dyspnoea on exertion | -168
bilateral lower extremity oedema | -168
rhinorrhea | -168
fever | -168
systolic murmur | 0
heart failure exacerbation | 0
erythematous non-tender macules | 0
methicillin-resistant Staphylococcus aureus positive | 0
amphetamine and opiate IVDU | 0
diastolic heart failure with preserved ejection fraction | 0
coronary artery disease | 0
coronary artery bypass graft | 0
aortic stenosis | 0
aortic valve replacement | 0
aortic valve thrombosis | 0
bioprosthetic valve replacement | 0
sick sinus syndrome | 0
dual-chamber pacemaker | 0
atrial fibrillation | 0
diabetes mellitus | 0
hypertension | 0
post-traumatic stress disorder | 0
chronic back pain | 0
septic shock | 72
broad-spectrum antibiotics | 72
vasopressors | 72
methicillin-susceptible Staphylococcus aureus | 120
C-reactive protein elevated | 120
white blood cell count elevated | 120
computed tomography of the head | 120
blood cultures | 120
intravenous antibiotics | 120
vancomycin | 120
rifampin | 120
gentamicin | 120
piperacillin-tazobactam | 120
transoesophageal echocardiogram | 192
three-valve endocarditis | 192
aortic root abscess | 192
pacemaker lead infection | 192
cardiovascular and thoracic surgery service evaluation | 192
hospice care | 216
expired | 336 
septic shock | 336
disseminated intravascular coagulation | 336