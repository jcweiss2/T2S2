22 years old | 0
male | 0
gastroesophageal reflux disease | 0
cholecystectomy | -17520
omeprazole | -17520
esophageal dysphagia | -17520
EGD | 0
propofol | 0
mild esophageal stricture | 0
esophageal mucosal changes | 0
ringed esophagus | 0
feline appearance | 0
longitudinal furrows | 0
eosinophilic esophagitis | 0
severe epigastric pain | 1.5
emesis | 1.5
elevated lipase | 1.5
leukocytosis | 1.5
normal triglycerides | 1.5
peripancreatic fluid | 1.5
hypoxia | 24
hemodynamic instability | 24
acute hypoxic respiratory failure | 24
ARDS | 24
septic shock | 24
pleural effusion | 24
acute kidney injury | 24
pancreatic necrosis | 240
retroperitoneal fluid collection | 240
ischemic colitis | 240
subtotal colectomy | 240
multiorgan failure | 24
intensive care admission | 24
vasopressor support | 24
broad-spectrum antibiotics | 24
antifungal agents | 24
thoracentesis | 24
chest tube placement | 24
percutaneous drain placement | 240
pancreatic necrosectomy | 240
prolonged hospitalization | 4320
rehabilitation | 4320
propofol-induced pancreatitis | 1.5
severe necrotizing pancreatitis | 1.5
no gallstone pancreatitis | 1.5
no alcohol use | 1.5
negative infectious workup | 1.5
negative autoimmune etiology | 1.5
normal serum triglyceride | 1.5
no trauma or toxin exposure | 1.5
negative cystic fibrosis | 1.5
negative myotonic dystrophy | 1.5
no vasculitis | 1.5
no drug allergies | 1.5
