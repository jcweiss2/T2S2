54 years old | 0
female | 0
admitted to the Emergency Department | 0
syncope | 0
hematemesis | 0
smoking habit | 0
alcohol consumption |.0
hemodynamically stable | 0
asymptomatic | 0
hemoglobin 10.2 mg/dl | 0
cranial CT scan | 0
initial EGD | 0
hiatal hernia | 0
no active bleeding | 0
in-hospital observation | 0
hemodynamic instability | -72
melenae | -72
hemoglobin stable | -72
EGD after 48 hours | 48
discharged | 72
readmitted | 120
syncope | 120
hypotension | 120
heart rate 92 bpm | 120
fluid replacement | 120
hemodynamic stability | 120
hemoglobin 8.4 mg/dl | 120
transfusion of 2 units PRBC | 120
melenae | 120
EGD pulsatile vessel | 120
aortic aneurysm | 120
duodenal AEF | 120
mural thrombus | 120
urgent laparotomy | 120
ligation of iliac arteries | 120
axilo-bifemoral bypass | 120
resection of fistula | 120
primary suture repair | 120
vasoactive drugs | 120
transfusion of 5 units PRBC | 120
admitted to ICU | 120
hemodynamically stable | 126
asymptomatic | 126
transferred to ward | 144
discharged | 264
stable hemoglobin | 264
no active bleeding | 264
pathology report | 264
gram positive aerobic flora | 264
Streptococcus viridians | 264
coagulase-negative Staphyloccocus | 264
Piperacillin/Tazobactam | 264
follow-up CT scan | 1080
no recurrent AEF | 1080
no further gastrointestinal bleeding | 1080
