26 years old | 0
female | 0
otherwise healthy | 0
referred to the department | 0
rising levels of human chorionic gonadotropin | 0
intermittent vaginal bleeding | 0
6 weeks after a legal medical abortion | -1008
intrauterine pregnancy | -1008
vaginal ultrasound scan | 0
placental remnants in the uterus | 0
surgical evacuation of the uterus | 0
discharged | 12
readmitted | 24
temperature of 39.5°C | 24
abdominal pain | 24
severe endometritis | 24
metronidazole administered | 24
benzylpenicillin administered | 24
gentamicin administered | 24
deteriorated | 48
saturation fell to 90% | 48
respiratory rate rose to around 40 breaths per minute | 48
oxygen given by mask | 48
temperature peaked at 40.7°C | 48
C-reactive protein rose to around 300 mg/L | 48
leukocytes to around 15 × 10^9/L | 48
moved to the intensive care unit | 48
intubated | 48
CT scan performed | 48
thrombophlebitis of the internal jugular vein | 48
hepatomegaly | 48
diagnosed with Lemierre's syndrome | 48
benzylpenicillin discontinued | 48
gentamicin discontinued | 48
tazocin administered | 48
clindamycin administered | 48
metronidazole continued | 48
heparin injections | 48
recovered | 360
discharged | 504
infection with F. necrophorum | 48
blood cultures showed infection with F. necrophorum | 48
F. necrophorum cultivated from the patient's cervix | 48
infection originated from the cervix | 48
no symptoms from the oropharyngeal tract | 0