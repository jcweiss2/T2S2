72 years old | 0
female | 0
known diabetic | -5760
admitted to the hospital | 0
unconsciousness | -12
poor glycemic control | 0
hypertensive | 0
on oral hypoglycemic drugs | -5760
on medication for hypertension | -5760
no history of convulsions | 0
no history of fever | 0
no history of vomiting | 0
no history of headache | 0
no history of trauma | 0
no neurodeficit | 0
Glasgow Coma scale 5/15 | 0
pulse 88/min | 0
blood pressure 140/80 mm Hg | 0
respiratory rate 16/min | 0
irregular bilateral vesicular breath sounds | 0
capillary blood glucose 28 mg/dL | 0
Total leukocyte count 16,200/mm3 | 0
neutrophil predominance | 0
serum alanine aminotransferase 31 IU/mL | 0
serum aspartate aminotransferase 71 IU/mL | 0
alkaline phosphatase 22 IU/L | 0
total protein 4.8 g/dL | 0
albumin 2.4 g/dL | 0
urea 54 mg/dL | 0
creatinine 1.2 mg/dL | 0
total bilirubin 0.6 mg/dL | 0
conjugated bilirubin 0.3 mg/dL | 0
focal ischemia on CT scan | 0
hypoglycemic encephalopathy | 0
hypoxic brain damage | 0
intubated | 0
ventilator support | 0
piperacillin + tazobactam | 0
uncontrolled blood sugar | 72
fluctuating blood sugar | 72
low grade fever | 72
endotracheal secretions sent for culture | 72
Acinetobacter baumanii isolated | 96
sensitive to netilmicin | 96
sensitive to polymixin B | 96
netilmicin started | 96
cefepime started | 96
high grade fever | 168
total leukocyte count 8400/mm3 | 168
neutrophilic predominance | 168
serum creatinine 2 mg/dL | 168
catheterized urine sample sent for culture | 168
blood sent for culture | 168
Escherichia coli isolated | 168
sensitive to meropenem | 168
sensitive to poymyxin B | 168
sensitive to cotrimoxazole | 168
sensitive to nitrofurantoin | 168
meropenem added to treatment | 168
general condition deteriorated | 168
total leukocyte counts dropped to 4000/mm3 | 168
E. faecium isolated from blood | 168
E. faecium resistant to linezolid | 168
MIC of E. faecium > 256 μg/mL | 168
MIC of E. faecium 1024 μg/mL | 168
vancomycin started | 192
condition further deteriorated | 360
declared dead | 360