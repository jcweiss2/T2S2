41 years old | 0
male | 0
admitted to the hospital | 0
fever | -72
fatigue | -72
weight loss | -72
disseminated skin lesions | -72
low urine output | -72
mental confusion | -72
thoracic herpes zoster | -504
HIV infection | -504
diagnosed with HIV | -504
decided not to initiate antiretroviral therapy | -504
afebrile | 0
dehydrated | 0
blood pressure 109/72 mmHg | 0
pulse rate 130 beats/min | 0
oxygen saturation 97% | 0
mental confusion | 0
Glasgow Coma Scale 14 | 0
lung sounds clear | 0
abdomen innocent | 0
no peripheral lymphadenopathy | 0
diffuse maculopapular and crusty skin lesions | 0
hemoglobin 13.9 g/dL | 0
white blood cell count 6,500/mm3 | 0
platelet count 82,000/mm3 | 0
C-reactive protein 26.1 mg/dL | 0
creatinine level 4.0 mg/dL | 0
sodium concentration 127 mg/dL | 0
lactate dehydrogenase 5,782 U/L | 0
aspartate aminotransferase 342 U/L | 0
alanine aminotransferase 340 U/L | 0
total bilirubin 3.9 mg/dL | 0
direct bilirubin 3.4 mg/dL | 0
international normalized ratio 1.71 | 0
triglycerides 324 mg/dL | 0
ferritin > 100,000 ng/mL | 0
serologic diagnosis of HIV-1 infection | 0
CD4 count 4 cells/mm3 | 0
HIV-1 viral load 1,749,163 copies/mL | 0
chest computed tomography unspecific | 0
brain CT scan normal | 0
cerebrospinal fluid normal | 0
abdominal CT scan no hepatosplenomegaly | 0
retroperitoneal, periaortic, and interaortocaval lymph node enlargement | 0
sequential organ failure assessment score 8 | 0
septic shock | 0
multiorgan dysfunction | 0
acute renal failure | 0
metabolic acidosis | 0
hepatic failure | 0
coagulopathy | 0
volemic expansion initiated | 0
ceftriaxone administered | 0
yeasts suggestive of Histoplasma spp. | 0
transferred to the ICU | 24
supplemental oxygen | 24
amphotericin B deoxycholate initiated | 24
reduced level of consciousness | 48
Glasgow Coma Scale 10 | 48
refractory septic shock | 48
high doses of vasopressors | 48
corticosteroids | 48
mechanical ventilation | 48
hemodialysis | 48
yeasts suggestive of Histoplasma spp. in bone marrow | 72
yeasts suggestive of Histoplasma spp. in skin samples | 168
hemophagocytosis not observed | 72
Histoplasma spp. cultures positive | 336
antiretroviral therapy initiated | 240
discharged from the hospital | 768
follow-up in the outpatient clinic | 768
creatinine level 1.3 mg/dL | 2304
CD4 count 180 cells/mm3 | 2304
HIV-1 viral load < 40 copies/mL | 2304
darunavir/ritonavir | 2304
dolutegravir | 2304
lamivudine | 2304
prophylactic trimethoprim-sulfamethoxazole | 2304
itraconazole | 2304