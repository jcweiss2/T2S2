38 years old | 0
male | 0
admitted to the hospital | 0
fever | 0
cough | 0
shortness of breath | 0
myalgia | 0
BMI 29.9 | 0
history of daily vaping | 0
CT angiogram | 0
no pulmonary embolism | 0
bilateral numerous multifocal ground glass opacities | 0
SARS COV2 PCR nasopharyngeal swab test | 0
COVID-19 positive | 0
droplet precautions | 0
contact isolation | 0
blood and sputum culture | 0
urine/sputum legionella testing | 0
mycoplasma IGM tests | 0
negative results | 0
subcutaneous Heparin | 0
elevated D-dimer | 0
intubated | 120
acute hypoxemic respiratory failure | 120
admitted to the intensive care unit | 120
Plaquenil | 120
supplemental oxygen | 120
albuterol sulfate | 120
tiotropium bromide | 120
Tocilizumab | 120
Zithromax | 120
multi organ failure | 144
acute renal failure | 144
sepsis | 816
toxic metabolic encephalopathy | 936
low white blood cell | 0
normal red blood cell | 0
high platelet | 0
high neutrophil percentage | 0
low lymphocyte percentage | 0
high C-reactive protein | 24
high creatinine | 24
high PTT | 24
high fibrinogen | 24
high pro-calcitonin | 24
high lactate dehydrogenase | 24
high alanine aminotransferase | 24
high aspartate aminotransferase | 24
low calcium | 24
high potassium | 240
high glucose | 240
insulin therapy | 240
continuous veno-venous hemofiltration | 240
intermittent hemodialysis | 240
high troponin-I | 240
high creatinine kinase | 240
anemic | 240
transfused | 240
Hemophagocytic lymphohistiocytosis syndrome | 480
toxic metabolic encephalopathy | 480
normal head CT | 480
second CT scan of the chest | 1104
scattered centrilobular ground glass opacities | 1104
new right hydropneumothorax | 1104
bilateral lower lobe consolidations | 1104
thick-walled cavity | 1104
superimposed E faecalis bacterial infection | 1104
pulmonary hypertension | 1104
high attenuation foci | 1104
bilateral symmetrical muscle calcification | 1104
rhabdomyolysis | 1104
discharge arrangements | 2160