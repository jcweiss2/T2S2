38 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
HBV-associated PAN | -156 | 0 | Factual
acute abdomen | 0 | 0 | Factual
septic shock | 0 | 0 | Factual
prednisolone | -4320 | 0 | Factual
cyclophosphamide | -4320 | 0 | Factual
Tenofovir | -4320 | -144 | Factual
chronic renal failure | -156 | 0 | Factual
diabetes mellitus Type II | -156 | 0 | Factual
free sub diaphragmatic air | 0 | 0 | Factual
peritonitis | 0 | 0 | Factual
three perforations of the small intestine | 0 | 0 | Factual
segmental enterectomy with anastomosis | 0 | 0 | Factual
mechanical ventilation | 0 | 72 | Factual
circulatory support | 0 | 72 | Factual
acute-on-chronic renal failure | 0 | 72 | Factual
weaned off the ventilator | 72 | 72 | Factual
haemodynamically stable | 72 | 168 | Factual
tenofovir orally | 72 | 168 | Factual
IV methylprednisolone | 72 | 168 | Factual
abdominal drain catheter presented enteric content | 168 | 168 | Factual
second explorative laparotomy | 168 | 168 | Factual
two new perforations | 168 | 168 | Factual
multiple areas of patchy necrosis | 168 | 168 | Factual
plasma exchanges | 168 | 360 | Factual
IV cyclophosphamide | 168 | 168 | Factual
IV methylprednisolone | 168 | 192 | Factual
IV prednisone | 192 | 360 | Factual
third laparotomy | 240 | 240 | Factual
three new necrotic lesions | 240 | 240 | Factual
necrotic lesion on the left lobe of the liver | 240 | 240 | Factual
fourth laparotomy | 336 | 336 | Factual
segmental enterectomy with anastomosis | 336 | 336 | Factual
cholecystectomy | 336 | 336 | Factual
anastomotic leak | 336 | 336 | Factual
gangrenous gallbladder | 336 | 336 | Factual
septic shock | 360 | 360 | Factual
multiple organ failure | 360 | 360 | Factual
death | 360 | 360 | Factual
weight loss | -8760 | -156 | Factual
myalgias | -8760 | -156 | Factual
fever | -8760 | -156 | Factual
skin erythema | -8760 | -156 | Factual
deterioration of renal function | -8760 | -156 | Factual
new onset of diabetes mellitus Type II | -8760 | -156 | Factual
hypertension | -8760 | -156 | Factual
HBsAg | 0 | 0 | Factual
HBeAg | 0 | 0 | Factual
Anti-HBcAb | 0 | 0 | Factual
absence of Anti-HBsAb | 0 | 0 | Factual
absence of Anti-HBeAb | 0 | 0 | Factual