76 years old | 0
male | 0
admitted to the hospital | 0
severe hyponatremia | 0
pancreatic adenocarcinoma | -672
metastasis to the liver | -672
diastolic heart failure | -672
atrial fibrillation | -672
coronary artery disease | -672
port placement for chemotherapy | -672
routine preoperative evaluation | -672
sodium level of 116 mmol/L | -672
pneumonia | -672
x-ray findings | -672
broad-spectrum antibiotics | -672
fluid for hyponatremia | -672
transferred to the intensive care unit | -672
jugular vein distention | -672
lower extremity pitting edema | -672
transthoracic echocardiogram | -672
normal left ventricular cavity size | -672
mildly reduced systolic function | -672
septal flattening | -672
left atrial enlargement | -672
suspected MV vegetation | -672
severe mitral regurgitation | -672
tricuspid regurgitation Doppler | -672
elevated RV systolic pressure | -672
type 2 and type 3 pulmonary arterial hypertension | -672
ill-defined thickening in the TV leaflets | -672
afebrile | -672
leukocytosis | -672
recent urethral instrumentation | -672
blood cultures | -672
consulted infectious disease specialist | -672
broad-spectrum antibiotics | -672
infective endocarditis | -672
day 1 | -672
valvular vegetations via echocardiography | -672
tricuspid valve (TV) and mitral valve (MV) | -672
transesophageal echocardiogram (TEE) | -24
normal left ventricular size and function | -24
normal RV size and function | -24
hypermobile interatrial septum | -24
no left atrial or left atrial appendage thrombus | -24
2 large vegetations on the atrial aspect of MV leaflets | -24
severe mitral regurgitation | -24
tricuspid regurgitation | -24
RVSP 47 mm Hg | -24
negative blood cultures | -24
polymerase chain reaction testing | -24
Coxiella urnetiid | -24
Legionella spp | -24
Brucella spp | -24
antiphospholipid syndrome | -24
discontinued apixaban | -24
low molecular weight heparin or unfractionated heparin | -24
computed tomography imaging of the head | -24
intracerebral hemorrhage | -24
observation of clinic course | -24
enoxaparin | -24
platelets recovered to above 50,000 10^9/L | -24
nonbacterial thrombotic endocarditis (NBTE) | -24
advanced malignancy | -24
systemic lupus erythematosus | -24
antiphospholipid syndrome | -24
rheumatoid arthritis | -24
sepsis | -24
burns | -24
echocardiogram | -24
infectious endocarditis | -24
valvular destruction | -24
unfractionated heparin | -24
vitamin K antagonists | -24
warfarin | -24
surgical intervention | -24
heart failure | -24
acute valve rupture | -24
prevention of recurrent embolization | -24
bivalvular involvement | -24
valvular dysfunction | -24
valvular regurgitation | -24
anticoagulation | -24
resolution of valvular dysfunction | -24
advanced pancreatic malignancy | -24
outpatient follow-up | -24
death | -24