39 years old | 0\
female | 0\
palpable mass on her right breast | 0\
Hodgkin lymphoma | -192 months\
chemotherapy | -192 months\
mantle field radiation | -192 months\
inflammatory colitis | -216 months\
mesalazine | -12 months\
invasive ductal carcinoma | 0\
triple-negative phenotype | 0\
MIB1 85% | 0\
neoadjuvant chemotherapy | 0\
paclitaxel | 0\
carboplatin | 0\
port-à-cath insertion | 48\
fever | 72\
subcutaneous cellulitis | 72\
colliquative necrosis | 72\
elevated white blood cell count | 72\
neutrophilia | 72\
elevated C-reactive protein | 72\
broad-spectrum i.v. antibiotic therapy | 72\
piperacillin/tazobactam | 72\
daptomycin | 72\
PORT rimotion | 72\
necrosectomy | 72\
defervescence | 96\
improvement in subcutaneous cellulitis | 96\
improvement in blood works | 96\
febrile seizure | 120\
WBC rise | 120\
worsening of skin lesion | 120\
second necrosectomy | 120\
peripheral blood cultures negative | 120\
skin plug negative | 120\
i.v. catheter tip positivity for Klebsiella pneumoniae | 120\
meropenem | 120\
levofloxacin | 120\
mediastinitis | 120\
bilateral pleural effusion | 120\
left pulmonary atelectasis | 120\
thoracoscopy | 120\
pleural and mediastinal drainage | 120\
sepsis | 120\
broad-spectrum antibiotic and antifungal therapy | 120\
hemodynamic support | 120\
non-invasive ventilation | 120\
intensive inflammatory infiltrate | 120\
neutrophils | 120\
systemic methylprednisolone | 120\
topical cyclosporine | 120\
progressive resolution of mediastinitis | 168\
progressive resolution of pleural effusion | 168\
wound improvement | 168\
scar | 168\
progressive normalization of blood count | 168\
progressive normalization of flogosis index | 168\
breast ultrasound | 168\
right mastectomy | 168\
axillary dissection | 168\
breast surgical wound healing | 168\
fibroelastosis | 168\
chronic inflammation | 168\
isolated neoplastic cells | 168\
negative axillary nodes | 168\
negative restaging brain/chest/abdomen CT | 168\
negative BRCA mutation test | 168\
negative p53 mutation test | 168\
autologous skin graft | 336\
PICC implant | 336\
chemotherapy with carboplatin and paclitaxel | 336\
dose reduction | 336\
completion of chemotherapy | 504\
follow-up | 504