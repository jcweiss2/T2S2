27 years old|0
male|0
presented at the emergency department|0
massive hemorrhage from the tracheostomy tube|0
multiple traumas due to a car accident|-5760
neck fracture|-5760
quadriplegic|-5760
operated (neck fracture)|-5760
nasogastric tube inserted|-5760
discharge of food from the foramen of tracheostomy tube after oral feeding|-5760
massive bleeding from tracheostomy stoma|0
vital signs became unstable|0
blood pressure below 80/60|0
peripheral pulse not palpable|0
urgent surgery performed|0
general anesthesia|0
rigid bronchoscopy performed|0
tracheal stenosis below the vocal cords|0
unclear view of trachea|0
tracheoesophageal fistula (TEF)|0
TEF located in membranous part of trachea|0
bleeding stopped during operation|0
pressure of tracheostomy cuff|0
dissection of tracheostomy stoma|0
division and ligature of innominate artery|0
separation of trachea from the divided artery|0
repair of tracheal defect|0
reinforcement with strap muscle|0
reinsertion of tracheostomy tube|0
insertion of jejunostomy tube due to TEF|0
vital signs stabilized post-operation|0
neurologic examination unchanged post-operation|0
weaker right radial pulse|0
discharged from hospital|312
readmitted for TEF repair|1752
endoscopy performed|1752
large foramen in anterior wall of esophagus|1752
deep vein thrombosis in left leg|1752
progression to inferior vena cava|1752
heparin administered|1752
colored Doppler sonography after 7 days|1752
deep vein thrombosis resolved|1752
severe purulent discharge from tracheostomy tube|1752
chest X-ray showed bronchiectasis|1752
chest X-ray showed pneumonia|1752
antibiotic treatment based on culture|1752
gradual deterioration|1752
septic shock|1752
unresponsive to medical treatment|1752
patient expired|1104
