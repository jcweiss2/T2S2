newborn female | 0
born at 24 weeks + 3 days | 0
breech presentation | 0
cord prolapse | 0
birth weight of 645 g | 0
HIV negative mother | 0
Apgar score of 4 | 0
Apgar score of 8 | 5
mechanical ventilation | 0
central umbilical catheters | 0
total parenteral nutrition | 0
empiric antibiotics | 0
skin sensors | 0
late-onset sepsis | 216
Escherichia coli bacteremia | 216
antimicrobial therapy with cefepime | 216
adhesive patch removal | 480
skin abrasion | 480
erythema | 480
induration | 480
plaque with necrotic center | 480
ulcer | 528
subcutaneous cell tissue extension | 528
necrotic area progression | 528
intensive treatment by wound care team | 480
thermic instability | 528
metabolic acidosis | 528
hyperglycemia | 528
hypotension | 528
cutaneous mucormicosis suspicion | 528
skin biopsy | 528
empiric antifungal treatment with liposomal amphotericin B | 528
fungal biomarkers | 528
refractory shock | 552
renal failure | 552
death | 564
fungal cultures | 528
Rhizopus spp. | 528
histopathology report | 528
broad aseptate hyphae | 528
Mucorales | 528
mass spectroscopy | 528
polymerase chain reaction | 528
Rhizopus arrhizus | 528
fungal blood cultures | 528 
negative fungal blood cultures | 528