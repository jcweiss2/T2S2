27 years old | 0
male | 0
admitted to the hospital | 0
pancytopenia | 0
neutrophils: 0.8×10^9/L | 0
hemoglobin: 9.4 gr/dl | 0
platelets: 4×10^9/L | 0
muco-cutaneous hemorrhages | 0
marrow aspiration | 0
trephine biopsy | 0
diagnosis of idiopathic severe aplastic anemia | 0
empirical broad spectrum antibiotherapy | 5
piperacillin–tazobactam | 5
amikacin | 5
febrile neutropenia | 5
fever resolved | 10
neutropenia worsened | 10
neutrophils: 0.3×10^9/L | 10
oral prednisone | 12
admitted to the intensive care unit (ICU) | 19
septic shock | 19
piperacillin-tazobactam restarted | 20
levofloxacin | 20
blood cultures returned positive for Streptococcus mitis | 20
blood cultures returned positive for Klebsiella pneumoniae | 20
patient recovered | 24
admitted to the hematology unit | 24
central venous catheter (CVC) inserted | 25
fever reappeared | 29
piperacillin–tazobactam and levofloxacin replaced by meropenem | 29
antifungal treatment by caspofungin | 29
fever persisted | 29
poor clinical condition | 29
diarrhea | 29
abdominal pain | 29
dry cough | 29
left thoracic pain | 29
peripheral and central venous blood cultures performed | 29
caspofungin replaced by liposomal amphotericin B | 31
voriconazole | 31
stool examination revealed rare colonies of S. clavata | 31
CT scan revealed a left pulmonary nodular lesion | 31
diffuse bowel thickening | 31
multiple nodular lesions of spleen, kidneys, and liver | 31
liver function tests were normal | 31
CVC removed | 31
left blurred vision | 31
cerebral CT scan and magnetic resonance imaging were normal | 31
ophtalmological examination revealed a left retinal hemorrhage | 31
echocardiogram excluded the diagnosis of fungal endocarditis | 31
patient remained severely neutropenic | 31
S. clavata identified from the first blood culture | 33
clinical condition rapidly improved | 33
daily blood cultures returned positive for S. clavata until day 34 | 33
weekly stool examinations and daily blood cultures returned negative | 34
fever persisted until day 42 | 42
weekly galactomannan antigenemia results were negative | 42
voriconazole blood levels were weekly checked | 42
antifungal susceptibility testing | 42
patient underwent a sibling allogeneic bone marrow transplantation | 42
conditioning regimen combining IV cyclophosphamide | 35
IV fludarabine | 35
IV alemtuzumab | 36
cyclosporine started | 41
granulocyte transfusions | 39
granulocyte transfusions | 40
granulocyte transfusions | 41
granulocyte transfusions | 48
granulocyte transfusions | 49
neutrophil counts reached 0.5 to 1×10^9 /L | 39
neutrophil counts returned below 0.1×10^9/L | 40
neutrophil counts reached 0.5×10^9/L | 68
voriconazole replaced by posaconazole | 84
liposomal amphotericine B discontinued | 84
abdominal ultrasound showed only small splenic residual lesions | 84
patient left the unit | 88
fever did not recur | 88
left vision progressively normalized | 88
no recurrence of infection or complication of transplantation | 120