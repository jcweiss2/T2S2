27 years old | 0
    man | 0
    mitochondrial neurogastrointestinal encephalopathy disease | 0
    central catheter line peripherally inserted | 0
    jejunal diverticulosis | 0
    partial small bowel resection | 0
    insulin-dependent type I diabetes mellitus | 0
    presented with fever | 0
    presented with vomiting | 0
    presented with abdominal pain | 0
    core temperature of 38.5°C | 0
    heart rate of 120 beat/min | 0
    blood pressure of 120/70 mmHg | 0
    rapid heart sounds | 0
    regular heart sounds | 0
    no additional heart sounds | 0
    no murmurs | 0
    no lung abnormalities | 0
    mild abdominal tenderness | 0
    no guarding | 0
    functioning percutaneous endoscopic gastrostomy | 0
    no signs of infection at gastrostomy | 0
    marked redness around central catheter line | 0
    pussy secretion around central catheter line | 0
    no stigmata of endocarditis | 0
    leukocytosis | 0
    C-reactive protein 25 mg/dL | 0
    acute kidney injury | 0
    creatinine 1.3 mg/dL | 0
    urea 50 mg/dL | 0
    diabetic ketoacidosis | 0
    serum glucose level 420 mg/dL | 0
    positive ketones in peripheral blood | 0
    metabolic acidosis | 0
    pH 7.2 | 0
    pCO2 32 mmHg | 0
    HCO3 11 mmHg |$