35 years old | 0
female | 0
gave birth to healthy twins | 0
cesarean section | 0
threatened preterm delivery | 0
first pregnancy | 0
in vitro fertilization | 0
facial nerve paresis | 0
no hypertension | 0
no cardiac diseases | 0
no vision abnormalities | 0
no seizures | 0
severe headache | 0
generalized tonic-clonic seizures | 0
loss of consciousness | 0
arterial blood pressure 195/110 mmHg | 0
heart rate 120 beats/min | 0
diagnosis of eclampsia | 0
transferred to intensive care unit | 0
antihypertensive therapy | 0
intravenous magnesium sulphate | 0
ebrantil | 0
20% manitol | 0
oral diazepam | 0
bilateral vision loss | 0
complete blood count normal | 0
liver function tests normal | 0
clotting parameters normal | 0
electrocardiogram normal | 0
proteinuria 2+ | 0
other system examinations normal | 0
seizures not repeated | 24
headache alleviated | 24
bilateral loss of vision | 0
light perception | 0
normal pupillary responses | 0
normal fundus findings | 0
diagnosis of cortical blindness | 0
mild right-sided facial nerve paresis | 0
no other neurological disorders | 0
MSCT scan hypodensity posterior white matter | 0
MRI T2 hyperintense signals | 0
MRI FLAIR hyperintense signals | 0
vasogenic edema | 0
PRES diagnosis | 0
blood pressure stabilized | 24
oral enalapril maleate | 24
oral methyldopa | 24
IV human albumin | 24
bilateral improvement of visual function | 120
best-corrected visual acuity 1.0 | 120
normal anterior eye segment | 120
normal fundus | 120
peripheral relative scotoma | 120
depressed sensitivity paracentral left visual field | 120
right-sided partial facial nerve paresis | 120
MRI regression of edema | 192
discrete residual changes posterior horns | 192
discharged | 216
oral antihypertensive therapy | 216
physical therapy for facial nerve paresis | 216
hypertension | 0
proteinuria | 0
PET | 0
eclampsia | 0
cortical blindness | 0
PRES | 0
status epilepticus | 0
intracranial hemorrhage | 0
cerebral ischemia | 0
neurological deficits | 0
complications | 0
seizures | 0
vision loss | 0
headache | 0
blood pressure elevation | 0
MSCT findings | 0
MRI findings | 0
antihypertensive treatment | 0
magnesium sulphate | 0
manitol | 0
diazepam | 0
enalapril | 0
methyldopa | 0
human albumin | 0
physical therapy | 0
visual improvement | 120
edema regression | 192
residual changes | 192
discharge | 216
oral enalapril continuation | 216
physical therapy continuation | 216
