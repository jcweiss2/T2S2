42 years old | 0
male | 0
hypertension | 0
shortness of breath | -120
subjective fever | -120
chills | -120
occasional cough productive of clear sputum | -120
generalized bone pain | -120
intermittent headache | -120
watery diarrhea | -120
anorexia | -120
home temperature recording of 105 °F | -120
no chest pain | -120
no abdominal pain | -120
no numbness | -120
no tingling | -120
no weakness | -120
no history of pulmonary embolism | -120
no history of deep vein thrombosis | -120
no recent travel | -120
denied use of tobacco | -120
denied use of drugs | -120
temperature: 38.6 °C | 0
heart rate: 109 beats per minute | 0
respiratory rate 39 breaths per minute | 0
SpO2: 57 | 0
blood pressure: 132/66 mm Hg | 0
dyspneic | 0
unable to speak in full sentences | 0
breath sounds equal | 0
symmetrical chest wall expansion | 0
regular rhythm | 0
strong and symmetrical peripheral pulses | 0
alert | 0
oriented | 0
no focal neurological deficits | 0
chest X-ray revealed scattered bilateral airspace opacities | 0
sodium: 120 mEq/L (L) | 0
potassium: 4 mEq/L | 0
blood urea nitrogen: 21 mg/dL (H) | 0
creatinine: 1.1 mg/dL (H) | 0
white blood cell: 13 900/µL (H) | 0
neutrophil %: 89.4 (H) | 0
lymphocyte %: 5.5 (L) | 0
hemoglobin: 13.3 g/dL | 0
platelets: 250 000/µL | 0
Dimer 2.74 (H) | 0
C-reactive protein: 29.32 mg/dL (H) | 0
ferritin: 826.30 ng/mL (H) | 0
lactate dehydrogenase: 1883 U/L (H) | 0
interleukin-6: 224.35 pg/mL (H) | 0
troponin <0.019 (ng/mL) | 0
RT-PCR positive for COVID | 0
managed on nonrebreather mask | 0
managed on nasal cannula | 0
received ceftriaxone | 0
received azithromycin | 0
received hydroxychloroquine | 0
received tocilizumab | 0
enrolled in remdesivir trial | 0
severe hypoxia on day 2 | 48
oxygen saturation in 60s | 48
removed non-rebreather mask | 48
rapidly intubated | 48
hypotension post-intubation | 48
vasopressor therapy | 48
no overt shock | 48
lactate remained below 2.5 | 48
serum creatinine remained below 0.8 mg/dL | 48
troponinemia worsened (0.194-0.682 ng/mL) | 48
concern for acute PE | 48
heparin drip initiated | 48
fluctuating hypoxia on ventilation | 48
receiving heparin (intravenous) | 48
receiving sedatives | 48
receiving occasionally paralytics | 48
continuously febrile | 48
required pressor support | 48
suboptimal blood pressures | 48
duplex study revealed no deep vein thrombosis | 48
transthoracic echocardiography without intracavitary thrombus | 48
diminished pupillary reflexes | 144
mid-dilated pupils | 144
no corneal reflexes | 144
no oculocephalic reflexes | 144
persisted after withdrawing sedation | 144
CT head revealed large ischemic infarcts | 144
CT chest with angiography disclosed multifocal dense ground-glass opacities | 144
no PE | 144
clinical deterioration | 144
no further workup | 144
pronounced dead | 168
