33 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
nausea | -24 | 0 | Factual
vomiting | -24 | 0 | Factual
abdominal pain | -24 | 0 | Factual
discharged | -36 | -36 | Factual
hospitalized | -36 | -36 | Factual
recurrent pericarditis | -36 | -36 | Factual
colchicine | -36 | -12 | Factual
febrile | 0 | 0 | Factual
hypotensive | 0 | 0 | Factual
leukocytosis | 0 | 0 | Factual
elevated serum lactate | 0 | 0 | Factual
acute kidney injury | 0 | 0 | Factual
acute transaminitis | 0 | 0 | Factual
severe coagulopathy | 0 | 0 | Factual
normal serum troponin | 0 | 0 | Factual
negative toxicology screen | 0 | 0 | Factual
normal sinus rhythm | 0 | 0 | Factual
normal biventricular function | 0 | 0 | Factual
no valvular disease | 0 | 0 | Factual
no pericardial effusion | 0 | 0 | Factual
sepsis suspected | 0 | 0 | Possible
fluid resuscitation | 0 | 24 | Factual
broad-spectrum antibiotics | 0 | 24 | Factual
vasopressor therapy | 0 | 24 | Factual
multisystem organ failure | 24 | 24 | Factual
intubated | 24 | 24 | Factual
paralyzed | 24 | 24 | Factual
intravascular volume repletion | 24 | 48 | Factual
intravenous vasopressors | 24 | 48 | Factual
stress-dose steroids | 24 | 48 | Factual
high-dose vitamin B12 | 24 | 48 | Factual
Swan-Ganz catheter | 24 | 24 | Factual
distributive shock | 24 | 24 | Factual
cardiac output | 24 | 24 | Factual
pulmonary artery diastolic pressure | 24 | 24 | Factual
systemic vascular resistance | 24 | 24 | Factual
cardiogenic shock | 48 | 48 | Factual
high filling pressures | 48 | 48 | Factual
low cardiac output | 48 | 48 | Factual
high systemic vascular resistance | 48 | 48 | Factual
elevated troponin | 48 | 48 | Factual
severe biventricular failure | 48 | 48 | Factual
left ventricular ejection fraction | 48 | 48 | Factual
intravenous milrinone | 48 | 72 | Factual
continuous renal replacement therapy | 48 | 72 | Factual
anuric renal failure | 48 | 72 | Factual
PRBC transfusion | 48 | 48 | Factual
normalized cardiac output | 72 | 72 | Factual
decreased troponin | 72 | 72 | Factual
improved multisystem organ failure | 72 | 72 | Factual
neutropenia | 96 | 96 | Factual
recovered left ventricular ejection fraction | 144 | 144 | Factual
weaned from vasopressors | 240 | 240 | Factual
taken off CRRT | 240 | 240 | Factual
extubated | 312 | 312 | Factual
hair loss | 576 | 576 | Factual
admitted to taking colchicine | 576 | 576 | Factual
elevated serum colchicine | 30 | 30 | Factual
elevated whole blood colchicine | 14 | 14 | Factual
hypertension | -36 | 0 | Factual
pulmonary emboli | -36 | 0 | Factual
polysubstance abuse | -36 | 0 | Factual
discharged | 720 | 720 | Factual