13 years old | 0
female | 0
admitted to the hospital | 0
difficult-to-control seizures | 0
worsening of handwriting | -72
involuntary, repetitive pill-rolling hand movements | -72
focal seizures | -72
GTCS | -72
facio-brachial dystonic seizures | -72
agitation | -72
unresponsiveness | -72
mutism | -72
lucid | -72
attempting to form words | -72
without speech production | -72
bruxism | -24
dystonic posturing | -24
full body rigidity | -24
opisthotonic posturing | -24
insomnia | -24
afraid | -24
agitated | -24
cried abnormally | -24
spontaneously | -24
brisk reflexes | -24
unsustained clonus | -24
bilateral | -24
waxy catatonia | -24
opsoclonus | -24
high-grade fever | 240
sensorium deteriorated | 240
orofacial dyskinesia | 240
autonomic instability | 240
irregular respiration | 240
sepsis | 240
urinary tract infection | 240
colitis | 240
mRS score 5 | 240
hemogram normal | 0
liver function tests normal | 0
renal function tests normal | 0
serum electrolytes normal | 0
thyroid function normal | 0
viral markers normal | 0
MRI Brain normal | 0
repeat MRI Brain normal | 336
EEG delta slowing | 0
left hemispheric regions | 0
CSF analysis normal | 0
cell count normal | 0
sugar normal | 0
protein normal | 0
Herpes Simplex negative | 0
Japanese Encephalitis negative | 0
ANA negative | 0
chest X-ray normal | 0
CECT abdomen normal | 0
thorax normal | 0
ultrasound pelvis normal | 0
skeletal survey normal | 0
tumor markers not done | 0
Acyclovir started | 0
AEDs started | 0
anti-NMDAR antibody detected | 240
methylprednisolone started | 240
intravenous immunoglobulins started | 240
oral prednisolone started | 240
symptoms improving | 480
mRS 4 | 672
AEDs tapered | 672
mRS 1 | 1152
amnesia | 1152
mild language disintegration | 1152
occasional agitation | 1152
follow-up advised | 1152
relapse after 8 years | -6720
subacute onset AED resistant seizures | -6720
abnormal behavior | -6720
abnormal body movements | -6720
routine investigations normal | -6720
CSF analysis unremarkable | -6720
MRI Brain normal | -6720
recovery after 3 months | -6390
fully functional | -6390