male | 0
2.98 kg | 0
born by emergency cesarean section | 0
bradycardia fetal distress | -1
gestational diabetes | -40
positive Group B streptococcus screen | -40
infection treatment | -40
sibling with undiagnosed skeletal dysplasia | -260
fetal anomaly scan | -10
bilateral bowing of the femur | -10
bilateral bowing of the tibia | -10
bilateral bowing of the fibula | -10
rocker-bottom feet | -10
mandible receding | -10
infant crying | 0
stable vital signs | 0
Apgar scores at 1 minute | 0
Apgar scores at 5 minutes | 5
dysmorphic features | 0
abnormal head trait | 0
micrognathia | 0
retrognathia | 0
short arms | 0
genu varum | 0
abnormally curved index | 0
camptodactyly | 0
pansystolic murmur | 0
grunting | 5
retractions | 5
fluctuating SpO2 | 5
respiratory distress | 5
nasal continuous positive airway pressure | 5
ground-glass opacity | 5
bilateral peribronchial cuffing | 5
bilateral pneumothorax | 10
hyperpyrexia | 10
mechanical ventilation | 10
nasogastric tube insertion | 10
inability to tolerate oral feeding | 10
hypertonic limbs | 10
fisting | 10
rhizomelia | 10
recurrent episodes of upper respiratory tract infections | 20
recurrent episodes of respiratory distress | 20
intolerance to oral feeding | 20
bronchoscopy | 20
laryngomalacia | 20
brain magnetic resonance imaging | 20
cranial ultrasound | 20
eye examination | 20
echocardiogram | 20
anterior muscular ventricular septal defect | 20
mild-to-moderate tricuspid regurgitation | 20
skeletal survey | 20
bilateral symmetric bowing of the femur | 20
bilateral symmetric bowing of the tibia | 20
diaphyseal cortical thickening | 20
skeletal dysplasia | 20
short stature | 20
severe joint contractures | 20
failure to thrive | 20
hypertonia | 20
swallowing difficulties | 20
genetic testing | 30
pathogenic variant in the LIFR gene | 30
c.1387_1390del p.(Asn463Phefs∗24) | 30
autosomal recessive SWS | 30
neonatal Schwartz-Jampel syndrome type 2 | 30
genetic counseling | 30
prenatal counseling | 30
gastrostomy tube insertion | 40
open Nissen fundoplication procedure | 40
pyloromyotomy | 40
discharge | 50
physiotherapy | 50
rehabilitation services | 50
dietary management | 50
recurrent episodes of chest infection | 100
respiratory distress | 100
fever | 1860
decreased activity | 1860
poor feeding | 1860
intubation | 1860
high frequency ventilation | 1860
inotropic support | 1860
antibiotics | 1860
multi-organ failure | 1860
septic shock | 1860
severe bronchopneumonia | 1860
acute respiratory distress syndrome | 1860
death | 1860