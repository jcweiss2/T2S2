65 years old | 0 | 0 
female | 0 | 0 
liver cirrhosis | -8760 | 0 
hepatocellular carcinoma | -8760 | 0 
scheduled for left lobe hepatectomy | 0 | 0 
administered intravenous glycopyrrolate | 0 | 0 
general anesthesia induced with propofol | 0 | 0 
general anesthesia induced with rocuronium | 0 | 0 
general anesthesia induced with remifentanil | 0 | 0 
general anesthesia maintained with sevoflurane | 0 | 300 
general anesthesia maintained with remifentanil | 0 | 300 
general anesthesia maintained with rocuronium | 0 | 300 
intubated and ventilated mechanically | 0 | 300 
monitored by electrocardiography | 0 | 300 
monitored by arterial blood pressure | 0 | 300 
monitored by central venous pressure | 0 | 300 
monitored by SpO2 | 0 | 300 
stable vital signs | 0 | 60 
sudden decrease in arterial blood pressure | 60 | 60 
sudden decrease in end-tidal carbon dioxide | 60 | 60 
sudden decrease in SpO2 | 60 | 60 
tachycardia | 60 | 60 
ST elevation on the EKG | 60 | 60 
resuscitation with colloid and catecholamines | 60 | 70 
intraoperative ultrasonography revealed massive air emboli | 60 | 60 
diagnosed with VAE and PAE | 60 | 60 
arterial blood gas analysis | 60 | 60 
catecholamine administration | 60 | 300 
systolic blood pressure maintained | 70 | 300 
heart rate maintained | 70 | 300 
central venous pressure maintained | 70 | 300 
end-tidal carbon dioxide restored | 70 | 300 
ABGA at 30 minutes after the occurrence of VAE | 90 | 90 
norepinephrine infusion | 70 | 300 
fluid resuscitation | 70 | 300 
air emboli in left heart disappeared | 130 | 130 
hepatectomy restarted | 130 | 300 
systolic pressure maintained | 130 | 300 
total anesthesia time | 0 | 300 
total fluid administered | 0 | 300 
total urinary output | 0 | 300 
total blood loss | 0 | 300 
intubated and ventilated mechanically in ICU | 300 | 744 
responded only to intense pain | 300 | 744 
systolic pressure maintained in ICU | 300 | 744 
norepinephrine infusion in ICU | 300 | 744 
postoperative laboratory findings | 300 | 300 
postoperative EKG | 300 | 300 
EKG findings recovered normally | 744 | 744 
trans-thoracic echocardiogram | 744 | 744 
vital signs stable | 744 | 744 
norepinephrine infusion tapered out | 744 | 744 
mental status unchanged | 744 | 744 
brain CT and MRI | 120 | 120 
multiple acute cerebral infarctions | 120 | 120 
weaned to spontaneous ventilation | 264 | 264 
extubated | 264 | 264 
vital signs became unstable | 360 | 360 
intravenous administration of catecholamines | 360 | 744 
panperitonitis confirmed | 360 | 744 
expired due to cardiac arrest | 744 | 744 
septic shock | 744 | 744 
cardiac arrest | 744 | 744