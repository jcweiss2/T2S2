35 years old|0
female|0
Hodgkin lymphoma|0
nodular sclerosis subtype|0
primary refractory HL|0
admitted to the hospital|0
generalized pruritus|0
atopic dermatitis|0
corticoid-based therapy|0
laterocervical lymphadenopathies|0
night fever|0
intense sweating|0
supra-diaphragmatic lymphadenopathies|0
infra-diaphragmatic lymphadenopathies|0
abdominal masses|0
lymphadenopathy biopsy|0
NS classic HL|0
stage IIIB HL|0
International Prognostic Score 2|0
ABVD chemotherapy regimen|0
partial response|-5520
early relapse|-5520
primary refractory to ABVD|-5520
ESHAP salvage chemotherapy regimen|-5520
no response|-5520
GemOx chemotherapy regimen|-5520
neutropenia grade 4|-5520
thrombocytopenia grade 4|-5520
dose-intensity failures|-5520
chemotherapy discontinuation|-5520
radiotherapy consolidation|-5520
HL progression|-5520
IFE chemotherapy regimen|-5520
stable disease|-5520
watch-and-wait policy|-5520
localized progression with radiotherapy|-5520
transient partial responses|-5520
new mass in D8–D9|-5520
medullar compression syndrome|-5520
HL relapse|-5520
radiotherapy|-5520
GemOx chemotherapy|-5520
new progression in left cervical nodes|-5520
new progression in axillary nodes|-5520
symptomatic disease progression|-5520
PET/CT confirmation|-5520
bendamustine 90 mg/m2|-5520
disease stability|-5520
significant B symptoms|-5520
worsening clinical status|-5520
celecoxib 200 mg every 12 hours|0
lenalidomide 20 mg|0
compassionate use treatment|0
unremarkable toxicity|0
excellent tolerance|0
complete response|0
interim CT/PET after three cycles|0
final CT/PET after six cycles|0
CT scan in August 2015|0
celecoxib maintenance 200 mg/12 hours|0
anemia due to gastrointestinal bleeding|0
celecoxib discontinuation|0
disease relapse|0
supra-abdominal adenopathies|0
infra-abdominal adenopathies|0
hepatic lesions|0
splenic lesions|0
negative biopsies|0
asymptomatic situation|0
celecoxib restarted 200 mg every 12 hours|0
disease progression to ascites|0
paracentesis|0
persistent HL|0
brentuximab vedotin|0
intensive care admission|0
sepsis|0
fatal outcome|0
