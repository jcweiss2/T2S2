51 years old | 0
male | 0
referred to the emergency room | 0
abdominal pain | -72
distended abdomen | 0
severe tenderness to palpation | 0
IV fluids started | 0
IV ondansetron | 0
morphine sulfate | 0
leukocytosis | 0
WBC count 14.5 thou/cm | 0
laparotomy | 0
normal small and large intestine | 0
normal vasculature | 0
discharged | 48
nausea | 0
abdominal pain | 48
dyspnea | 48
came back to ER | 72
tachypnea | 72
tachycardia | 72
low-grade fever | 72
lung CT | 72
abdominopelvic CT | 72
intubated | 72
Covid-19 RT-PCR | 72
WBC 17000 per microliter | 72
Hb 12:8.7 g/dL | 72
Plt 350000 per microliter | 72
urea 170 mg/dL | 72
Cr 4.2 mg/dL | 72
LDH 504 U/L | 72
CRP 47mg/L | 72
negative viral disease | 72
treated with hydroxychloroquine sulfate | 72
lopinavir/ritonavir | 72
ribavirin | 72
β interferon | 72
fecaloid discharged | 168
sepsis | 168
WBC 24000 per microliter | 168
Hb 12 g/dL | 168
Plt 347000 per microliter | 168
urea 206 mg/dL | 168
Cr 3.2 mg/dL | 168
amylase 67 U/L | 168
re-laparotomy | 168
serosanguinous secretions | 168
necrotic changes in small intestine | 168
130 cm resected | 168
leakage from anastomosis site | 192
smaller bowel necrosis | 192
100 cm resected | 192
ileostomy | 192
intravascular thrombosis | 192
necrotic margin | 192
RT-PCR positive | 192
treated with heparin infusion | 192
broad-spectrum antibiotics | 192
extubated | 240
hemodynamic stable | 240
platelet count decrease | 240
gastrointestinal bleeding | 240
WBC 7100 per microliter | 240
Hb 8.7 g/dL | 240
plt 162000 per microliter | 240
Cr 1.3 mg/dL | 240
amylase 65 U/L | 240
plt 69000 per microliter | 264
Cr 1.1 mg/dL | 264
heparin discontinued | 264
D-dimer 2500 ng/mL | 264
fibrinogen 150 mg/dL | 264
PT 44 sec | 264
PTT 44 sec | 264
INR 1.7 | 264
no schistocyte | 264
treatment-resistant sepsis | 264
DIC | 264
died | 264
