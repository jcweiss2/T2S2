newborn female | 0 | 0 
24 weeks + 3 days | 0 | 0 
breech presentation | 0 | 0 
cord prolapse | 0 | 0 
birth weight of 645 g | 0 | 0 
36-year-old mother | 0 | 0 
HIV negative | 0 | 0 
Apgar score of 4 | 0 | 0 
Apgar score of 8 | 0 | 5 
mechanical ventilation | 0 | 216 
central umbilical catheters | 0 | 216 
total parenteral nutrition | 0 | 216 
empiric antibiotics | 0 | 216 
skin sensors | 0 | 216 
late-onset sepsis | -216 | -216 
Escherichia coli bacteremia | -216 | -216 
cefepime | -216 | -96 
adhesive patch removal | -192 | -192 
skin abrasion | -192 | -192 
erythema | -168 | -168 
induration | -168 | -168 
plaque with necrotic center | -168 | -168 
ulcer | -144 | -144 
subcutaneous cell tissue extension | -144 | -144 
necrotic area progression | -144 | -144 
intensive treatment | -144 | -72 
wound care | -144 | -72 
healings | -144 | -72 
hydrating dermal wound dressings | -144 | -72 
sodium alginate | -144 | -72 
carboxymethylcellulose | -144 | -72 
hydrocolloids | -144 | -72 
thermic instability | -72 | -72 
metabolic acidosis | -72 | -72 
hyperglycemia | -72 | -72 
hypotension | -72 | -72 
clinical deterioration | -72 | -72 
cutaneous mucormicosis suspicion | -72 | -72 
skin biopsy | -72 | -72 
empiric antifungal treatment | -72 | 0 
liposomal amphotericin B | -72 | 0 
fungal biomarkers | -72 | -72 
serum galactomannan | -72 | -72 
1,3 beta-D-glucan | -72 | -72 
refractory shock | 0 | 36 
metabolic acidosis progression | 0 | 36 
renal failure | 0 | 36 
death | 36 | 36 
fungal cultures | -72 | -72 
Rhizopus spp. | -72 | -72 
histopathology | -72 | -72 
broad aseptate hyphae | -72 | -72 
right angle branching | -72 | -72 
Mucorales | -72 | -72 
mass spectroscopy | -72 | -72 
MALDI-TOF MS | -72 | -72 
polymerase chain reaction | -72 | -72 
PCR | -72 | -72 
Rhizopus arrhizus | -72 | -72 
fungal blood cultures | -216 | -216 
negative fungal blood cultures | -216 | -216 
necrotizing cellulitis | -144 | 36 
primary cutaneous mucormycosis | -192 | 36 
gangrenous form | -144 | 36 
necrotic eschar | -144 | 36 
skin abscesses | -144 | 36 
surgical debridement | 0 | 36 
anti-fungal treatment | -72 | 36 
L-AmB | -72 | 36 
ischemic necrosis | 0 | 36 
leukocytes | 0 | 36 
anti-fungal agents | 0 | 36 
infection control | 0 | 36 
traditional diagnostic methods | -72 | -72 
microbiology | -72 | -72 
histopathology | -72 | -72 
mass spectrometry | -72 | -72 
molecular studies | -72 | -72 
etiological diagnosis | -72 | -72 
infection site | -192 | 36 
left arm | -192 | 36 
cellulitis | -144 | 36 
ulcer | -144 | 36 
tissue necrosis | -144 | 36 
primary skin infection | -192 | 36 
secondary skin involvement | -192 | 36 
disseminated infection | -192 | 36 
autopsy | 36 | 36 
vesicle | -168 | -168 
pustule | -168 | -168 
erythematous plaque | -168 | -168 
necrotic plaque | -168 | -168 
papule | -144 | -144 
necrotizing cellulitis | -144 | 36 
distant tissues | -144 | 36 
skin abscesses | -144 | 36 
R. microsporus | -72 | -72 
R. arrhizus | -72 | -72 
R. oryzae | -72 | -72 
Lichtheimia corymbifera | -72 | -72 
Absidia corymbifera | -72 | -72 
cutaneous aspergillosis | -72 | -72 
hyalohyphomycosis | -72 | -72 
Fusarium | -72 | -72 
necrotizing fasciitis | -72 | -72 
clostridial gas gangrene | -72 | -72 
sepsis-associated purpura fulminans | -72 | -72 
bacterial cellulitis | -72 | -72 
pyoderma gangrenosum | -72 | -72 
broad hyaline hyphae | -72 | -72 
aseptate hyphae | -72 | -72 
vascular invasion | -72 | -72 
necrotic tissue | -72 | -72 
MALDI-TOF MS | -72 | -72 
PCR assays | -72 | -72 
mass spectrometry tests | -72 | -72 
fungal identification | -72 | -72 
species level | -72 | -72 
traditional methods | -72 | -72 
microbiology | -72 | -72 
histopathology | -72 | -72 
surgical debridement | 0 | 36 
anti-fungal treatment | -72 | 36 
L-AmB | -72 | 36 
underlying disease | 0 | 36 
predisposing factors | 0 | 36 
disease severity | 0 | 36 
ischemic necrosis | 0 | 36 
leukocytes | 0 | 36 
anti-fungal agents | 0 | 36 
infection control | 0 | 36 
Francis JR | -72 | -72 
pediatric patients | -72 | -72 
mucormycosis | -72 | -72 
antifungal therapy | -72 | -72 
surgical debridement | 0 | 36 
death risk | 0 | 36 
pooled data | -72 | -72 
children | -72 | -72 
antifungal therapy | -72 | -72 
surgical debridement | 0 | 36 
infection control | 0 | 36 
high suspicion | 0 | 36 
prompt recognition | 0 | 36 
aggressive approach | 0 | 36 
traditional diagnostic methods | -72 | -72 
microbiology | -72 | -72 
histopathology | -72 | -72 
mass spectrometry | -72 | -72 
molecular studies | -72 | -72 
etiological diagnosis | -72 | -72 
Álvaro Hoyos | 0 | 0 
María Adelaida Mejía | 0 | 0 
Verónica Herrera | 0 | 0 
Andrés Soto | 0 | 0 
Clara Rico | 0 | 0 
Alejandro Díaz-Díaz | 0 | 0 
Institutional Ethics Committee | 0 | 0 
Clínica Universitaria Bolivariana | 0 | 0 
Universidad Pontificia Bolivariana | 0 | 0 
CRediT authorship | 0 | 0 
conceptualization | 0 | 0 
writing | 0 | 0 
review | 0 | 0 
editing | 0 | 0 
supervision | 0 | 0 
formal analysis | 0 | 0 
investigation | 0 | 0 
validation | 0 | 0 
visualization | 0 | 0 
funding | 0 | 0 
grant | 0 | 0 
public | 0 | 0 
commercial | 0 | 0 
not-for-profit | 0 | 0 
sectors | 0 | 0 
consent | 0 | 0 
case report | 0 | 0 
approval | 0 | 0 
declaration | 0 | 0 
competing interest | 0 | 0 
authors | 0 | 0 
conflicting interests | 0 | 0 
acknowledgements | 0 | 0 
critical review | 0 | 0