44 years old | 0
male | 0
admitted to the hospital | 0
bronchobiliary fistula | -720
pneumonia | -720
pancreaticoduodenectomy | -4032
transarterial embolization | -672
dilation of the bile duct | -720
multiple bilomas | -720
poor oral intake | -720
fluctuating fever | -720
jaundice | -720
intravenous antibiotic treatment | -720
repeated drainage | -720
endoscopic retrograde biliary drainage | -720
percutaneous transhepatic biliary drainage | -720
recurrent biliary stent obstruction | -168
acute dyspnea | -168
yellowish sputum | -168
bilirubin in sputum | -168
preoperative chest X-ray | 0
progressive consolidation | 0
pleural effusion | 0
abdominal computed tomography | 0
dilated bile duct | 0
bilomas | 0
chest computed tomography | 0
subdiaphragmatic abscess | 0
pneumonic consolidation | 0
necrotizing change | 0
bilateral pleural effusion | 0
tubogram | 0
fistulous communication | 0
fiberoptic bronchoscopy | 0
copious bile | 0
preoperative arterial blood gas analysis | 0
leukocytosis | 0
total bilirubin | 0
direct bilirubin | 0
alkaline phosphatase | 0
γ-glutamyl transferase | 0
albumin | 0
lactate | 0
international normalized ratio | 0
Staphylococcus aureus | 0
Escherichia coli | 0
Enterococcus faecium | 0
Pseudomonas aeruginosa | 0
surgical treatment | 0
percutaneous transhepatic biliary drainage | 0
preoperative biliary decompression | 0
electrocardiogram | 0
pulse oximetry | 0
invasive arterial blood pressure | 0
oxygen saturation | 0
heart rate | 0
preoxygenation | 0
rapid sequence induction | 0
etomidate | 0
rocuronium | 0
left-sided double-lumen endobronchial tube | 0
auscultation | 0
visualization | 0
fiberoptic bronchoscopy | 0
ventilation | 0
target-controlled infusion | 0
propofol | 0
remifentanil | 0
bispectral index | 0
central venous pressure | 0
cannulation | 0
esophageal temperature | 0
urine output | 0
bile-stained secretions | 0
trachea | 0
carina | 0
right bronchus | 0
one-lung ventilation | 0
tidal volume | 0
respiratory rate | 0
positive end-expiratory pressure | 0
lateral decubitus position | 0
oxygenation | 0
repeated bronchial lavage | 0
resection of the fistula | 0
bilobectomy | 0
perforated diaphragm | 0
subphrenic drain | 0
two-lung ventilation | 0
recruit maneuver | 0
oxygenation | 0
anesthesia | 445
operation | 340
estimated blood loss | 0
crystalloid | 0
packed red blood cells | 0
dopamine | 0
urine output | 0
hypokalemia | 0
potassium repletion | 0
single-lumen endotracheal tube | 0
postoperative mechanical ventilation | 0
sedation | 0
dexmedetomidine | 0
remifentanil | 0
controlled mandatory ventilation | 0
postoperative chest X-ray | 0
decreased effusion | 0
extubation | 96
follow-up examination | 720
no sign of BBF recurrence | 720
progressive sepsis | 4032
wound infection | 4032
hepatic failure | 4032
necrotizing pneumonia | 4032
repeated biliary stent stricture | 4032