80 years old | 0
female | 0
hypertension | 0
asthma | 0
hypothyroidism | 0
presented to the Emergency Department | 0
erythematous right lower extremity | 0
edematous right lower extremity | 0
ecchymosis | 0
superficial erosions | 0
clear drainage | 0
laceration to the affected leg | -96
remained in wet pants for multiple hours | -96
increased edema | -72
increased erythema | -72
increased pain | -72
bullae developed | -72
drained the lesions | -48
expression of clear fluid | -48
sloughing of the epidermis | -48
vital signs within normal limits | 0
WBC count 7400 cells/mcL | 0
50% band neutrophils | 0
elevated lactate 3.0 mmol/L | 0
blood cultures obtained | 0
ceftriaxone IVPB 1g | 0
admitted to the hospital | 0
cellulitis of the right lower extremity | 0
bandemia | 0
lactic acidosis | 0
acute hypoxic respiratory failure | 24
altered mentation | 24
hypotension | 24
transferred to the Intensive Care Unit | 24
severe sepsis | 24
cefepime started | 24
metronidazole started | 24
returned to the medical floor | 72
blood cultures grew Plesiomonas shigelloides | 72
antimicrobial susceptibilities sensitive to ceftriaxone | 72
antimicrobial susceptibilities sensitive to ciprofloxacin | 72
antimicrobial susceptibilities sensitive to ertapenem | 72
antimicrobial susceptibilities sensitive to meropenem | 72
ciprofloxacin added | 72
changes in stool | 168
ciprofloxacin discontinued | 168
concerns for Clostridium difficile infection | 168
general surgery consulted | 168
wound debridement performed | 168
condition continued to improve | 336
discharged to inpatient rehab | 336
metronidazole 500 mg TID | 336
ceftriaxone IVPB 2g daily | 336
discharged from inpatient rehab | 504
instructions to follow up with family doctor | 504
