75 years old | 0
female | 0
admitted to the emergency department | 0
unconscious | 0
productive cough | -96
fever | -96
high blood pressure | -672
paroxysmal atrial fibrillation | -672
type 2 diabetes | -672
bisoprolol | -672
propafenone | -672
atorvastatin | -672
metformin | -672
aspirin | -672
nonsmoker | 0
no occupational exposures | 0
tachypnoea | 0
tachycardia | 0
atrial fibrillation | 0
normal blood pressure | 0
transcutaneous arterial oxygen saturation decreased | 0
diffuse wheezing | 0
diminished breath sounds | 0
mild dullness at the right base of the lung | 0
severe inflammation | 0
white blood cell count 20.9×10^9 cells per L | 0
neutrophils 17.2×10^9 cells per L | 0
C-reactive protein 326.1 mg·L−1 | 0
elevated liver transaminases | 0
alanine aminotransferase 3216 U·L−1 | 0
aspartate aminotransferase 4359 U·L−1 | 0
decreased kidney function | 0
creatinine 313 µmol·L−1 | 0
urea 26.2 mmol·L−1 | 0
severe hypercapnic respiratory failure | 0
carbon dioxide tension 107 mmHg | 0
oxygen tension 63 mmHg | 0
pH 7.04 | 0
HCO3− 28.9 mmol·L−1 | 0
chest radiography | 0
computed tomography (CT) | 0
pulmonary oedema | 0
right-sided infiltrates | 0
aspiration pneumonia | 0
antibiotic therapy with intravenous piperacillin/tazobactam | 0
intubated | 0
mechanically ventilated | 0
transferred to the intensive care unit (ICU) | 0
regained consciousness | 24
laboratory tests returned to normal | 24
cultures from bronchoalveolar lavage were positive for Haemophilus influenzae | 24
persistent hypercapnic respiratory failure | 48
tracheostomy | 48
mechanical ventilation discontinued | 360
breathing spontaneously through the tracheostomy tube | 360
dyspnoea | 360
mild weakness | 360
severe shortness of breath | 360
stridor | 360
acute respiratory insufficiency | 360
tracheal dyskinesia | 360
bilateral vocal cord paresis | 360
neuromuscular pathology suspected | 360
slight muscular weakness in the proximal leg muscles | 360
fatigability of the extraocular muscles | 360
myasthenia gravis suspected | 360
critical illness polyneuropathy | 360
Guillain–Barré syndrome | 360
nerve conduction studies with repetitive nerve stimulation (RNS) | 360
single-fibre electromyography (SFEMG) | 360
acetylcholine receptor (AChR) antibodies | 360
antibodies against muscle-specific kinase (MuSK) | 360
AChR antibodies negative | 360
RNS studies showed a decremental muscle electrical response | 360
myasthenia gravis diagnosed | 360
pyridostigmine 150 mg·day−1 | 360
prednisolone 5 mg·day−1 | 360
dyspnoea and difficulty breathing disappeared | 384
hypercapnia resolved | 384
permanent tracheostomy tube placed | 504
discharged | 504