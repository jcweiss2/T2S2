35 years old | 0
male | 0
Samoan American | 0
congenital deafness | 0
hypertension | 0
asthma | 0
admitted to the hospital | 0
night sweats | -144
rash | -144
productive cough | -144
shortness of breath | -144
fevers | -144
intermittent back pain | -144
enlarging neck nodule | -144
diagnosed with Valley Fever | -1440
fluconazole | -1440
scaling plaques to the right forehead | 0
small ulcerated lesions to the right lower mouth and posterior neck | 0
coarse breath sounds in the left upper lung fields | 0
nontender lymph node to the left anterior neck | 0
leukocytosis with predominant neutrophilia | 0
elevated erythrocyte sedimentation rate | 0
elevated C-reactive protein | 0
elevated liver enzymes | 0
total protein of 10.0 g/dL | 0
albumin of 1.7 g/dL | 0
corrected calcium of 11.0 mg/dL | 0
elevated alkaline phosphatase of 167 U/L | 0
elevated lactic acid of 2.7 mmol/L | 0
elevated lactate dehydrogenase of 341 U/L | 0
ferritin of 3366 ng/mL | 0
anemia of chronic disease | 0
respiratory viral panel positive for respiratory syncytial virus | 0
disseminated fungal diseases | 0
histoplasmosis | 0
blastomycosis | 0
tuberculosis | 0
secondary hemophagocytic lymphohistiocytosis | 0
HIV | 0
malignancy | 0
Infectious Diseases consulted | 0
serum coccidioides IgG ELISA | 0
serum coccidioides IgM ELISA | 0
direct microscopy of the sputum revealed spherules resembling coccidioides | 0
magnetic resonance imaging of the spine | 24
magnetic resonance imaging of the pelvis | 24
computed tomography–guided biopsy of the right iliac crest | 48
computed tomography–guided biopsy of the cervical lymph node | 48
lumbar puncture | 48
high-flow nasal cannula | 24
intravenous fluids | 24
itraconazole | 24
liposomal amphotericin B | 24
supplemental oxygen | 24
transferred to the intensive care unit | 48
intubated | 48
vasopressors | 48
chest X-ray | 72
computed tomography scan of the chest | 96
ceftriaxone | 96
azithromycin | 96
acute kidney injury | 120
paralytic ileus | 120
right internal jugular deep vein thrombosis | 120
gluteal hematoma | 120
voriconazole | 168
mechanical ventilation | 168
discharged | 1008
intensive inpatient rehabilitation program | 1008
severe physical deconditioning | 1008