72 years old | 0
woman | 0
cough | -168
shortness of breath | -168
weakness | -168
hypoxic | 0
oxygen saturation of 80% | 0
admitted for COVID-19 pneumonia | 0
superimposed bacterial pneumonia | 0
sepsis | 0
hypertension | 0
hypothyroidism | 0
obesity | 0
dexamethasone | 0
albuterol | 0
nasal cannula oxygen | 0
therapeutic dosing of enoxaparin |C0
gram-positive cocci in clusters | 0
vancomycin | 0
meropenem | 0
doxycycline | 0
intravenous piggyback | +48
doxycycline infiltration | +48
mild swelling | +48
pain | +48
worsening respiratory failure | +96
endotracheal intubation | +96
transfer to intensive care unit | +96
norepinephrine | +96
hypotension | +96
pronEd periodically | +96
gradual improvement of respiratory status | +96
triple lumen central catheter | +96
no peripheral intravenous catheters | +96
poor peripheral venous access | +96
left hand swelling | +432
dorsal purplish bulla | +432
responsive | +432
pain in hand | +432
pain in distal forearm | +432
unable to flex fingers | +432
denied numbness | +432
vascular surgery consultation | +432
no signs of arterial insufficiency | +432
computed tomography demonstrated hematoma | +432
no evidence of venous thrombosis | +432
nonsurgical management | +432
local wound care | +432
hand surgery consultation | +504
hematoma evacuation | +504
worsened swelling | +504
worsened pain | +504
faint ulnar Doppler signal | +504
faint radial Doppler signal | +504
cool fingers | +504
blistering | +504
mottling | +504
intrinsic minus posturing | +504
passive extension pain | +504
limited active range of motion | +504
compartment pressures elevated | +504
delta pressures | +504
decompressive fasciotomy | +504
thenar muscle edema | +504
hypothenar muscle edema | +504
dorsal incisions | +504
compartments released | +504
dorsal fasciotomies closed | +504
improved pain | +552
limited range of motion | +552
improved swelling | +552
superficial necrosis | +744
eschar ulnarly | +744
discharged | +744
continued recovery through physical therapy | +1248
composite fist formation | +1248
full finger extension | +1248
necrotic eschar debridement | +1248
wound fully healed | +4872
mild scar contracture | +4872
wrist flexion limitation | +4872
full wrist extension | +4872
full range of motion | +4872
Disabilities of the Arm, Shoulder, and Hand score 60 | +4872
very satisfied | +4872
resolution of neuropathic pain | +4872
