68 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
type 1 diabetic | 0 | 0 | Factual
hypertensive | 0 | 0 | Factual
on amlodipine | 0 | 0 | Factual
operated for treatment of right inguinal hernia | -7200 | -7200 | Factual
admitted to the emergency room | 0 | 0 | Factual
abdominal pain | -72 | 0 | Factual
ketoacidosis decompensation | -72 | 0 | Factual
uremic syndrome | -72 | 0 | Factual
conscious patient | 0 | 0 | Factual
hemodynamically stable | 0 | 0 | Factual
dyspneic | 0 | 0 | Factual
febrile at 39,6 °C | 0 | 0 | Factual
right lumbar tenderness | 0 | 0 | Factual
oliguric | 0 | 0 | Factual
diuresis at 300 ml/24h | 0 | 0 | Factual
altered renal function | 0 | 0 | Factual
creatinine at 92 mg/l | 0 | 0 | Factual
urea at 3,1 g/l | 0 | 0 | Factual
K+ at 6.9 mmol/l | 0 | 0 | Factual
Na+ at 123 mmol/l | 0 | 0 | Factual
blood sugar at 6.5 g/l | 0 | 0 | Factual
alkaline reserves at 8 mEq/l | 0 | 0 | Factual
infectious syndrome | 0 | 0 | Factual
CRP at 418 mg/l | 0 | 0 | Factual
white blood cells at 26000/ml | 0 | 0 | Factual
hemoglobin at 12,3 g/dl | 0 | 0 | Factual
leucocyturia 320,000 | 0 | 0 | Factual
hematuria at 120,000 | 0 | 0 | Factual
single anatomical right kidney | 0 | 0 | Factual
emphysematous pyelonephritis | 0 | 0 | Factual
renal abscess | 0 | 0 | Factual
pneumoperitoneum | 0 | 0 | Factual
admitted to intensive care | 0 | 0 | Factual
dialysis sessions | 0 | 72 | Factual
insulin therapy | 0 | 240 | Factual
antibiotic therapy | 0 | 240 | Factual
ceftriaxone | 0 | 48 | Factual
metronidazole | 0 | 48 | Factual
surgical drainage of abscesses | 48 | 48 | Factual
right double J stent | 48 | 336 | Factual
favorable evolution | 72 | 240 | Factual
decrease of the infectious syndrome | 72 | 240 | Factual
apyrexia | 48 | 48 | Factual
chronic renal failure | 240 | 240 | Factual
creatinine plateau of 20 mg/l | 240 | 240 | Factual
discharged | 240 | 240 | Factual
oral antibiotics | 240 | 672 | Factual
abdominopelvic CT | 672 | 672 | Factual
clear regression of the bubbles of air | 672 | 672 | Factual
double J catheter removed | 1008 | 1008 | Factual