35-year-old woman | 0
    gravid 3 | 0
    para 2 | 0
    referred to radiology department | 0
    second-trimester ultrasonography | -1680
    omphalocele | -1680
    prior normal vaginal delivery | -1440
    healthy offspring | -1440
    no history of smoking | 0
    no medical illness | 0
    no specific medications | 0
    no congenital anomalies | 0
    23rd week of gestation | -1680
    small fetal chest | -1680
    loss of anterior chest wall | -1680
    heart exposed outside | -1680
    cardiac chambers with slight loss of configuration | -1680
    cardiac anomalies not excluded | -1680
    Pentalogy of Cantrell | -1680
    supra/umbbilical omphalocele | -1680
    bowel loops | -1680
    liver | -1680
    amniocentesis not performed | -1680
    MRI revealed extra-thoracic heart | -1680
    anterior to chest cavity | -1680
    herniation of left lung | -1680
    herniated liver through anterior abdominal wall | -1680
    dilated bowel | -1680
    stenosis possibility | -1680
    atresia possibility | -1680
    spinal deformity | -1680
    ectopia cordis | -1680
    33rd gestational week | -432
    male gender | -432
    diagnosis of Pentalogy of Cantrell | -432
    caesarian section | 0
    newborn length 46 cm | 0
    weight 2100 g | 0
    head circumference 30 cm | 0
    thoracic perimeter 25 cm | 0
    Apgar score 3/10 (first minute) | 0
    Apgar score 6/10 (fifth minute) | 0
    bulky omphalocele | 0
    liver out of abdomen | 0
    bowel loops out of abdomen | 0
    thick membranous covering | 0
    maldevelopment of distal sternum | 0
    diaphragmatic hernia | 0
    heart located outside chest | 0
    cardiac abnormalities | 0
    admitted to NICU | 0
    mechanical ventilation | 0
    progressive respiratory failure | 0
    severe respiratory acidosis | 0
    electrolyte imbalance | 0
    general condition deteriorated | 24
    died | 48
    septicemia | 48
    respiratory failure | 48
    <|eot_id|>
    