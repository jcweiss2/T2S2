68 years old | 0
male | 0
transferred to hospital | 0
dyspnea | -2160
femoral neck fracture | -2160
radiation therapy for tonsil cancer | -87600
recurrent aspiration | -87600
refused nasogastric tube | -2160
refused percutaneous endoscopic gastrostomy feeding | -2160
admitted to secondary hospital for nutritional support | -2160
malnutrition | -2160
slipped and broke femur | -2160
refused femur operation | -2160
dyspnea aggravation | -2160
aspiration pneumonia | 0
recommended nothing per oral | 0
mother gave vegetable soup with solid materials | 120
respiratory failure | 120
shock | 120
intubated | 120
transferred to ICU | 120
ventilator care | 120
monitoring | 120
bronchoscopy | 120
extracted vegetables (carrot, potato) | 120
recovered from pneumonia | 120
difficulty liberating from ventilator | 120
recommended tracheostomy | 120
family refused tracheostomy | 120
sustained persuasion over 2 months | 120
family agreed to tracheostomy | 120
percutaneous dilatational tracheostomy | 120
discharged to nursing hospital with home ventilator | 432
visited ER with fever and dyspnea | 4320
transferred to another hospital | 4320
chest CT showing pneumonia | 4320
visited ER due to secretion resembling enteral feeding materials | 6480
chest CT revealed TEF | 6480
continuous leakage of ventilator circuit | 6480
changed T-tube to endotracheal tube | 6480
inflated balloon to maximum | 6480
bronchoscopy revealed TEF | 6480
oval-shaped TEF 2 cm in diameter | 6480
TEF located on left side of proximal trachea | 6480
NG tube visible through TEF | 6480
consulted radiologist | 6480
consulted gastroenterologist | 6480
consulted pulmonary interventionist | 6480
consulted chest surgeon | 6480
radiologist: esophageal stent impossible | 6480
gastroenterologist: endosponge and vacuum therapy impossible | 6480
pulmonary interventionist: no stent available | 6480
thoracic surgeon: recommended primary closure after PEG and liberation from ventilator | 6480
intensivists: liberation from ventilator impossible due to muscle weakness | 6480
family refused PEG | 6480
gave up primary treatment of TEF | 6480
discharged to nursing hospital | 6480
family agreed to withdraw life-sustaining treatment | 6480
patient and family changed mind, wanted PEG | 65520
admitted to ICU | 65520
planned esophagogastroscopy and PEG | 65520
routine scope could not enter esophagus due to stenosis | 65520
complication from radiation therapy | 65520
PEG impossible | 65520
thinner scope investigated esophagus | 65520
balloon of endotracheal tube in esophagus | 65520
discussed jejunostomy | 65520
malnutrition | 65520
pneumonia | 65520
septic shock | 65520
died | 65520
