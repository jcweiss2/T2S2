75 years old | 0
female | 0
hypertension | 0
hyperlipidemia | 0
leukocytosis | -730
weight loss | -730
fatigue | -90
admitted to the hospital | 0
T-PLL | 0
alemtuzumab | 0
pentostatin | 0
rash | 196
facial swelling | 196
sore throat | 196
dysphagia | 196
conjunctivitis | 196
anasarca | 200
respiratory distress | 200
intubation | 216
mechanical ventilation | 216
sepsis | 220
death | 240
WBC count of 461 × 10^9/L | 0
Hgb of 6.9 gm/dL | 0
flow cytometry of the peripheral blood showed T-PLL | 0
bone marrow biopsy | 0
cytogenetic analysis | 0
inversion at chromosome 14 | 0
trisomy 8 | 0
karyotype analysis | 0
clonal T-cell gene rearrangement | 0
computed tomography chest, abdomen, and pelvis | 0
splenomegaly | 0
lymphadenopathy | 0
hepatomegaly | 0
skin lesions | 196
cutaneous manifestations | 196
diffuse skin rash | 196
edema | 200
lymphocytic infiltration | 200
tumor lysis syndrome | 200
uric acid elevated | 200
creatinine elevated | 200
rasburicase | 200
alemtuzumab and pentostatin therapy | 200
CMV and PCP prophylaxis | 200
valganciclovir | 200
Bactrim | 200
peripheral blood smear | 200
flow cytometry | 200
skin biopsy | 200
atypical perivascular lymphocytic infiltrate | 200
CD7+, CD2+, CD3+, CD4+, and CD5+ | 200
CD8, CD30, and CD56 negative | 200
lymphadenopathy in the mediastinal and cervical chains | 208
tachypnea | 216
oxygen saturation dropped | 216
hypotension | 216
shock | 216
racemic epinephrine | 216
Benadryl | 216
methylprednisolone | 216
intubation | 216
ventilation | 216
intravenous pressor support | 216
lactate increased | 220
creatinine increased | 220
infectious workup | 220
sepsis suspected | 220
medical intensive care unit | 220
death | 240