72 years old | 0
female | 0
gravida 2 | 0
para 2 | 0
hypothyroidism | -6720
hyperlipidemia | -6720
hypertension | -6720
osteoarthritis | -6720
bilateral oophorectomy | -1440
bilateral knee replacements | -240
colonoscopy | -480
severe abdominal pain | -8
vaginal bleeding | -8
nausea | -8
vomiting | -8
chills | -8
severe distress | 0
tympanic abdomen | 0
distended abdomen | 0
tender to palpation | 0
rebound tenderness | 0
moderate leukocytosis | 0
anion gap metabolic acidosis | 0
azotemia | 0
minimal urine output | 0
given 2 L of normal saline | 0
catheterized with a Foley catheter | 0
uterine prolapse | 0
mild vaginal bleeding | 0
computed tomography scan | 0
pneumoperitoneum | 0
pneumobilia | 0
colonic perforation | 0
enterofistula | 0
taken to the operating room | 2
emergent exploratory laparotomy | 2
foul-smelling gas | 2
spontaneous rupture of the posterior fundus | 2
intrauterine malignancy | 2
total abdominal hysterectomy | 2
salpingectomy | 2
appendectomy | 2
peritoneal cavity irrigated | 2
antibiotic solution | 2
peritoneal-cavity fluid cultures | 2
uterine myometrial tissue sent for pathology | 2
abdomen closed with retention sutures | 2
Jackson-Pratt drain placed | 2
severe end organ damage | 4
multi end organ failure | 4
intubated | 4
transferred to surgical intensive care unit | 4
pathologic report | 24
advanced high-grade serous adenocarcinoma | 24
blood gram stain | 24
C. perfringens | 24
broad-spectrum antibiotics | 24
norepinephrine | 24
pressure support | 24
piperacillin/tazobactam | 24
vancomycin | 24
metronidazole | 24
blood and peritoneal fluid cultures | 48
antibiotic regimen changed | 48
vancomycin | 48
intravenous penicillin G | 48
abdomen tense and distended | 96
worsening multiorgan failure | 96
reexploration of abdominal cavity | 96
necrosis of distal half of small bowel | 96
necrosis of entire colon | 96
ileectomy | 96
total colectomy | 96
resection of proximal rectum | 96
washout of peritoneal cavity | 96
bowel left in discontinuity | 96
wound vacuum in place | 96
ileostomy creation | 144
focal areas of patchy necrosis | 144
multiple resections | 144
ileostomy created | 144
necrosis at site of ileostomy | 144
hemodynamic instability | 144
advance directives revisited | 144
comfort care with terminal wean | 144
died | 144