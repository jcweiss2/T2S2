47 years old | 0
female | 0
hypothyroidism | -6480
Hashimoto’s thyroiditis | -6480
iron deficiency anemia | -6480
lymphadenopathy | -6480
ITP | -6480
Pfizer-BioNTech mRNA vaccine | 0
mild arm soreness | 0
easy bruising | 432
gum bleeding | 432
epistaxis | 432
ecchymosis | 432
petechiae | 432
thrombocytopenia | 432
platelet count 1000/mcL | 432
prothrombin time 16.2 seconds | 432
international normalized ratio 1.5 mg/dL | 432
reticulocyte count 2.2% | 432
lactate dehydrogenase 310 U/L | 432
atypical lymphocytes | 432
alkaline phosphatase 109 U/L | 432
antinuclear antibody screen negative | 432
dexamethasone | 432
admitted to ICU | 432
platelet transfusion | 432
IVIG | 432
CT scans | 432
Sjogren’s SS-A antibody positive | 432
ANA positive | 432
Epstein-Barr virus DNA positive | 432
hepatitis C negative | 432
hepatitis B negative | 432
HIV negative | 432
thyroid-stimulating hormone negative | 432
discharged | 456
ITP diagnosed | -6480
platelets 4000/mcL | -6480
prednisone | -6480
complete remission | -6480
ITP flare-up | -4320
platelets 3000/mcL | -4320
human immune globulin | -4320
dexamethasone | -4320
direct platelet antibody level 1962 | -4320
rheumatoid factor 20.7 IU/mL | -4320
bone marrow biopsy | -4320
karyotyping 46XX | -4320
enlarged left axillary lymph node | -1092
left axillary and retroperitoneal adenopathy | -1092
biopsy of left axillary lymph node | -1092
follicular hyperplasia | -1092
flow cytometry negative | -1092
fine needle aspirate negative | -1092
excisional biopsies negative | -1092
COVID-19 vaccine administration | 0 
first dose | 0 
Pfizer-BioNTech COVID mRNA vaccine | 0 
mild arm soreness | 48 
easy bruising | 432 
gum bleeding | 432 
epistaxis | 432 
ecchymosis | 432 
petechiae | 432 
thrombocytopenia | 432 
platelet count 1000/mcL | 432 
prothrombin time 16.2 seconds | 432 
international normalized ratio 1.5 mg/dL | 432 
reticulocyte count 2.2% | 432 
lactate dehydrogenase 310 U/L | 432 
atypical lymphocytes | 432 
alkaline phosphatase 109 U/L | 432 
antinuclear antibody screen negative | 432 
dexamethasone | 432 
admitted to ICU | 432 
platelet transfusion | 432 
IVIG | 432 
CT scans | 432 
Sjogren’s SS-A antibody positive | 432 
ANA positive | 432 
Epstein-Barr virus DNA positive | 432 
hepatitis C negative | 432 
hepatitis B negative | 432 
HIV negative | 432 
thyroid-stimulating hormone negative | 432 
discharged | 456 
ITP diagnosed | -6480 
platelets 4000/mcL | -6480 
prednisone | -6480 
complete remission | -6480 
ITP flare-up | -4320 
platelets 3000/mcL | -4320 
human immune globulin | -4320 
dexamethasone | -4320 
direct platelet antibody level 1962 | -4320 
rheumatoid factor 20.7 IU/mL | -4320 
bone marrow biopsy | -4320 
karyotyping 46XX | -4320 
enlarged left axillary lymph node | -1092 
left axillary and retroperitoneal adenopathy | -1092 
biopsy of left axillary lymph node | -1092 
follicular hyperplasia | -1092 
flow cytometry negative | -1092 
fine needle aspirate negative | -1092 
excisional biopsies negative | -1092 
COVID-19 vaccine administration | 0 
first dose | 0 
Pfizer-BioNTech COVID mRNA vaccine | 0 
mild arm soreness | 48 
easy bruising | 432 
gum bleeding | 432 
epistaxis | 432 
ecchymosis | 432 
petechiae | 432 
thrombocytopenia | 432 
platelet count 1000/mcL | 432 
prothrombin time 16.2 seconds | 432 
international normalized ratio 1.5 mg/dL | 432 
reticulocyte count 2.2% | 432 
lactate dehydrogenase 310 U/L | 432 
atypical lymphocytes | 432 
alkaline phosphatase 109 U/L | 432 
antinuclear antibody screen negative | 432 
dexamethasone | 432 
admitted to ICU | 432 
platelet transfusion | 432 
IVIG | 432 
CT scans | 432 
Sjogren’s SS-A antibody positive | 432 
ANA positive | 432 
Epstein-Barr virus DNA positive | 432 
hepatitis C negative | 432 
hepatitis B negative | 432 
HIV negative | 432 
thyroid-stimulating hormone negative | 432 
discharged | 456 
ITP diagnosed | -6480 
platelets 4000/mcL | -6480 
prednisone | -6480 
complete remission | -6480 
ITP flare-up | -4320 
platelets 3000/mcL | -4320 
human immune globulin | -4320 
dexamethasone | -4320 
direct platelet antibody level 1962 | -4320 
rheumatoid factor 20.7 IU/mL | -4320 
bone marrow biopsy | -4320 
karyotyping 46XX | -4320 
enlarged left axillary lymph node | -1092 
left axillary and retroperitoneal adenopathy | -1092 
biopsy of left axillary lymph node | -1092 
follicular hyperplasia | -1092 
flow cytometry negative | -1092 
fine needle aspirate negative | -1092 
excisional biopsies negative | -1092 
COVID-19 vaccine administration | 0 
first dose | 0 
Pfizer-BioNTech COVID mRNA vaccine | 0 
mild arm soreness | 48 
easy bruising | 432 
gum bleeding | 432 
epistaxis | 432 
ecchymosis | 432 
petechiae | 432 
thrombocytopenia | 432 
platelet count 1000/mcL | 432 
prothrombin time 16.2 seconds | 432 
international normalized ratio 1.5 mg/dL | 432 
reticulocyte count 2.2% | 432 
lactate dehydrogenase 310 U/L | 432 
atypical lymphocytes | 432 
alkaline phosphatase 109 U/L | 432 
antinuclear antibody screen negative | 432 
dexamethasone | 432 
admitted to ICU | 432 
platelet transfusion | 432 
IVIG | 432 
CT scans | 432 
Sjogren’s SS-A antibody positive | 432 
ANA positive | 432 
Epstein-Barr virus DNA positive | 432 
hepatitis C negative | 432 
hepatitis B negative | 432 
HIV negative | 432 
thyroid-stimulating hormone negative | 432 
discharged | 456 
ITP diagnosed | -6480 
platelets 4000/mcL | -6480 
prednisone | -6480 
complete remission | -6480 
ITP flare-up | -4320 
platelets 3000/mcL | -4320 
human immune globulin | -4320 
dexamethasone | -4320 
direct platelet antibody level 1962 | -4320 
rheumatoid factor 20.7 IU/mL | -4320 
bone marrow biopsy | -4320 
karyotyping 46XX | -4320 
enlarged left axillary lymph node | -1092 
left axillary and retroperitoneal adenopathy | -1092 
biopsy of left axillary lymph node | -1092 
follicular hyperplasia | -1092 
flow cytometry negative | -1092 
fine needle aspirate negative | -1092 
excisional biopsies negative | -1092 
COVID-19 vaccine administration | 0 
first dose | 0 
Pfizer-BioNTech COVID mRNA vaccine | 0 
mild arm soreness | 48 
easy bruising | 432 
gum bleeding | 432 
epistaxis | 432 
ecchymosis | 432 
petechiae | 432 
thrombocytopenia | 432 
platelet count 1000/mcL | 432 
prothrombin time 16.2 seconds | 432 
international normalized ratio 1.5 mg/dL | 432 
reticulocyte count 2.2% | 432 
lactate dehydrogenase 310 U/L | 432 
atypical lymphocytes | 432 
alkaline phosphatase 109 U/L | 432 
antinuclear antibody screen negative | 432 
dexamethasone | 432 
admitted to ICU | 432 
platelet transfusion | 432 
IVIG | 432 
CT scans | 432 
Sjogren’s SS-A antibody positive | 432 
ANA positive | 432 
Epstein-Barr virus DNA positive | 432 
hepatitis C negative | 432 
hepatitis B negative | 432 
HIV negative | 432 
thyroid-stimulating hormone negative | 432 
discharged | 456 
ITP diagnosed | -6480 
platelets 4000/mcL | -6480 
prednisone | -6480 
complete remission | -6480 
ITP flare-up | -4320 
platelets 3000/mcL | -4320 
human immune globulin | -4320 
dexamethasone | -4320 
direct platelet antibody level 1962 | -4320 
rheumatoid factor 20.7 IU/mL | -4320 
bone marrow biopsy | -4320 
karyotyping 46XX | -4320 
enlarged left axillary lymph node | -1092 
left axillary and retroperitoneal adenopathy | -1092 
biopsy of left axillary lymph node | -1092 
follicular hyperplasia | -1092 
flow cytometry negative | -1092 
fine needle aspirate negative | -1092 
excisional biopsies negative | -1092 
COVID-19 vaccine administration | 0 
first dose | 0 
Pfizer-BioNTech COVID mRNA vaccine | 0 
mild arm soreness | 48 
easy bruising | 432 
gum bleeding | 432 
epistaxis | 432 
ecchymosis | 432 
petechiae | 432 
thrombocytopenia | 432 
platelet count 1000/mcL | 432 
prothrombin time 16.2 seconds | 432 
international normalized ratio 1.5 mg/dL | 432 
reticulocyte count 2.2% | 432 
lactate dehydrogenase 310 U/L | 432 
atypical lymphocytes | 432 
alkaline phosphatase 109 U/L | 432 
antinuclear antibody screen negative | 432 
dexamethasone | 432 
admitted to ICU | 432 
platelet transfusion | 432 
IVIG | 432 
CT scans | 432 
Sjogren’s SS-A antibody positive | 432 
ANA positive | 432 
Epstein-Barr virus DNA positive | 432 
hepatitis C negative | 432 
hepatitis B negative | 432 
HIV negative | 432 
thyroid-stimulating hormone negative | 432 
discharged | 456 
ITP diagnosed | -6480 
platelets 4000/mcL | -6480 
prednisone | -6480 
complete remission | -6480 
ITP flare-up | -4320 
platelets 3000/mcL | -4320 
human immune globulin | -4320 
dexamethasone | -4320 
direct platelet antibody level 1962 | -4320 
rheumatoid factor 20.7 IU/mL | -4320 
bone marrow biopsy | -4320 
karyotyping 46XX | -4320 
enlarged left axillary lymph node | -1092 
left axillary and retroperitoneal adenopathy | -1092 
biopsy of left axillary lymph node | -1092 
follicular hyperplasia | -1092 
flow cytometry negative | -1092 
fine needle aspirate negative | -1092 
excisional biopsies negative | -1092 
COVID-19 vaccine administration | 0 
first dose | 0 
Pfizer-BioNTech COVID mRNA vaccine | 0 
mild arm soreness | 48 
easy bruising | 432 
gum bleeding | 432 
epistaxis | 432 
ecchymosis | 432 
petechiae | 432 
thrombocytopenia | 432 
platelet count 1000/mcL | 432 
prothrombin time 16.2 seconds | 432 
international normalized ratio 1.5 mg/dL | 432 
reticulocyte count 2.2% | 432 
lactate dehydrogenase 310 U/L | 432 
atypical lymphocytes | 432 
alkaline phosphatase 109 U/L | 432 
antinuclear antibody screen negative | 432 
dexamethasone | 432 
admitted to ICU | 432 
platelet transfusion | 432 
IVIG | 432 
CT scans | 432 
Sjogren’s SS-A antibody positive | 432 
ANA positive | 432 
Epstein-Barr virus DNA positive | 432 
hepatitis C negative | 432 
hepatitis B negative | 432 
HIV negative | 432 
thyroid-stimulating hormone negative | 432 
discharged | 456 
ITP diagnosed | -6480 
platelets 4000/mcL | -6480 
prednisone | -6480 
complete remission | -6480 
ITP flare-up | -4320 
platelets 3000/mcL | -4320 
human immune globulin | -4320 
dexamethasone | -4320 
direct platelet antibody level 1962 | -4320 
rheumatoid factor 20.7 IU/mL | -4320 
bone marrow biopsy | -4320 
karyotyping 46XX | -4320 
enlarged left axillary lymph node | -1092 
left axillary and retroperitoneal adenopathy | -1092 
biopsy of left axillary lymph node | -1092 
follicular hyperplasia | -1092 
flow cytometry negative | -1092 
fine needle aspirate negative | -1092 
excisional biopsies negative | -1092 
COVID-19 vaccine administration | 0 
first dose | 0 
Pfizer-BioNTech COVID mRNA vaccine | 0 
mild arm soreness | 48 
easy bruising | 432 
gum bleeding | 432 
epistaxis | 432 
ecchymosis | 432 
petechiae | 432 
thrombocytopenia | 432 
platelet count 1000/mcL | 432 
prothrombin time 16.2 seconds | 432 
international normalized ratio 1.5 mg/dL | 432 
reticulocyte count 2.2% | 432 
lactate dehydrogenase 310 U/L | 432 
atypical lymphocytes | 432 
alkaline phosphatase 109 U/L | 432 
antinuclear antibody screen negative | 432 
dexamethasone | 432 
admitted to ICU | 432 
platelet transfusion | 432 
IVIG | 432 
CT scans | 432 
Sjogren’s SS-A antibody positive | 432 
ANA positive | 432 
Epstein-Barr virus DNA positive | 432 
hepatitis C negative | 432 
hepatitis B negative | 432 
HIV negative | 432 
thyroid-stimulating hormone negative | 432 
discharged | 456 
ITP diagnosed | -6480 
platelets 4000/mcL | -6480 
prednisone | -6480 
complete remission | -6480 
ITP flare-up | -4320 
platelets 3000/mcL | -4320 
human immune globulin | -4320 
dexamethasone | -4320 
direct platelet antibody level 1962 | -4320 
rheumatoid factor 20.7 IU/mL | -4320 
bone marrow biopsy | -4320 
karyotyping 46XX | -4320 
enlarged left axillary lymph node | -1092 
left axillary and retroperitoneal adenopathy | -1092 
biopsy of left axillary lymph node | -1092 
follicular hyperplasia | -1092 
flow cytometry negative | -1092 
fine needle aspirate negative | -1092 
excisional biopsies negative | -1092 
COVID-19 vaccine administration | 0 
first dose | 0 
Pfizer-BioNTech COVID mRNA vaccine | 0 
mild arm soreness | 48 
easy bruising | 432 
gum bleeding | 432 
epistaxis | 432 
ecchymosis | 432 
petechiae | 432 
thrombocytopenia | 432 
platelet count 1000/mcL | 432 
prothrombin time 16.2 seconds | 432 
international normalized ratio 1.5 mg/dL | 432 
reticulocyte count 2.2% | 432 
lactate dehydrogenase 310 U/L | 432 
atypical lymphocytes | 432 
alkaline phosphatase 109 U/L | 432 
antinuclear antibody screen negative | 432 
dexamethasone | 432 
admitted to ICU | 432 
platelet transfusion | 432 
IVIG | 432 
CT scans | 432 
Sjogren’s SS-A antibody positive | 432 
ANA positive | 432 
Epstein-Barr virus DNA positive | 432 
hepatitis C negative | 432 
hepatitis B negative | 432 
HIV negative | 432 
thyroid-stimulating hormone negative | 432 
discharged | 456 
ITP diagnosed | -6480 
platelets 4000/mcL | -6480 
prednisone | -6480 
complete remission | -6480 
ITP flare-up | -4320 
platelets 3000/mcL | -4320 
human immune globulin | -4320 
dexamethasone | -4320 
direct platelet antibody level 1962 | -4320 
rheumatoid factor 20.7 IU/mL | -4320 
bone marrow biopsy | -4320 
karyotyping 46XX | -4320 
enlarged left axillary lymph node | -1092 
left axillary and retroperitoneal adenopathy | -1092 
biopsy of left axillary lymph node | -1092 
follicular hyperplasia | -1092 
flow cytometry negative | -1092 
fine needle aspirate negative | -1092 
excisional biopsies negative | -1092 
COVID-19 vaccine administration | 0 
first dose | 0 
Pfizer-BioNTech COVID mRNA vaccine | 0 
mild arm soreness | 48 
easy bruising | 432 
gum bleeding | 432 
epistaxis | 432 
ecchymosis | 432 
petechiae | 432 
thrombocytopenia | 432 
platelet count 1000/mcL | 432 
prothrombin time 16.2 seconds | 432 
international normalized ratio 1.5 mg/dL | 432 
reticulocyte count 2.2% | 432 
lactate dehydrogenase 310 U/L | 432 
atypical lymphocytes | 432 
alkaline phosphatase 109 U/L | 432 
antinuclear antibody screen negative | 432 
dexamethasone | 432 
admitted to ICU | 432 
platelet transfusion | 432 
IVIG | 432 
CT scans | 432 
Sjogren’s SS-A antibody positive | 432 
ANA positive | 432 
Epstein-Barr virus DNA positive | 432 
hepatitis C negative | 432 
hepatitis B negative | 432 
HIV negative | 432 
thyroid-stimulating hormone negative | 432 
discharged | 456 
ITP diagnosed | -6480 
platelets 4000/mcL | -6480 
prednisone | -6480 
complete remission | -6480 
ITP flare-up | -4320 
platelets 3000/mcL | -4320 
human immune globulin | -4320 
dexamethasone | -4320 
direct platelet antibody level 1962 | -4320 
rheumatoid factor 20.7 IU/mL | -4320 
bone marrow biopsy | -4320 
karyotyping 46XX | -4320 
enlarged left axillary lymph node | -1092 
left axillary and retroperitoneal adenopathy | -1092 
biopsy of left axillary lymph node | -1092 
follicular hyperplasia | -1092 
flow cytometry negative | -1092 
fine needle aspirate negative | -1092 
excisional biopsies negative | -1092 
COVID-19 vaccine administration | 0 
first dose | 0 
Pfizer-BioNTech COVID mRNA vaccine | 0 
mild arm soreness | 48 
easy bruising | 432 
gum bleeding | 432 
epistaxis | 432 
ecchymosis | 432 
petechiae | 432 
thrombocytopenia | 432 
platelet count 1000/mcL | 432 
prothrombin time 16.2 seconds | 432 
international normalized ratio 1.5 mg/dL | 432 
reticulocyte count 2.2% | 432 
lactate dehydrogenase 310 U/L | 432 
atypical lymphocytes | 432 
alkaline phosphatase 109 U/L | 432 
antinuclear antibody screen negative | 432 
dexamethasone | 432 
admitted to ICU | 432 
platelet transfusion | 432 
IVIG | 432 
CT scans | 432 
Sjogren’s SS-A antibody positive | 432 
ANA positive | 432 
Epstein-Barr virus DNA positive | 432 
hepatitis C negative | 432 
hepatitis B negative | 432 
HIV negative | 432 
thyroid-stimulating hormone negative | 432 
discharged | 456 
ITP diagnosed | -6480 
platelets 4000/mcL | -6480 
prednisone | -6480 
complete remission | -6480 
ITP flare-up | -4320 
platelets 3000/mcL | -4320 
human immune globulin | -4320 
dexamethasone | -4320 
direct platelet antibody level 1962 | -4320 
rheumatoid factor 20.7 IU/mL | -4320 
bone marrow biopsy | -4320 
karyotyping 46XX | -4320 
enlarged left axillary lymph node | -1092 
left axillary and retroperitoneal adenopathy | -1092 
biopsy of left axillary lymph node | -1092 
follicular hyperplasia | -1092 
flow cytometry negative | -1092 
fine needle aspirate negative | -1092 
excisional biopsies negative | -1092 
COVID-19 vaccine administration | 0 
first dose | 0 
Pfizer-BioNTech COVID mRNA vaccine | 0 
mild arm soreness | 48 
easy bruising | 432 
gum bleeding | 432 
epistaxis | 432 
ecchymosis | 432 
petechiae | 432 
thrombocytopenia | 432 
platelet count 1000/mcL | 432 
prothrombin time 16.2 seconds | 432 
international normalized ratio 1.5 mg/dL | 432 
reticulocyte count 2.2% | 432 
lactate dehydrogenase 310 U/L | 432 
atypical lymphocytes | 432 
alkaline phosphatase 109 U/L | 432 
antinuclear antibody screen negative | 432 
dexamethasone | 432 
admitted to ICU | 432 
platelet transfusion | 432 
IVIG | 432 
CT scans | 432 
Sjogren’s SS-A antibody positive | 432 
ANA positive | 432 
Epstein-Barr virus DNA positive | 432 
hepatitis C negative | 432 
hepatitis B negative | 432 
HIV negative | 432 
thyroid-stimulating hormone negative | 432 
discharged | 456 
ITP diagnosed | -6480 
platelets 4000/mcL | -6480 
prednisone | -6480 
complete remission | -6480 
ITP flare-up | -4320 
platelets 3000/mcL | -4320 
human immune globulin | -4320 
dexamethasone | -4320 
direct platelet antibody level 1962 | -4320 
rheumatoid factor 20.7 IU/mL | -4320 
bone marrow biopsy | -4320 
karyotyping 46XX | -4320 
enlarged left axillary lymph node | -1092 
left axillary and retroperitoneal adenopathy | -1092 
biopsy of left axillary lymph node | -1092 
follicular hyperplasia | -1092 
flow cytometry negative | -1092 
fine needle aspirate negative | -1092 
excisional biopsies negative | -1092 
COVID-19 vaccine administration | 0 
first dose | 0 
Pfizer-BioNTech COVID mRNA vaccine | 0 
mild arm soreness | 48 
easy bruising | 432 
gum bleeding | 432 
epistaxis | 432 
ecchymosis | 432 
petechiae | 432 
thrombocytopenia | 432 
platelet count 1000/mcL | 432 
prothrombin time 16.2 seconds | 432 
international normalized ratio 1.5 mg/dL | 432 
reticulocyte count 2.2% | 432 
lactate dehydrogenase 310 U/L | 432 
atypical lymphocytes | 432 
alkaline phosphatase 109 U/L | 432 
antinuclear antibody screen negative | 432 
dexamethasone | 432 
admitted to ICU | 432 
platelet transfusion | 432 
IVIG | 432 
CT scans | 432 
Sjogren’s SS-A antibody positive | 432 
ANA positive | 432 
Epstein-Barr virus DNA positive | 432 
hepatitis C negative | 432 
hepatitis B negative | 432 
HIV negative | 432 
thyroid-stimulating hormone negative | 432 
discharged | 456 
ITP diagnosed | -6480 
platelets 4000/mcL | -6480 
prednisone | -6480 
complete remission | -6480 
ITP flare-up | -4320 
platelets 3000/mcL | -4320 
human immune globulin | -4320 
dexamethasone | -4320 
direct platelet antibody level 1962 | -4320 
rheumatoid factor 20.7 IU/mL | -4320 
bone marrow biopsy | -4320 
karyotyping 46XX | -4320 
enlarged left axillary lymph node | -1092 
left axillary and retroperitoneal adenopathy | -1092 
biopsy of left axillary lymph node | -1092 
follicular hyperplasia | -1092 
flow cytometry negative | -1092 
fine needle aspirate negative | -1092 
excisional biopsies negative | -1092 
COVID-19 vaccine administration | 0 
first dose | 0 
Pfizer-BioNTech COVID mRNA vaccine | 0 
mild arm soreness | 48 
easy bruising | 432 
gum bleeding | 432 
epistaxis | 432 
ecchymosis | 432 
petechiae | 432 
thrombocytopenia | 432 
platelet count 1000/mcL | 432 
prothrombin time 16.2 seconds | 432 
international normalized ratio 1.5 mg/dL | 432 
reticulocyte count 2.2% | 432 
lactate dehydrogenase 310 U/L | 432 
atypical lymphocytes | 432 
alkaline phosphatase 109 U/L | 432 
antinuclear antibody screen negative | 432 
dexamethasone | 432 
admitted to ICU | 432 
platelet transfusion | 432 
IVIG | 432 
CT scans | 432 
Sjogren’s SS-A antibody positive | 432 
ANA positive | 432 
Epstein-Barr virus DNA positive | 432 
hepatitis C negative | 432 
hepatitis B negative | 432 
HIV negative | 432 
thyroid-stimulating hormone negative | 432 
discharged | 456 
ITP diagnosed | -6480 
platelets 4000/mcL | -6480 
prednisone | -6480 
complete remission | -6480 
ITP flare-up | -4320 
platelets 3000/mcL | -4320 
human immune globulin | -4320 
dexamethasone | -4320 
direct platelet antibody level 1962 | -4320 
rheumatoid factor 20.7 IU/mL | -4320 
bone marrow biopsy | -4320 
karyotyping 46XX | -4320 
enlarged left axillary lymph node | -1092 
left axillary and retroperitoneal adenopathy | -1092 
biopsy of left axillary lymph node | -1092 
follicular hyperplasia | -1092 
flow cytometry negative | -1092 
fine needle aspirate negative | -1092 
excisional biopsies negative | -1092 
COVID-19 vaccine administration | 0 
first dose | 0 
Pfizer-BioNTech COVID mRNA vaccine | 0 
mild arm soreness | 48 
easy bruising | 432 
gum bleeding | 432 
epistaxis | 432 
ecchymosis | 432 
petechiae | 432 
thrombocytopenia | 432 
platelet count 1000/mcL | 432 
prothrombin time 16.2 seconds | 432 
international normalized ratio 1.5 mg/dL | 432 
reticulocyte count 2.2% | 432 
lactate dehydrogenase 310 U/L | 432 
atypical lymphocytes | 432 
alkaline phosphatase 109 U/L | 432 
antinuclear antibody screen negative | 432 
dexamethasone | 432 
admitted to ICU | 432 
platelet transfusion | 432 
IVIG | 432 
CT scans | 432 
Sjogren’s SS-A antibody positive | 432 
ANA positive | 432 
Epstein-Barr virus DNA positive | 432 
hepatitis C negative | 432 
hepatitis B negative | 432 
HIV negative | 432 
thyroid-stimulating hormone negative | 432 
discharged | 456 
ITP diagnosed | -6480 
platelets 4000/mcL | -6480 
prednisone | -6480 
complete remission | -6480 
ITP flare-up | -4320 
platelets 3000/mcL | -4320 
human immune globulin | -4320 
dexamethasone | -4320 
direct platelet antibody level 1962 | -4320 
rheumatoid factor 20.7 IU/mL | -4320 
bone marrow biopsy | -4320 
karyotyping 46XX | -4320 
enlarged left axillary lymph node | -1092 
left axillary and retroperitoneal adenopathy | -1092 
biopsy of left axillary lymph node | -1092 
follicular hyperplasia | -1092 
flow cytometry negative | -1092 
fine needle aspirate negative | -1092 
excisional biopsies negative | -1092 
COVID-19 vaccine administration | 0 
first dose | 0 
Pfizer-BioNTech COVID mRNA vaccine | 0 
mild arm soreness | 48 
easy bruising | 432 
gum bleeding | 432 
epistaxis | 432 
ecchymosis | 432 
petechiae | 432 
thrombocytopenia | 432 
platelet count 1000/mcL | 432 
prothrombin time 16.2 seconds | 432 
international normalized ratio 1.5 mg/dL | 432 
reticulocyte count 2.2% | 432 
lactate dehydrogenase 310 U/L | 432 
atypical lymphocytes | 432 
alkaline phosphatase 109 U/L | 432 
antinuclear antibody screen negative | 432 
dexamethasone | 432 
admitted to ICU | 432 
platelet transfusion | 432 
IVIG | 432 
CT scans | 432 
Sjogren’s SS-A antibody positive | 432 
ANA positive | 432 
Epstein-Barr virus DNA positive | 432 
hepatitis C negative | 432 
hepatitis B negative | 432 
HIV negative | 432 
thyroid-stimulating hormone negative | 432 
discharged | 456 
ITP diagnosed | -6480 
platelets 4000/mcL | -6480 
prednisone | -6480 
complete remission | -6480 
ITP flare-up | -4320 
platelets 3000/mcL | -4320 
human immune globulin | -4320 
dexamethasone | -4320 
direct platelet antibody level 1962 | -4320 
rheumatoid factor 20.7 IU/mL | -4320 
bone marrow biopsy | -4320 
karyotyping 46XX | -4320 
enlarged left axillary lymph node | -1092 
left axillary and retroperitoneal adenopathy | -1092 
biopsy of left axillary lymph node | -1092 
follicular hyperplasia | -1092 
flow cytometry