73 years old | 0
    male | 0
    inoperable adenocarcinoma of the right lung | -8760
    concurrent chemoradiotherapy | -8760
    Salmonella Group D necrotising pneumonia | -6720
    empyema necessitans | -6720
    hospital admission for haemoptysis | 0
    purulent discharge | 0
    invasive pulmonary aspergillosis (IPA) suspected | 0
    persistent cavitation on CT thorax | 0
    elevated serum ß-D-glucan titre | 0
    positive serum galactomannan assay | 0
    Aspergillus niger growth in sputum | 0
    voriconazole 400 mg/day | 0
    cefoperazone-sulbactam | 0
    metronidazole | 0
    vancomycin | 0
    piperacillin-tazobactam | 0
    meropenem | 0
    acetaminophen (APAP) 4 g/day | 0
    intractable pain | 0
    acidotic breathing | 960
    severe metabolic acidosis | 960
    raised anion gap | 960
    no lactic acidosis | 960
    normal serum osmolal gap | 960
    no exposure to salicylate | 960
    no exposure to toxic alcohols | 960
    no exposure to glycols | 960
    moderately raised creatinine | 960
    moderately raised beta-hydroxybutyrate | 960
    elevated urine anion gap | 960
    pyroglutamic acidosis (PGA) suspected | 960
    APAP discontinued | 960
    intravenous N-acetylcysteine (NAC) infusion | 960
    transferred to ICU | 960
    acid–base imbalance improved | 960
    discharged from ICU | 1032
    urine pyroglutamic acid hyper-excretion confirmed | 1032
    massive haemoptysis | 1464
    death | 1464
    