78 years old | 0
male | 0
high-grade T1 urothelial carcinoma | -672
transurethral resection of bladder tumor | -672
intravesical BCG instillation | -336
fever | -24
rigors | -24
altered mental status | -24
shortness of breath | -24
denies cough | -24
denies chest pain | -24
no urinary symptoms | -24
no gastrointestinal symptoms | -24
BCG instillation | -24
temperature of 102.8 F | 0
pulse rate of 92/min | 0
respiratory rate of 40/min | 0
blood pressure 78/45 mmHg | 0
oxygen saturation of 93% | 0
toxic appearance | 0
dehydrated | 0
respiratory distress | 0
asymmetric chest expansion | 0
dullness to percussion | 0
decreased tactile fremitus | 0
reduced air entry on auscultation | 0
unremarkable cardiovascular examination | 0
leukocytosis | 0
white cell count of 27,200/microliter | 0
hemoglobin of 11.5 g/dL | 0
lactate of 7.8 meq/L | 0
high anion gap metabolic acidosis | 0
creatinine of 2.31 mg/dL | 0
blood urea nitrogen of 28 mg/dL | 0
normal oral flora on sputum culture | 0
negative urinary streptococcal and legionella antigens | 0
left basilar pneumonia | 0
small left pleural effusion | 0
no acute intracranial abnormalities on CT head | 0
negative preliminary blood culture | 0
intubation | 0
ventilation | 0
vasopressors | 0
intravenous Vancomycin | 0
intravenous Piperacillin-Tazobactam | 0
septic shock | 0
low-grade pyrexia | 24
failure to improve clinically | 24
suspicion for systemic BCG dissemination | 24
positive blood cultures for acid-fast bacilli | 48
discontinuation of broad-spectrum antibiotics | 48
triple therapy with Isoniazid, Ethambutol, and Rifampicin | 48
clinical improvement | 72
discharge | 120
planned follow-up with infectious disease team | 120
completion of 2 months of triple therapy | 2880
maintenance therapy with Rifampicin and Isoniazid | 4320