63 years old | 0
male | 0
recurrent abdominal adhesions | 0
multiple surgeries | 0
Abcarian stoma | 0
mucus fistula | 0
abdominal pain | -unknown
fever | -unknown
body temperature 36.8°C | 0
blood pressure 109/54 mmHg | 0
pulse rate 109 beats/min | 0
respiratory rate 18 breaths/min | 0
coarse breathing sounds | 0
regular heartbeats without murmur | 0
soft abdomen | 0
tenderness in right upper quadrant | 0
positive Murphy sign | 0
no palpable mass | 0
no hepatosplenomegaly | 0
mild anemia | 0
hemoglobin 10.6g/dl | 0
neutrophilic leukocytosis | 0
white blood cell count 28,000/ml | 0
C-reactive protein 100 mg/L | 0
troponin I 48 ng/L | 0
creatinine 176 umol/L | 0
urea 19 mmol/L | 0
normal electrolytes | 0
normal liver function tests | 0
normal serology | 0
normal urinalysis | 0
unremarkable chest X-ray | 0
unremarkable initial ECG | 0
thick gallbladder wall >3mm | 0
pericholecystic fluid | 0
gallbladder sludge | 0
cholelithiasis | 0
admission for sepsis secondary to acute cholecystitis | 0
antibiotics started | 0
supportive measures started | 0
continued fever | 24
hypotension | 24
ICU admission | 24
inotropic support | 24
retrosternal chest pain | 48
profuse sweating | 48
ST-segment elevation V2–V4 | 48
troponin-T 781 ng/L | 48
diagnosis of anterior wall ST-segment elevation myocardial infarction considered | 48
emergent coronary angiography | 48
nonobstructive CAD | 48
dilated left ventricular cavity | 48
apical dyskinesis | 48
preservation of basal to midseptal and basal-lateral wall contraction | 48
left ventricular ejection fraction 25% | 48
sepsis-induced Takotsubo cardiomyopathy diagnosis | 48
antibiotics continued | 48
conservative therapies | 48
recovery | 672
discharge | 240
repeated echocardiogram | 672
complete resolution of left ventricular systolic function | 672
ejection fraction >55% | 672
no obstructive coronary artery disease | 48
no acute plaque rupture | 48
no recent heart trauma | 48
no intracranial bleeding | 48
no pheochromocytoma | 48
no myocarditis | 48
no hypertrophic cardiomyopathy | 48
normotensive | 0
no palpitations | 0
no excessive diaphoresis | 0
no recent viral illness | 0
no cardiogenic shock | 48
no malignant arrhythmias | 48
intravenous hydration | 48
noradrenaline infusion | 48
empiric antibiotics | 48
uneventful hospital stay | 240
left ventricular function recovery within 4 weeks | 672
In the assistant's answer, they listed "abdominal pain | -unknown" and "fever | -unknown", which might be incorrect per the problem's instructions, which require approximation. Therefore, perhaps the correct approach is to assign these to 0, as they are part of the admission presentation.
