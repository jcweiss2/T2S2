39 years old | 0
male | 0
diabetes mellitus | -8760
dyslipidemia | -8760
admitted to the hospital | 0
abdominal pain | -24
nausea | -24
vomiting | -24
heart rate 81 per minute | 0
blood pressure 151/82 mmHg | 0
respiratory rate 20 per minute | 0
oxygen saturation 100% | 0
temperature 37.1°C | 0
distension in the epigastrium | 0
tenderness in the epigastrium | 0
elevated white cell count | 0
hyponatremia | 0
hyperglycemia | 0
lactic acidosis | 0
elevated creatinine | 0
lipase level 3500 U/L | 0
triglyceride level 3531 mg/dL | 0
denies binge drinking | 0
denies abdominal trauma | 0
denies recent change in medications | 0
denies recent procedures | 0
diffuse pancreatitis on CT scan | 0
hepatic steatosis on ultrasound | 0
no evidence of gall stones | 0
started on intravenous fluid resuscitation | 0
started on electrolyte management | 0
started on intravenous insulin drip | 0
intubated for respiratory failure | 72
tachypnea | 72
altered mental status | 72
worsening acidosis | 72
plasmapheresis initiated | 48
triglycerides improved | 96
initiated on hemodialysis | 96
renal failure | 96
elevated bladder pressures | 120
peak airway pressures | 120
emergent decompressive laparotomy | 120
serous ascitic fluid drained | 120
areas of saponification noted | 120
sepsis | 144
delirium | 144
renal function improved | 240
hemodialysis stopped | 240
discharged to home | 240
started on icosapent ethyl | 240
started on omega 3 fatty acids | 240
started on fenofibrate | 240