47 years old | 0
male | 0
admitted to ICU | 0
confirmed COVID-19 | -144
six-days history of shortness of breath | -144
hospitalization in COVID-19 ICU | -144
typical anginal pain | -48
hypertension | -672
fever | -288
six days of non-productive cough | -288
dyspnea | -288
progressive oxygen desaturation | -168
thorax CT revealed diffuse bilateral infiltrates | -168
ground glass opacities | -168
crazy paving with thickened interlobular septa | -168
consolidation in lower lobes | -168
treatment with enoxaparin sodium | -168
treatment with prednisolon | -168
treatment with moxifloksasin | -168
treatment with amlodipin | -168
treatment with favirapiravir | -240
treatment with ceftriaxone | -168
HFNO support | -48
blood pressure 135/68 mmHg | -48
heart rate 73 bpm | -48
oxygen saturation 88-93% | -48
body temperature 36.7°C | -48
normal cardiac examination | -48
inferior STEMI | -48
treatment with acetylsalicylic acid | -48
treatment with ticagrelor | -48
treatment with heparin | -48
cardiac symptoms decreased | -48
cardiac symptoms disappeared within 30 minutes | -48
coronary angiography showed 30-40% stenosis in LAD | -48
normal LMCA | -48
normal LCA | -48
normal RCA | -48
ST segment elevation regressed | -48
no ischemic cardiac symptoms after intervention | -48
hs-cTnI 0.012 ng/mL | -48
hs-cTnI 0.056 ng/mL | -48
normal kidney function tests | -48
normal liver function tests | -48
increased d-dimer | -48
increased fibrinogen | -48
increased ferritin | -48
increased lactate dehydrogenase | -48
increased C-reactive protein | -48
normal pro-brain natriuretic peptide | -48
CTPA no pulmonary embolism | -48
MINOCA diagnosis | -48
cardiogoniometry showed septal inferior myocardial ischemia | 24
medical treatment started | -48
transferred to normal medical ward | 72
discharged | 240
