49 years old | 0
male | 0
admitted to the hospital | 0
dry cough | -168
shortness of breath | -168
nausea | -168
vomiting | -168
tachypneic | 0
tachycardiac | 0
normotensive | 0
hypoxic | 0
oxygen saturation 64% | 0
tested positive for COVID-19 | 0
nasal cannula | 0
non-rebreather mask | 0
prone positioning | 0
oxygen saturation improved | 0
D-dimer level high | 0
subcutaneous enoxaparin | 0
therapeutic clinical trial of sarilumab | 0
methylprednisolone | 0
persistent tachycardia | 264
chest pain | 264
pulmonary embolism | 264
RV thrombus | 264
transferred to ICU | 264
dry cough | 336
increased work of breathing | 336
spiking fevers | 336
re-admitted to ICU | 480
respiratory condition worsened | 576
transferred to tertiary referral center | 576
COVID-19 pneumonia | 0
secondary bacterial infection | 336
reactivation | 480
relapse | 480
reinfection | 480
reverse transcription-polymerase chain reaction | 0
chest X-ray | 0
diffuse patchy bilateral pulmonary opacities | 0
repeat CXR | 240
extensive bilateral airspace disease | 240
CTPA | 264
right lower lobe PE | 264
echocardiogram | 264
dilated right ventricle | 264
mobile echo density | 264
thrombolytic therapy | 264
repeat echocardiogram | 336
resolution of RV thrombus | 336
CTPA and venous duplex ultrasound | 336
no evidence of new thrombus | 336
deteriorated clinically | 480
repeat echocardiogram | 480
second RV thrombus | 480
left gastrocnemius vein DVT | 480
empiric broad-spectrum antibiotics | 504
cytokine storm | 504
tocilizumab | 504
transferred to advanced care facility | 576
venovenous extracorporeal membrane oxygenation | 576
respiratory condition worsened | 600
percutaneous thrombectomy | 600
tracheostomy | 912
decannulated | 1368
septic shock | 1692
percutaneous endoscopic gastrostomy tube placement | 2232
discharged | 2976
passed away | 3000