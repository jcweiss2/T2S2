38 years old | 0
male | 0
admitted to the hospital | 0
warm, swollen, painful right knee | -1314
redness | -1314
car accident | -1344
craniocerebral trauma | -1344
coma | -1344
intracranial hypertension | -1344
temporary ventricular drainage | -1344
sepsis with Klebsiella Pneumoniae | -1344
sepsis with Pseudomonas Aeruginosa | -1344
multi-organ failure | -1344
swelling of the right knee | -728
rehabilitation | -728
no evidence of infection in the synovial fluid | -728
referred for further diagnosis | -728
warm, swollen, painful right knee | 0
no redness | 0
no other joints involved | 0
normal body temperature | 0
normal clinical examination | 0
arthrocentesis of the knee | 0
white blood cell count (WBC) of 57000 | 0
90% neutrophils | 0
negative cultures | 0
no crystals in the fluid | 0
elevated C-reactive protein (CRP 43 mg/L) | 0
elevated blood WBC of 11.500 /mm³ | 0
negative rheumatoid factor | 0
negative anti-CCP antibodies | 0
negative anti-nuclear factor | 0
negative Borellia antibodies | 0
negative Chlamydia Trachomatis PCR | 0
negative Neisseria Gonorrhoeae PCR | 0
magnetic resonance imaging of the knee | 0
no major cartilage problems | 0
no meniscal or ligamental lesions | 0
bony infarctions in femur and tibia | 0
needle arthroscopy | 24
hyperemic and very hypertrophic synovium | 24
white film | 24
biopsies of synovial tissue | 24
important inflammation | 24
high amount of neutrophils | 24
direct cultures of the synovial tissue | 24
Staphylococcus Warneri | 24
resistant only to penicillin | 24
negative PCR for Borrelia | 24
negative PCR for mycobacteria genus | 24
negative PCR for mycobacterium complex | 24
treatment with Levofloxacin | 24
clear improvement | 408
persisting swelling of the knee | 408
repeated needle arthroscopy | 408
decreased inflammatory infiltrate | 408
synovial fluid | 408
3.810 WBC | 408
38% neutrophils | 408
CRP dropped | 408
discharged | 504