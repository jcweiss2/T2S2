48 years old | 0
male | 0
admitted to the emergency department | 0
cough | -96
dyspnea | -96
fever | -48
highest temperature of 39.3°C | -48
yellowish sputum | -48
chills | -48
sweats | -48
denied hemoptysis | -48
oral cefixime | -48
diclofenac sodium | -48
no effect | -48
good health | 0
no history of hypertension | 0
no history of diabetes | 0
no history of stroke | 0
no history of myocardial infarction | 0
no prior illnesses | 0
no hospitalizations | 0
no known drug allergies | 0
living in Chengdu | 0
no tobacco | 0
no alcohol | 0
no drug abuse | 0
married | 0
three healthy daughters | 0
family history negative for genetic disease | 0
body temperature 40.0°C | 0
heart rate 130 beats/min | 0
breathing rate 41 breaths/min | 0
blood pressure 111/59 mmHg | 0
oxygen saturation (SpO2) of 93% | 0
Chest computed tomography (CT) | 0
diffuse, bilateral, and interstitial infiltrates | 0
white blood cell (WBC) count of 6.88×10^9/L | 0
neutrophil percentage was 85.4% | 0
lymphocyte percentage 11.0% | 0
erythrocyte sedimentation rate (ESR) 23 mm/h | 0
concentration of procalcitonin (PCT) 0.12 ng/mL | 0
prothrombin time (PT) 12.5 s | 0
international normalized ratio (INR) 1.16 | 0
fibrinogen (Fbg) 7.01 g/L | 0
thrombin time (TT) 148 s | 0
D-dimer (D2) 1.66 µg/mL | 0
fibrin degradation products (FDP) 6.80 µg/mL | 0
blood gas analysis | 0
pH 7.492 | 0
PCO2 36 mmHg | 0
PO2 60.4 mmHg | 0
oxygenation index of 234 mmHg | 0
electrolytes | 0
renal function | 0
myocardial injury markers | 0
tumor markers | 0
infection markers | 0
Chlamydia pneumoniae | 0
Mycoplasma pneumoniae | 0
respiratory failure | 24
transferred to the intensive care unit | 24
mechanical ventilation | 24
supportive care | 24
moxifloxacin | 24
piperacillin tazobactam | 24
oseltamivir | 24
fever continued | 48
pulmonary infection | 48
repeat CT scan | 48
moxifloxacin replaced with linezolid | 72
meropenem | 72
fever subsided | 96
other symptoms and signs persisted | 96
WBC count | 96
PCT | 96
inflammatory activity | 96
inspiratory crackles | 96
C-reactive protein (CRP) | 120
ESR | 120
PCT | 120
all of the tests for viruses were negative | 120
influenza A and B virus | 120
cytomegalovirus | 120
Toxoplasma | 120
Epstein–Barr virus | 120
rubella virus | 120
herpes simplex virus | 120
Cryptococcal antigen | 120
galactomannan test | 120
β-D-glucan test | 120
anti-nuclear antibody | 120
anti-extractable nuclear antigen antibody | 120
anti-neutrophilic cytoplasmic antibody | 120
peripheral blood cultures | 120
contact with domestic pigeons | 120
unbiased metagenomic next-generation sequencing (mNGS) | 120
bronchoalveolar lavage fluid (BALF) | 120
C. psittaci infection | 120
doxycycline | 168
moxifloxacin | 168
meropenem | 168
empirical antiviral agents ceased | 168
PCT and WBC count continued to decline | 168
fever finally returned to normal | 360
acrocyanosis of both lower extremities | 72
palpable purpura | 72
left dorsalis pedis artery occlusion | 72
right peroneal vein thrombosis | 72
amputation of both legs | 360
multiple organ failure | 360
repatriated for further rehabilitation | 360
one-year follow-up | 8760
doing well | 8760
no further symptoms | 8760