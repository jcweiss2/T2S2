54 years old | 0
male | 0
admitted to the hospital | 0
fever | -168
cough | -168
dyspnea | -168
syncope | -168
nausea | -168
vomiting | -168
diarrhea | -168
smoking history | -8760
exposure to SARS-CoV-2 | -168
COVID-19 diagnosis | 0
SARS-CoV-2 positive | 0
lymphopenia | 0
elevated lactate dehydrogenase | 0
elevated ferritin | 0
elevated D-dimer | 0
elevated inter-leukin-6 | 0
elevated troponin-I | 0
bilateral alveolar infiltrates | 0
S1Q3T3 pattern on electrocardiogram | 0
ARDS | 1
septic shock | 1
intubation | 1
mechanical ventilation | 1
norepinephrine | 1
tricuspid valve thrombus | 1
right ventricle thrombus | 1
LMWH | 1
enoxaparin | 1
hydroxychloroquine | 1
azithromycin | 1
tocilizumab | 1
tracheostomy | 336
percutaneous endoscopic gastrostomy tube placement | 336
discharged | 624
apixaban | 624
follow-up transthoracic echocardiogram | 168
thrombus dissolution | 168