48 years old | 0
    man | 0
    presented to hospital | 0
    transpelvic gunshot wound | 0
    right lower quadrant of the abdomen | 0
    hemodynamically unstable | 0
    blood pressure 82/63 mm Hg | 0
    heart rate 120 bpm | 0
    exploratory laparotomy | 0
    small bowel injury | 0
    rectosigmoid injury | 0
    multiple areas of hemorrhage | 0
    resection of affected small bowel and rectosigmoid | 0
    small bowel anastomosed | 0
    colostomy created | 0
    rectal stump created | 0
    admitted to intensive care unit | 0
    ongoing medical care | 0
    day 13 | 312
    coffee-ground output from nasogastric tube | 312
    hemoglobin drop from 8.9 to 7.1 g/dL | 312
    transfusion of 2 units packed red blood cells | 312
    esophagogastroduodenoscopy performed | 312
    large ulcer at stomach body and fundus | 312
    irregular ulcer borders | 312
    vessel at ulcer edge | 312
    greyish coating in ulcer bed | 312
    exudate in ulcer bed | 312
    tissue biopsy obtained | 312
    intravenous pantoprazole initiated | 312
    oral sucralfate initiated | 312
    36 hours later | 336
    tissue pathology results revealed necrotic exudate with fungal aseptate hyphae | 336
    diagnosis of invasive gastric mucormycosis | 336
    intravenous liposomal amphotericin initiated | 336
    no further bleeding | 336
    stabilization of hemoglobin | 336
    no surgical intervention | 336
    day 15 | 360
    necrotic area at open left flank wound | 360
    sepsis development | 360
    white blood cell count 23,000/µL | 360
    heart rate 120 bpm | 360
    lactic acid level 4.4 mmol/L | 360
    broad-spectrum intravenous antibiotics initiated | 360
    vancomycin initiated | 360
    piperacillin-tazobactam initiated | 360
    repeat exploratory laparotomy | 360
    multifocal necrotic bowel around small bowel anastomosis and rectal stump | 360
    areas of perforation around anastomotic site | 360
    debridement of areas | 360
    resection of necrotic bowel | 360
    histopathological evaluation of resected specimen revealed fungal aseptate hyphae | 360
    day 17 | 408
    bloody output from nasogastric tube | 408
    bloody output from abdominal surgical drains | 408
    hemorrhagic shock development | 408
    refractory to blood transfusion | 408
    refractory to intravenous hydration | 408
    refractory to inotrope therapy | 408
    immediate laparotomy performed | 408
    8x4 cm perforation with necrosis at gastric ulcer site | 408
    active bleeding | 408
    unsuccessful control of bleeding | 408
    patient died | 408

    48 years old | 0
    man | 0
    presented to hospital | 0
    transpelvic gunshot wound | 0
    right lower quadrant of the abdomen | 0
    hemodynamically unstable | 0
    blood pressure 82/63 mm Hg | 0
    heart rate 120 bpm |6
    exploratory laparotomy |0
    small bowel injury |0
    rectosigmoid injury |0
    multiple areas of hemorrhage |0
    resection of affected small bowel and rectosigmoid |0
    small bowel anastomosed |0
    colostomy created |0
    rectal stump created |0
    admitted to intensive care unit |0
    ongoing medical care |0
    day 13 |312
    coffee-ground output from nasogastric tube |312
    hemoglobin drop from 8.9 to 7.1 g/dL |312
    transfusion of 2 units packed red blood cells |312
    esophagogastroduodenoscopy performed |312
    large ulcer at stomach body and fundus |312
    irregular ulcer borders |312
    vessel at ulcer edge |312
    greyish coating in ulcer bed |312
    exudate in ulcer bed |312
    tissue biopsy obtained |312
    intravenous pantoprazole initiated |312
    oral sucralfate initiated |312
    36 hours later |336
    tissue pathology results revealed necrotic exudate with fungal aseptate hyphae |336
    diagnosis of invasive gastric mucormycosis |336
    intravenous liposomal amphotericin initiated |336
    no further bleeding |336
    stabilization of hemoglobin |336
    no surgical intervention |336
    day 15 |360
    necrotic area at open left flank wound |360
    sepsis development |360
    white blood cell count 23,000/µL |360
    heart rate 120 bpm |360
    lactic acid level 4.4 mmol/L |360
    broad-spectrum intravenous antibiotics initiated |360
    vancomycin initiated |360
    piperacillin-tazobactam initiated |360
    repeat exploratory laparotomy |360
    multifocal necrotic bowel around small bowel anastomosis and rectal stump |360
    areas of perforation around anastomotic site |360
    debridement of areas |360
    resection of necrotic bowel |360
    histopathological evaluation of resected specimen revealed fungal aseptate hyphae |360
    day 17 |408
    bloody output from nasogastric tube |408
    bloody output from abdominal surgical drains |408
    hemorrhagic shock development |408
    refractory to blood transfusion |408
    refractory to intravenous hydration |408
    refractory to inotrope therapy |408
    immediate laparotomy performed |408
    8x4 cm perforation with necrosis at gastric ulcer site |408
    active bleeding |408
    unsuccessful control of bleeding |408
    patient died |408