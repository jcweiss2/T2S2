44 years old | 0
male | 0
admitted to the emergency room | 0
weakness | -48
physical deconditioning | -48
type I diabetes mellitus | 0
peptic ulcer disease | 0
depression |: 0
seizure disorder | 0
Charcot foot of the left foot | 0
mild developmental delay | 0
insulin detemir | 0
escitalopram | 0
depakote | 0
clonazepam | 0
gabapentin | 0
levetiracetam | 0
lisinopril | 0
finasteride | 0
non-compliance to medications | 0
previous hospital admissions for diabetic ketoacidosis | 0
substance abuse with tobacco | 0
seven pack-years of smoking | 0
alcohol consumption | 0
occasional use of marijuana | 0
diabetic ketoacidosis | 0
acute kidney injury | 0
drug-induced acute tubular necrosis | 0
dehydration | 0
hyperkalemia | 0
intravenous fluids | 0
insulin infusion | 0
DKA resolved | 0
blood culture positive for MSSA | 0
vancomycin | 0
renal adjusted dose of piperacillin/tazobactam | 0
persistent positive blood cultures with MSSA | 0
chronic fracture of left humerus proximally | 0
non-union fracture for 1 year | 0
limited range of movements | 0
orthopedic consultation | 0
CT scan of upper extremity | 0
osteomyelitis | 0
large septated fluid collections in subcutaneous soft tissues and muscles | 0
seromas related to old hemorrhage | 0
incision and drainage | 0
drains placed | 0
culture of fluid drained grew MSSA | 0
septicemia | 0
localized abscess | 0
cardiac transthoracic echo | 0
transesophageal echocardiography | 0
benzocaine | 0
lidocaine | 0
persistent hypoxemia | 0
oxygen saturation 85-87% on 100% non-rebreather mask | 0
arterial blood gas pH 7.43 | 0
arterial blood gas PCO2 41 | 0
arterial blood gas PO2 249 | 0
oxygen saturation 85% | 0
no cyanosis | 0
arterial blood color not noted | 0
chest X-ray no abnormalities | 0
CT angiogram of chest no evidence of pulmonary embolism | 0
probable diagnosis of methemoglobinemia | 0
methemoglobin level 28.6% | 0
methylene blue 2 mg/kg IV | 0
oxygen saturation 92-94% on 2 L nasal cannula | 2
repeat methemoglobin levels 8.2% | 2
hypoxia improved | 2
good saturation on room air | 2
repeat blood cultures negative | 48
medical condition improved | 0
discharged | 0
IV antibiotics | 0
skilled nursing facility | 0
