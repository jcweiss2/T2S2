71 years old | 0
male | 0
admitted to the hospital | 0
rectal bleeding | 0
denied abdominal pain | 0
denied nausea | 0
denied vomiting | 0
denied hematemesis | 0
denied previous history of gastrointestinal bleeding | 0
cirrhosis of the liver | -672
alcohol use | -672
hypertension | -672
coronary artery disease | -672
atrial fibrillation | -672
systolic congestive heart failure | -672
coronary artery bypass surgery | -168
not taking warfarin | 0
pallor | 0
hemodynamically stable | 0
nasogastric aspiration clear | 0
rectal examination revealed maroon-colored blood | 0
admitted to the intensive care unit | 0
initial hematocrit 11% | 0
received more than 6 units of packed red blood cells | 0
hematocrit 18% | 0
emergency endoscopy | 2
emergency colonoscopy | 2
bowel cleansing with polyethylene glycol | 1
upper gastrointestinal endoscopy revealed two clean based cratered ulcers in the duodenal bulb | 2
no blood in the upper gastrointestinal tract | 2
colonoscopy revealed large amount of fresh and altered blood with clots in the entire colon | 2
no lesion identified to explain the bleeding | 2
exploratory laparotomy | 4
two irregular appearing areas in the ascending colon | 4
right hemicolectomy | 4
MALT lymphoma | 4
marginal zone cells infiltrating the lamina propria | 4
immunohistochemical stains showed cells reactive to CD20, CD43 and BCL-2 antibodies | 4
nonreactive to cyclin D1, CD3, CD5, CD10, and BCL-6 antibodies | 4
H. pylori negative | 4
hematology/oncology team evaluated the patient | 8
staging work-up planned | 8
developed sepsis | 120
expired two weeks after surgery | 336