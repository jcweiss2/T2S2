52 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
body mass index 23.6 kg/m2 | 0 | 0 | Factual
no comorbidities | 0 | 0 | Factual
open modified Scopinaro procedure | -7440 | -7440 | Factual
initial weight 216 kg | -7440 | -7440 | Factual
BMI 57.4 kg/m2 | -7440 | -7440 | Factual
weight reganance | -2400 | 0 | Factual
incisional hernia | -2400 | 0 | Factual
bariatric revisional surgery | -168 | -168 | Factual
hernia repair | -168 | -168 | Factual
weight 170 kg | -168 | -168 | Factual
BMI 45.1 | -168 | -168 | Factual
gastric pouch leak | -168 | -168 | Factual
intra-abdominal collections | -168 | -168 | Factual
sepsis | -168 | -168 | Factual
conservative management | -168 | 0 | Factual
open abdomen | -168 | 0 | Factual
negative wound pressure therapy | -168 | 0 | Factual
parenteral nutrition | -168 | 0 | Factual
intravenous antibiotics | -168 | 0 | Factual
epithelized gastrocutaneous fistula | -72 | 0 | Factual
controlled but persistent drainage | -72 | 0 | Factual
upper endoscopy | -72 | -72 | Factual
fistulous orifice | -72 | -72 | Factual
extraluminal extravasation | -72 | -72 | Factual
recurrent left subphrenic abscess | -72 | -72 | Factual
endoscopic treatment | -72 | 0 | Factual
argon plasma coagulation | -72 | -72 | Factual
internal and external drainages | -72 | -72 | Factual
clipping | -72 | -72 | Factual
fibrin sealants | -72 | -72 | Factual
e-vac therapy | -72 | -72 | Factual
stenting | -72 | -72 | Factual
multidisciplinary team discussion | 0 | 0 | Factual
decision to proceed with innovative endoscopic technique | 0 | 0 | Factual
placement of CSDO | 0 | 0 | Factual
Occlutech muscular VSD occluder | 0 | 0 | Factual
procedure performed in catheterization laboratory | 0 | 0 | Factual
intravenous sedation | 0 | 0 | Factual
topic anesthesia | 0 | 0 | Factual
fistula cannulated | 0 | 0 | Factual
extraluminal leakage documented | 0 | 0 | Factual
Amplatz extra stiff guidewire | 0 | 0 | Factual
delivery system introduced | 0 | 0 | Factual
CSDO deployed | 0 | 0 | Factual
no immediate adverse events | 0 | 0 | Factual
contrast study | 0 | 0 | Factual
no extravasation of contrast material | 0 | 0 | Factual
restricted oral intake | 0 | 24 | Factual
liquid diet | 24 | 240 | Factual
regular diet | 240 | 240 | Factual
10-15cc remaining daily drainage | 240 | 432 | Factual
pigtail displaced | 432 | 432 | Factual
systemic signs of sepsis | 432 | 432 | Factual
computed tomography | 432 | 432 | Factual
fluoroscopy | 432 | 432 | Factual
recurrence of abscess | 432 | 432 | Factual
partial dislodgment of CSDO | 432 | 432 | Factual
second attempt with oversized disc | 432 | 432 | Factual
Occlutech Figulla Flex II UNI 24-mm | 432 | 432 | Factual
device sealed fistulous orifice | 432 | 432 | Factual
6-month clinical and imaging follow-up | 1296 | 1296 | Factual
upper endoscopy | 1296 | 1296 | Factual
contrast-enhanced CT scan | 1296 | 1296 | Factual
device engrafted | 1296 | 1296 | Factual
significant reduction of chronic abscess | 1296 | 1296 | Factual
no signs of fistula recurrence | 1296 | 1296 | Factual
pigtail removed | 1296 | 1296 | Factual
no drainage observed | 1296 | 1296 | Factual