67 years old | 0
female | 0
admitted to the intensive care unit | 0
chronic back pain | -2160
obesity | 0
hypertension | 0
gastritis | 0
HSV1 | 0
tobacco use | 0
prednisone | -2160
desaturated to SpO2 of 85% | 24
oxygenation improved with continuous positive airway pressure | 24
chest X-ray bilateral lower lobe infiltrates | 24
glucocorticoid taper with dexamethasone and hydrocortisone | 0
hydrocortisone 100 mg | 0
dexamethasone 10 mg twice daily | 24
dexamethasone 8 mg twice daily | 48
dexamethasone 6 mg | 24
hydrocortisone 50 mg every 6 hours | 72
hydrocortisone 25 mg every 6 hours | 96
acute kidney injury | 48
febrile episodes | 48
vancomycin initiated | 48
piperacillin–tazobactam initiated | 48
hemodynamically unstable | 120
hypercapnic respiratory failure | 120
intubated | 120
norepinephrine initiated | 120
hemodialysis initiated | 120
white blood cell count doubled | 144
procalcitonin elevated | 144
repeat cultures sent | 144
vancomycin continued | 144
meropenem initiated | 144
chest X-ray acute respiratory distress syndrome | 144
Candida albicans in blood | 144
Candida albicans in urine | 144
Candida albicans in sputum | 144
fluconazole initiated | 144
immunosuppression concerns | 144
β-D-Glucan not performed | 144
sputum negative for Pneumocystis jirovecii | 144
immunostaining HSV positive | 144
disseminated HSV1 infection confirmed | 144
acyclovir initiated | 144
history of oral HSV1 | 144
recurrent oral infections | 144
bloody output from orogastric tube | 360
esophagogastroduodenoscopy performed | 360
diffuse esophageal ulcerations | 360
gastric ulcerations | 360
HSV esophagitis | 360
improving clinically | 360
vasopressors discontinued | 360
extubated | 360
transferred out of ICU | 672
renal function improvement | 672
dialysis discontinued | 672
discharged | 936
