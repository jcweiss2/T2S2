81 years old | 0  
    woman | 0  
    transferred to Neurocritical Care Unit | 0  
    severe encephalopathy | 0  
    right frontal mass | 0  
    coronary artery disease | -8760  
    stent placement | -8760  
    type 2 diabetes mellitus | 0  
    endometrial carcinoma | -262080  
    hysterectomy | -262080  
    chemotherapy | -262080  
    aseptic meningitis | -175200  
    syncope | -168  
    seizure | -168  
    dysarthria | -168  
    runny nose | -168  
    nausea | -168  
    diarrhea | -168  
    ciprofloxacin | -168  
    rapid deterioration of neurological status | -168  
    profound lethargy | -168  
    bilateral weakness | -168  
    right-sided weakness | -168  
    left-sided weakness | -168  
    cranial nerve abnormalities | -168  
    viral encephalitis | -168  
    acyclovir | -168  
    brain CT | -168  
    chest CT | -168  
    abdomen CT | -168  
    pelvis CT | -168  
    afebrile | 0  
    stable vital signs | 0  
    stuporous | 0  
    opens eyes to painful stimuli | 0  
    attempts to localize with left upper extremity | 0  
    not following commands | 0  
    nonverbal | 0  
    left gaze preference | 0  
    anisocoric pupils | 0  
    left pupil 6 mm | 0  
    right pupil 4 mm | 0  
    reactive pupils | 0  
    right upper extremity flaccid | 0  
    right lower extremity flaccid | 0  
    no response to painful stimuli | 0  
    minimal withdrawal in left lower extremity | 0  
    hyponatremia | 0  
    sodium level 131 | 0  
    hyperglycemia | 0  
    glucose 248 | 0  
    mild anemia | 0  
    Hgb 11 | 0  
    brain MRI | 0  
    high FLAIR signal | 0  
    tubular/lobulated/ring enhancement | 0  
    bifrontal regions | 0  
    left anterior midbrain | 0  
    multicentric glioma | 0  
    multicentric primary CNS lymphoma | 0  
    lumbar puncture | 0  
    CSF studies | 0  
    bacterial etiology | 0  
    viral etiology | 0  
    fungal etiology | 0  
    normal CSF chemical profile | 0  
    mildly elevated protein level 78 | 0  
    brain abscesses | 0  
    empiric antimicrobial treatment | 0  
    ampicillin | 0  
    meropenem | 0  
    vancomycin | 0  
    voriconazole | 0  
    pyrimethane/sulfadiazine | 0  
    intravenous dexamethasone | 0  
    open brain biopsy | 72  
    Gram-positive rods | 72  
    L. monocytogenes infection | 72  
    antibiotics discontinued | 72  
    steroids tapered off | 240  
    transferred to regular floor | 240  
    percutaneous endoscopic gastrostomy | 240  
    unable to swallow safely | 240  
    transferred to rehabilitation facility | 768  
    neurological examination improvement | 768  
    eye opening to verbal stimuli | 768  
    command-following with left upper extremity | 768  
    incomprehensible sounds | 768  
    pupils 4 mm bilaterally | 768  
    reactive pupils | 768  
    partial left third cranial nerve palsy | 768  
    left nasolabial fold flattening | 768  
    persistent right upper extremity weakness | 768  
    persistent right lower extremity weakness | 768  
    persistent left lower extremity weakness | 768  
    minimal withdrawal to pain | 768  
    <|eot_id|>
    