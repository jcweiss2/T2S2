32 years old | 0
female | 0
fever | -720
cough | -216
hoarseness of voice | -168
odynophagia | -168
ectopic pregnancy | -280
ruptured ectopic pregnancy | -274
admitted to the hospital | -274
laparoscopic exploration | -274
Mycobacterium tuberculosis | -274
sepsis | -274
adult respiratory distress syndrome | -274
central line placed | -274
Pseudomonas aeruginosa | -274
Enterobacter cloacae | -274
pulmonary tuberculosis | -274
antibiotics started | -274
anti-TB medications started | -274
discharged home | -264
vomiting | -128
headache | -128
exertional dyspnea | -128
inability to talk | -128
difficulty opening left eye | -128
weight loss | -128
disseminated central nervous system TB | -128
anti-TB regimen adjusted | -128
left-sided hemiparesis | -128
recovered | -126
discharged home | -126
hoarseness of voice | 0
odynophagia | 0
superior mediastinal mass | 0
CT scan | 0
large subclavian artery pseudoaneurysm | 0
CT angiogram | 0
compression effects on trachea, esophagus, and recurrent laryngeal nerves | 0
radial artery blood pressures on the right side higher than that on the left | 0
preoperative diagnosis | 0
left subclavian artery pseudoaneurysm | 0
repair of the aneurysm | 24
left posterolateral thoracotomy incision | 24
pleural adhesions excised | 24
pericardial patch used | 24
histopathology | 24
chronic granulomatous inflammation | 24
necrosed tissue | 24
uneventful recovery | 168
discharged | 168
followed for 2 months | 216
doing well | 216