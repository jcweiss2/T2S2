48 years old | 0
    male | 0
    admitted to the Emergency Service | 0
    toothache | -96
    dyspnea | -96
    chest pain | -96
    sweating | -96
    tachyarrhythmia | -96
    sore throat | -96
    fever (38.2°C) | -96
    gross swelling of the lower right cheek | 0
    swelling of the submandibular region | 0
    swelling of the mental region | 0
    erythematous and warm on palpation | 0
    difficulties in opening the jaw | 0
    inflammatory changes of the oral cavity mucous membrane | 0
    treatment with ceftriaxone-steroids-based 3 g once daily | -96 (assuming started at the beginning of the 4-day history)
    ineffective treatment | -72 (assuming treatment started 24 hours after onset)
    condition worsened | -72
    dyspnea | -72
    chest pain | -72
    increase in white blood cells (WBC = 17 × 10^9/L) | 0
    increase in neutrophils (88%) | 0
    increase in C-reactive protein (4 mg/L) | 0
    urgent orotracheal intubation | 0
    chest and neck CT scan showing left pleural effusion | 0
    mediastinitis | 0
    right parapharyngeal abscess | 0
    possible complication of odontogenic infection | 0
    drainage of the right neck by cervicotomy | 0
    placement of left chest drain on the left sixth intercostal space | 0
    initiation of intravenous piperacillin sodium plus tazobactam sodium (4 × 500 mg die) | 0
    clinical condition worsened | 48 (after 2 days from admission)
    transfer to Intensive Care Unit | 48
    chest and neck CT scan demonstrating air collections in right submandibular, left carotid, retroesophageal, and pretracheal spaces | 48
    air and fluid collections in upper, anterior, and posterior mediastinum | 48
    diagnosis of cervical necrotizing fasciitis with DNM | 48
    insertion of additive pleural drain on the right side | 48
    chest and neck CT angiography showing abscesses in cervical spaces | 72 (after 1 day from previous CT)
    extensive mediastinal empyema | 72
    left pleural effusion | 72
    right hydropneumothorax | 72
    aggressive mediastinal debridement | 72
    VATS performed | 72
    incision and drainage of neck abscesses | 72
    insertion of 2 surgical drains | 72
    oral tooth extraction (48th) | 72
    drainage and packing of purulent fluid by maxillofacial surgical team | 72
    microscopy and culture revealing Streptococcus anginosus | 72
    microscopy and culture revealing Gemella morbillorum | 72
    microscopy and culture revealing Staphylococcus lugdunensis | 72
    initiation of amoxicillin 1000 mg intravenously 6 hourly | 72
    initiation of metronidazole 500 mg intravenously 12 hourly | 72
    dismissal in better health conditions | 168 (1 week later)
    