62 years old | 0
woman | 0
primary progressive multiple sclerosis | 0
acute altered level of consciousness | 0
hypoxemia | 0
shock | 0
tested positive for severe acute respiratory syndrome coronavirus-2 | -168
blood pressure 55/32 mm Hg | 0
heart rate 120 beats/min | 0
respiratory rate 32 breaths/min | 0
oxygen saturation 95% on 100% oxygen | 0
dense airspace opacities in the right lung | 0
ground-glass opacity in the left lung | 0
sinus tachycardia | 0
diffuse anterolateral ST-elevation | 0
high-sensitivity cardiac Troponin T 4986 ng/L | 0
N-terminal pro-B-type natriuretic peptide 51,439 ng/L | 0
ferritin 3067 U/L | 0
C-reactive protein 68.2 mg/L | 0
D-dimer 6920 ng/mL |"0
lactate dehydrogenase 1094 U/L | 0
lactate 2.4 mmol/L | 0
creatinine 252 umol/L | 0
blood cultures negative | 0
sputum cultures negative | 0
resuscitated with intravenous fluids | 0
intravenous dexamethasone | 0
ceftriaxone | 0
azithromycin | 0
no intubation | 0
no inotropes | 0
severe left ventricular dysfunction | 0
lung ultrasound findings consistent with pneumonia | 0
urgent cardiac magnetic resonance imaging | 24
global hypokinesia | 24
relative sparing of the basal segments | 24
extensive sub-epicardial late gadolinium enhancement in the anterolateral and inferolateral left ventricular walls | 24
elevation in tissue mapping-based markers of inflammatory injury | 24
elevated native T1 | 24
elevated native T2 | 24
marked expansion of the extracellular volume | 24
left ventricular ejection fraction 24% | 24
anakinra administered intravenously 100 mg twice daily | 24
rapid clinical improvement during the following 72 hours | 72
reduced oxygen requirements | 72
improved blood pressure | 72
reduction in heart rate | 72
anakinra treatment continued for 5 days | 24
renal function improved | 72
progressive reduction in inflammatory markers | 72
alert | 72
hemodynamically stable | 72
required 1 liter of supplemental oxygen | 72
repeat CMR imaging on day 14 | 336
left ventricular ejection fraction improved from 24% to 54% | 336
reduction in late gadolinium enhancement signal intensity | 336
global reductions in myocardial T1 | 336
global reductions in myocardial T2 | 336
reduction in extracellular volume | 336
small pericardial effusion | 336
enhancement of the parietal pericardium | 336
pericarditis | 336
resolution of pulmonary consolidation | 336
resolution of pleural effusions | 336
discharged | 360
