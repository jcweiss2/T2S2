79 years old | 0
male | 0
admitted to the hospital | 0
fever | -1176
fatigue | -1176
anorexia | -1176
body temperature reaching 38.5 °C | -1176
body temperature fluctuating between 36.5 °C and 38 °C | -1176
pulmonary bacterial infection | 0
respiratory failure | 0
co-morbid diseases | 0
poor nutrition | 0
nasogastric tube insertion | 0
cerebral infarction | 0
coronary atherosclerotic heart disease | 0
COVID-19 | 0
anti-infection treatment | 0
antiviral treatment | 0
treatments for improving cardiac function | 0
blood transfusions | 0
symptomatic treatments | 0
brain computed tomography scan showing multiple small punctate hypodense foci | 0
chest computed tomography scan showing scattered patches and cloudy fuzzy shadows | 0
ischemic changes | 0
acute ischemic stroke | 0
nasogastric tube placement using ultrasound | 0
gastric juice extraction failure | 0
auscultation failure due to stethoscope unavailability | 0
no bubble overflow in normal saline solution | 0
ultrasonic probe identification of nasogastric tube | 0
comet tail sign through cross-section after esophageal inlet | 0
parallel transparent hyperechoic images in the shape of "=" | 0
100 mL nutrient solution injected | 0
no discomfort | 0
vital signs stable | 0
no adverse reactions | 0
severe COVID-19 | 0
malnutrition | 0
enteral nutritional support | 0
nasal feeding feasibility assessment | 0
nasal septum deviation investigation | 0
nasal inflammation investigation | 0
obstruction investigation | 0
cerebrospinal fluid rhinorrhea investigation | 0
no contact with COVID-19 patients | -1176
no history of COVID-19 in family | 0
recovery from cerebral infarction | 0
no impairment of action or speech | 0
Level 3 protection requirements | 0
X-ray radiation avoidance | 0
decreased oxygen saturation risk | 0
tube slippage risk | 0
inadvertent aspiration risk | 0
viral exposure risk reduction | 0
clinical workload reduction | 0
immediate accurate results | 0
prognosis improvement | 0
treatment success potential improvement | 0
informed consent provided | 0
no conflicts of interest | 0
CARE Checklist compliance | 0
peer-reviewed | 0
single blind peer-review | 0
Grade C peer-review | 0
Grade D peer-review | 0
no shortness of breath | 0
denies chest pain | 0
co-morbid diseases |7 0
