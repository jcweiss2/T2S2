31 years old|0
male|0
presented to his general practitioner| -24
bilateral joint pains|-24
joint swelling|-24
ankle joint involvement|-24
wrist joint involvement|-24
polyarthralgia| -48
coryzal symptoms| -72
sore throat| -72
fever| -72
no headache|0
no photophobia|0
no neck stiffness|0
alert and orientated|0
temperature 36.9°C|0
heart rate 101 bpm|0
blood pressure 125/85 mmHg|0
respiratory rate 16 breaths per minute|0
oxygen saturations 99%|0
qSOFA score of zero|0
bilateral swelling in small joints of hands|0
wrist joint pain|0
knee joint swelling|0
knee joint pain|0
mild purpuric rash on limbs|0
metabolic acidosis|0
raised lactate 9.29 mmol/L|0
cryptic shock|0
C reactive protein 223 mg/L|0
erythrocyte sedimentation rate 45 mm/h|0
white cell count 4.9 × 10^9/L|0
international normalized ratio 2|0
prothrombin time 24.9 s|0
D-dimer 42,011 ng/mL|0
alanine aminotransferase 58 U/L|0
alkaline phosphatase 81 U/L|0
haematuria|0
proteinuria|0
sepsis of unknown source with DIC|0
blood cultures taken|0
commenced intravenous piperacillin/tazobactam|0
commenced intravenous fluids|0
intravenous vitamin K 10 mg|0
ankle joint aspiration|0
negative joint fluid cultures|0
negative ANCA|0
negative ANA|0
negative ASOT|0
negative rheumatoid factor|0
negative lupus anticoagulant|0
negative HIV|0
negative hepatitis B|0
negative hepatitis C|0
mildly raised rheumatoid factor|0
mildly raised lupus anticoagulant|0
urine total protein:creatinine ratio 164.2 mg/mmol|0
blood cultures grew Neisseria meningitidis group W135|48
switched to benzylpenicillin|48
household contacts received ciprofloxacin prophylaxis|48
remained febrile after 9 days|216
inflammatory markers rising CRP 354 mg/L|216
developed extensive ecchymosis|216
purpuric macules|216
large bullous lesions|216
soft tissue induration|216
cutaneous lesions on limbs|216
ankle and wrist joint swelling persisted|216
vasculitic element|216
purpura fulminans|216
CT chest, abdomen, pelvis normal|216
transthoracic echocardiogram normal|216
skin necrosis evolved|240
MRI of four limbs performed|240
failure to defervesce|240
daily fevers up to 39.5°C|240
non-resolving inflammatory response|240
new skin lesions|240
immune-driven complications|240
immune-complex formation|240
ibuprofen 400 mg TID ineffective|240
pulsed intravenous methylprednisolone 500 mg|240
fever lysis post methylprednisolone|240
clinical improvement|240
biochemical improvement|240
antibiotics stopped after 14 days|336
recrudescence of fever|336
reintroduced intravenous meropenem|336
reintroduced oral prednisolone|336
majority cutaneous lesions regressed|336
tissue loss over right foot dorsum|336
CT angiogram excluded macrovascular ischemia|336
repeat MRI right foot showed soft tissue collection|336
referred to plastic surgeons|336
surgical debridement|336
attempted flap cover unsuccessful|336
right above-knee amputation|336
convalescence complicated|336
