88 years old | 0
female | 0
admitted to the hospital | 0
hypertension | -672
atrial fibrillation | -672
unstable angina | -672
left-side motor weakness | -168
right-side eyeball deviation | -168
right middle cerebral artery (MCA) infarction | -168
tissue plasminogen activator (tPA) | -168
dyspnea | -120
unstable vital signs | -120
blood pressure 80/40 mmHg | -120
heart rate 150 beats/min | -120
respiration 44 breaths/min | -120
body temperature 39.1℃ | -120
O2 saturation 94% | -120
intubated | -120
left subclavian venous catheterization | -120
lidocaine injection | -120
left subclavian vein identified | -120
Seldinger-type central venous catheter set used | -120
guidewire passed through introducer needle | -120
guidewire advanced 30 cm | -120
guidewire could not be advanced further | -120
guidewire could not be withdrawn | -120
chest X-ray showed knotted and kinked guidewire | -120
transferred to hospital | -120
admitted to hospital | 0
portable chest X-ray | 0
subclavian venogram | 0
guidewire knotted and kinked in left clavicle area | 0
guidewire folded back on itself | 0
guidewire entered mediastinum | 0
subclavian vein intact | 0
surgical exploration decided | 0
general anesthesia | 12
etomidate injection | 12
rocuronium injection | 12
arterial catheter placed | 12
femoral venous catheter applied | 12
incision made | 12
guidewire found beneath subclavian vein | 12
guidewire cut and removed | 12
patient transferred to surgical intensive care unit | 24
patient discharged to ward | 48