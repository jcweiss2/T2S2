11 years old | 0
    female | 0
    repetitive focal to bilateral tonic-clonic seizures | 0
    febrile illness | -48
    abdominal pain | -48
    vomiting | -48
    normal neurodevelopment | 0
    unremarkable personal and family medical history | 0
    serial seizures began with right version | 0
    status epilepticus (SE) | 0
    refractory to first-line antiseizure treatment | 0
    refractory to second-line antiseizure treatment | 0
    transferred to intensive care unit (ICU) | 0
    sedated | 0
    intubated | 0
    mechanically ventilated | 0
    EEG on day 2 showed slow background with extreme delta brushes | 48
    extensive diagnostic work-up performed | 0
    hyperproteinorrachy identified | 0
    rhinovirus DNA isolated in PCR panel on nasal exudate | 0
    clinical picture critical on day 23 | 552
    escalation of anesthetics | 552
    continuous convulsive seizures with focal clonic jerks of the right hemibody | 552
    bilateral clonic jerking | 552
    EEG monitoring from day 18 to day 48 | 432
    seizure burden peaked on day 26 with abundant epileptiform EEG activity | 624
    focal to bilateral tonic-clonic seizures for >90% of recording time | 624
    seizures arose from left occipital region | 624
    temporal left seizures | 624
    central left seizures | 624
    occipital right seizures | 624
    brain MRI negative on first day of seizure recurrence | 24
    T2-FLAIR bilateral hyperintensity of claustra on day 7 | 168
    T2-FLAIR hyperintensity less marked on day 13 | 312
    T2-FLAIR hyperintensity in left cuneus on day 34 | 816
    failure of midazolam | 0
    failure of thiopental | 0
    failure of propofol | 0
    failure of ketamine | 0
    failure of topiramate | 0
    failure of cannabidiol | 0
    failure of valproate | 0
    failure of ospolot | 0
    failure of phenobarbital | 0
    failure of phenytoin | 0
    failure of lacosamide | 0
    failure of brivaracetam | 0
    failure of methylprednisone 1 g/day for 5 days | 0
    failure of IgIV for 5 days | 0
    failure of plasmapheresis for 5 days | 0
    ketogenic diet started on day 32 | 768
    target ketonemia (>2.5 mmol/L) achieved after one week | 768
    anakinra administration delayed by fever | 0
    anakinra administration delayed by raised inflammatory biomarkers | 0
    anakinra started on day 34 at 200 mg/day | 816
    anakinra increased to 400 mg/day on day 40 | 960
    seizures reduced by 50% after 3 days of anakinra | 888
    seizures stopped after 10 days of anakinra | 960
    focal seizures persisted on day 48 | 1152
    discharged from ICU on day 48 | 1152
    anakinra stopped on day 56 due to candida albicans sepsis | 1344
    continuous IV midazolam for subtle focal seizures | 1152
    eye deviation to the right | 1152
    IV midazolam stopped on day 90 | 2160
    regained awareness on day 90 | 2160
    focal seizures became less frequent | 2160
    transferred to rehabilitation on day 137 | 3288
    relapse of seizures during febrile illness due to gastroenteritis on day 217 | 5208
    IV midazolam controlled seizures | 5208
    discharged home on day 270 | 6480
    lacosamide 400 mg/day | 6480
    phenobarbital 100 mg/day | 6480
    clobazam 25 mg/day | 6480
    no clinical seizures at thirteen months | 9480
    no motor disability | 9480
    moderate intellectual disability | 9480
    milder impact on verbal functioning | 9480
    ketogenic diet weaned due to compliance issues | 9480
    low carbohydrate diet continued | 9480
