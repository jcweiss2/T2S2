49 years old | 0  
    male | 0  
    obese | 0  
    BMI-33.9 | 0  
    ethanol related decompensated liver cirrhosis | 0  
    recurrent life threatening variceal bleeds | 0  
    mild ascites | 0  
    jaundice | 0  
    CTP score −9 | 0  
    Child: B | 0  
    MELD Na: 17 | 0  
    referred for liver transplant | 0  
    no hypertension | 0  
    no diabetes | 0  
    no asthma | 0  
    wife evaluated as donor | 0  
    first nasopharyngeal swab for COVID-19 RT-PCR | -720  
    subsequent two swabs 48 hours apart | -720  
    negative COVID-19 RT-PCR | -720  
    informed consent for nosocomial COVID-19 risk | 0  
    live donor liver transplant | 0  
    partial MHV right lobe graft | 0  
    splenic artery ligation | 0  
    GRWR-0.70 | 0  
    right graft weight-635 gms | 0  
    intraoperative high portal pressure 16 mmHg | 0  
    intraoperative course uneventful | 0  
    extubated on POD1 | 24  
    post-operative doppler showed high portal blood flows 2000 ml/min | 168  
    pharmacological modulation with octreotide infusion | 168  
    intravenous methylprednisolone 10 mg/kg during anhepatic phase | 0  
    methylprednisolone tapered to 100 mg on POD1 | 24  
    methylprednisolone tapered to 80 mg on POD2 | 48  
    methylprednisolone tapered to 60 mg on POD3 | 72  
    methylprednisolone tapered to 40 mg on POD4 | 96  
    switched to oral wysolone 20 mg from POD5 | 120  
    tacrolimus started on POD2 | 48  
    tacrolimus trough level 8-10 ng/ml | 48  
    unable to start MMF in first post-operative week | 0  
    low platelet count | 0  
    low total leucocyte count | 0  
    low dose MMF 250 mg/12 hr started on POD8 | 192  
    rising aminotransferases | 192  
    serum AST and ALT rising trend in 2nd post-operative week | 336  
    methylprednisolone pulse therapy | 336  
    response to methylprednisolone | 336  
    percutaneous liver biopsy not performed | 336  
    thrombocytopenia | 336  
    four fold rise of aminotransferases | 336  
    absence of sepsis | 336  
    normal doppler study | 336  
    cirrhosis ethanol related | 336  
    acute cellular rejection suggested | 336  
    satisfactory hospital course | 0  
    discharge planned on POD20 | 480  
    developed fever on POD20 | 480  
    temperature 101°F | 480  
    heart rate 110 per minute | 480  
    respiratory rate 26 per minute | 480  
    saturation drop to 88% on ambient air | 480  
    RT-PCR positive for SARS‐CoV‐2 on day 2 of fever | 504  
    nasopharyngeal aspirate negative for other respiratory viruses | 504  
    immunosuppression modified | 504  
    MMF stopped | 504  
    oral steroid switched to intravenous hydrocortisone | 504  
    tacrolimus continued in low dose | 504  
    oxygen saturation 94-96% with high-flow nasal cannula | 504  
    day 3 of fever (POD22) | 528  
    tachypnoeic (RR-37/min) | 528  
    chest x-ray showed bilateral patchy parenchymal opacities | 528  
    shifted to intensive care isolation | 528  
    blood tests for inflammatory markers | 528  
    septic screening | 528  
    remdesivir 200 mg on first day | 528  
    remdesivir 100 mg once daily for next five days | 528  
    enoxaparin 60 mg once daily | 528  
    non-invasive ventilation continued | 528  
    clinical deterioration on day 6 of fever (POD25) | 600  
    IL-6-253.9 pg/ml | 600  
    CRP-106.04 mg/L | 600  
    NT-ProBNP%1426 pg/ml | 600  
    ferritin-108.62 ng/ml | 600  
    hypoxia worsened | 600  
    PF ratio-143 | 600  
    additional 3rd plasma aliquot transfused | 600  
    convalescent plasma aliquots from different donors | 600  
    IgG antibody titres >1:1000 | 600  
    deterioration halted | 600  
    no endotracheal intubation | 600  
    good recovery | 600  
    inflammatory markers improved | 600  
    off oxygen therapy on POD40 | 960  
    absolute lymphocyte count 1.42×103 per microliter | 960  
    radiological resolution of lung opacities | 960  
    aminotransferases improved | 960  
    total bilirubin improved | 960  
    repeat nasopharyngeal swabs positive | 960  
    discharged on 6th August 2020 | 960  
    doing well | 960  
    telephonic follow-up | 960  
