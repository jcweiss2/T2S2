27 years old | 0
female | 0
admitted to the emergency department | 0
ingestion of venlafaxine | -12
ingestion of alcohol | -12
hallucinations | 0
hyperreflexia | 0
mydriasis | 0
trism | 0
opsoclonus | 0
myoclonus | 0
serotonergic syndrome | 0
body temperature 37.0° C | 0
blood pressure 115/80 mmHg | 0
pulse 145 bpm | 0
sinus-tachycardia | 0
prolonged corrected QT-interval (QTc) of 513ms | 0
blood-alcohol level 2.32 ‰ | 0
glucose level 238 mg/dL | 0
symptomatic therapy | 0
given 2000 ml Sterofundin | 0
given 12 mg of midazolam | 0
transferred to the hospital’s intensive care unit | 0
severe intoxication | 0
high risk for hemodynamic failure | 0
glucose 200 ml of 20% glucose solution | 2
recurring severe hypoglycaemia | 2
invasive ventilation | 12
induction of anaesthesia | 12
given 5 mg of midazolam | 12
given 50 μg of sufentanil | 12
given 50 mg of rocuronium | 12
vasopressors | 12
noradrenaline up to 10 mg/h | 12
dobutamine up to 30 mg/h | 12
progressive lactic acidosis | 12
transthoracic echocardiography (TTE) | 13
severe left-ventricular dysfunction | 13
left ventricular ejection fraction (LVEF) of 10-15 % | 13
global left-ventricular hypokinesia | 13
veno-arterial extracorporeal life support (ECLS) | 17
diffuse bleeding | 17
acute liver failure | 17
disseminated intravascular coagulation | 17
venlafaxine serum concentration > 720 μg/L | 17
acute kidney failure | 17
slow low-efficiency dialysis | 17
systemic heparin | 17
septic shock | 96
serum procalcitonin (PCT) levels 11.6mmols/L | 96
serum lactate 5.6 mmol/L | 96
increase noradrenaline | 96
fluid replacement | 96
ventilator-associated pneumonia | 96
antibiotic therapy | 96
meropenem | 96
vancomycin | 96
anisocoria | 96
distorted pupils | 96
cranial imaging | 96
high doses of sedative medication | 96
midazolam | 96
sufentanil | 96
two-dimensional echocardiogram | 168
gradually recovering left ventricular function | 168
LVEF of 45% | 168
ECLS weaned | 168
extubated | 336
pneumonia improved | 336
transferred to a general ward | 336
transferred to rehabilitation | 336
clinically apparent lesion of the N. peroneus | 336