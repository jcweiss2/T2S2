47 years old | 0
male | 0
admitted to the hospital | 0
diarrhea | -336
nausea | -336
vomiting | -336
acute kidney injury | -336
kidney transplant | -6048
type two diabetes | 0
hypertension | 0
hyperlipidemia | 0
endocarditis | 0
coronary artery disease | 0
heart failure with reduced ejection fraction | 0
coronary artery bypass surgery | -7776
mitral valve replacement | -7776
aspirin | 0
atorvastatin | 0
carvedilol | 0
clopidogrel | 0
sacubitril-valsartan | 0
warfarin | 0
insulin | 0
tacrolimus | 0
mycophenolic acid | 0
no shortness of breath | 0
no cough | 0
no fever | 0
no chills | 0
no recent travel | 0
no known contact with sick person | 0
temperature 36.6 °C | 0
blood pressure 90/58 mm Hg | 0
heart rate 103 beats per minute | 0
respiratory rate 16 breaths per minute | 0
oxygen saturation 98% | 0
body-mass index 42.2 | 0
normal heart sounds | 0
clear lungs | 0
blood creatinine level 6.7 mg/dL | 0
blood potassium level 5.7 mMol/L | 0
blood urea nitrogen 175 mg/dL | 0
bicarbonate level 14 mMol/L | 0
white-cell count 2.9 K/CUMM | 0
lymphocytes count 0.2 K/CUMM | 0
INR 2.75 | 0
hypotension resolved | 0
insulin administered | 0
beta-agonists administered | 0
calcium administered | 0
polystyrene sulfonates administered | 0
nasopharyngeal swab tested positive for SARS-CoV-2 RNA | 0
no evidence of pulmonary infiltrates | 0
vital signs stable | 24
no respiratory symptoms | 24
oxygen saturation 96% | 24
diarrhea resolved | 24
nausea resolved | 24
vomiting resolved | 24
soft diet tolerated | 24
acute kidney injury unresolved | 72
hyperkalemia | 72
metabolic acidosis | 72
leukopenia | 72
mild thrombocytopenia | 72
oliguric | 72
transplant nephrology consultation | 72
renal ultrasonography normal | 72
urinary sediment examination normal | 72
intravenous fluid administered | 72
immunosuppressive therapy discontinued | 72
INR monitored | 72
warfarin administered | 24
INR increased | 48
productive cough | 96
shortness of breath | 96
oxygen saturation decreased | 96
oxygen administered | 96
filgrastim administered | 96
shortness of breath worsened | 102
oxygen saturation decreased | 102
high-flow nasal cannula initiated | 102
transferred to ICU | 102
blood and sputum specimen obtained | 102
chest radiograph obtained | 102
multifocal air-space opacities | 102
prominent pulmonary vascular markings | 102
enlarged cardiac silhouette | 102
intravenous furosemide administered | 102
vancomycin administered | 102
cefepime administered | 102
intubation and mechanical ventilation | 120
blood pressure decreased | 120
norepinephrine administered | 120
vasopressin administered | 120
CRRT initiated | 120
white blood cell count increased | 120
c-reactive protein increased | 120
ferritin increased | 120
lactate dehydrogenase increased | 120
creatine phosphokinase increased | 120
repeated chest radiograph | 120
bilateral opacities worsened | 120
prosthetic mitral valve normal | 120
left ventricular ejection fraction 20% | 120
atrial fibrillation | 144
amiodarone administered | 144
hypotension worsened | 144
CRRT held | 144
death | 216