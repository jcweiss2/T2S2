32 years old | 0
male | 0
Turkish | 0
obese | 0
body mass index 30kg/m2 | 0
admitted to ICU | 0
lymphoma with plasmablastic differentiation | -720
tumor lysis syndrome | -720
septic shock | -720
HIV diagnosis | -720
dolutegravir/abacavir/lamivudine treatment | -720
dolutegravir/abacavir/lamivudine administration by nasogastric tube | 0
Cp-DTG measurement | 96
meropenem concentration measurement | 96
linezolid concentration measurement | 96
anidulafungin concentration measurement | 96
undetectable Cp-DTG | 96
detectable meropenem concentration | 96
detectable linezolid concentration | 96
detectable anidulafungin concentration | 96
inflammation | -720
immunosuppression | -720
ferritin elevation | -720
C-Reactive protein elevation | -720
D-dimer elevation | -720
procalcitonin elevation | -720
enteric malabsorption | -720
mesenteric hypoperfusion | -720
hyperlactatemia | -720
high norepinephrine requirements | -720
trophic enteral feeding | 0
EF intolerance | 0
atrophy of the intestinal mucosa | 0
decreased dolutegravir absorption | 96
drug distribution alterations | 0
severe hypoalbuminemia | -720
hyperbilirubinemia | -720
increased dolutegravir clearance | 96
fever | -720
high and persistent fever | -720
haematological malignancies | -720
lymphoma impact on dolutegravir pharmacokinetics | 0
NT drug administration | 0
sedoanalgesia drugs | 0
delay in gastric emptying | 0
prokinetic drugs | 96
drug-drug interactions | 0
rifampin treatment | -168
rifampin suspension | -24
double dose dolutegravir reduction | -24
continuous venovenous hemodialysis | 0
minimal dolutegravir removal by hemodialysis | 96
no specific dolutegravir dosage adjustments required | 96
discharge | unknown