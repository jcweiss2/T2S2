63 years old| 0
    male | 0
    admitted to the hospital (initial diagnosis with SRCC) | 0
    signet ring cell carcinoma (SRCC) in the gastric corpus | 0
    neoadjuvant chemotherapy | 0
    gastrectomy with Roux-en-Y reconstruction | 0
    postoperative period with full recovery | 0
    infrarenal AAA (4.1 cm diameter) diagnosed | 0
    assigned follow-up for AAA | 0
    admitted due to urosepsis | -14,560
    admitted due to pyelonephritis | -14,560
    admitted due to anaemia (Hb 85 g/L) | -14,560
    previous antibiotic therapy | -14,560
    high inflammation markers (WBC 33.3 × 10^9/L; CRP 87 mg/L; PCT 3.3 ng/mL) | -14,560
    CTA scan detected AAA enlargement to 54 mm | -14,560
    thrombosed intramural haematoma (9 mm) in right aortic wall | -14,560
    no extravasation | -14,560
    assigned fatal rupture risk monitoring | -14,560
    hospitalization for 10 days | -14,560
    nonspecific symptoms (subfebrile fever, constipation) | -14,560
    condition worsened | -14,560
    severe fatigue | -14,560
    anaemia (Hb 78 g/L, Hct 23 %, CRP 123 g/L, PCT 6.5 ng/mL) | -14,560
    negative FOBT | -14,560
    absent GI tract bleeding symptoms | -14,560
    diagnostic delay | -14,560
    second CTA scan detected ruptured AAA (rAAA) | -14,560
    anteriorly located pseudoaneurysm (44x43mm) | -14,560
    urgent operation admission | -14,560
    total laparotomy performed | -14,560
    enlarged pulsating inflammatory conglomerate without active blood leakage | -14,560
    PAEF (2 cm defect in duodenum) | -14,560
    duodenal compression | -14,560
    inadequate perfusion | -14,560
    entire pars ascendens appeared necrotic | -14,560
    infrarenal AAA resected | -14,560
    replaced with 16 mm linear silver-coated Dacron graft | -14,560
    complete resection of pars horizontalis and pars ascendens | -14,560
    no severe postoperative complications | -14,560
    readmitted after 40 months | 40,320
    recurrent fainting episodes | 40,320
    pain in the abdomen | 40,320
    haematemesis (Hb 98 g/L) | 40,320
    severe idiopathic hypoglycaemia (1.7 mmol/L) | 40,320
    received RBC transfusions | 40,320
    underwent CT scans | 40,320
    underwent CTA scans | 40,320
    underwent gastroscopies | 40,320
    underwent coloscopies | 40,320
    no clinically significant findings | 40,320
    capsule-endoscopy detected jejunal ulcer | 40,320
    PET scan visualized metabolically active regions in distal jejunum and aortic graft | 40,320
    no definite diagnosis from PET scan | 40,320
    preoperative diagnostic hypotheses: tumor or SAEF | 40,320
    total laparotomy performed | 40,320
    stapler-lined jejuno-jejunal anastomosis adhered to Dacron graft | 40,320
    SAEF confirmed (between distal anastomosis of Dacron prosthesis and jejunum) | 40,320
    infrarenal aortic cross-clamping | 40,320
    Dacron graft removed | 40,320
    microbiological analysis (no malignancy or infection) | 40,320
    replaced with new linear xenograft | 40,320
    intravenous antibiotic therapy for 4 weeks postoperatively | 40,320
    per os acetylsalicylic acid initiated | 40,320
    follow-up CTA confirmed intact aortic graft after 30 months | 40,320
    no signs of inflammation or fistulisation | 40,320
