70 years old | 0
female | 0
Caucasian | 0
admitted to the hospital | 0
complaints of worsening shortness of breath | 0
productive cough | -72
nasal congestion | -72
diarrhea | -72
vomiting | -72
hypertension | -6720
tobacco use | -6720
oxygen saturation of 77% | 0
blood pressure of 94/53 mmHg | 0
heart rate of 122 bpm | 0
temperature of 36.8 °C | 0
poor air movement | 0
diminished breath sounds | 0
no audible wheezing | 0
no audible crackles | 0
pH of 7.30 | 0
pCO2 of 43 mmHg | 0
pO2 of 48 mmHg | 0
lactic acid 4.4 mmol/L | 0
leukocyte count of 25,000/mm3 | 0
bandemia | 0
hemoglobin 13.2 g/dL | 0
hematocrit 40.2% | 0
platelet count of 199,000/mm3 | 0
hazy bibasilar opacities | 0
no pleural effusion | 0
no pneumothorax | 0
full face noninvasive bi-level ventilation | 0
oxygen saturation increased to 93% | 0
shortness of breath improved | 0
desire not to be intubated | 0
desire not to be resuscitated | 0
blood cultures obtained | 0
urine cultures obtained | 0
respiratory virus panel | 0
influenza panel | 0
urine streptococcal antigens | 0
urine legionella antigens | 0
piperacillin-tazobactam | 0
vancomycin | 0
admitted to the medical intensive care unit | 0
antimicrobial coverage changed to ceftriaxone and azithromycin | 0
blood cultures grew Pasteurella multocida | 24
sensitive to all antibiotics tested | 24
de-escalated to monotherapy with ceftriaxone | 24
all other cultures and viral panels returned negative | 24
owns sixteen indoor cats | -6720
no recent scratches or bites | -6720
skin fully inspected | 0
no evidence of scratches or bites | 0
no tetanus shot administered | 0
noninvasive ventilation weaned | 72
transitioned to venturi mask | 72
hemodynamics remained stable | 72
off vasopressor support | 72
leukocytosis significantly improved | 72
lactic acidosis had resolved | 72
bilateral pleural effusions visualized | 72
diagnostic thoracentesis performed | 72
removal of 1000 mL of straw-colored fluid | 72
transudate by Light's criteria | 72
gram stain returned negative | 72
culture returned negative | 72
CT angiogram performed | 144
multifocal pneumonia | 144
right middle lobe | 144
right lower lobe | 144
left lower lobe | 144
moderate sized right pleural effusion | 144
no pulmonary embolism | 144
discharged home | 144
home oxygen | 144
IV ceftriaxone | 144
complete 14 days of treatment | 168