60 years old | 0
male | 0
insulin dependent diabetes mellitus | -7200
failed renal allograft | -7200
maintenance hemodialysis | -7200
fever | -72
diffuse abdominal pain | -72
elevated white blood cell count | -72
air in failed renal allograft | -72
focal segmental glomerulosclerosis | -9360
end-stage renal disease | -9360
dilated cardiomyopathy | -9360
bilateral radical nephrectomies | -9360
kidney cancer | -9360
deceased donor renal transplant | -7200
worsening left ventricular function | -7200
ejection fraction of 25% | -7200
severe mitral regurgitation | -7200
acute renal failure | -5760
transplant ureteric stricture | -5760
balloon dilatation | -5760
insertion of a stent | -5760
transplant ureterectomy | -5760
pyelovesicostomy of allograft | -5760
psoas hitch of the bladder | -5760
myocardial infarction | -4320
medical therapy | -4320
no revascularization | -4320
transplant failure | -3600
anuric | -3600
started on hemodialysis | -3600
put on deceased donor transplant wait list | -3600
admitted to ICU | -2160
hypoglycemia | -2160
non-ST-elevation myocardial infarction | -2160
in-hospital arrest | -2160
hepatomegaly | -2160
venous congestion | -2160
right-sided heart failure | -2160
elevated white blood cell count | -2160
blood culture grew Bacteroids | -2160
ciprofloxacin | -2160
metronidazole | -2160
CT scan of abdomen and pelvis | -2160
locules of gas in failed renal transplant | -2160
piperacillin-tazobactam | -2160
broaden antibiotic coverage | -2160
transferred to tertiary care institution | -1440
allograft nephrectomy | 0
hemodynamic stabilization | 0
emergent subcapsular nephrectomy | 0
necrotic kidney with pus | 0
no significant blood loss | 0
postoperatively transferred to ICU | 0
stable over next few days | 0
died on 4th postoperative day | 96
myocardial infarction | 96
histopathology | 96
necrotic kidney with acute inflammation | 96
total effacement of kidney architecture | 96