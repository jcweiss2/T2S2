67 years old | 0
male | 0
African American | 0
admitted to the hospital | 0
shortness of breath | -24
generalized weakness | -24
nausea | -24
diarrhea | -24
history of schizophrenia | 0
hypertension | 0
no history of splenectomy | 0
nonsmoker | 0
no use of illicit drugs | 0
no heavy alcohol consumption | 0
lived in a group home | 0
denied sick contacts | 0
refused pneumococcal vaccination | 0
refused influenza vaccination | 0
no sickle cell disease | 0
hypotension | 0
fever | 0
heart rate within normal range | 0
respiratory rate within normal range | 0
ill-appearing male patient | 0
alert and oriented | 0
lungs clear to auscultation | 0
heart sounds regular | 0
no tachycardia | 0
no murmurs | 0
abdominal examination normal | 0
neurologic examination normal | 0
no meningeal signs | 0
denied headache | 0
denied cough | 0
denied chest pain | 0
watery diarrhea | 0
elevated WBC count | 0
neutrophils | 0
low hemoglobin | 0
low platelet count | 0
elevated BUN | 0
elevated creatinine | 0
low bicarbonate | 0
elevated anion gap | 0
elevated lactic acid | 0
elevated alkaline phosphatase | 0
elevated AST | 0
elevated total bilirubin | 0
elevated direct bilirubin | 0
elevated CK | 0
elevated LDH | 0
elevated D-dimer | 0
microangiopathic hemolytic anemia | 0
CT scan negative for pulmonary infiltrates | 0
CT scan negative for colitis | 0
CT scan negative for intraabdominal source of infection | 0
diagnosed with severe sepsis | 0
treated with fluid resuscitation | 0
treated with broad-spectrum antibiotics | 0
developed retiform violaceous patches | 12
developed central dusky necrosis | 12
developed gangrene | 24
required norepinephrine infusion | 12
blood cultures grew Gram positive cocci | 48
identified as S. pneumoniae | 48
treated with ceftriaxone | 48
treated with clindamycin | 48
hemodialysis initiated | 72
echocardiogram normal | 72
repeat blood cultures negative | 72
weaned off norepinephrine | 72
renal function improved | 168
liver function improved | 168
weaned off hemodialysis | 168
rash nearly resolved | 168
discharged | 168