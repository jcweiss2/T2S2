69 years old | 0
female | 0
nonischemic dilated cardiomyopathy | -672
left ventricular ejection fraction (LVEF) of 35% | -672
guideline-directed medical therapy | -672
cardiac resynchronization therapy | -672
recovered LVEF | -168
fever | -168
chills | -168
diarrhea | -168
worsening dyspnea | -168
signs and symptoms of shock | -168
end-organ hypoperfusion | -168
admitted to the hospital | 0
negative result of SARS CoV-2 polymerase chain reaction testing | 0
elevated Coxsackie B virus titer to 1:320 | 0
transthoracic echocardiogram | 0
LVEF of 20% | 0
severe right ventricular (RV) dysfunction | 0
severe mitral regurgitation | 0
right heart catheterization | 0
right atrial (RA) pressure of 6 mm Hg | 0
RV pressure of 32/9 mm Hg | 0
pulmonary artery (PA) pressure of 30/20/25 mm Hg | 0
pulmonary capillary wedge pressure of 22 mm Hg | 0
V waves of 30 mm Hg | 0
left ventricular end diastolic pressure of 32 mm Hg | 0
cardiac output of 3.3 L/min | 0
cardiac index of 1.95 L/min/m2 | 0
electrocardiogram | 0
markedly low voltage | 0
ventricular paced rhythm | 0
coronary angiogram | 0
nonobstructive coronary artery disease | 0
cardiac biopsy | 12
nondiagnostic endomyocardial biopsy results | 12
empiric high-dose steroids with 1 g methylprednisolone | 12
worsening shock | 14
acute kidney and liver injury | 14
incessant ventricular tachycardia/fibrillation | 14
intravenous lidocaine | 14
amiodarone | 14
procainamide drips | 14
axillary LV-aortic microaxial pump | 14
venoarterial-ECMO | 14
RA of 11 mm Hg | 14
PA of 22/18/19 mm Hg | 14
pulmonary capillary wedge pressure of 20 mm Hg | 14
mixed venous saturation of 78% | 14
4 L of ECMO flow | 14
1.4 L of LV-aortic pump flow | 14
P4 setting | 14
refractory cardiogenic shock | 15
continued electrical instability | 15
transfer to hospital for consideration of durable mechanical support or OHT | 15
preliminary evaluation for OHT | 15
no major contraindications to heart transplantation | 15
temporary mechanical circulatory support | 15
PA outflow cannula | 15
refractory arrhythmias | 15
progressive multiorgan system dysfunction | 15
surgical temporary biventricular assist device | 15
oxygenator | 15
drainage cannulas in RA and LV apex | 15
reinfusion cannula in the ascending aorta | 15
expedited evaluation for durable mechanical circulatory support and OHT | 18
urgently listed for OHT | 18
cardiogenic shock | 18
surgically implanted VAD support | 18
OHT | 20
dobutamine 10 μg/kg/min | 20
norepinephrine 2 μg/min | 20
inhaled nitric oxide 20 ppm | 20
no mechanical circulatory support | 20
vasopressors weaned | 72
inotropes weaned | 72
inhaled nitric oxide weaned | 72
extubated | 96
pathologic examination of the explanted heart | 120
consistent with GCM | 120
massive myocarditis | 120
infiltrate predominantly of lymphocytes | 120
numerous mononuclear cells | 120
scattered eosinophils | 120
multinucleate giant cells | 120
extensive healing fibrosis | 120