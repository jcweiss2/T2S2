7 years old | 0\
male | 0\
admitted to the hospital | 0\
pre-B-ALL | -672\
relapse of pre-B-ALL | -672\
allogeneic HSCT | -672\
hemoglobin 8.5 g/dl | 0\
thrombocytes 13.000/μl | 0\
WBC 940/μl | 0\
neutrophils 50/μl | 0\
CRP 6.83 mg/dl | 0\
ferritin 182 μg/dl | 0\
cachexia | 0\
dry skin | 0\
pallor | 0\
multiple hematomas | 0\
hepatosplenomegaly | 0\
antibiotic, antiviral, and antifungal chemoprophylaxis | 0\
ceftriaxone | 0\
teicoplanin | 0\
acyclovir | 0\
caspofungin | 0\
pain in the left flank | 0\
morphine | 0\
blinatumomab treatment | 0\
somnolent and sleepy | 144\
delayed reaction | 144\
cerebral side effect of blinatumomab | 144\
cerebral CT scan | 144\
MRI scan | 144\
multiple cerebral hemorrhages | 144\
cardio-respiratory decompensation | 144\
mechanical ventilation | 144\
catecholamine therapy | 144\
blinatumomab treatment stopped | 144\
hemoglobin 6.7 g/dl | 144\
thrombocytes 49.000/μl | 144\
WBC 120/μl | 144\
neutrophils 20/μl | 144\
CRP 23.13 mg/dl | 144\
ferritin 1439 μg/dl | 144\
multiple thrombi in the left and right ventricle | 144\
thromboembolic events | 144\
endocarditis | 144\
septic embolisms | 144\
meropenem | 144\
gentamicin | 144\
CT scans of the thorax, abdomen and pelvis | 168\
multiple, systemic thromboembolic lesions | 168\
ischemia | 168\
bleeding | 168\
infarction | 168\
bone marrow aspiration | 168\
bone marrow aplasia | 168\
lymphatic blasts | 168\
cerebral pressure rising | 168\
cerebral herniation | 168\
death | 168\
invasive mycosis of R. pusillus | 168\
autopsy | 168\
R. pusillus identified via PCR-based methods | 168