65 years old | 0  
    man | 0  
    presented to emergency room | 0  
    muscular pain in the back of the neck | -144  
    generalized fatigue | 0  
    weakness | 0  
    received nonsteroidal anti-inflammatory drugs | -144  
    poor oral intake | 0  
    no weight loss | 0  
    loose motion | 0  
    no significant gastrointestinal symptoms | 0  
    no significant cardiorespiratory symptoms | 0  
    general physical examination | 0  
    dehydration | 0  
    jaundice | 0  
    normal heart sounds | 0  
    no added murmurs | 0  
    temperature of 39.7 C | 0  
    increased creatine kinase | 0  
    high sensitivity troponin T | 0  
    aspartate aminotransferase elevation | 0  
    alanine aminotransferase elevation | 0  
    total bilirubin elevation | 0  
    direct bilirubin elevation | 0  
    white blood count | 0  
    no clear consolidation on chest X-ray | 0  
    normal sinus heart rate | 0  
    left axis deviation | 0  
    no ischemic changes on ECG | 0  
    hypertension | 0  
    diabetes mellitus | 0  
    chronic renal impairment | 0  
    obesity | 0  
    metabolic syndrome | 0  
    obstructive sleep apnea | 0  
    cervical spondylosis | 0  
    lumbar spondylosis | 0  
    G6PD deficiency | 0  
    admitted as fever with jaundice | 0  
    infection-related hepatic dysfunction | 0  
    hemolytic episode | 0  
    virology screen negative | 0  
    autoimmune screens negative | 0  
    started on Ceftriaxone | 0  
    blood culture taken | 0  
    no more high temperatures after admission | 0  
    became unconscious | 48  
    unresponsive | 48  
    no seizure activity | 48  
    normal heart rate | 48  
    normal rhythm | 48  
    normal blood pressure | 48  
    normal blood glucose | 48  
    left hemispheric syndrome | 48  
    severe hemiparesis on the right | 48  
    gaze deviation to the left | 48  
    global aphasia | 48  
    hemianopia | 48  
    hypoesthesia | 48  
    NIHSS score 18 | 48  
    urgent CT brain | 48  
    no acute changes on CT | 48  
    left MCA ischemic stroke | 48  
    informed consent collected | 48  
    IV r-tPA administered | 48  
    onset to needle 30 min | 48  
    kept in ICU | 48  
    follow-up CT brain | 72  
    new ischemic infarct | 72  
    no hemorrhagic changes | 72  
    blood culture positive | 72  
    Gentamicin added | 72  
    TTE performed | 96  
    TEE performed | 96  
    vegetation on mitral valve | 96  
    mild to moderate mitral regurgitation | 96  
    Streptococcus agalactiae in blood culture | 120  
    Gentamycin for 2 weeks | 120  
    Vancomycin for 6 weeks | 120  
    follow-up TEE | 1344  
    no fresh vegetations | 1344  
    no abscess | 1344  
    follow-up CT brain | 1344  
    no hemorrhage | 1344  
    no mycotic aneurysms | 1344  
    speech difficulties | 1344  
    right hemiparesis | 1344  
    requiring cane to ambulate | 1344  

  