85 years old | 0
male | 0
Caucasian | 0
admitted to the hospital | 0
history of prior THA | -27648
elevated cobalt and chromium ions | -27648
head and liner exchange | -27648
atrial fibrillation | 0
congestive heart failure | 0
peripheral vascular disease | 0
abdominal aortic aneurysm | 0
renal artery stenosis | 0
chronic kidney disease | 0
hypertension | 0
chronic obstructive pulmonary disease | 0
prostate cancer | 0
anticoagulated with rivaroxaban | 0
abdominal aortic aneurysm repair | -27648
aortobifemoral bypass | -27648
hospitalized with E. coli sepsis | -144
E. coli sepsis secondary to pneumonia | -144
urinary tract infection | -144
right hip pain | -144
readmitted with worsening right hip pain | -72
swelling | -72
transferred to our institution | -72
diagnosed with right THA PJI | -72
cultures grew E. coli | -72
irrigation and debridement | -72
removal of the THA | -72
extended trochanteric osteotomy | -72
placement of an antibiotic-impregnated cement spacer | -72
treated with 6 weeks of intravenous antibiotics | -72
treated with 6 weeks of oral antibiotics | -36
antibiotic holiday | -14
fluoroscopically guided aspiration of his right hip | -14
serologic markers demonstrated a significant downward trend | -14
synovial fluid cell count and differential normalized | -14
alpha defensin testing | -14
bacterial cultures were found to be negative | -14
cleared his infection | -14
second stage of his reimplantation was scheduled | -14
physical examination revealed a well-healed posterolateral scar | -14
no pain with passive range of motion of the hip | -14
flex to 110° | -14
20° of internal rotation | -14
40° of external rotation | -14
no appreciable leg length discrepancy | -14
feet were warm and well perfused clinically | -14
palpable dorsalis pedis and posterior tibial pulses | -14
radiographs revealed the cement spacer remained in appropriate position | -14
fracture of the greater trochanter with significant displacement | -14
evaluated by his vascular surgeon and cardiologist | -14
optimized as much as possible before reimplantation | -14
rivaroxaban was discontinued 72 hours before the second-stage surgery | -3
revision right THA via posterior approach | 0
irrigation and debridement | 0
removal of the antibiotic impregnated spacer | 0
reimplantation of the right THA | 0
noncemented acetabular component | 0
2 screws for secondary fixation | 0
proximal femoral replacement | 0
no intraoperative complications | 0
estimated blood loss of 500 cubic centimeters | 0
transferred to the postanesthesia care unit | 0
transferred to the floor in stable condition | 0
palpable dorsalis pedis and posterior tibial pulses | 0
postoperative hemoglobin (Hgb) in the postanesthesia care unit was 7.4 | 0
preoperative anticoagulation, rivaroxaban was reinitiated at noon of postoperative day one (POD 1) | 12
at a lower dose (10 mg daily instead of 20 mg) | 12
given his low Hgb | 12
Hgb was found to be 5.8 on POD 2 | 48
transfused 2 units of packed red blood cells | 48
appropriate response | 48
systolic blood pressure was consistently in the 100s-140s | 48
without any periods of hypotension | 48
white blood cell count had increased from 15 on POD 1 to 25 | 48
loose bowel movements | 48
Clostridioides difficile testing was found to be positive | 48
started on oral vancomycin | 48
right lower extremity was found to be cool to the touch | 48
distal pulses which were palpable on morning rounds were now no longer palpable | 48
denied any significant discomfort or pain | 48
denied any weakness or changes in sensation from baseline | 48
stat computed tomography (CT) angiography was obtained | 48
revealed an occlusion in the right limb of his aortobifemoral graft | 48
taken emergently to the interventional vascular suite | 48
attempted percutaneous thrombectomy via the left brachial artery | 48
aborted after an arterial injury was noted in the brachial artery | 48
taken to the operating room | 48
underwent an open repair of his left brachial artery | 48
open groin exploration with open balloon thrombectomy of the right aortobifemoral graft | 48
intraoperative angiogram confirmed restoration of blood flow to the right lower extremity | 48
extubated and taken to the intensive care unit postoperatively | 48
started on a heparin drip | 48
rivaroxaban was held | 48
heparin drip was stopped | 72
restarted on the rivaroxaban | 72
vascular examination remained stable | 72
compartments remained soft | 72
recovered well and was discharged from the hospital 2 weeks later | 336
transferred to a skilled nursing facility | 336
doing well at his most recent clinic visit, 8 months postoperatively | 5376
pain-free | 5376
ambulating with the use of a walker and an ankle-foot orthosis | 5376
some residual weakness in the right foot | 5376
no complaints | 5376
no signs of recurrent infection or compromised blood flow to his right lower extremity | 5376
remains on chronic anticoagulation, currently on warfarin | 5376