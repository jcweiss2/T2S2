45 years old | 0
    woman | 0
    admitted to the heart center | 0
    severe mitral stenosis | 0
    left atrial clot | 0
    shortness of breath on minimal exertion | -168
    no cerebral symptoms | 0
    no headache | 0
    no dizziness | 0
    no transient ischemic attacks | 0
    no strokes | 0
    fully conscious | 0
    alert | 0
    oriented | 0
    stable vital signs | 0
    blood pressure 110/80 mmHg | 0
    diastolic murmur audible over the mitral area | 0
    intact cranial nerves | 0
    motor power intact | 0
    sensation intact | 0
    no evidence of vasculitis | 0
    no Osler’s nodes | 0
    no Jane way pad | 0
    no palmer erythema | 0
    no cyanosis of fingers | 0
    erythrocyte sedimentation rate 4 mm | 0
    no leukocytosis | 0
    white blood cell 10,000 mm3 | 0
    electrolytes within normal limits | 0
    kidney function within normal limits | 0
    liver function within normal limits | 0
    chest X-ray showing prominence of the left cardiac border | 0
    electrocardiography indicative of no change | 0
    two-dimensional echocardiography revealing large bulky non-mobile thrombosis in the left atrium | 0
    severe mitral stenosis | 0
    mitral valve area 0.6 cm2 | 0
    other cardiac valves normal | 0
    negative antinuclear antibodies | 0
    negative rheumatoid factor | 0
    elevation of C4 & C3 components of complement | 0
    negative HBS Antigen | 0
    underwent open heart surgery | 0
    ascending aorta cannulation | 0
    bicaval cannulation | 0
    aorta cross-clamped | 0
    heart arrested with cold cardioplegia | 0
    systemic hypothermia at 30 °C | 0
    cardiopulmonary bypass | 0
    stenotic mitral valve found with bulky clot | 0
    diseased mitral valve excised | 0
    left atrial clot excised | 0
    left atrial cavity irrigated with normal saline | 0
    valve implanted | 0
    left ventricle filled with saline and blood | 0
    left ventricle deaired | 0
    weaned off cardiopulmonary bypass | 0
    inotropic support initiated | 0
    transferred to intensive care unit | 0
    blood pressure dropped | 6
    central venous pressure elevated | 6
    extremity became cool | 6
    cyanotic | 6
    inotropic support with dobutamine | 6
    inotropic support with adrenaline | 6
    inotropic drugs tapered | 72
    blood pressure stabilized | 72
    cyanosis changed to gangrene | 72
    acral part of the extremity amputated | 288
    histopathological examination showed non-specific vasculitis with thrombosis | 288
    did not regain full consciousness | 24
    quadriplegic | 24
    non-voluntary movements of four limbs | 24
    non-voluntary movements of face | 24
    eyes could move only on vertical plane | 24
    pupils became small and fixed | 24
    managed to respond by blinking | 72
    managed to respond by moving eyes vertically | 72
    brain MRI revealed multiple infarction of the brainstem | 72
    prolonged ventilatory support | 72
    tracheostomy performed | 72
    acute renal failure | 72
    anemia | 72
    kidneys recovered | 72
    locked-in state for 4 weeks | 672
    no neurological improvement | 672
    expired from hepatic failure | 672
    generalized sepsis | 672
<|eot_id|>
