69 years old | 0
    primary arterial hypertension | 0
    dyslipidemia | 0
    ischemic heart disease | 0
    severe heart ejection fraction 15–20% | 0
    mechanical aortic valve | 0
    stage 4 chronic kidney disease | 0
    early-stage Alzheimer’s dementia | 0
    middle-class art teacher | 0
    living in an urban environment | 0
    no history of recent travel | 0
    no dairy intake | 0
    admitted to the emergency department | 0
    non-bloody diarrhea | -96
    diffuse abdominal pain | -96
    dyspnoea | -96
    unquantified fever | -96
    prostrated | 0
    hypotensive | 0
    chest X-ray | 0
    homogeneous opacity | 0
    pleural effusion | 0
    protein C-reactive protein 27 mg/dL | 0
    serum creatinine 6 mg/dl | 0
    hypoxemic respiratory failure | 0
    lactate level 1.37 mmol/L | 0
    septic shock | 0
    multiorgan dysfunction | 0
    empirical antibiotic therapy with ceftriaxone | 0
    admitted to the ICU | 0
    fluid filling | 0
    vasopressor support | 0
    invasive mechanical ventilation | 0
    continuous renal function replacement technique | 0
    early escalation antibiotic therapy for meropenem | 0
    early escalation antibiotic therapy for linezolid | 0
    L. monocytogenesis identified in blood cultures | 0
    L. monocytogenesis identified in pleural fluid | 0
    HIV negative | 0
    delay invasive diagnostic investigation | 0
    family denied consumption of contaminated food | 0
    no additional cases of listeria infection | 0
    chest CT scan | 0
    extensive multiloculated right pleural effusion | 0
    attempt for pleural decortication | 0
    hemothorax | 0
    linezolid changed to ampicillin | 0
    meropenem maintained | 0
    decrease in inflammatory parameters | 0
    treated with 12 days of meropenem | 0
    treated with 21 days of ampicillin | 0
    meningeal doses despite absence of CNS involvement | 0
    day 13 of ampicillin | 312
    increase in inflammatory parameters | 312
    worsening of pleural imaging | 312
    piperacillin-tazobactam added | 312
    new laboratory worsening | 312
    new clinical worsening | 312
    co-morbidities | 0
    suspension of invasive measures | 600
    patient died | 720
    