69 years old | 0
female | 0
admitted to the hospital | 0
general myalgia | -72
fever | -72
nausea | -72
picking ginkgo nuts in the mountains | -240
resided in an urban area | 0
right upper abdominal tenderness | 0
enlarged cervical lymph nodes | 0
rebound tenderness | 0
no eschar found | 0
blood pressure 110/90 mm Hg | 0
pulse rate 78/min | 0
respiratory rate 24/min | 0
body temperature 38.5℃ | 0
white blood cell count 4,510/mm3 | 0
segmented neutrophils 70.6% | 0
hemoglobin 14.0 g/dL | 0
platelet count 57 × 10^3/mm3 | 0
C-reactive protein 17.51 mg/dL | 0
aspartate aminotransferase 374 IU/L | 0
alanine aminotransferase 254 IU/L | 0
alkaline phosphatase 982 IU/L | 0
lactate dehydrogenase 1,141 IU/L | 0
total protein 7.0 g/dL | 0
albumin 3.8 g/dL | 0
total bilirubin 1.2 mg/dL | 0
abdominal computed tomography showed edematous change in the GB wall with GB stones | 0
intravenous ceftriaxone 2 g/d initiated | 0
percutaneous cholecystostomy performed | 0
sustained symptoms | 0
nausea persisted | 0
abdominal pain persisted | 0
progressive shortness of breath | 96
increasing sputum production | 96
hypoxemia | 96
confusion | 96
oxygen delivered at 5 L/min via nasal cannula | 96
arterial blood gas analysis pH 7.45 | 96
PaCO2 36 mm Hg | 96
PaO2 67 mm Hg | 96
HCO3- 25 | 96
extensive airspace consolidation in both lungs | 96
endotracheal intubation performed | 96
admitted to the intensive care unit | 96
maculopapular rash on her trunk and face | 120
sputum and blood cultures negative | 120
oral doxycycline 200 mg/d initiated | 120
intravenous piperacillin 4.5 g/d initiated | 120
serologic test for Orientia tsutsugamushi positive | 120
multi-organ function returned to normal state | 216
mental alertness improved | 216
follow-up chest radiography showed resolved abnormalities | 216
discharged | 312
percutaneous cholecystostomy catheter removed | 312
elective cholecystectomy performed | 312
three black pigment stones found | 312