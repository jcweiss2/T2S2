31 years old | 0
    female | 0
    cesarean section | -408
    cesarean section | -48
    presented 17 days post delivery | -408
    suprapubic abdominal pain | -72
    bilateral flank pain | -72
    dysuria | -72
    nausea | -72
    vomiting | -72
    diarrhea | -72
    afebrile | -72
    subjective rigors | -72
    chills | -72
    hypotension | 0
    leukocytosis 23,000 WBC/μl | 0
    left shift | 0
    elevated serum lactate 4.1 mmol/L | 0
    intravenous fluid resuscitation | 0
    empiric broad spectrum IV antibiotics | 0
    admitted to ICU | 0
    sepsis without established source | 0
    unremarkable urologic exam | 0
    unremarkable radiologic exam | 0
    clean urinalysis | 0
    suction D&C | 0
    laparoscopic intra-abdominal exam | 0
    white blood cell count rose to 42,000/μl | 24
    septic shock worsened | 24
    leukemoid reaction 112,000 WBC/μl | 24
    disseminated intravascular coagulation (DIC) | 24
    consideration of Clostridium sordellii infection | 24
    supra-cervical hysterectomy | 48
    bilateral salpingectomy | 48
    abdominal compartment syndrome | 48
    acute and chronic endo-myometritis | 48
    necrotic features | 48
    acute salpingitis | 48
    omental fat necrosis and hemorrhage | 48
    IV immunoglobulin | 48
    exploratory laparotomy | 120
    abdominal washout | 120
    vacuum-assisted closure (VAC) device | 120
    abdominal washout | 168
    Wittmann temporary abdominal fascia patch | 168
    exploratory laparotomy | 288
    abdominal washout | 288
    Wittmann patch tightening | 288
    abdominal washout | 336
    fascial closure | 336
    white blood cell count normalized | 144
    discharged | 600
    walker for ambulation | 600
    physical therapy home visits | 600
    de-conditioned | 600
    doing well at follow-up | 720
