56 years old | 0
male | 0
admitted to the hospital | 0
fever | -168
difficulty breathing | -168
diabetes | 0
hypertension | 0
hyperlipidaemia | 0
tested positive for COVID-19 | -168
intubated | -168
ventilation | -168
persistent temperature spikes | -504
fatigue symptoms | -504
blood culture isolated coagulase-negative Staphylococcus | -504
echocardiogram showed mitral valve vegetation | -504
received antibiotic combinations | -504
meropenem | -504
levofloxacin | -504
teicoplanin | -504
no resolution of fever | -504
no resolution of mitral valve vegetation | -504
referred to the current centre | -504
complained of right leg pain | 0
calf swelling | 0
pulse of 90 bpm | 0
blood pressure of 122/77 mmHg | 0
respiratory rate of 20 breaths/minute | 0
temperature of 38.5 oC | 0
pansystolic murmur over the mitral valve area | 0
bilateral coarse inspiratory crepitations | 0
right calf was swollen | 0
could not move his ankle due to pain and weakness | 0
left leg pulses were normal | 0
right foot pulses were impalpable | 0
elevated inflammatory parameters | 0
white blood cell count of 13 x 10^9/L | 0
C reactive protein of 341 mg/L | 0
haemoglobin level of 7.1 g/dL | 0
antibiotic therapy was changed | 0
vancomycin | 0
ceftriaxone | 0
pre-operative full body computed tomography angiography | 0
right 7 x 7.5 cm tibioperoneal trunk aneurysm | 0
transoesophageal echocardiogram examination | 0
posterior mitral valve leaflet vegetation | 0
moderate eccentric mitral regurgitation | 0
open surgical repair | 0
lung and cardiac assessment | 0
considered fit for surgery | 0
combined one stage operation | 0
cardiac surgery | 0
heparin | 0
activated clotting time of >400 seconds | 0
heart-lung machine | 0
extended vertical transatrial-septal approach | 0
mitral valve replacement | 0
bioprosthesis | 0
Edwards Magna | 0
size 29 | 0
heparin was reversed with protamine | 0
peripheral aneurysm repair | 0
harvest of the right saphenous vein | 0
exposure of the distal superficial femoral artery | 0
posterior tibial artery was exposed | 0
proximal control was obtained | 0
aneurysm was approached | 0
aneurysm was opened | 0
organised thrombus without pus was observed | 0
thrombus was evacuated | 0
aneurysm was ligated | 0
distal popliteal artery was ligated | 0
vascular reconstruction | 0
reversed saphenous vein graft | 0
end to side proximal anastomosis | 0
distal anastomosis | 0
intra-operative handheld Doppler examination | 0
no microorganisms were recovered | 0
aspirin | 24
atorvastatin | 24
cardiac surgery stage took 3 hours and 31 minutes | 0
vascular surgery took 3 hours 30 minutes | 0
total blood loss was 300 mL | 0
extubated on post-operative day two | 48
discharged from ICU on day seven | 168
discharged from hospital on day 31 | 744
echocardiography showed a normal functioning mitral valve at five months | 1140
free of symptoms at six months | 1344
palpable right PTA pulse at the ankle | 1344
advised to remain on 75 mg aspirin once daily | 1344