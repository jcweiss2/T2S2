73 years old | 0
female | 0
admitted to the ICU | -72
abdominal pain | -72
dizziness | -48
decompensated cirrhosis | -72
abdominal infection | -72
spontaneous peritonitis | -72
hypoproteinemia | -72
acute respiratory distress syndrome (ARDS) | -72
septic shock | -72
noninvasive ventilation | -48
oral and perioral herpes infection | -48
large wound around the lips and in the mouth | -48
consciousness intact | 0
no ongoing abdominal pain | 0
no distension | 0
no chest tightness | 0
no asthma | 0
perioral wound progressed to exhibit local bleeding with crusting of blood | 0
wound measured approximately 10 cm × 10 cm | 0
Prothrombin time 15.9 sec | 0
partial thromboplastin time 34.5 sec | 0
albumin 27.9 g/L | 0
alanine aminotransferase 56 U/L | 0
total bilirubin 129.4 μmol/L | 0
neutrophils 79.2% | 0
hemoglobin 87 g/L | 0
platelet count 48 × 10^9/L | 0
high sensitivity C-reactive protein 77 mg/L | 0
multidisciplinary consultation | 0
treatment with oral antiviral drugs | 0
intramuscular injection of nutritious nerve drugs | 0
application of topical penciclovir and mupirocin | 0
wet application of topical nitrocilin | 0
oral and topical antiviral and antibiotic administration | 24
nutritional and symptomatic supportive care | 24
anti-inflammatory effect of furacilin | 24
hemostasis with local epinephrine injection | 24
application of topical thrombin lyophilized powder | 24
wet wound healing approach | 24
wound fully healed | 168
discharged from the hospital | 168