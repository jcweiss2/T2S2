66 years old | 0
female | 0
unconscious | 0
previous suicide attempts | -87600
rheumatologist check-ups | -87600
blood laboratory findings in reference range | 0
last psychiatrist consultation 10 years ago | -87600
rare alcohol consumption | -87600
general good physical condition | 0
regular medication: enalapril | 0
methotrexate | 0
folic acid | 0
diclofenac | 0
lansoprazole | 0
Vit D3 | 0
cholecalciferol | 0
calcium-carbonate | 0
5-hydroxytryptophane | 0
occasional Alprazolam use | 0
coma | 0
blood pressure 115/70 mmHg | 0
heart rate 85/min | 0
oxygen saturation 97% on room air | 0
temperature 36.0°C | 0
tachypnoeic | 0
bilateral miosis | 0
fingers in ulnar deviation | 0
absent reflexes | 0
discrete pretibial edema bilateral | 0
no clonus | 0
no extrapyramidal signs |0
hypotension 70/50 mmHg |0
SaO2 decrease to 85% |0
pulmonary edema |0
miosis |0
no pupillary reflexes on light |0
no nuchal rigidity |0
absent limb reflexes |0
GCS 3 |0
pulmonary crackles bilaterally |0
respiration rate 25-30/min |0
non-invasive monitoring |0
laboratory findings: serum glucose deviation |0
sodium deviation |0
potassium deviation |0
urine ketones |0
urine proteins |0
GFR 92.9 mL/min/1.73 m² |0
D-dimer 3254.36 ng/mL |0
ECG HR 80/min |0
normal ECG axis |0
WBC 7.9 109/L |0
platelets 339 109/L |0
Hb 148 g/L |0
RBC 4.7 1012/L |0
Hct 0.42 |0
CRP 2.5 mg/L |0
glycemia 12.2 mmol/L |0
BUN 4.3 mol/L |0
creatinine 59.6 µmol/L |0
Na 136 mmol/L |0
K 3.76 mmol/L |0
Ca 2.3 mmol/L |0
AST 17.9 U/L |0
ALT 12.1 U/L |0
GGT 15.3 U/L |0
AF 85.5 U/L |0
myoglobin 49.6 ng/mL |0
troponin 11.1 ng/L |0
urine ketones + |0
urine proteins 30 |0
ethanol 526 mg/dL |0
PT 10.67 s |0
aTPP 26.37 s |0
TT 20 s |0
ABGA pH 7.26 |0
pCO2 3.5 kPa |0
SaO2 94% with O2 support |0
HCO3 14 mmol/L |0
BE -15.4 mmol/L |0
anion gap 21.7 mmol/L |0
lactates >2 mmol/L |0
symptomatic treatment: pulmonary aspiration |0
intravenous colloids 500 mL |0
NaCl 0.9% 500 mL |0
oxygen support 4-5 L/min |0
amp furosemide 10 mg IV |0
stabilized hemodynamic condition |0
BP increased to 110/70 mmHg |0
HR 110-120/min |0
urine output 3.5 mL/min |0
coma persistence |0
reflexes absence |0
toxicological screening: low benzodiazepines 477 ng/mL |0
opiates excluded |0
tramadol excluded |0
methadone excluded |0
cannabis excluded |0
5-HTP not assessed |0
hypotensive reaction 80/60 mmHg |0
SaO2 drop to 85% |0
tachypnea 35-40/min |0
shallow respirations |0
family report of 250 mL 70% ethanol disinfectant missing |0
BAC 526 mg/dL |0
ABGA metabolic acidosis confirmed |0
osmolality 403-421 mOsm/kg |0
D-dimer 3254 ng/mL |0
anaesthesiology consultant recommended monitoring without mechanical ventilation |0
treatment: D5 NS 100 mL/h |0
potassium 10 mmol/h |0
thiamine 100 mg IV |0
oxygen 4-5 L/min |0
BP average 90/60 mmHg |0
PCR SARS-COV-2 negative |0
hemodynamic instability |0
age-related reduced biotransformation |0
risk of fluid overload |0
immunocompromised condition |0
decision to perform hemodialysis |0
hemodialysis via femoral catheter |0
HD discontinued after 2.5 hours due to coagulation |2.5
nadroparin 0.6 mL administered |2.5
stuporous state |2.5
reflexes restoration |2.5
post-HD BAC 250 mg/dL |2.5
ABGA corrected |2.5
D-dimer increased to 8098 ng/mL |2.5
glycemia 6.4 mmol/L |2.5
BUN 5.5 mol/L |2.5
creatinine 64 µmol/L |2.5
Na 138 mmol/L |2.5
K 4.2 mmol/L |2.5
Ca 2.05 mmol/L |2.5
AST 50 U/L |2.5
ALT 26 U/L |2.5
GGT 17 U/L |2.5
AF 83 U/L |2.5
myoglobin 10 ng/mL |2.5
troponin 12.2 ng/L |2.5
D-dimer 8098 ng/mL |2.5
urine ketones - |2.5
proteins - |2.5
ethanol 200.107 mg/dL |2.5
treatment: D5NS 100 mL/h |12
ceftriaxone 2.0 g |12
famotidine 20 mg IV tid |12
nadroparin 0.6 mL tid |12
LOC improved to mild somnolence |12
depressed mood |12
BAC 104 mg/dL |12
no gastric discomfort |12
no hematemesis |12
no haemogram reduction |12
denial of excessive 5-HTP intake |12
RA therapy discontinued for 48 hours |12
transfer to psychiatric clinic |24
stable hemodynamic status |24
stable mental status |24
LMWH recommended for 7 days |24
haemostatic parameters control |24
continue regular therapy |24
PCR test for SARS-COV-2 negative |0
ethanol poisoning diagnosis |0
decision to use hemodialysis |0
coagulopathy due to metabolic acidosis |0
D-dimer increase post-HD |2.5
serotonin syndrome excluded |0
RA-related immunocompromise |0
risk of infections |0
proinflammatory cytokine activation |0
renal impairment risk due to enalapril and diclofenac |0
hypovolemia risk from furosemide |0
tartrazine exposure excluded |0
thrombotic complications monitoring |24
differential diagnosis of coma |0
suicidal poisoning confirmed |0
monitoring of haemostasis |24
avoidance of severe hypocalcemia |2.5
discontinuation of NSAID and ACE inhibitors during treatment |0
hypocalcemia post-HD |2.5
coagulopathy management |0
psychiatric follow-up |24
acute alcohol poisoning management |0
hemodialysis efficacy |2.5
fluids overload prevention |0
infection risk mitigation |0
thrombotic risk mitigation |24
enhanced monitoring post-HD |2.5
controlled glycemia |0
alcohol elimination monitoring |0
