29 years old|0
female|0
referred to the emergency department|0
vomiting|-96
general malaise|-96
atypical chest pain|-96
epigastric pain|-96
polyuria|-720
polydipsia|-720
mild eczema|0
3 pack-year smoking history|0
normotensive|0
blood pressure 141/100 mmHg|0
sinus tachycardia 127 b.p.m.|0
temperature 34.6°C|0
oxygen saturation 98% on room air|0
respiratory rate 22 breaths/min|0
normal lung examination|0
normal heart examination|0
normal lower limb examination|0
severe high anion gap metabolic acidosis|0
arterial pH 6.87|0
hyperglycaemia 31.6 mmol/L|0
capillary ketones 4.6 mmol/L|0
bicarbonate 2.9 mmol/L|0
PO2 11.7 kPa|0
PCO2 1.5 kPa|0
normal CXR|0
sinus tachycardia on ECG|0
hypokalaemia 3.2 mmol/L|0
white cell count 33.09 ×10^9/L|0
neutrophils 28.43 ×10^9/L|0
CRP 13.9 mg/L|0
normal plasma sodium|0
normal serum creatinine|0
diagnosed with new-onset type 1 DM|0
commenced treatment for DKA|0
potassium replacement|0
fixed rate insulin infusion|0
volume expansion with crystalloids|0
empiric intravenous amoxicillin/clavulanic acid|0
pH 7.07|0
capillary ketones 4.1 mmol/L|0
hypothermia resolved|0
desaturated to 88% on room air|24
commenced on supplemental oxygen|24
ABG on 3 L of oxygen|24
PaO2 6.4 kPa|24
PCO2 2.3 kPa|24
pH 7.24|24
bicarbonate 7.5 mmol|24
suspected case of SARS-CoV2|24
nasopharyngeal swab taken|24
desaturated further with type 1 respiratory failure|24
bilateral infiltrates on CXR|24
ARDS-like picture|24
deterioration with fall in pO2 to 5.3 kPa|24
high flow oxygen via AIRVO|24
diuretic treatment|24
continuation of antibiotics|24
transferred to ICU|24
intubated and ventilated|24
FiO2 100%|24
peak end expiratory pressure 15 cm H2O|24
PaO2 10.3 kPa|24
haemodynamic support with noradrenaline 40 µg/min|24
vasopressin 2.4 units/h|24
ECMO|24
CVVH|24
negative SARS-CoV2 swabs|72
troponin rose from 38 to 2869 ng/L|48
normal creatine kinase 84 U/L|48
TTE showed reduced ejection fraction 45%|48
discontinue ECMO after 4 days|96
extubated|168
PaO2 16.7 kPa on FiO2 30%|168
troponin 401 ng/L|168
ejection fraction 50-55% on echo|168
minimally thickened trileaflet aortic valve|168
insulin infusion discontinued|192
commenced subcutaneous insulin|192
negative cultures|192
normal CXR|192
no cardiomegaly|192
no mediastinal lymphadenopathy|192
discharged to endocrine ward|264
discharged home|384
HbA1c 58 mmol/mol|0
positive GAD antibodies|0
normal cardiac function|0
troponin <14 ng/L|0
no shortness of breath|0
clear chest examination|0
oxygen saturation 99% on room air|0
diagnosis of ARDS in association with severe DKA|0
type 1 DM|0
no significant sequels|0
