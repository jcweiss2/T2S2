10 years old | 0
male | 0
referred to hospital | -504
persistent fever | -504
cough | -504
weight loss | -504
chest X-ray | -504
treatment for acute bronchitis | -504
thiamphenicol | -504
clavulanic acid | -504
amoxicillin | -504
conscious | 0
respiratory distress | 0
dyspnoea | 0
polypnea | 0
heart rate | 0
temperature | 0
hepatomegaly | 0
distended neck veins | 0
muffled heart sounds | 0
admitted to paediatric intensive care unit | 0
thoracoabdominal sonogram | 0
left liver lobe abscess | 0
chest and abdominal CT scan | 0
bilateral pleuropneumopathy | 0
diaphragmatic collection | 0
hepatosplenomegaly | 0
minor ascites | 0
amoebic serology | 0
IV antibiotic | 0
amoxicillin | 0
clavulanic acid | 0
gentamicin | 0
pericardial effusion | 0
mediastinal abscess | 0
mediastinal drainage | 0
evacuated 500ml pus | 0
no improvement | 0
antibiotic changed | 0
ceftriaxone | 0
metronidazole | 0
blood transfusion | 0
severe anaemia | 0
no improvement after 3 days | 72
ASA class V | 72
thoracotomy | 96
pericardiectomy | 96
removed 2 litres pus | 96
drains left in place | 96
febrile | 120
culture of pus grew Staphylococcus aureus | 120
HIV serology positive | 120
gentamicin stopped | 120
ciprofloxacin started | 120
temperature subsided | 216
hemodynamic parameters improved | 216
persistent purulent drainage | 216
stable | 312
corticotherapy introduced | 312
drains removed | 312
chest radiograph | 312
bilateral lower lobe infiltrate | 312
mild cardiomegaly | 312
cardiac sonogram | 312
thickened pericardium | 312
no pericardial effusion | 312
no valvular anomaly | 312
discharged home | 576
per os ciprofloxacin | 576
iron treatment | 576
steroids stopped | 576
seen in out-patient department 1 week after | 672
doing well | 672
seen 1 month after discharge | 1344
confirmation HIV testing positive | 1344
CD4 count 14 cells/ml | 1344
antiretroviral drugs | 1344
cotrimoxazole | 1344
referred back to hospital | 1344
mother admitted antiretroviral treatment | 1344
sepsis | 0
cardiac tamponade | 0
HIV infection transmitted by mother | -504
massive purulent pericarditis | 0
severe sepsis | 0
life-threatening empyema | 0
cardiomegaly | 0
immune depression | 0
amoebic liver abscess differential diagnosis | 0
HIV testing requested | 0
pericardiostomy recommended | 0
pericardial effusion confused with liver abscess | 0
pericardiectomy necessary | 96
thick pus | 96
massive pus | 96
cardiac failure | 0
high mortality | 0
infection spread hematogenously | 0
contiguous spread | 0
secondary to foreign body | 0
pneumonia | 0
empyema | 0
Streptococcus | 0
Staphylococcus | 0
chronic pericarditis | 0
tuberculosis infection | 0
HIV positive | 0
pericardial collection | 0
immune depressed | 0
amoebic infection | 0
frank thick pus | 0
decortication | 0
purulent drainage | 216
fibrosis | 312
lower lobe infiltrate | 312
antiretroviral treatment | 1344
cotrimoxazole prophylaxis | 1344
cardiac tamponade signs | 0
immunosuppression | 0
pericarditis diagnosis | 0
liver abscess differential | 0
CT scan misread | 0
left liver lobe | 0
Larrey's aperture | 0
immune depressed patients | 0
pericardiostomy | 0
HIV infected children | 0
sepsis presentation | 0
cardiac tamponade presentation | 0
purulent pericarditis suspicion | 0
