48 years old | 0
male | 0
admitted to the hospital | 0
transpelvic gunshot wound | 0
hemodynamically unstable | 0
blood pressure 82/63 mm Hg | 0
heart rate 120 bpm | 0
exploratory laparotomy | 0
small bowel injury | 0
rectosigmoid injury | 0
multiple areas of hemorrhage | 0
small bowel resected | 0
rectosigmoid resected | 0
small bowel anastomosed | 0
colostomy created | 0
intensive care unit | 0
coffee-ground output from nasogastric tube | -312
drop in hemoglobin from 8.9 to 7.1 g/dL | -312
transfused with 2 units of packed red blood cells | -312
esophagogastroduodenoscopy | -312
large ulcer at the body and fundus of the stomach | -312
irregular borders along with a vessel at the ulcer edge | -312
greyish coating and a large amount of exudate | -312
tissue biopsy from the ulcer | -312
intravenous pantoprazole | -312
oral sucralfate | -312
tissue pathology results revealed necrotic exudate containing fungal aseptate hyphae | -276
invasive gastric mucormycosis | -276
intravenous liposomal amphotericin | -276
no further bleeding | -276
stabilization of hemoglobin | -276
necrotic area at the open wound on the left flank | -288
development of sepsis | -288
white blood cell count of 23,000/µL | -288
heart rate of 120 bpm | -288
lactic acid level of 4.4 mmol/L | -288
broad-spectrum intravenous antibiotics | -288
vancomycin | -288
piperacillin-tazobactam | -288
repeat exploratory laparotomy | -288
multifocal necrotic bowel | -288
perforation around the anastomotic site | -288
necrotic bowel resected | -288
histopathological evaluation of resected specimen | -288
fungal aseptate hyphae consistent with the diagnosis of invasive GIM | -288
bloody output from the nasogastric tube | -264
abdominal surgical drains | -264
hemorrhagic shock | -264
refractory to blood transfusion | -264
refractory to intravenous hydration | -264
refractory to inotrope therapy | -264
immediate laparotomy | -264
perforation with necrosis at the previously seen gastric ulcer site | -264
active bleeding | -264
attempts to control the bleeding remained unsuccessful | -264
patient died in the operating room | -264