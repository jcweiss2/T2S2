43 years old | 0
male | 0
uncontrolled diabetes mellitus | -336
chronic kidney disease | -336
infected post-amputation surgical wound | -336
admitted to the hospital | 0
infected surgical wound on the right foot | 0
purulent discharge | 0
cellulitis | 0
decreased urination | 0
Foley catheter | 0
plain X-rays | 0
blood analysis | 0
white blood cells | 0
neutrophils | 0
lymphocytes | 0
hemoglobin | 0
hematocrit | 0
platelets | 0
fasting blood sugar | 0
creatinine | 0
blood urea nitrogen | 0
C-reactive protein | 0
bilirubin | 0
venous blood gas | 0
pH | 0
PCO2 | 0
HCO3 | 0
broad-spectrum intravenous antibiotics | 0
Vancomycin | 0
Piperacillin/Tazobactam | 0
Imipenem | 0
wound irrigation | 0
fever | 168
systolic hypotension | 168
confusion | 168
Guillotine Ankle Amputation | 168
sepsis under control | 336
necrotic ulcer | 336
IV injections | 336
extensive debridement | 336
necrotic tissue | 336
pathological evaluation | 336
skin | 336
underlying fat | 336
non-septate broad fungal hyphae | 336
cutaneous mucormycosis | 336
liposomal amphotericin B | 336
pulseless radial and ulnar arteries | 360
Color-Doppler ultrasound | 360
occlusive clot formation | 360
proximal brachial artery | 360
acute deep vein thrombosis | 360
axillary vein | 360
surgical embolectomy | 360
severe sepsis | 432
multi-organ failure | 432
death | 432