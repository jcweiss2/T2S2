85 years old | 0
severe valvular cardiopathy | 0
ischaemic-hypertensive cardiopathy | 0
slight chronic renal failure | 0
chronic venous leg ulcers | 0
plunged legs in seawater | -336
first clinical evaluation | 0
no fever | 0
pain on distal left lower limb | 0
ulcer left lateral ankle | 0
fibrinous coating | 0
greenish coating | 0
smelly coating | 0
ulcers on right leg | 0
pretibial ulcers | 0
perimalleolar ulcers | 0
chronic venous insufficiency | 0
varicose veins | 0
stasis dermatitis | 0
lipodermatosclerosis | 0
elevated CRP | 0
no leucocytosis | 0
ankle-brachial pressure index 0.9 | 0
X-ray no involvement of joints | 0
X-ray no involvement of bones | 0
admitted to hospital | 0
intravenous antibiotic therapy | 0
amoxicillin | 0
clavulanic acid | 0
fever | 0
increased inflammatory parameters | 0
cellulitis left leg | 12
hypotension | 12
acute renal failure | 12
septic shock | 12
changed antibiotic to imipenem | 12
treated with intravenous catecholamines | 12
blood cultures growth Vibrio parahaemolyticus | 12
diagnosed septic shock Vibrio parahaemolyticus | 12
bacteriological smear wounds growth Vibrio parahaemolyticus | 12
bacteriological smear wounds growth Pseudomonas aeruginosa | 12
bacteriological smear wounds growth Morganella morganii | 12
bacteriological smear wounds growth Streptococcus mitis | 12
bacteriological smear wounds growth Enterococcus spp | 12
stopped imipenem | 12
started ciprofloxacin | 12
started doxycycline | 12
normalization of haemodynamics | 336
return to usual renal parameters | 336
chronic hepatitis B infection | 336
no virulence detected in blood | 336
hepatic function intact | 336
sonography showed cardiac liver | 336
portal hypertension | 336
daily curettage | 0
topical sulphonamide | 0
pressure bandage lower limbs | 0
negative pressure wound treatment | 0
stopped negative pressure wound treatment | 0
discharged from hospital | 336
outpatient clinic visits | 2880
satisfactory granulation | 2880
split-thickness skin graft | 2880
complete wound healing | 2880
