62 years old | 0
    man | 0
    febrile neutropenia | 0
    dry cough | 0
    dyspnea | 0
    autologous bone marrow transplant | -384
    mantle cell lymphoma | -384
    chest CT | 0
    diffuse tracheobronchial thickening | 0
    densification of adjacent mediastinal fat | 0
    empirical antibiotic therapy | 0
    coverage for fungal infections with amphotericin B | 0
    persistence of cough | 24
    hemoptysis | 24
    CT performed one month and ten days after first CT | 912
    worsening of tracheal and bronchial walls thickening | 912
    increased densification of adjacent mediastinal fat | 912
    laryngotracheobronchoscopy | 504
    attached whitish plaques | 504
    detachable whitish plaques | 504
    friable mucosa | 504
    segmental ostial obstruction | 504
    bronchoalveolar lavage | 504
    endobronchial biopsy | 504
    presence of bifurcated hyphae at 45° | 504
    Aspergillus sp | 504
    chest CT two days after laryngotracheobronchoscopy | 528
    progression of disease | 528
    bronchoalveolar lavage culture positive for Aspergillus sp | 504
    discharged | 504
    outpatient follow-up | 504
    prescribed oral voriconazole | 504
    new admission | 576
    abdominal pain | 576
    diarrhea | 576
    hypotension | 576
    febrile peak | 576
    septic shock from abdominal origin | 576
    intensive care unit admission | 576
    death | 720
    <|eot_id|>

    