22 years old | 0
man | 0
presented to emergency department | 0
diagnosed with mild COVID-19 illness | -1032
sore throat | -1032
loss of sense of smell | -1032
positive COVID-19 PCR | -1032
full recovery | -1032
negative PCR | -1032
received first dose of inactivated SARS-CoV-2 vaccine | -1008
remained asymptomatic and well | -1008
received second dose of inactivated SARS-CoV-2 vaccine | -336
started to experience headache | -336
started to experience fatigue | -336
started to develop fever | -312
started to develop sore throat | -312
started to develop abdominal pain | -312
illness progressed over the following 4 days | -264
high-grade fever | 0
myalgia | 0
nausea | 0
vomiting | 0
diarrhoea | 0
faint erythematous non'itchy rash over torso | 0
dry irritant cough | 0
no shortness of breath | 0
no chest discomfort | 0
no urinary symptoms | 0
no pain | 0
no swelling of joints | 0
no history of recent travel | 0
no sick contacts | 0
no animal exposure | 0
no consumption of raw dairy products | 0
not on chronic medications | 0
no known allergies | 0
reported taking ibuprofen | 0
reported taking one dose of antibiotic | 0
non-smoker | 0
did not use recreational drugs | 0
temperature of 39°C | 0
systolic blood pressure of 110 mm Hg | 0
tachycardia | 0
dry mucous membranes | 0
congested throat | 0
bilateral conjunctival injection | 0
left conjunctival haemorrhage | 0
generalised erythematous maculopapular rash | 0
peripheral lymph nodes not enlarged | 0
no audible cardiac murmurs | 0
chest clear to auscultation | 0
abdomen examination unremarkable | 0
WBC 15 | 0
platelet 122 | 0
creatinine 115 | 0
AST 53 | 0
ALT 81 | 0
direct bilirubin 35 | 0
albumin 16 | 0
C reactive protein 249 | 0
ferritin 4357 | 0
D-dimer 14 | 0
procalcitonin 9 | 0
interleukin-6 90 | 0
SARS-CoV-2 PCR negative | 0
SARS-CoV-2 IgG strongly positive | 0
throat swab negative for group A streptococcus | 0
sputum culture showed mixed flora | 0
bacterial blood cultures negative | 0
urinalysis showed significant proteinuria | 0
ANA negative | 0
dsDNA negative | 0
c-ANCA negative | 0
p=ANCA negative | 0
C3 reduced | 0
C4 reduced | 0
admitted to intensive care unit | 0
hypotension | 0
diagnosis of probable sepsis | 0
diagnosis of vaccine-related illness | 0
treated with ceftriaxone | 0
treated with levofloxacin | 0
intravenous fluids | 0
intravenous hydrocortisone | 0
hydrocortisone stopped | 48
blood pressure stabilised | 0
fever initially improved | 0
fever remained persistent | 0
started to develop facial puffiness | 0
started to develop generalised body oedema | 0
remained tachycardic | 0
diarrhoea persisted | 0
difficult to mobilise | 0
renal impairment | 0
significant proteinuria | 0
ECG showed sinus tachycardia | 0
ECG showed non-specific T-wave abnormalities | 0
troponin-I raised | 0
pro-BNP over 8000 pg/mL | 0
transthoracic echocardiogram showed severe tricuspid regurgitation | 0
transthoracic echocardiogram showed normal tricuspid valve structure | 0
pulmonary hypertension | 0
PASP 46 mm Hg | 0
right atrium moderately dilated | 0
right ventricle moderately dilated | 0
normal systolic function | 0
left ventricle cavity size normal | 0
mildly reduced ejection fraction | 0
thin rim of pericardial effusion | 0
computed tomography scan negative for pulmonary embolism | 0
bilateral moderate pleural effusion | 0
basal atelectasis | 0
hydrocortisone discontinued | 48
shifted to medical ward | 48
high-level fever began to recur | 48
all cultures negative | 0
other workup unrevealing | 0
multisystem inflammatory syndrome in adults | 0
multisystem involvement | 0
cardiac involvement | 0
renal involvement | 0
haematologic involvement | 0
dermatologic involvement | 0
ophthalmologic involvement | 0
raised inflammatory markers | 0
therapy with intravenous dexamethasone | 168
condition improved | 168
generalised oedema subsided | 168
skin rash resolved | 168
conjunctivitis resolved | 168
white blood cell count normalised | 168
renal function improved | 168
inflammatory markers normalised | 168
repeat transthoracic echocardiography showed trace tricuspid regurgitation | 168
marked improvement in right ventricular systolic function | 168
normal size of right atrium | 168
normal size of right ventricle | 168
pulmonary artery systolic pressure normalised | 168
dexamethasone continued | 168
switched to oral prednisolone | 192
discharged home | 192
tapering dose of prednisolone | 192
symptoms resolved | 432
some general weakness | 432
fatigue | 432
repeat echocardiogram completely normal | 432
