60 years old | 0
male | 0
admitted to the hospital | 0
fever | -48
abdominal pain | -48
edema of the scrotum | -48
edema of the penis | -48
edema of the perineum | -48
edema of the right gluteal region | -48
hypertension | -672
osteoporosis | -672
hemorroids | -672
high degree of inflammation | 0
white blood cell count 13.11/μL | 0
C-reactive protein level 61.4 mg/dL | 0
serum creatinine 4.3 mg/dL | 0
blood urea 157 mg/dL | 0
blood sugar 142 mg/dL | 0
procalcitonin 8.53 ng/mL | 0
SARS-CoV-2 infection suspected | 0
SARS-CoV-2 infection confirmed | 0
CT of the abdomen and the pelvis | 0
inflammatory infiltration of the subcutaneous tissues of the hypogastrium | 0
liquefaction, and presence of gas in the subcutaneous tissues of the scrotum, the perineum, and the right gluteal region | 0
Fournier's gangrene | 0
meropenem | 0
metronidazole | 0
linezolid | 0
resection of the necrotic tissues | 0
bilateral orchiectomy | 0
excision of the penile and scrotal skin | 0
mechanical ventilation | 12
broad-spectrum antibiotics | 12
supportive and nutritional therapies | 12
colostomy | 12
wound debridement | 12
negative pressure wound therapy | 12
Escherichia coli | 24
Pseudomonas aeruginosa | 24
cephazolin | 24
catheterization | 24
free-skin grafts | 24
testosterone supplementation | 24
colostomy reversal | 48
continous nursing care | 48
free-skin graft care | 48
regular dressing changes | 48
physiotherapy | 48
urological and surgical clinic | 48