18 years old | 0
male | 0
fever | -672
rash | -672
acne | -672
minocycline | -672
increased WBC count | 0
eosinophilia | 0
systemic involvement | 0
diffuse erythematous or maculopapular eruption | 0
pruritis | 0
DRESS syndrome | 0
fever persisted | 0
rash persisted | 0
discharged | 24
admitted to the hospital | 0
right upper quadrant pain | -168
abdominal fullness and distention | -168
abdominal tenderness | -168
fever | -168
abdominal distension | -48
mild bellyache | -48
extreme thirst | -48
temperature of 36.8 °C | -48
fulvous fluid | -48
abdominal and pelvic computed tomography (CT) scan | -48
irregular, slightly low-density lesion in the right posterior hepatic lobe | -48
gas density shadow inside | -48
liquid density shadow and high-density drainage tube shadow | -48
round-like low-density lesion of about 0.8 cm in diameter | -48
thickened appendix | -48
structure of the ascending colon near the ileocecal region became disorganised | -48
multiple gas accumulation and dilation in the bowel | -48
air-fluid levels inside the abdomen | -48
hepatic abscesses | -48
ileus | -48
mild ascites | -48
appendicitis | -48
liver cyst | -48
abdominal infection | -48
peritonitis | -48
surgical exploration | -48
fulvous purulent exudate and necrotic tissue | -48
partial postnecrotic defect in the peritoneum | -48
massive epiploon adhesion in the right upper abdomen | -48
ileocecal resection | -48
partial resection of the ascending colon | -48
ileostomy and drainage of hepatic, abdominal and extraperitoneal abscesses | -48
orotracheal intubation | -24
hypotension | -24
anemia | -24
fever | -24
transferred to the intensive care unit (ICU) | -24
noradrenaline | -24
ventilator | -24
intravenous hydration | -24
nutritional support therapy | -24
blood transfusion | -24
blood cultures and drainage fluids | -24
tigecycline and piperacillin/tazobactam | -24
body temperature | -24
routine blood count | -24
procalcitonin level | -24
C-reactive protein (CRP) level | -24
elevated leukocyte count | -24
electrocardiogram monitor | -24
pulse rate of 130 beats/minute | -24
positive anaerobic blood culture vials | -24
Gram stain revealed short Gram-positive bacillus without spores | -24
MALDI-TOF MS | -24
E. lenta | -24
antimicrobial susceptibility testing | -24
tigecycline was replaced by teicoplanin | -24
piperacillin/tazobactam was discontinued | -24
ertapenem was added to teicoplanin | -24
cultures of the drainage fluid were obtained | -24
Escherichia coli | -24
ertapenem and teicoplanin | -24
fever, leukocytosis, PCT level and CRP level promptly improved | -24
transferred to the general ward | -24
ertapenem and teicoplanin | -24
debridement, dressing change and symptomatic supportive treatment | -24
repeated blood cultures | -24
negative | -24
repeat CT | -24
size of the hepatic abscess and the amount of ascites decreased | -24
intravenous ertapenem and teicoplanin | -24
symptoms achieved further alleviation | -24
discharged from the hospital | -24
oral antibiotics (clindamycin) | -24
follow-up with a six-week course of intravenous ertapenem | -24
electronic search on PubMed/MEDLINE | 0
Eggerthella lenta | 0
Eubacterium lentum | 0
key words | 0
case studies | 0
English language | 0
published from 1970 through 2020 | 0
E. lenta bacteremia | 0
liver abscess | 0
hepatic puncture and drainage | -1
admitted to our hospital | 0
complaints of right upper quadrant pain and discomfort | 0
right upper quadrant pain | 0
abdominal fullness and distention | 0
abdominal tenderness | 0
fever | 0
abdominal distension | 0
mild bellyache | 0
extreme thirst | 0
temperature of 36.8 °C | 0
fulvous fluid | 0
abdominal and pelvic computed tomography (CT) scan | 0
irregular, slightly low-density lesion in the right posterior hepatic lobe | 0
gas density shadow inside | 0
liquid density shadow and high-density drainage tube shadow | 0
round-like low-density lesion of about 0.8 cm in diameter | 0
thickened appendix | 0
structure of the ascending colon near the ileocecal region became disorganised | 0
multiple gas accumulation and dilation in the bowel | 0
air-fluid levels inside the abdomen | 0
hepatic abscesses | 0
ileus | 0
mild ascites | 0
appendicitis | 0
liver cyst | 0
abdominal infection | 0
peritonitis | 0
surgical exploration | 0
fulvous purulent exudate and necrotic tissue | 0
partial postnecrotic defect in the peritoneum | 0
massive epiploon adhesion in the right upper abdomen | 0
ileocecal resection | 0
partial resection of the ascending colon | 0
ileostomy and drainage of hepatic, abdominal and extraperitoneal abscesses | 0
orotracheal intubation | 0
hypotension | 0
anemia | 0
fever | 0
transferred to the intensive care unit (ICU) | 0
noradrenaline | 0
ventilator | 0
intravenous hydration | 0
nutritional support therapy | 0
blood transfusion | 0
blood cultures and drainage fluids | 0
tigecycline and piperacillin/tazobactam | 0
body temperature | 0
routine blood count | 0
procalcitonin level | 0
C-reactive protein (CRP) level | 0
elevated leukocyte count | 0
electrocardiogram monitor | 0
pulse rate of 130 beats/minute | 0
positive anaerobic blood culture vials | 0
Gram stain revealed short Gram-positive bacillus without spores | 0
MALDI-TOF MS | 0
E. lenta | 0
antimicrobial susceptibility testing | 0
tigecycline was replaced by teicoplanin | 0
piperacillin/tazobactam was discontinued | 0
ertapenem was added to teicoplanin | 0
cultures of the drainage fluid were obtained | 0
Escherichia coli | 0
ertapenem and teicoplanin | 0
fever, leukocytosis, PCT level and CRP level promptly improved | 0
transferred to the general ward | 0
ertapenem and teicoplanin | 0
debridement, dressing change and symptomatic supportive treatment | 0
repeated blood cultures | 0
negative | 0
repeat CT | 0
size of the hepatic abscess and the amount of ascites decreased | 0
intravenous ertapenem and teicoplanin | 0
symptoms achieved further alleviation | 0
discharged from the hospital | 0
oral antibiotics (clindamycin) | 0
follow-up with a six-week course of intravenous ertapenem | 0
electronic search on PubMed/MEDLINE | 0
Eggerthella lenta | 0
Eubacterium lentum | 0
key words | 0
case studies | 0
English language | 0
published from 1970 through 2020 | 0
E. lenta bacteremia | 0
liver abscess | 0
hepatic puncture and drainage | -1
admitted to our hospital | 0
complaints of right upper quadrant pain and discomfort | 0
right upper quadrant pain | 0
abdominal fullness and distention | 0
abdominal tenderness | 0
fever | 0
abdominal distension | 0
mild bellyache | 0
extreme thirst | 0
temperature of 36.8 °C | 0
fulvous fluid | 0
abdominal and pelvic computed tomography (CT) scan | 0
irregular, slightly low-density lesion in the right posterior hepatic lobe | 0
gas density shadow inside | 0
liquid density shadow and high-density drainage tube shadow | 0
round-like low-density lesion of about 0.8 cm in diameter | 0
thickened appendix | 0
structure of the ascending colon near the ileocecal region became disorganised | 0
multiple gas accumulation and dilation in the bowel | 0
air-fluid levels inside the abdomen | 0
hepatic abscesses | 0
ileus | 0
mild ascites | 0
appendicitis | 0
liver cyst | 0
abdominal infection | 0
peritonitis | 0
surgical exploration | 0
fulvous purulent exudate and necrotic tissue | 0
partial postnecrotic defect in the peritoneum | 0
massive epiploon adhesion in the right upper abdomen | 0
ileocecal resection | 0
partial resection of the ascending colon | 0
ileostomy and drainage of hepatic, abdominal and extraperitoneal abscesses | 0
orotracheal intubation | 0
hypotension | 0
anemia | 0
fever | 0
transferred to the intensive care unit (ICU) | 0
noradrenaline | 0
ventilator | 0
intravenous hydration | 0
nutritional support therapy | 0
blood transfusion | 0
blood cultures and drainage fluids | 0
tigecycline and piperacillin/tazobactam | 0
body temperature | 0
routine blood count | 0
procalcitonin level | 0
C-reactive protein (CRP) level | 0
elevated leukocyte count | 0
electrocardiogram monitor | 0
pulse rate of 130 beats/minute | 0
positive anaerobic blood culture vials | 0
Gram stain revealed short Gram-positive bacillus without spores | 0
MALDI-TOF MS | 0
E. lenta | 0
antimicrobial susceptibility testing | 0
tigecycline was replaced by teicoplanin | 0
piperacillin/tazobactam was discontinued | 0
ertapenem was added to teicoplanin | 0
cultures of the drainage fluid were obtained | 0
Escherichia coli | 0
ertapenem and teicoplanin | 0
fever, leukocytosis, PCT level and CRP level promptly improved | 0
transferred to the general ward | 0
ertapenem and teicoplanin | 0
debridement, dressing change and symptomatic supportive treatment | 0
repeated blood cultures | 0
negative | 0
repeat CT | 0
size of the hepatic abscess and the amount of ascites decreased | 0
intravenous ertapenem and teicoplanin | 0
symptoms achieved further alleviation | 0
discharged from the hospital | 0
oral antibiotics (clindamycin) | 0
follow-up with a six-week course of intravenous ertapenem | 0
electronic search on PubMed/MEDLINE | 0
Eggerthella lenta | 0
Eubacterium lentum | 0
key words | 0
case studies | 0
English language | 0
published from 1970 through 2020 | 0
E. lenta bacteremia | 0
liver abscess | 0
hepatic puncture and drainage | -1
admitted to our hospital | 0
complaints of right upper quadrant pain and discomfort | 0
right upper quadrant pain | 0
abdominal fullness and distention | 0
abdominal tenderness | 0
fever | 0
abdominal distension | 0
mild bellyache | 0
extreme thirst | 0
temperature of 36.8 °C | 0
fulvous fluid | 0
abdominal and pelvic computed tomography (CT) scan | 0
irregular, slightly low-density lesion in the right posterior hepatic lobe | 0
gas density shadow inside | 0
liquid density shadow and high-density drainage tube shadow | 0
round-like low-density lesion of about 0.8 cm in diameter | 0
thickened appendix | 0
structure of the ascending colon near the ileocecal region became disorganised | 0
multiple gas accumulation and dilation in the bowel | 0
air-fluid levels inside the abdomen | 0
hepatic abscesses | 0
ileus | 0
mild ascites | 0
appendicitis | 0
liver cyst | 0
abdominal infection | 0
peritonitis | 0
surgical exploration | 0
fulvous purulent exudate and necrotic tissue | 0
partial postnecrotic defect in the peritoneum | 0
massive epiploon adhesion in the right upper abdomen | 0
ileocecal resection | 0
partial resection of the ascending colon | 0
ileostomy and drainage of hepatic, abdominal and extraperitoneal abscesses | 0
orotracheal intubation | 0
hypotension | 0
anemia | 0
fever | 0
transferred to the intensive care unit (ICU) | 0
noradrenaline | 0
ventilator | 0
intravenous hydration | 0
nutritional support therapy | 0
blood transfusion | 0
blood cultures and drainage fluids | 0
tigecycline and piperacillin/tazobactam | 0
body temperature | 0
routine blood count | 0
procalcitonin level | 0
C-reactive protein (CRP) level | 0
elevated leukocyte count | 0
electrocardiogram monitor | 0
pulse rate of 130 beats/minute | 0
positive anaerobic blood culture vials | 0
Gram stain revealed short Gram-positive bacillus without spores | 0
MALDI-TOF MS | 0
E. lenta | 0
antimicrobial susceptibility testing | 0
tigecycline was replaced by teicoplanin | 0
piperacillin/tazobactam was discontinued | 0
ertapenem was added to teicoplanin | 0
cultures of the drainage fluid were obtained | 0
Escherichia coli | 0
ertapenem and teicoplanin | 0
fever, leukocytosis, PCT level and CRP level promptly improved | 0
transferred to the general ward | 0
ertapenem and teicoplanin | 0
debridement, dressing change and symptomatic supportive treatment | 0
repeated blood cultures | 0
negative | 0
repeat CT | 0
size of the hepatic abscess and the amount of ascites decreased | 0
intravenous ertapenem and teicoplanin | 0
symptoms achieved further alleviation | 0
discharged from the hospital | 0
oral antibiotics (clindamycin) | 0
follow-up with a six-week course of intravenous ertapenem | 0
electronic search on PubMed/MEDLINE | 0
Eggerthella lenta | 0
Eubacterium lentum | 0
key words | 0
case studies | 0
English language | 0
published from 1970 through 2020 | 0
E. lenta bacteremia | 0
liver abscess | 0
hepatic puncture and drainage | -1
admitted to our hospital | 0
complaints of right upper quadrant pain and discomfort | 0
right upper quadrant pain | 0
abdominal fullness and distention | 0
abdominal tenderness | 0
fever | 0
abdominal distension | 0
mild bellyache | 0
extreme thirst | 0
temperature of 36.8 °C | 0
fulvous fluid | 0
abdominal and pelvic computed tomography (CT) scan | 0
irregular, slightly low-density lesion in the right posterior hepatic lobe | 0
gas density shadow inside | 0
liquid density shadow and high-density drainage tube shadow | 0
round-like low-density lesion of about 0.8 cm in diameter | 0
thickened appendix | 0
structure of the ascending colon near the ileocecal region became disorganised | 0
multiple gas accumulation and dilation in the bowel | 0
air-fluid levels inside the abdomen | 0
hepatic abscesses | 0
ileus | 0
mild ascites | 0
appendicitis | 0
liver cyst | 0
abdominal infection | 0
peritonitis | 0
surgical exploration | 0
fulvous purulent exudate and necrotic tissue | 0
partial postnecrotic defect in the peritoneum | 0
massive epiploon adhesion in the right upper abdomen | 0
ileocecal resection | 0
partial resection of the ascending colon | 0
ileostomy and drainage of hepatic, abdominal and extraperitoneal abscesses | 0
orotracheal intubation | 0
hypotension | 0
anemia | 0
fever | 0
transferred to the intensive care unit (ICU) | 0
noradrenaline | 0
ventilator | 0
intravenous hydration | 0
nutritional support therapy | 0
blood transfusion | 0
blood cultures and drainage fluids | 0
tigecycline and piperacillin/tazobactam | 0
body temperature | 0
routine blood count | 0
procalcitonin level | 0
C-reactive protein (CRP) level | 0
elevated leukocyte count | 0
electrocardiogram monitor | 0
pulse rate of 130 beats/minute | 0
positive anaerobic blood culture vials | 0
Gram stain revealed short Gram-positive bacillus without spores | 0
MALDI-TOF MS | 0
E. lenta | 0
antimicrobial susceptibility testing | 0
tigecycline was replaced by teicoplanin | 0
piperacillin/tazobactam was discontinued | 0
ertapenem was added to teicoplanin | 0
cultures of the drainage fluid were obtained | 0
Escherichia coli | 0
ertapenem and teicoplanin | 0
fever, leukocytosis, PCT level and CRP level promptly improved | 0
transferred to the general ward | 0
ertapenem and teicoplanin | 0
debridement, dressing change and symptomatic supportive treatment | 0
repeated blood cultures | 0
negative | 0
repeat CT | 0
size of the hepatic abscess and the amount of ascites decreased | 0
intravenous ertapenem and teicoplanin | 0
symptoms achieved further alleviation | 0
discharged from the hospital | 0
oral antibiotics (clindamycin) | 0
follow-up with a six-week course of intravenous ertapenem | 0
electronic search on PubMed/MEDLINE | 0
Eggerthella lenta | 0
Eubacterium lentum | 0
key words | 0
case studies | 0
English language | 0
published from 1970 through 2020 | 0
E. lenta bacteremia | 0
liver abscess | 0
hepatic puncture and drainage | -1
admitted to our hospital | 0
complaints of right upper quadrant pain and discomfort | 0
right upper quadrant pain | 0
abdominal fullness and distention | 0
abdominal tenderness | 0
fever | 0
abdominal distension | 0
mild bellyache | 0
extreme thirst | 0
temperature of 36.8 °C | 0
fulvous fluid | 0
abdominal and pelvic computed tomography (CT) scan | 0
irregular, slightly low-density lesion in the right posterior hepatic lobe | 0
gas density shadow inside | 0
liquid density shadow and high-density drainage tube shadow | 0
round-like low-density lesion of about 0.8 cm in diameter | 0
thickened appendix | 0
structure of the ascending colon near the ileocecal region became disorganised | 0
multiple gas accumulation and dilation in the bowel | 0
air-fluid levels inside the abdomen | 0
hepatic abscesses | 0
ileus | 0
mild ascites | 0
appendicitis | 0
liver cyst | 0
abdominal infection | 0
peritonitis | 0
surgical exploration | 0
fulvous purulent exudate and necrotic tissue | 0
partial postnecrotic defect in the peritoneum | 0
massive epiploon adhesion in the right upper abdomen | 0
ileocecal resection | 0
partial resection of the ascending colon | 0
ileostomy and drainage of hepatic, abdominal and extraperitoneal abscesses | 0
orotracheal intubation | 0
hypotension | 0
anemia | 0
fever | 0
transferred to the intensive care unit (ICU) | 0
noradrenaline | 0
ventilator | 0
intravenous hydration | 0
nutritional support therapy | 0
blood transfusion | 0
blood cultures and drainage fluids | 0
tigecycline and piperacillin/tazobactam | 0
body temperature | 0
routine blood count | 0
procalcitonin level | 0
C-reactive protein (CRP) level | 0
elevated leukocyte count | 0
electrocardiogram monitor | 0
pulse rate of 130 beats/minute | 0
positive anaerobic blood culture vials | 0
Gram stain revealed short Gram-positive bacillus without spores | 0
MALDI-TOF MS | 0
E. lenta | 0
antimicrobial susceptibility testing | 0
tigecycline was replaced by teicoplanin | 0
piperacillin/tazobactam was discontinued | 0
ertapenem was added to teicoplanin | 0
cultures of the drainage fluid were obtained | 0
Escherichia coli | 0
ertapenem and teicoplanin | 0
fever, leukocytosis, PCT level and CRP level promptly improved | 0
transferred to the general ward | 0
ertapenem and teicoplanin | 0
debridement, dressing change and symptomatic supportive treatment | 0
repeated blood cultures | 0
negative | 0
repeat CT | 0
size of the hepatic abscess and the amount of ascites decreased | 0
intravenous ertapenem and teicoplanin | 0
symptoms achieved further alleviation | 0
discharged from the hospital | 0
oral antibiotics (clindamycin) | 0
follow-up with a six-week course of intravenous ertapenem | 0
electronic search on PubMed/MEDLINE | 0
Eggerthella lenta | 0
Eubacterium lentum | 0
key words | 0
case studies | 0
English language | 0
published from 1970 through 2020 | 0
E. lenta bacteremia | 0
liver abscess | 0
hepatic puncture and drainage | -1
admitted to our hospital | 0
complaints of right upper quadrant pain and discomfort | 0
right upper quadrant pain | 0
abdominal fullness and distention | 0
abdominal tenderness | 0
fever | 0
abdominal distension | 0
mild bellyache | 0
extreme thirst | 0
temperature of 36.8 °C | 0
fulvous fluid | 0
abdominal and pelvic computed tomography (CT) scan | 0
irregular, slightly low-density lesion in the right posterior hepatic lobe | 0
gas density shadow inside | 0
liquid density shadow and high-density drainage tube shadow | 0
round-like low-density lesion of about 0.8 cm in diameter | 0
thickened appendix | 0
structure of the ascending colon near the ileocecal region became disorganised | 0
multiple gas accumulation and dilation in the bowel | 0
air-fluid levels inside the abdomen | 0
hepatic abscesses | 0
ileus | 0
mild ascites | 0
appendicitis | 0
liver cyst | 0
abdominal infection | 0
peritonitis | 0
surgical exploration | 0
fulvous purulent exudate and necrotic tissue | 0
partial postnecrotic defect in the peritoneum | 0
massive epiploon adhesion in the right upper abdomen | 0
ileocecal resection | 0
partial resection of the ascending colon | 0
ileostomy and drainage of hepatic, abdominal and extraperitoneal abscesses | 0
orotracheal intubation | 0
hypotension | 0
anemia | 0
fever | 0
transferred to the intensive care unit (ICU) | 0
noradrenaline | 0
ventilator | 0
intravenous hydration | 0
nutritional support therapy | 0
blood transfusion | 0
blood cultures and drainage fluids | 0
tigecycline and piperacillin/tazobactam | 0
body temperature | 0
routine blood count | 0
procalcitonin level | 0
C-reactive protein (CRP) level | 0
elevated leukocyte count | 0
electrocardiogram monitor | 0
pulse rate of 130 beats/minute | 0
positive anaerobic blood culture vials | 0
Gram stain revealed short Gram-positive bacillus without spores | 0
MALDI-TOF MS | 0
E. lenta | 0
antimicrobial susceptibility testing | 0
tigecycline was replaced by teicoplanin | 0
piperacillin/tazobactam was discontinued | 0
ertapenem was added to teicoplanin | 0
cultures of the drainage fluid were obtained | 0
Escherichia coli | 0
ertapenem and teicoplanin | 0
fever, leukocytosis, PCT level and CRP level promptly improved | 0
transferred to the general ward | 0
ertapenem and teicoplanin | 0
debridement, dressing change and symptomatic supportive treatment | 0
repeated blood cultures | 0
negative | 0
repeat CT | 0
size of the hepatic abscess and the amount of ascites decreased | 0
intravenous ertapenem and teicoplanin | 0
symptoms achieved further alleviation | 0
discharged from the hospital | 0
oral antibiotics (clindamycin) | 0
follow-up with a six-week course of intravenous ertapenem | 0
electronic search on PubMed/MEDLINE | 0
Eggerthella lenta | 0
Eubacterium lentum | 0
key words | 0
case studies | 0
English language | 0
published from 1970 through 2020 | 0
E. lenta bacteremia | 0
liver abscess | 0
hepatic puncture and drainage | -1
admitted to our hospital | 0
complaints of right upper quadrant pain and discomfort | 0
right upper quadrant pain | 0
abdominal fullness and distention | 0
abdominal tenderness | 0
fever | 0
abdominal distension | 0
mild bellyache | 0
extreme thirst | 0
temperature of 36.8 °C | 0
fulvous fluid | 0
abdominal and pelvic computed tomography (CT) scan | 0
irregular, slightly low-density lesion in the right posterior hepatic lobe | 0
gas density shadow inside | 0
liquid density shadow and high-density drainage tube shadow | 0
round-like low-density lesion of about 0.8 cm in diameter | 0
thickened appendix | 0
structure of the ascending colon near the ileocecal region became disorganised | 0
multiple gas accumulation and dilation in the bowel | 0
air-fluid levels inside the abdomen | 0
hepatic abscesses | 0
ileus | 0
mild ascites | 0
appendicitis | 0
liver cyst | 0
abdominal infection | 0
peritonitis | 0
surgical exploration | 0
fulvous purulent exudate and necrotic tissue | 0
partial postnecrotic defect in the peritoneum | 0
massive epiploon adhesion in the right upper abdomen | 0
ileocecal resection | 0
partial resection of the ascending colon | 0
ileostomy and drainage of hepatic, abdominal and extraperitoneal abscesses | 0
orotracheal intubation | 0
hypotension | 0
anemia | 0
fever | 0
transferred to the intensive care unit (ICU) | 0
noradrenaline | 0
ventilator | 0
intravenous hydration | 0
nutritional support therapy | 0
blood transfusion | 0
blood cultures and drainage fluids | 0
tigecycline and piperacillin/tazobactam | 0
body temperature | 0
routine blood count | 0
procalcitonin level | 0
C-reactive protein (CRP) level | 0
elevated leukocyte count | 0
electrocardiogram monitor | 0
pulse rate of 130 beats/minute | 0
positive anaerobic blood culture vials | 0
Gram stain revealed short Gram-positive bacillus without spores | 0
MALDI-TOF MS | 0
E. lenta | 0
antimicrobial susceptibility testing | 0
tigecycline was replaced by teicoplanin | 0
piperacillin/tazobactam was discontinued | 0
ertapenem was added to teicoplanin | 0
cultures of the drainage fluid were obtained | 0
Escherichia coli | 0
ertapenem and teicoplanin | 0
fever, leukocytosis, PCT level and CRP level promptly improved | 0
transferred to the general ward | 0
ertapenem and teicoplanin | 0
debridement, dressing change and symptomatic supportive treatment | 0
repeated blood cultures | 0
negative | 0
repeat CT | 0
size of the hepatic abscess and the amount of ascites decreased | 0
intravenous ertapenem and teicoplanin | 0
symptoms achieved further alleviation | 0
discharged from the hospital | 0
oral antibiotics (clindamycin) | 0
follow-up with a six-week course of intravenous ertapenem | 0
electronic search on PubMed/MEDLINE | 0
Eggerthella lenta | 0
Eubacterium lentum | 0
key words | 0
case studies | 0
English language | 0
published from 1970 through 2020 | 0
E. lenta bacteremia | 0
liver abscess | 0
hepatic puncture and drainage | -1
admitted to our hospital | 0
complaints of right upper quadrant pain and discomfort | 0
right upper quadrant pain | 0
abdominal fullness and distention | 0
abdominal tenderness | 0
fever | 0
abdominal distension | 0
mild bellyache | 0
extreme thirst | 0
temperature of 36.8 °C | 0
fulvous fluid | 0
abdominal and pelvic computed tomography (CT) scan | 0
irregular, slightly low-density lesion in the right posterior hepatic lobe | 0
gas density shadow inside | 0
liquid density shadow and high-density drainage tube shadow | 0
round-like low-density lesion of about 0.8 cm in diameter | 0
thickened appendix | 0
structure of the ascending colon near the ileocecal region became disorganised | 0
multiple gas accumulation and dilation in the bowel | 0
air-fluid levels inside the abdomen | 0
hepatic abscesses | 0
ileus | 0
mild ascites | 0
appendicitis | 0
liver cyst | 0
abdominal infection | 0
peritonitis | 0
surgical exploration | 0
fulvous purulent exudate and necrotic tissue | 0
partial postnecrotic defect in the peritoneum | 0
massive epiploon adhesion in the right upper abdomen | 0
ileocecal resection | 0
partial resection of the ascending colon | 0
ileostomy and drainage of hepatic, abdominal and extraperitoneal abscesses | 0
orotracheal intubation | 0
hypotension | 0
anemia | 0
fever | 0
transferred to the intensive care unit (ICU) | 0
noradrenaline | 0
ventilator | 0
intravenous hydration | 0
nutritional support therapy | 0
blood transfusion | 0
blood cultures and drainage fluids | 0
tigecycline and piperacillin/tazobactam | 