55 years old | 0
female | 0
Saudi | 0
admitted to the hospital | 0
end-stage liver disease | -720
cryptogenic cirrhosis | -720
type 2 diabetes mellitus | -720
oral metformin | -720
hypertension | -720
oral amlodipine | -720
non-smoker | 0
no alcohol consumption | 0
no history of drug abuse | 0
fever | -24
cough | -24
progressive lower limb edema | -24
abdominal distention | -24
admitted to hospital for one week | -168
liver transplantation team | -168
temperature 37.7°C | 0
heart rate 111 beats per minute | 0
respiratory rate 26 breaths per minute | 0
normal blood pressure | 0
oxygen saturation on breathing room air | 0
mild peripheral blood leukocytosis | 0
platelets 41×10^9/L | 0
albumin 26 g/L | 0
bilirubin 47 µmol/L | 0
creatinine 59 µmol/L | 0
screen for infection | 0
blood examination | 0
sputum examination | 0
urine examination | 0
ascitic fluid examination | 0
chest X-ray | 0
right-sided pleural effusion | 0
hydrothorax | 0
possible consolidation | 0
empirically on antibiotics | 0
diuretics dosage increased | 0
ascitic and pleural fluid drained | 0
urine culture positive for Streptococcus agalactiae | 0
sensitive to antimicrobials | 0
clinical condition improved | 24
repeated chest X-ray | 24
reduction in right hydrothorax | 24
discharged home | 168
oral ciprofloxacin | 168
oral lasix | 168
multivitamin tablets | 168
admitted to hospital for liver transplant | 720
live organ donation | 720
total hepatectomy | 720
transplantation using full right lobe graft | 720
three biliary anastomoses | 720
arterial anastomosis repeated twice | 720
transfusion of 12 units packed red blood cells | 720
transferred to ICU | 720
extubated after 24 hours | 744
re-intubated for 24 hours | 768
ARDS | 768
immunosuppressive therapy | 816
oral tacrolimus | 816
oral mycophenolate mofetil | 816
oral prednisolone | 816
anastomotic biliary stricture | 1008
bile leak | 1008
PTC | 1008
PTBD | 1008
internal-external biliary catheter | 1008
pigtail catheter | 1008
drains kept in place for few weeks | 1008
pigtail catheter removed | 1056
internal-external PTBD catheter left in place | 1056
right upper quadrant abdominal pain | 1344
no fever | 1344
no vomiting | 1344
no change in peripheral blood leukocyte count | 1344
no change in bilirubin | 1344
no change in ALT | 1344
no change in alkaline phosphatase | 1344
CRP increased | 1344
ultrasound of abdomen | 1344
right-sided sub-diaphragmatic collection | 1344
septic screen | 1344
blood sampling | 1344
urine sampling | 1344
biliary drain fluid sampling | 1344
abdominal collection sampling | 1344
IV meropenem | 1344
culture from PTBD catheter positive for E. meningoseptica | 1344
multidrug-resistant organism | 1344
IV meropenem changed to IV ciprofloxacin | 1392
metronidazole | 1392
repeat cultures from PTBD catheter | 1440
repeat culture results positive for E. meningoseptica | 1440
clinical condition improved | 1440
abdominal pain resolved | 1440
decision to continue antibiotics for two weeks | 1440
asymptomatic | 1560
normal peripheral blood leukocyte count | 1560
CRP dropped | 1560
repeat fluid cultures from PTBD catheter negative | 1560
no complications from antibiotic treatment | 1560