40 years old | 0
male | 0
businessman | 0
admitted to ICU | 0
fever with chills | -480
vomiting | -96
seizures | -96
decreased urine output | -96
shock | 0
intubated | 0
mechanical ventilation | 0
icteric | 0
acute kidney injury | 0
dengue antigen non-structural (NS1) positive | -480
malaria negative | -480
enteric fever negative | -480
hematocrit 35.2% | 0
total leukocyte count 9600/mm3 | 0
coagulopathy | 0
endotracheal bleed | 0
anuria | 0
liver function deteriorating | 0
septic shock | 0
lung protective mechanical ventilation | 0
slow low efficiency daily dialysis | 0
vasopressors (noradrenaline) | 0
broad spectrum antibiotics (ceftriaxone) | 0
artesunate | 0
dengue IgM positive | 0
Leptospira IgM positive | 0
HEV IgM positive | 0
malaria test negative | 0
enteric fever test negative | 0
hepatitis A test negative | 0
hepatitis B test negative | 0
hepatitis C test negative | 0
human immunodeficiency virus test negative | 0
serum procalcitonin rising | 0
no growth of organisms from blood | 0
no growth of organisms from endotracheal samples | 0
no growth of organisms from urine samples | 0
condition deteriorated | 120
died | 144
renal biopsy not done | 144
liver biopsy not done | 144
thrombocytopenia | 0
endothelial dysfunction | 0
cytokine expression | 0
chemokines expression | 0
adhesion molecules expression | 0
T-lymphocytes activation | 0
hemostatic system dysfunction | 0
co-infection detected | 0
triple co-infection | 0
rapid urbanization | 0
increasing population density | 0
frequent travel | 0
poor water drainage infrastructure | 0
inadequate vector control measures | 0
high mortality | 0
high morbidity | 0
endothelial dysfunction related mortality | 0
antibodies against NS proteins | 0
cross-reactivity with endothelial cells | 0
tumor necrosis factor alpha-α production | 0
interleukin-8 production | 0
nitric oxide production | 0
renal dysfunction | 0
cerebral edema | 0
disseminated intravascular coagulation | 0
microscopic agglutination test not available | 0
IgM ELISA test for leptospira | 0
IgM ELISA test for HEV | 0
RT-PCR testing not done | 0
HEV RNA viremia not demonstrated | 0
early treatment initiation | 0
early detection of co-infection | 0
early endothelial involvement | 0
favorable outcome | 0