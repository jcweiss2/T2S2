38 years old | 0
female | 0
gravida 2 | 0
para 1 | 0
admitted to the Department of Obstetrics | 0
difficulty walking | -672
pain in right inguinal region | -672
pain in lower back | -672
low-lying placenta | -672
elective Caesarean section scheduled | -672
body temperature 36.3°C | -24
pulse rate 83 beats/min | -24
blood pressure 116/50 mmHg | -24
respiratory rate 15 breaths/min | -24
SpO2 98% | -24
lower abdominal pain | -24
massive vaginal bleeding | -24
emergency Caesarean section | 0
dramatically deteriorating dyspnea | 0
transferred to ICU | 0
chest X-ray showed cardiac dilatation and opacity | 0
anemia | 0
Hb level 6.1 g/dL | 0
bilateral pleural effusions | 24
multiple lung nodules | 24
multiple liver masses | 24
multiple osteolytic changes | 24
thrombi in splenic vein | 24
thrombi in abdominal inferior vena cava | 24
thrombi in left common iliac vein | 24
no signs of pulmonary embolism | 24
SpO2 deteriorated to 94% | 24
non-invasive positive-pressure ventilation | 24
diuretic | 24
resolution of respiratory distress | 48
transferred to Division of General Medicine | 72
left hip pain | 72
body temperature 37.1°C | 72
pulse rate 93 beats/min | 72
blood pressure 126/82 mmHg | 72
respiratory rate 25 breaths/min | 72
SpO2 96% | 72
conjunctiva anemic and icteric | 72
lymph nodes palpated on left side of neck | 72
lymph nodes palpated superior to left clavicle | 72
respiratory sounds attenuated | 72
bilateral breast engorgement | 72
Caesarean operation scar | 72
white blood cell count 11,470/μL | 72
normocytic normochromic anemia | 72
hypoalbuminemia | 72
elevated lactate dehydrogenase | 72
elevated alkaline phosphatase | 72
elevated tumor markers | 72
pleural fluid cytology revealed adenocarcinoma | 120
sputum cytology revealed adenocarcinoma | 120
stopped breastfeeding | 120
oxygen therapy changed to nasal high-flow oxygen | 168
cell block cytology of pleural effusion revealed adenocarcinoma | 168
immunostaining positive for CK7 | 168
immunostaining positive for TTF-1 | 168
immunostaining positive for napsin A | 168
immunostaining negative for CK20 | 168
estrogen receptor 1-5% positive | 168
EGFR mutation detected | 216
gefitinib therapy initiated | 216
transferred to Division of Respiratory Medicine | 240
pleural effusion reduced | 240
SpO2 improved | 240
discharged | 360
continued treatment on outpatient basis | 360