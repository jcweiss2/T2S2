54 years old | 0
male | 0
type 2 diabetes mellitus | 0
acute abdominal pain | -48
fever | 0
blood pressure 82/45 mmHg | 0
pulse rate 135/min | 0
distended abdomen | 0
tight abdomen | 0
no jaundice | 0
diabetic ketoacidosis | 0
elevated white blood cells 24000/mm³ | 0
high C-reactive protein 270 mg/l | 0
normal liver function tests | 0
massive ascites | 0
increased gallbladder wall thickness | 0
resolved gallbladder distention | 0
no pneumoperitoneum | 0
no choledocholithiasis | 0
diagnostic paracentesis | 0
bile ascites | 0
exploratory laparotomy | 0
diffuse biliary peritonitis | 0
retroperitoneal cavity bile staining | 0
peritoneal lavage | 0
no duodenal perforation | 0
no gallbladder perforation | 0
cholecystectomy | 0
intraoperative cholangiography | 0
common bile duct extravasation | 0
perforation repair over T-tube | 0
Salem tube drainage | 0
discharged | 360
T-tube removal | 768
normal cholangiogram | 768
no biliary leakage | 768
no pancreaticobiliary junction | 768
no distal stricture | 768
symptoms not recurred | 768
ulcerous acalculous cholecystitis | 0
