63 years old | 0
male | 0
admitted to the hospital | 0
hypertension | -6720
chronic back pain | -6720
spinal stenosis | -6720
lower extremity edema | -6720
oxycodone | -6720
losartan | -6720
furosemide started | -6720
watery diarrhea | -336
hematochezia | -336
abdominal pain | -336
diffuse maculopapular rash | -168
itch | -168
dry cough | -168
nonproductive cough | -168
fever up to 38.6°C | -168
furosemide discontinued | -168
moderate distress | 0
temperature 38.6°C | 0
blood pressure 126/59 mm Hg | 0
heart rate 103 bpm | 0
respiratory rate 22 bpm | 0
oxygen saturation 95% | 0
diffuse erythematous maculopapular rash | 0
no conjunctival injection | 0
no mucosal involvement | 0
tachycardia | 0
normal cardiovascular exam | 0
clear lungs | 0
soft abdomen | 0
nontender abdomen | 0
no hepatosplenomegaly | 0
no focal neurological deficits | 0
leukocytosis 11.8×10^9/L | 0
elevated eosinophil count 1.29×10^9/L | 0
normal hemoglobin | 0
normal platelets | 0
normal creatinine | 0
normal electrolytes | 0
normal liver enzymes | 0
CRP 229 | 0
ESR 31 | 0
hypoxemia | 0
partial oxygen 66 mm Hg | 0
hilar lymphadenopathy | 0
interstitial changes | 0
pneumonitis | 0
levofloxacin | 0
IV fluids | 0
rash worsened | 24
cough persisted | 24
fever persisted | 24
thrombocytopenia | 24
doxycycline | 24
afebrile | 48
cough persisted | 48
eosinophilic leukocytosis persisted | 48
furosemide resumed | 72
rash worsened | 72
hypoxia | 72
dyspnea | 72
fever up to 39.4°C | 72
leukocytosis worsened | 72
eosinophilia worsened | 72
acute kidney injury | 72
atrial fibrillation | 72
rapid ventricular response | 72
DRESS syndrome suspected | 72
negative infectious workup | 96
negative autoimmune workup | 96
hematuria | 96
proteinuria | 96
skin biopsy consistent with drug reaction | 96
normal LV ejection fraction | 120
no pericardial effusion | 120
no wall motion abnormalities | 120
negative troponin | 120
negative CK-MB | 120
negative TSH | 120
amiodarone | 120
steroids initiated | 120
prednisone 1 mg/kg daily | 120
levofloxacin discontinued | 120
doxycycline discontinued | 120
clinical improvement | 144
discharged | 144
prednisone taper | 144
atovaquone prophylaxis | 144
spironolactone | 144
fatigue | 1008
mild shortness of breath | 1008
insomnia | 1008
normalized labs | 1008
