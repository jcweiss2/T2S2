64 years old | 0
    male | 0
    type 2 diabetes | 0
    hypertension | 0
    kidney transplant recipient | 0
    tacrolimus | 0
    mycophenolic acid | 0
    prednisone | 0
    progressive shortness of breath | -96
    recurrent fever | -96
    cough | -96
    admitted to the emergency department | 0
    serum creatinine 0.7 mg/dL | 0
    GFR >60 ml/min/1.73 m2 | 0
    chest radiography showing diffuse interstitial and airspace opacities | 0
    gram stain negative | 0
    rapid influenza test negative | 0
    pneumococcal urinary antigen test negative | 0
    legionella urinary antigen test negative | 0
    SARS-CoV-2 positive | 0
    admitted to the intensive care unit | 0
    electively intubated | 0
    hydroxychloroquine | 0
    azithromycin | 0
    cefepime | 0
    mycophenolic acid suspension | 0
    tacrolimus reduction | 0
    prednisone continuation | 0
    low tidal volume lung-protective strategy | 0
    prone positioning | 0
    neuromuscular blockade (atracurium) | 0
    high positive end-expiratory pressure therapy | 0
    day 3 sputum sample redrawn | 72
    increased endotracheal secretions | 72
    worsening CXR | 72
    hypoxemia | 72
    high dose corticosteroids (60 mg IV methylprednisolone) | 72
    sputum positive for gram-negative bacilli | 96
    S. maltophilia identified | 120
    TMP/SMX initiated | 120
    cefepime discontinued | 120
    AKI developed | 168
    serum creatinine 2.1 mg/dL | 168
    oliguria | 168
    TMP/SMX discontinued | 192
    levofloxacin initiated | 192
    serum creatinine 3.4 mg/dL | 192
    GFR 18 ml/min/1.73 m2 | 192
    hyperkalemia (6.1 mmol/L) | 192
    hemodialysis initiated | 192
    urinalysis no eosinophiluria | 192
    urinalysis no white cell casts | 192
    steroids continued | 192
    tacrolimus levels therapeutic | 192
    kidney biopsy considered unsafe | 192
    remdesivir unavailable | 192
    convalescent plasma unavailable | 192
    supportive therapy continued | 192
    oxygenation declined | 264
    clinical status declined | 264
    comfort care measures | 264
    death | 288
    