7 years old | 0
male | 0
admitted to the hospital | 0
generalized convulsive status epilepticus | 0
fever | -96
diffuse skin rash | -96
right tibia fracture | -336
maculopapular rash | 0
nonpurulent conjunctivitis | 0
cracked, fissured lips | 0
cervical lymphadenopathy | 0
fever of 39°C | 0
meningeal signs were negative | 0
Glasgow Coma Scale (GCS) score was 7 | 0
seizure treated and stopped with administration of one dose of midazolam and phenobarbital | 0
treated with phenobarbital, ceftriaxone, acyclovir, and osmotic therapy with mannitol | 0
intubated with initiation of mechanical ventilation | 24
respiratory failure | 24
urgent brain magnetic resonance imaging (MRI) | 24
cerebral vasculitis | 24
severe encephalitis | 24
treated with IVIG as a single infusion of 2 g/kg along with acetylsalicylic acid (50 mg/kg/day) | 48
fever resolved | 48
disappearance of skin rash | 48
mild improvement in the level of consciousness | 48
successfully extubated | 72
acyclovir treatment was discontinued | 72
confused, occasionally extremely irritable and delirious | 72
persistence of GCS score in the range of 8–10 | 72
recurrence of fever | 72
brain MRI showed progression of initially noted changes | 120
intravenous steroid pulse therapy (methylprednisolone 30 mg/kg/day for 5 days) | 216
oral prednisolone (2 mg/kg/day) | 216
response to steroid therapy was excellent | 216
significant improvement in neurological status | 216
full motor function recovery | 360
improvement of cognitive function | 360
periungual desquamation of the fingers | 504
repeated echocardiogram was normal | 504
discharged | 1080
follow-up brain MRI, 2 months after the onset of the disease, did not reveal areas with restricted water diffusion | 1440
T2W image showed parenchymal atrophy | 1440
3D-TOF MR angiography confirmed normalization of the cerebral circulation | 1440
dosage of corticosteroids was gradually decreased and then stopped completely | 2160