29 years old | 0
female | 0
admitted to the hospital | 0
history of chronic ulcerative pancolitis | -8760
history of autoimmune hepatitis | -8760
history of cirrhosis | -8760
treated with azathioprine | -8760
treated with corticosteroids | -8760
fever | -96
left leg pain | -96
diarrhoea | -96
septic shock | 10
temperature 39.4°C | 10
heart rate 120 beats per minute | 10
blood pressure 70/50 mm Hg | 10
oxygen saturation 50% | 10
acute respiratory distress | 10
Glasgow Coma Score 8 | 10
purpuric erythema | 10
mechanical ventilation | 10
large-volume expansion | 10
cathecholaminergic support by adrenaline | 10
cardiac arrest | 10
low-flow time 5 minutes | 10
acute renal failure | 10
increased creatinine kinase level | 10
disseminated intravascular coagulation | 10
leucopenia | 10
hepatocellular failure | 10
lactate level 16 mmol/L | 10
C-reactive protein 13.4 mg/L | 10
broad-spectrum antibiotic therapy with piperacillin–tazobactam | 10
broad-spectrum antibiotic therapy with vancomycin | 10
broad-spectrum antibiotic therapy with amikacin | 10
clindamycin | 12
bullae | 12
superficial excoriations | 12
erythema | 12
leg and abdomen computed tomography | 12
subcutaneous fat infiltration | 12
diagnosis of NSTI | 12
surgery | 14
extensive debridement of cutaneous and subcutaneous tissues | 14
necrotizing fascia | 14
continuous renal replacement therapy | 14
haemorrhagic shock | 14
massive transfusions | 14
second surgery debridement | 38
skin lesions extensive | 38
subcutaneous crackles | 38
lake of bleeding | 38
necrotizing fascia | 38
death | 38
E. coli strain belonged to phylogenetic group C | 0
E. coli strain carried genes encoding yersiniabactin | 0
E. coli strain carried genes encoding aerobactin | 0
E. coli strain carried genes encoding salmochelin | 0
E. coli strain carried genes encoding hemolysin | 0
E. coli strain carried genes encoding cytotoxic necrotizing factor 1 | 0
E. coli strain carried genes encoding adhesin/invasin Hra | 0
E. coli strain carried genes encoding P fimbriae pilin PapC | 0