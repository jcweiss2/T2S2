69 years old | 0
male | 0
admitted to the hospital | 0
cough | -72
sputum | -72
fever | -72
drowsy mental status | -72
traumatic intracranial hemorrhage | -504
epidural hemorrhage | -504
subdural hemorrhage | -504
accidental fall | -504
right craniectomy | -504
ventriculoperitoneal shunt | -504
posttraumatic hydrocephalus | -504
intensive rehabilitation treatment | -128
antipsychotic medication | -168
drowsiness | -168
aspiration event | -168
respiratory symptoms | -168
deteriorating mental status | -168
focal infiltrate at left lower lung field | 0
consolidation with air bronchogram | 0
aspirated materials at left upper lobe bronchus | 0
aspirated materials at LLL segmental bronchus | 0
food particles in esophagus | 0
pneumonia | 0
aspiration-induced pneumonia | 0
brain CT scan | 0
no notable findings | 0
previously inserted VP shunt | 0
focal encephalomalacic changes in right frontal lobe | 0
mental change due to pneumonia-induced sepsis | 0
oxygen partial pressure 43.9 mm Hg | 0
oxygen saturation 79.4% | 0
respiratory rate 24 breaths/minute | 0
high-flow nasal oxygen therapy | 0
fraction of inspired oxygen 0.5 | 0
flow 50 L/minute | 0
oxygen saturation 93-97% | 0
respiratory rate 22-26 breaths/minute | 0
comfortable respiration | 0
repeated sudden desaturation | 24
endotracheal intubation | 24
mechanical ventilation | 24
desaturation due to airway secretion | 24
attempted weaning from MV | 48
unable to effectively expectorate airway secretions | 48
alert mental status | 48
extubation | 48
high-flow nasal cannula | 48
FiO2 0.4 | 48
flow 50 L/minute | 48
oxygen saturation 93-100% | 48
transferred to general ward | 72
high-flow nasal cannula setting changed | 72
flow 40 L/minute | 72
FiO2 0.4 | 72
mentation became drowsy | 100
stupor | 100
brain CT scan | 100
pneumocephalus | 100
midline shifting | 100
near-collapse of left ventricle | 100
Mount Fuji sign | 100
tension pneumocephalus | 100
high-flow nasal cannula stopped | 100
simple nasal cannula | 100
follow-up brain CT scan | 112
pneumocephalus slightly decreased | 112
facial bone CT scan | 112
skull base fractures | 112
right frontal sinus | 112
ethmoidal sinuses | 112
positive pressure ventilation | 112
mental status improved | 168
follow-up brain CT | 168
pneumocephalus markedly decreased | 168
midline shifting improved | 168
left ventricle structure improved | 168
tracheostomy | 240
difficulties in expectorating airway secretions | 240
mental status improved | 280
sudden decline in mental status | 320
stupor | 320
intracranial infection | 320
craniotomy for drainage | 320
mental status did not fully recover | 320