80 years old | 0
    male | 0
    admitted to the hospital | 0
    suspected urinary tract infection | -120
    progressive fever | -120
    dysuria | -120
    clean catch urine specimen collected | -120
    empirically started on cephalexin | -120
    urine analysis positive for large leukocyte esterase | -120
    urine analysis positive for bacteria | -120
    culture grew Escherichia coli | -120
    resistance to ampicillin | -120
    resistance to levofloxacin | -120
    resistance to trimethoprim | -120
    resistance to sulfamethoxazole | -120
    intermediate sensitivity to ampicillin/sulbactam | -120
    sensitivity to cefazolin | -120
    sensitivity to gentamicin | -120
    sensitivity to nitrofurantoin | -120
    prescribed cephalexin 500 mg three times daily | -120
    extensive erythematous rash | -48
    sloughing of the skin | -48
    continued progression of severe reaction | -24
    cephalexin discontinued | 0
    transferred to BICU | 0
    chronic obstructive pulmonary disease | 0
    type 2 diabetes mellitus | 0
    coronary artery disease | 0
    hypertension | 0
    hypothyroidism | 0
    depression | 0
    end-stage renal disease | 0
    hemodialysis | 0
    multiple myocardial infarctions | 0
    ischemic cardiomyopathy | 0
    atrial fibrillation | 0
    home medications included hydrocodone/acetaminophen | 0
    home medications included levothyroxine | 0
    home medications included escitalopram | 0
    home medications included carvedilol | 0
    home medications included guaifenesin | 0
    home medications included docusate | 0
    home medications included calcitriol | 0
    home medications included albuterol | 0
    home medications included amiodarone | 0
    pulmonary infiltrates | 0
    respiratory failure | 0
    intubated | 0
    difficulty swallowing | 0
    endotracheal tube placed | 0
    diagnosed with toxic epidermal necrolysis syndrome | 0
    56% total body surface area involvement | 0
    blood pressure 81/45 mmHg | 0
    respiratory rate 12 breaths/min | 0
    temperature 36.8°C | 0
    WBC count 1.5 × 10³/mm³ | 0
    73% neutrophils | 0
    platelet count 77,000/µL | 0
    serum creatinine 2.12 mg/dL | 0
    venous serum lactate 3.1 mmol/L | 0
    oxygen saturation 99% on 6 L O₂ | 0
    advanced to 15 L O₂ via non-rebreather mask | 0
    pain assessed at 9/10 | 0
    peripheral blood cultures obtained | 0
    skin surveillance cultures of nares | 0
    skin surveillance cultures of axilla | 0
    skin surveillance cultures of groin | 0
    urine culture from Foley catheter | 0
    chest radiograph revealed right pleural effusion | 0
    right lower and left basilar opacities | 0
    marked respiratory distress | 0
    intubated | 0
    norepinephrine and vasopressin drips | 0
    continuous infusion of albumin 25% | 0
    lactated Ringer’s given at 300 mL/h | 0
    tetanus-diphtheria toxoids vaccine administered | 0
    single IV dose of gentamicin 120 mg | 0
    single IV dose of fluconazole 100 mg | 0
    WBC 5.4 × 10³/mm³ | 24
    serum creatinine 1.98 mg/dL | 24
    venous serum lactate 1.8 mmol/L | 24
    random serum gentamicin level 2.4 mg/dL | 24
    redosed with gentamicin 120 mg | 24
    supportive continuous renal replacement therapy | 24
    fluconazole continued at 200 mg IV | 24
    urine culture showed >100,000 cfu/mL Candida species | 24
    Gram’s stain showed Gram-negative rods | 24
    Gram’s stain showed Gram-positive rods | 24
    wide complex tachycardia | 96
    amiodarone restarted | 96
    gentamicin held | 96
    random gentamicin level 2.2 mg/dL | 96
    sloughing of skin over back, chest, upper extremities, abdomen, bilateral thighs, buttocks | 120
    Pseudomonas aeruginosa cultured | 120
    sensitive to anti-pseudomonal beta-lactams | 120
    sensitive to gentamicin | 120
    sensitive to tobramycin | 120
    sensitive to amikacin | 120
    sensitive to colistin | 120
    resistant to doripenem | 120
    resistant to quinolones | 120
    another 120 mg dose of gentamicin | 120
    patient continued to decline | 144
    expired | 144
    cause of death cardiac arrest | 144
    multisystem organ failure | 144
    autopsy reported TEN involving 80% body surface area | 144
    necrotizing bronchopneumonia | 144
    SCORTEN predicted mortality 62% | 144
