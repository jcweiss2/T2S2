65 years old | 0
female | 0
liver cirrhosis | -6720
chronic hepatitis B | -6720
hepatocellular carcinoma | 0
admitted to the hospital | 0
intravenous glycopyrrolate | 0
general anesthesia | 0
propofol | 0
rocuronium | 0
remifentanil | 0
sevoflurane | 0
mechanical ventilation | 0
electrocardiography | 0
arterial blood pressure | 0
central venous pressure | 0
SpO2 | 0
stable vital signs | 0
sudden decrease in arterial blood pressure | 1
tachycardia | 1
ST elevation on EKG | 1
resuscitation | 1
colloid administration | 1
catecholamines administration | 1
intraoperative ultrasonography | 1
massive air emboli | 1
VAE diagnosis | 1
PAE diagnosis | 1
arterial blood gas analysis | 1
catecholamine administration | 1.17
systolic blood pressure maintained | 1.17
heart rate maintained | 1.17
central venous pressure maintained | 1.17
end-tidal carbon dioxide restored | 1.17
ABGA | 1.5
norepinephrine infusion | 1.5
fluid resuscitation | 1.5
air emboli disappeared | 2.17
hepatectomy restarted | 2.17
surgery completed | 5
intensive care unit | 5
mechanical ventilation | 5
norepinephrine infusion | 5
abnormal PT/PTT | 5
fibrinogen | 5
d-dimer | 5
antithrombin III | 5
CK-MB | 5
troponin-T | 5
ST elevation on EKG | 5
EKG findings recovered | 24
trans-thoracic echocardiogram | 24
vital signs stable | 24
norepinephrine infusion tapered out | 24
mental status unchanged | 120
brain CT | 120
brain MRI | 120
multiple acute cerebral infarctions | 120
weaned to spontaneous ventilation | 264
extubated | 264
vital signs unstable | 360
intravenous administration of catecholamines | 360
panperitonitis | 360
gram (+) cocci on peritoneal culture | 360
cardiac arrest | 744
septic shock | 744
expired | 744