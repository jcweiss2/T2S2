74 years old | 0
male | 0
unconscious state | -672
asthma | -8760
nephritic syndrome | -8760
prednisolone | -8760
steroid-induced DM | -672
obesity | -50400
found in unconscious state | 0
transported to hospital | 0
Glasgow Coma Scale, E2V1M4 | 0
blood pressure, no measurable but positive pulsation on carotid artery | 0
heart rate, 110 beats per minute | 0
respiratory rate, 24 breaths per minute | 0
body temperature, 35.2°C | 0
body mass index, 28 | 0
obesity | 0
near obstruction of the airway | 0
left conjugated deviated ocular position | 0
right hemiparesis | 0
hematemesis | 0
double incontinence | 0
complete phimosis with hypogonadism | 0
rapid fluid resuscitation | 0
tracheal intubation | 0
mechanical ventilation | 0
indwelling nasogastric tube placement | 0
infusion of noradrenaline | 0
infusion of vasopressin | 0
sinus tachycardia with complete right bundle branch block | 0
atrophic liver | 0
multiple pancreatic cysts | 0
excess visceral fat | 0
penis buried under a layer of subcutaneous fat | 0
septic shock of unknown focus | 0
acute respiratory failure | 0
renal failure with hyperkalemia | 0
cerebral ischemia | 0
liver cirrhosis | 0
rhabdomyolysis | 0
DM | 0
upper gastrointestinal bleeding | 0
infusion of calcium chloride | 0
insulin therapy | 0
zirconium for hyperkalemia and hyperglycemia | 0
administration of broad-spectrum antibiotics | 0
mineral corticoid for septic shock | 0
emergency circumcision | 0
insertion of balloon catheter | 0
admitted to intensive care unit | 0
circulation stabilized without cardiopressor treatment | 72
PaO2/FiO2 reached >300 | 72
extubated | 72
blood culturing revealed Staphylococcus capitis | 72
steroid dose rapidly decreased | 72
circulation became unstable | 72
steroid dose gradually tapered | 72
adrenal insufficiency suspected | 72
ACTH level, 5 pg/mL | 72
cortisol level, 7.0 μg/dL | 72
adrenal insufficiency confirmed | 72
blood tests for hepatitis B, hepatitis C, and autoimmune antibodies conducted | 72
all tests negative | 72
M2BPGI: Mac-2 binding protein (M2BP) value, 2+ | 72
NAFLD fibrosis score, 2.0 points | 72
FIB-4 index, 9.45 | 72
liver cirrhosis confirmed | 72
burn-out NASH diagnosed | 72
ascites observed on abdominal CT | 144
no fresh ischemic lesions | 144
pituitary gland had normal appearance on cerebral magnetic resonance imaging | 144
initial neurological deficits judged to be due to transient ischemic attack or Todd's paralysis | 144
hypogonadism judged to be induced by NASH | 144
testosterone level, low | 144
estradiol level, high | 144
could feed himself but required assistance for transfer | 168
severe lower extremity muscle weakness due to disuse or critical illness myopathy | 168
respiratory function temporally deteriorated | 360
thrombosis in right pulmonary artery and right common iliac vein | 360
heparinization | 360
renal function returned to normal range | 360
rhabdomyolysis resolved | 360
liver dysfunction, coagulopathy, and anemia remained | 360
left leg phlegmon | 432
treated with antibiotics | 432
esophagogastroscopy showed only atrophic gastritis | 648
transferred to another hospital for rehabilitation | 816