61 years old | 0
male | 0
South Asian | 0
farmer | 0
admitted to the emergency treatment unit | 0
abdominal pain | -72
distension | -72
vomiting | -72
constipation | -72
diagnosed with type 2 diabetes mellitus | -13140
diagnosed with hypertension | -13140
treated with Metformin | -13140
treated with gliclazide | -13140
treated with amlodipine | -13140
febrile | 0
confused | 0
Glasgow coma scale of 10 | 0
low volume and thready pulse | 0
pulse rate of 130 per min | 0
noninvasive blood pressure of 70/40 mmHg | 0
rapid breathing | 0
peripheral oxygen saturation of 88% | 0
abdomen grossly distended with gas | 0
flank dullness | 0
diffuse tenderness | 0
guarding | 0
rigidity | 0
bowel sounds not audible | 0
presumptive diagnosis of septic shock | 0
arterial blood gas analysis | 0
septic screening | 0
broad-spectrum antibiotics | 0
30 mL/kg intravenous fluid bolus | 0
subclavian central venous line inserted | 0
noradrenaline infusion | 0
adrenaline infusion | 0
invasive arterial pressure monitoring | 0
elective intubation of the trachea | 0
inferior vena cava distensibility of 35% | 0
left ventricular volume status in the 2d echocardiogram | 0
hypovolaemia | 0
moderately impaired cardiac contractility | 0
dobutamine infusion | 0
left lateral decubitus X-ray abdomen | 0
grossly distended small bowel loops | 0
no air under the diaphragm | 0
ultrasound of the abdomen | 0
moderate ascites | 0
features suggestive of acute kidney injury | 0
nasogastric tube inserted | 0
mildly bilious drainage of 500 mL | 0
random blood sugar of 250 mg/dL | 0
urine ketone body absent | 0
subcutaneous soluble insulin 0.1 U/kg | 0
variable-rate intravenous insulin infusion | 0
blood urea of 8.4 mmol/L | 0
serum creatinine of 2 mg/dL | 0
liver and clotting profiles normal | 0
hemodynamics stabilized | 0
emergency exploratory laparotomy | 0
midline laparotomy | 0
four-quadrant gross faecal peritonitis | 0
grossly distended small bowel | 0
hooked fishbone in the distal ileal mesenteric border | 0
sealed 5 mm perforation | 0
surrounding purulent exudate | 0
10 cm portion of the distal ileum resected | 0
proximal and distal ends taken out as end stomas | 0
peritoneal lavage | 0
pelvic drainage inserted | 0
vasopressor and inotropic requirements increased | 0
fourth vasopressor | 0
no urine output for 4 hours | 0
serum lactate rose to 20 mmol/L | 0
severe metabolic acidosis | 0
intravenous sodium bicarbonate infusion | 0
intravenous sedation and analgesia | 0
condition deteriorated | 2
cardiac arrest | 8
passed away | 8