Here is the extracted table of clinical events and timestamps:

62 years old | 0
male | 0
admitted to the hospital | 0
bilateral otalgia | -120
Glasgow Coma Scale (GCS) score 8 | -120
CRS with nasal polyposis | -672
functional endoscopic sinus surgery (FESS) with nasal polypectomy | -672
chronic obstructive pulmonary disease | 0
hypertension | 0
glaucoma | 0
right sided keratoconus treated with a previous corneal graft | 0
hypercholesterolaemia | 0
beclomethasone/formoterol inhaler | 0
salbutamol inhaler | 0
amlodipine | 0
simvastatin | 0
beclometasone dipropionate nasal spray | 0
tachypnoeic | 0
tachycardic | 0
pyrexial | 0
Glasgow Coma Scale (GCS) score 11 | 0
bilateral green purulent rhinorrhea | 0
bilateral proptosis | 0
right sided chemosis | 0
flexible nasendoscopy (FNE) | 0
raised CRP | 0
raised white cell count | 0
raised neutrophil count | 0
low lymphocyte count | 0
raised lactate | 0
pus aspirates collected from both nasal cavities | 0
Streptococcus pneumoniae isolated | 0
contrast-enhanced computed tomography (CT) of the head and sinuses | 1
opacification of the paranasal sinuses | 1
bony erosion of the lateral walls of both ethmoid sinuses | 1
soft tissue bulging into the right orbit | 1
bilateral proptosis | 1
no intracranial abnormality | 1
increasingly combative | 2
confused | 2
aversion to light | 2
lumbar puncture | 2
pale cloudy fluid | 2
extremely cellular specimen | 2
high protein | 2
low glucose | 2
Streptococcus pneumoniae isolated | 2
treatment for sepsis and presumed meningitis initiated | 2
intravenous ceftriaxone | 2
fluticasone nasal spray | 2
xylometazoline hydrochloride nasal spray | 2
regular saline nasal irrigation | 2
admitted to the critical care unit (CCU) | 2
intubated and ventilated | 12
extubated | 192
completed 10-day course of intravenous antibiotics | 240
discharged home | 312
follow-up with the critical care and ENT teams | 312
prescribed betamethasone nasal drops | 312
prescribed fluticasone nasal spray | 312
regular saline nasal irrigation | 312
recovered well | 744
returned to work full time | 744
vivid memories of stay on CCU | 744
no signs of post-traumatic stress disorder | 744
managed medically as an outpatient by the ENT team | 744
contrast-enhanced magnetic resonance imaging (MRI) of the brain, orbits and postnasal space | 1032
extensive bilateral ethmoid polyposis | 1032
hypertrophied inferior turbinates | 1032
left sided smooth dural enhancement | 1032
Aspergillus and Alternaria specific IgE levels within normal range | 1032