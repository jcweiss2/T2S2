62 years old | 0
    male | 0
    hypertension | -109248
    smoking | -109248
    AICD implant | -113688
    ventricular fibrillation arrest | -113688
    scheduled for AICD generator box change | 0
    general anesthesia | 0
    good ventricular function on echocardiogram | 0
    attempted removal of AICD generator box | 0
    break in insulation of AICD lead component | 0
    generator box removed | 0
    leads left in situ | 0
    plan for laser extraction | 0
    laser extraction of leads attempted | 48
    monitoring included standard and invasive arterial pressures | 48
    pericardial tamponade | 48
    linear tear in free wall of right ventricle | 48
    emergency surgery | 48
    extubated in ICU | 48
    central venous pressure 18-22 cm H2O | 48
    intermittent hypoxemic | 72
    PaO2 6.8-13.3 kPa | 72
    high inspired oxygen via CPAP mask | 72
    central venous pressure 13-15 cm H2O | 72
    clinical examination | 72
    chest X-ray showed left basal collapse | 72
    transthoracic echocardiogram inconclusive | 72
    normal hemodynamics | 72
    normal metabolic parameters | 72
    CTPA showed small right solitary pulmonary embolism | 72
    small left pleural effusion | 72
    atelectasis | 72
    started on heparin infusion | 72
    remained hypoxemic despite anticoagulation and oxygen | 72
    aneurysmal interatrial septum on CTPA review | 72
    transesophageal echocardiography performed | 72
    flail tricuspid valve | 72
    severe eccentric tricuspid regurgitation | 72
    large PFO with bidirectional shunt | 72
    dilatation of right atrial and right ventricular | 72
    mild RV dysfunction | 72
    preserved left ventricular function | 72
    extubated | 72
    discussed with cardiothoracic surgeon | 72
    consented for surgical closure of PFO | 72
    tricuspid valve replacement | 72
    next day | 96
    tricuspid valve replacement | 96
    bovine pericardial patch closure of PFO | 96
    good postoperative recovery | 96
    discharged home | 120
    follow-up at 6 weeks | 1344
    well seated functioning tricuspid prosthesis | 1344
    no residual shunt across interatrial septum | 1344
    
