52 years old | 0
    male | 0
    presented to the Emergency Department | 0
    septic shock | 0
    right sided abdominal pain | 0
    witnessed cardiac arrest | 0
    cardiopulmonary resuscitation | 0
    return of spontaneous circulation | 10
    physiologic resuscitation | 10
    broad spectrum intravenous antibiotics | 10
    cefuroxime | 10
    metronidazole | 10
    intubation | 10
    ventilation | 10
    computer tomography scan of the abdomen | 10
    moderate volume of free fluid | 10
    locules of gas within the pelvis | 10
    hollow viscus perforation | 10
    calcified structure within the appendix | 10
    foreign body causing perforated appendicitis | 10
    laparotomy | 20
    perforated appendicitis | 20
    four-quadrant purulent peritonitis | 20
    healthy caecum | 20
    appendicectomy | 20
    perforation in the mid-point | 20
    firm foreign body causing luminal obstruction | 20
    decaying tooth | 20
    metallic filling | 20
    washout with copious irrigation | 20
    abdomen closure | 20
    transfer to intensive care unit | 20
    passed away | 56
    multi-organ failure | 56
    sepsis | 56