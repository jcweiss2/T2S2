62 years old | 0
female | 0
presented to the neurologic clinic | 0
headache | -120
fever | -120
rigor | -120
received the second dose of COVID-19 Pfizer vaccine | -120
acute confessional state | 0
inability to talk | 0
known case of ceftriaxone allergy | 0
conscious | 0
disoriented | 0
did not obey commands | 0
no aphasia | 0
dysarthria could not be evaluated | 0
positive meningeal irritation signs | 0
pupils were isocor bilaterally | 0
light reaction was positive | 0
no evidence of ophthalmoplegia | 0
Babinski sign was negative | 0
not able to stand up and walk | 0
on wheelchair | 0
body temperature elevated | 0
temp 38C | 0
SPO2 98% | 0
Pulse rate 105 bpm | 0
Blood pressure 125/80 mmHg | 0
mild leukocytosis | 0
agranulocytosis | 0
C reactive protein elevated | 0
normal serum electrolyte | 0
normal renal and liver function tests | 0
random blood sugar 185mg/dl | 0
brain CT scan was normal | 0
brain MRI performed | 12
brain MRI showed normal brain parenchyma | 12
lumbar puncture was clear CSF macroscopically | 12
lymphocytic pleocytosis of 170 cells | 12
Protein 802mg/dl | 12
Glucose 71mg/dl | 12
Lactate 19.61mg/dl | 12
negative gram stain | 12
viral polymerase chain reaction for Herpes simplex virus negative | 12
meropenem IV 1 gm twice daily started | -12
Dexamethasone IV 4 mg once daily started | -12
Acyclovir vial IV 750 mg three times daily started | 0
responded well to the acyclovir | 48
became conscious again and oriented | 48
discharged from the hospital | 336
no focal neurological deficit | 336