weight loss | -8760
myalgias | -8760
fever | -8760
skin erythema | -8760
deterioration of renal function | -8760
new onset of diabetes mellitus Type II | -8760
hypertension | -8760
diagnosis of PAN | -4320
diagnosis of HBV infection | -4320
treatment with prednisolone | -4320
treatment with cyclophosphamide | -4320
stopped taking Tenofovir | -1440
admission | 0
acute abdomen | 0
septic shock | 0
free sub diaphragmatic air | 0
peritonitis | 0
three perforations of the small intestine | 0
segmental enterectomy with anastomosis | 0
mechanical ventilation | 0
circulatory support | 0
acute-on-chronic renal failure | 0
weaned off the ventilator | 72
haemodynamically stable | 72
treatment with tenofovir | 72
treatment with IV methylprednisolone | 72
abdominal drain catheter presented enteric content | 168
second explorative laparotomy | 168
two new perforations | 168
multiple areas of patchy necrosis | 168
plasma exchanges | 168
treatment with IV cyclophosphamide | 168
treatment with IV methylprednisolone | 168
treatment with IV prednisone | 168
third laparotomy | 240
three new necrotic lesions | 240
necrotic lesion on the left lobe of the liver | 240
fourth laparotomy | 336
segmental enterectomy with anastomosis | 336
cholecystectomy | 336
anastomotic leak | 336
gangrenous gallbladder | 336
death | 360
septic shock | 360
multiple organ failure | 360