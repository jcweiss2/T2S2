74 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
low-grade fever | -48 | 0 | Factual
dry cough | -48 | 0 | Factual
shortness of breath | -48 | 0 | Factual
elective right total knee replacement | -168 | -168 | Factual
post-operative course uneventful | -168 | -168 | Factual
pain in the right knee | -168 | 0 | Factual
redness in the right knee | -168 | 0 | Factual
swelling in the right knee | -168 | 0 | Factual
essential hypertension | 0 | 0 | Factual
obesity | 0 | 0 | Factual
myasthenia gravis in remission | 0 | 0 | Factual
osteoarthritis | 0 | 0 | Factual
body temperature 37.3°C | 0 | 0 | Factual
blood pressure 121/82 | 0 | 0 | Factual
pulse 87 beats per minute | 0 | 0 | Factual
respiratory rate 16 breaths per minute | 0 | 0 | Factual
oxygen saturation 87% | 0 | 0 | Factual
bilateral rhonchi with rales | 0 | 0 | Factual
patchy air space opacity in the right upper lobe | 0 | 0 | Factual
rapid nucleic acid amplification test for influenza A and B negative | 0 | 0 | Factual
nasopharyngeal swab specimen obtained | 0 | 0 | Factual
broad-spectrum antibiotics with cefepime and levofloxacin | 0 | 96 | Factual
supportive care with 2 L of supplemental oxygen | 0 | 96 | Factual
mild diarrhea | 72 | 72 | Factual
generalized weakness | 72 | 72 | Factual
fatigue | 72 | 72 | Factual
intravenous immunoglobulin | 72 | 120 | Factual
mild MG exacerbation | 72 | 120 | Factual
pending MG crises | 72 | 120 | Factual
arterial blood gases monitored | 0 | 384 | Factual
complete blood count monitored | 0 | 384 | Factual
basic metabolic profile studies monitored | 0 | 384 | Factual
mild absolute lymphopenia | 0 | 0 | Factual
anemia | 0 | 0 | Factual
pH 7.46 | 0 | 0 | Factual
pCO2 44.6 mmHg | 0 | 0 | Factual
pO2 94.7 mmHg | 0 | 0 | Factual
bicarbonate 31.4 mmol/L | 0 | 0 | Factual
creatinine kinase normal | 144 | 144 | Factual
lactic acid normal | 144 | 144 | Factual
lactate dehydrogenase elevated | 144 | 144 | Factual
ferritin elevated | 144 | 144 | Factual
interleukin-6 elevated | 144 | 144 | Factual
progressively increasing shortness of breath | 24 | 96 | Factual
oxygen requirements increased | 24 | 96 | Factual
nasopharyngeal swab results positive for SARS-CoV-2 | 96 | 96 | Factual
hydroxychloroquine | 96 | 240 | Factual
azithromycin | 96 | 240 | Factual
zinc sulfate | 96 | 240 | Factual
oral vitamin C | 96 | 240 | Factual
blood and sputum cultures did not grow any organisms | 96 | 96 | Factual
broad-spectrum antibiotics discontinued | 96 | 96 | Factual
shortness of breath worsened | 144 | 144 | Factual
oxygen requirements increased | 144 | 144 | Factual
drowsy | 144 | 144 | Factual
moderate distress | 144 | 144 | Factual
unable to protect the airways | 144 | 144 | Factual
blood pressure 78/56 mmHg | 144 | 144 | Factual
heart rate 112 beats per minute | 144 | 144 | Factual
temperature 38°C | 144 | 144 | Factual
respiratory rate 28 breaths per minute | 144 | 144 | Factual
bilateral alveolar infiltrates | 144 | 144 | Factual
interstitial edema | 144 | 144 | Factual
intubated | 144 | 144 | Factual
mechanical ventilation | 144 | 240 | Factual
norepinephrine | 144 | 192 | Factual
colchicine | 144 | 240 | Factual
high-dose vitamin C | 168 | 384 | Factual
clinical condition improved | 192 | 384 | Factual
norepinephrine support stopped | 192 | 192 | Factual
CXR showed significant improvement | 240 | 240 | Factual
spontaneous breathing trial | 240 | 240 | Factual
extubated | 240 | 240 | Factual
breathing status continued to improve | 240 | 384 | Factual
oxygen saturation 92% | 384 | 384 | Factual
CXR revealed almost complete resolution | 384 | 384 | Factual
discharged from the hospital | 384 | 384 | Factual
inpatient physical and occupational rehabilitation | 240 | 384 | Factual
quarantine | 384 | 398 | Factual