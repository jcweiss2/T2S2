40 years old | 0
male | 0
admitted to the hospital | 0
fever | -24
diarrhea | -24
dyspnea | -24
confusion | -24
shock | -24
bleeding spots on the chest and abdomen | -24
florid spots on the lower limbs | -24
oxygen saturation of 60% | -24
hypertension | -672
fatty liver | -672
HFRS | -24
septic shock | 0
decompensated metabolic acidosis | 0
AKI | 0
multiple organ failure | 0
ventilator-assisted ventilation | 0
fluid replacement | 0
norepinephrine | 0
CRRT | 0
sedation and analgesia | 0
plasma and platelet transfusions | 0
nasal cavity filled with an expanded sponge | 24
left nasal alar became purple and swollen | 48
massive nasal necrotic lesions | 72
Rhizopus oryzae complex | 72
Aspergillus fumigatus | 72
pulmonary aspergillosis | 72
rhinomucormycosis | 72
caspofungin | 72
voriconazole | 72
local treatment with amphotericin B | 72
nasal cavity rinsed with saline | 72
nasal cavity filled with sterile dressing containing amphotericin B | 72
nasal cavity filled with sterile dressing containing sodium bicarbonate | 78
left nasal scab fell off | 288
large tissue defect remained | 288
computed tomography revealed no orbitocerebral involvement | 288
bronchoalveolar lavage fluid culture revealed no fungal growth | 264
lung imaging findings returned to normal | 264
urine output recovered | 264
renal function recovered | 264
weaning from the ventilator | 264
discontinuation of caspofungin | 312
discontinuation of voriconazole | 336
recovered | 672
discharged | 672