77 years old | 0
    male | 0
    presented to the emergency department | 0
    syncope | 0
    hypertension | 0
    hyperlipidemia | 0
    uncontrolled diabetes mellitus type two | 0
    recurrent diabetic foot ulcers | 0
    osteomyelitis | 0
    peripheral vascular disease | 0
    coronary artery disease | 0
    five-vessel coronary artery bypass grafting | -149520
    pacemaker/defibrillator implantation | -149520
    systolic heart failure | 0
    ischemic cardiomyopathy | 0
    dizziness | 0
    dyspnea | 0
    fevers 101°F to 102°F | -72
    elevated blood glucose readings | -72
    lethargy | -72
    rigors | -72
    chills | -72
    malaise | -72
    unwitnessed time | 0
    elevated troponin levels | 0
    NT-proBNP 24000 pg/mL | 0
    leukocyte count 16000/uL | 0
    wide complex tachycardia | 0
    tachypneic | 0
    hypertensive 157/136 mm Hg | 0
    cardioversion | 0
    right bundle branch block | 0
    left anterior fascicular block | 0
    QTc 445 msec | 0
    normal axis | 0
    Levophed initiated | 0
    empiric antibiotic therapy | 0
    vancomycin | 0
    piperacillin/tazobactam | 0
    blood cultures obtained | 0
    agonal breathing | 0
    intubated | 0
    transferred to ICU | 0
    hypotensive | 0
    dopamine started | 0
    cardiac catheterization | 0
    cardiogenic shock considered | 0
    septic shock considered | 0
    severe native vessel disease | 0
    PCI | 0
    stent deployment | 0
    pseudoaneurysm identified | 0
    intra-aortic balloon pump inserted | 0
    sustained ventricular tachycardia | 0
    lidocaine infusion | 0
    amiodarone infusion | 0
    defibrillator reprogrammed | 0
    blood cultures positive for MSSA | 48
    elevated liver function tests | 48
    elevated creatinine | 48
    IABP removed | 48
    gram-positive bacteremia | 48
    lactic acidosis resolved | 48
    persistent fevers | 48
    worsening leukocytosis | 48
    IV linezolid | 48
    extubated | 72
    BiPAP | 72
    volume overloaded | 72
    monitored diuresis | 72
    oral amiodarone | 72
    ventricular tachycardia episodes | 72
    amiodarone bolus infusions | 72
    amiodarone maintenance infusions reinstated | 72
    Infectious Disease Service consulted | 72
    transitioned to cefazolin | 72
    rifampin | 72
    leukocytosis resolved | 72
    defervesce | 72
    ventricular tachycardia runs | 72
    AICD discharges | 72
    oxygen via nasal cannula | 72
    Precedex initiated | 72
    disorientation | 72
    repeat blood cultures no growth | 72
    pacemaker interrogation | 72
    lidocaine infusion resumed | 72
    VT zone 140–150 seconds | 72
    anti-tachycardia pacing identified | 72
    mexiletine triggered V-tach | 72
    pacemaker EOL imminent | 72
    TEE recommended | 72
    transcutaneous pacer pads placed | 72
    Palliative care considered | 72
    Diuril started | 72
    Precedex discontinued | 72
    lidocaine transitioned to amiodarone | 72
    seven VT runs | 96
    mexiletine started | 96
    amiodarone infusion continued | 96
    TTE obtained | 96
    dilated LV | 96
    segmental wall motion abnormalities | 96
    LVEF 35% | 96
    moderate concentric LV hypertrophy | 96
    left atrial enlargement | 96
    pacemaker leads in right heart | 96
    mitral annular calcification | 96
    mild mitral regurgitation | 96
    TEE performed | 96
    fibrinous lead vegetations | 96
    right atrial abscess | 96
    moderate LV dysfunction | 96
    moderate mitral regurgitation | 96
    moderate tricuspid regurgitation | 96
    tertiary care transfer proposed | 96
    Gentamicin initiated | 96
    transfer declined | 96
    no VT episodes | 96
    lidocaine discontinued | 96
    amiodarone discontinued | 96
    mexiletine continued | 96
    oral amiodarone continued | 96
    defibrillator inhibited | 96
    pacemaker function intact | 96
    IV antibiotics for 15 days | 96
    rifampin 300 mg daily | 96
    Keflex 750 mg twice daily | 96
    discharged home with hospice | 96
    outpatient follow-up | 96
    negative blood cultures | 96
    <|eot_id|>
    