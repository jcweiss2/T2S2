54 years old | 0
    woman | 0
    height 170 cm | 0
    weight 68 kg | 0
    no drug allergy | 0
    heavy smoker | 0
    no coronary risk factors | 0
    bilateral cataract extraction | -17280
    local anesthesia | -17280
    breast augmentation | -17280
    abdominoplasty | -17280
    general anesthesia | -17280
    screening gastroscopy | 0
    colonoscopy under sedation | 0
    occult anemia | 0
    no premedication | 0
    anticholinergic medications not used | 0
    standard parameter monitoring | 0
    noninvasive blood pressure monitoring | 0
    SPO2 monitoring | 0
    EKG monitoring | 0
    oxygen supplementation | 0
    nasal cannula 4 L/min | 0
    baseline vital signs normal | 0
    NIBP 112/65 | 0
    heart rate 72 beats/min | 0
    respiratory rate 12 per minute | 0
    SPO2 100% | 0
    sedated with meperidine 50 mg | 0
    sedated with midazolam 2 mg | 0
    sedated with propofol 40 mg | 0
    gastroscopy started | 0
    bradycardia | 600
    SPO2 97% | 600
    asystole | 600
    premature ventricular contraction | 600
    bizarre QRS wave | 600
    undetectable blood pressure | 600
    no skin rash | 600
    received xylocaine 60 mg | 600
    received atropine 2 mg | 600
    received epinephrine 0.01 mg | 600
    received hydrocortisone 250 mg | 600
    face mask ventilation 100% | 600
    sinus tachycardia | 600
    heart rate 112 beats/min | 600
    NIBP 70/42 mmHg | 600
    spontaneous breathing | 600
    no dyspnea | 600
    regained consciousness | 600
    acute chest pain | 600
    pulmonary edema | 600
    dyspnea | 600
    hypoxia SPO2 60% | 600
    procedure aborted | 600
    transferred to intensive care unit | 600
    EKG not indicative | 600
    chest X-ray diffuse bilateral infiltrations | 600
    transthoracic echocardiography | 600
    global hypokinesia | 600
    ejection fraction 20-29% | 600
    respiratory acidosis | 600
    PH 7.31 | 600
    PO2 43.5 | 600
    PCO2 51.5 | 600
    SBE 0.5 | 600
    HCO3 23.2 | 600
    acute LV dysfunction | 600
    pulmonary edema confirmed | 600
    Lasix 80 mg intravenous | 600
    dobutamine 15 mcg/kg/min | 600
    clinical improvement | 720
    saturation 95% | 720
    BiPAP ventilation | 720
    complete improvement | 1440
    weaning dobutamine | 1440
    troponin 0.08 | 0
    troponin 0.54 | 432
    troponin 0.58 | 1080
    serial EKGs no evolving changes | 1440
    coronary angiography | 17280
    no significant coronary stenosis | 17280
    fully recovered | 17280
    no cardiac symptoms | 17280
    weaned from BiPAP | 17280
    discontinued inotropic support | 17280
    echocardiography improved LV function | 17280
    no regional wall motion abnormality | 17280
    EF 68% | 17280
    chest x-ray no pulmonary edema | 17280
    discharged | 17280
    carvedilol | 17280
    rabeprazole sodium | 17280
    doing well at three months follow-up | 17280
    