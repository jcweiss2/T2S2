35 years old | 0  
    gravida 3 para 1–0-1–1 | 0  
    referred to maternal-fetal medicine office | 0  
    diagnosis of early midtrimester oligohydramnios | 0  
    oligohydramnios incidentally found | 0  
    routine anatomical survey ultrasound examination at 18 weeks of gestation | -432  
    evaluated for preterm prelabor rupture of membranes | 0  
    pooling of amniotic fluid in posterior vaginal fornix | 0  
    arborization ferning testing | 0  
    nitrazine testing | 0  
    initial evaluation negative | 0  
    two subsequent assessments showed no evidence of rupture of amniotic membranes | 0  
    offered intra-amniotic dye infusion testing | 0  
    declined intra-amniotic dye infusion testing | 0  
    ultrasound at 20 6/7 weeks of gestation | -168  
    single live fetus | -168  
    amniotic fluid index of 2.8 cm | -168  
    ultrasound evidence of membrane separation | -168  
    possible membrane rupture distal to the cervical opening | -168  
    fetal kidneys seen | -168  
    fetal bladder seen | -168  
    gestational diabetes | 0  
    history of loop electrical excision procedure | 0  
    herpes simplex type 2 | 0  
    maternal obesity | 0  
    prepregnancy BMI 34 kg/m2 | 0  
    episode of domestic violence | 0  
    early genetic screening with cell free fetal DNA | 0  
    appropriate fetal fraction | 0  
    sex chromosomes XY | 0  
    low risk for trisomy 13 | 0  
    low risk for trisomy 18 | 0  
    low risk for trisomy 21 | 0  
    second trimester maternal serum α-fetoprotein 2.16 MoM | 0  
    prenatal counseling with neonatology | 0  
    prenatal counseling with maternal-fetal medicine | 0  
    expressed wishes for full neonatal resuscitation at 22 weeks | 0  
    understanding of prognosis | 0  
    offered amnioinfusion | 0  
    offered intra-amniotic dye instillation testing | 0  
    proceeded with amnioinfusion | 0  
    proceeded with intra-amniotic dye installation at 21 6/7 weeks of gestation | -168  
    ultrasound guidance | -168  
    22-gauge needle inserted into intra-amniotic cavity | -168  
    15 mL clear yellow fluid removed | -168  
    genetic testing | -168  
    infection testing | -168  
    40 mL warmed 0.9% sodium chloride solution infused | -168  
    1000 mg/L oxacillin infused | -168  
    5 mL indigo carmine added | -168  
    intra-amniotic dye instillation test | -168  
    400 mL warmed 0.9% sodium chloride solution infused | -168  
    patient ambulated for 30 minutes | -168  
    tampon testing confirmed rupture of fetal membranes | -168  
    admitted to the hospital | 0  
    latency antibiotics | 0  
    serial intra-amniotic infusions | 0  
    acyclovir prophylaxis started | 0  
    clinical exam confirmed no active herpes lesions | 0  
    completed 7-day course of latency antibiotics | 168  
    ampicillin | 168  
    azithromycin | 168  
    betamethasone administered at 23 weeks of gestation | 168  
    second amnioinfusion at 22 6/7 weeks of gestation | 24  
    800 mL warmed 0.9% sodium chloride solution infused | 24  
    1000 mg/L oxacillin infused | 24  
    normal maximum vertical pocket obtained | 24  
    plan for serial intra-amniotic infusions until 26 weeks of gestation | 24  
    denied continued leakage of fluid at 23 6/7 weeks | 168  
    MVP normal at 23 6/7 weeks | 168  
    suspected amnion resealed | 168  
    decision to cease further intra-amniotic infusions | 168  
    amniotic fluid testing returned no evidence of intra-amniotic infection | 168  
    genetic testing with karyotype confirmed no genetic abnormalities | 168  
    genetic testing with microarray confirmed no genetic abnormalities | 168  
    developed gestational hypertension at 27 weeks of gestation | 264  
    no clinical evidence for preeclampsia | 264  
    no laboratory evidence for preeclampsia | 264  
    expectantly managed in the hospital | 264  
    fetal status remained reassuring | 264  
    appropriate fetal growth on serial ultrasounds | 264  
    MVP remained normal | 264  
    second course of betamethasone at 33 0/7 weeks | 648  
    external cephalic version performed at 34 weeks | 768  
    breech presentation | 768  
    successful induction of labor at 34 2/7 weeks | 776  
    given penicillin in labor | 776  
    group B streptococcus prophylaxis | 776  
    delivered vigorous male infant | 776  
    birth weight 2160 g | 776  
    Apgar score 9 at 1 minute | 776  
    Apgar score 9 at 5 minutes | 776  
    placenta weighed 390 g | 776  
    evidence of moderate acute inflammation at the chorion | 776  
    no evidence of inflammation elsewhere on the amnion | 776  
    no evidence of inflammation on umbilical cord | 776  
    newborn's initial white blood cell count 11.7 × 1000 μL | 776  
    ampicillin given | 776  
    gentamycin given | 776  
    negative blood cultures | 776  
    neonatal intensive care protocol | 776  
    newborn stayed in hospital for 9 days | 776  
    no immediate complications | 776  
    
