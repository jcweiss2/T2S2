51 years old | 0
male | 0
admitted to the hospital | 0
abdominal pain | -72
vomiting | -72
intestinal obstruction | -72
ate persimmon | -168
previous abdominal operation | -7200
small bowel perforation | -7200
leukocytosis | 0
hemoglobin concentration 18.3 g/d | 0
C-reactive protein 0.07 mg/dL | 0
body temperature 36.5 | 0
abdominal distension | 0
mild tenderness over the epigastric area | 0
HIV antibody negative | 0
mechanical obstruction in the ileum | 0
bezoar | 0
mild splenomegaly | 0
decrease of leukocytosis | 96
increase for C-reactive protein | 96
bezoar removal operation | 120
small bowel dilatation | 120
no signs of small bowel ischemia | 120
bezoar extracted | 120
decompression of the dilated bowel | 120
fever | 48
postoperative atelectasis | 48
pass flatus | 120
started on a progressive diet | 120
dyspnea | 168
diffuse ground glass opacity | 168
ARDS | 168
mechanical ventilation | 168
blood cultures collected | 96
yeast | 96
empiric therapy of fluconazole | 96
C. famata | 120
C. parapsilosis | 144
fever persisted | 144
leukocytosis persisted | 144
antifungal treatment for tinea pedis | -8760
changed to amphotericin B | 144
methylprednisolone | 144
stool culture collected | 288
Candida glabrata | 288
changed to caspofugin | 432
nephrotoxicity | 432
afebrile | 504
clinical improvement | 504
blood cultures sterile | 504
discharged | 888