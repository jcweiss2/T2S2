54 years old | 0
female | 0
admitted to the hospital | 0
acute abdomen | 0
possible diagnosis intestinal obstruction | 0
central line insertion | 0
USG guidance | 0
right subclavian vein | 0
irritation near right ear | 0
guidewire inserted | 0
right IJV visualized | 0
hyperechoic object seen | 0
guidewire confirmed | 0
guidewire taken out | 0
reattempts done | 0
catheter inserted | 0
guidewire removed | 0
venous aspiration | 0
saline flushed | 0
turbulence in right atrium | 0
catheter tip in superior vena cava | 0 
central venous catheterization | -24
malpositioning | -24
blind procedures | -24
anatomical landmarks | -24
ultrasound guidance | -24
complications | -24
catheter malposition | -24
internal jugular vein | -24
subclavian vein | -24
catheterization | -24
ASA practice guidelines | -120
USG examination | -120
central line malposition | -120
X-ray confirmation | -120
guidewire malposition | -120
catheter malposition | -120
thoracic cavity | -120
mediastinum | -120
electrocardiographic guidance | -120
p-wave size | -120
pericardial reflection | -120
arterial placement | -120
venous placement | -120
real-time acoustic shadow | -120
USG for CVC insertion | -120
anatomy of vessel | -120
thrombus within vessel | -120
needle piercing vessel | -120
guidewire going within vessel | -120
guidewire in other vessels | -120
CVC going in vessel | -120
turbulence in right atrium | -120
saline in distal port | -120
pleural damage | -120
hematoma | -120
hemothorax | -120
catheter pierces wall | -120
mediastinal space | -120
pleural cavity | -120
color of blood | -120
pulsating blood flow | -120
backflow of blood | -120 
discharged | 24