36-year-old man | 0
transferred to ICU | 0
intubated | 0
ventilated | 0
worsening type 1 respiratory failure | 0
COVID-19 diagnosis | 0
1-week history of persistent fever | -168
dry cough | -168
3 days of coryzal symptoms | -72
radiographic features of COVID-19 | 0
SARS-CoV-2 PCR swab positive | 48
raised CRP (320 mg/L) | 0
raised ferritin (2020 µg/L) | 0
raised D-dimer (2262 ng/mL) | 0
lymphocytopaenia (0.7×10^9/L) | 0
concurrent neutrophilia | 0
normal HbA1c | 0
normal lipid profile | 0
serum vitamin D insufficiency (34 nmol/L) | 336
nutritional assessment | 0
initial estimated weight (75 kg) | 0
initial estimated height (1.75 m) | 0
BMI 24.5 kg/m² | 0
corrected weight (80-85 kg) | 0
nasogastric tube placement | 0
enteral tube feeding | 0
Penn State protocol (1631 kcal/day) | 0
ESPEN recommendations (1125-1500 kcal/day) | 0
protein requirements (906-112.5 g/day) | 0
propofol use (≥350 kcal/day) | 0
sepsis | 0
prolonged ICU admission (52 days) | 0
ventilatory support (50 days) | 0
poor lung compliance | 0
brittle ventilation | 0
oxygenation issues | 0
protracted ventilator wean | 0
tracheostomy wean | 0
pulmonary embolism | 168
CT pulmonary angiogram | 168
COVID-19 pneumonitis | 0
fibrotic lung changes | 0
multiple antibiotic therapies | 0
prone positioning (196 hours) | 0
low volume feeding during proning | 0
nasogastric tube feeding interruptions | 0
feed composition adjustments | 0
high energy/protein feeds | 0
concentrated feed (2 kcal/mL) | 0
energy deficit | 0
protein deficit | 0
fasting for investigations | 0
tube removal due to agitation | 0
delays in feed provision | 0
mild/moderate gastrointestinal symptoms | 0
loose bowels | 0
constipation | 0
abdominal distension | 0
laxatives/enemas | 0
minimal gastric aspirates | 0
severe weight loss (19 kg) | 0
deconditioning | 0
reduced subcutaneous fat | 0
muscle wasting | 0
reduced appetite | 0
poor oral intake | 0
modified texture diet | 0
enteral tube feeding continuation | 0
oral nutritional supplements | 0
tube removal request | 0
hospital stay post ICU (10 days) | 0
physiotherapy | 0
speech and language therapy | 0
dietetic support | 0
fortified diets | 0
virtual clinic | 0
malnutrition | 0
cachexia | 0
sarcopenia | 0
metabolic dysregulation | 0
hypermetabolic state | 0
vitamin D deficiency | 336
hypocaloric feeding | 0
hypocaloric feeding adjustment | 0
underfeeding | 0
parenteral nutrition consideration | 0
micronutrient supplementation | 0
Pabrinex supplementation | 0
vitamin D replacement advice | 0
logistical challenges | 0
remote assessments | 0
PPE preservation | 0
staff redeployment | 0
anthropometric data issues | 0
feed delivery protocols | 0
nursing staff shortages | 0
nutritional interventions | 0
patient-reported weight loss | 0
appetite improvement | 0
sleep improvement | 0
protein requirements (90-112.5 g/day) | 0
