61 years old | 0
female | 0
end-stage renal disease | 0
adult polycystic kidney disease | 0
living-related kidney transplant | 0
fever | -120
diarrhea | -120
nausea | -120
attended a funeral | -240
denied cough | 0
denied shortness of breath | 0
denied chest pain | 0
denied abdominal pain | 0
denied vomiting | 0
denied fatigue | 0
denied myalgia | 0
denied headache | 0
hypertension | 0
gout | 0
histoplasmosis | 0
tacrolimus | 0
mycophenolate mofetil (MMF) | 0
prednisone | 0
itraconazole | 0
allopurinol | 0
labetalol | 0
hydralazine | 0
febrile | 0
pulse rate 87 beats per minute | 0
blood pressure 151/85 mm Hg | 0
respiratory rate 24 breaths per minute | 0
oxygen saturation 92% to 97% | 0
respiratory distress | 0
decreased breath sounds on left chest | 0
unremarkable physical exam | 0
hemoglobin 13.3 g/dL | 0
WBC 4.7 103/µL | 0
lymphocytes 24.4% | 0
neutrophils 67% | 0
sodium 135 mmol/L | 0
potassium 4.1 mmol/L | 0
bicarbonate 21 mEq | 0
BUN 13 mg/dL | 0
creatinine 1.3 mg/dL | 0
magnesium 1.6 mg/dL | 0
creatine kinase 83 U/L | 0
ferritin 734.4 ng/mL | 0
CRP 5.3 mg/L | 0
tacrolimus trough level 7 µg/L | 0
COVID-19 positive | 0
chest X-ray mid to lower lung infiltrates | 0
CT chest ground glass opacities | 0
ceftriaxone | 0
azithromycin | 0
intravenous fluids | 0
antipyretics | 0
MMF held | 0
tacrolimus continued | 0
prednisone continued | 0
oxygen 2-3 L | 0
fever resolved | 48
discharged | 120
MMF restarted | 120
doing well after discharge | 264
