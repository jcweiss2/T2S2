54 years old | 0
    male | 0
    admitted to the emergency department | 0
    progressive pain (right lower extremity) | -168
    swelling (right lower extremity) | -168
    permanent redness (right lower extremity) | -168
    petechial haemorrhage (right lower extremity) | -168
    hit leg | -168
    septic shock | 0
    tachycardia | 0
    dyspnoea | 0
    arterial hypotension | 0
    blood pressure 81/42 mmHg | 0
    heart rate 128 bpm | 0
    temperature 39.2°C | 0
    respiratory rate 38 breaths per minute | 0
    SpO2 96% on 6 L/min oxygen | 0
    paO2 114 mmHg | 0
    moderately impaired left ventricular ejection fraction (40%) | 0
    well-functioning heart valves | 0
    no endocarditis | 0
    no pericardial effusion | 0
    elevated white blood cell count (20.23 × 109/L) | 0
    elevated C-reactive protein (3362 nmol/L) | 0
    elevated procalcitonin (43.5 µg/L) | 0
    elevated lactate (8.8 mmol/L) | 0
    platelet count 160 × 109/L | 0
    elevated total bilirubin (42.75 µmol/L) | 0
    elevated aspartate aminotransferase (950 nmol/s*L) | 0
    elevated alanine aminotransferase (850 nmol/s*L) | 0
    elevated blood glucose (20.8 mmol/L) | 0
    suspected necrotising fasciitis | 0
    severe sepsis with multiple organ failure | 0
    liver failure | 0
    renal failure | 0
    elevated creatinine (382 µmol/L) | 0
    elevated urea (18.8 mmol/L) | 0
    absent urine output | 0
    elevated myoglobin (125 nmol/L) | 0
    continuous veno;venous haemodialysis | 0
    calcium-citrate anticoagulation | 0
    somnolent | 0
    Richmond Agitation and Sedation Scale score -2 | 0
    intubated | 2
    acidosis | 2
    paO2 179 mmHg | 2
    FiO2 70% | 2
    Horowitz Index 256 mmHg | 2
    mild ARDS | 2
    wound debridement | 6
    excision of the fascia | 6
    microbiological biopsy sampling | 6
    haemodynamic deterioration | 24
    excessive volume therapy (4 L crystalloids) | 24
    catecholamine therapy (1.2 mg/h norepinephrine) | 24
    whole-body CT scan | 24
    subcutaneous fluid retention (right thigh) | 24
    small air bubbles along the fascia | 24
    transfemoral amputation | 24
    increased catecholamine requirement (1.6 mg/h norepinephrine) | 24
    temperature 39.1°C | 24
    leukocytes 25.8 × 109/L | 24
    CRP 4067 nmol/L | 24
    PCT 60.40 µg/L | 24
    IL-6 2532 U/L | 24
    LBP 91 U/L | 24
    HLA-DR 27.3% | 24
    amputation | 24
    stump revision | 96
    wound closure | 216
    severe necrotising florid inflammation | 216
    empiric antimicrobial therapy (piperacillin/tazobactam) | 0
    clindamycin administration | 0
    Streptococcus pyogenes detected (wound swab and blood cultures) | 24
    antibiotic therapy changed to penicillin G | 24
    immunoglobulin therapy (Pentaglobin) | 48
    gradual weaning from mechanical ventilation | 168
    extubated | 168
    temperature 36.8°C | 168
    leukocytes 15.8 × 109/L | 168
    CRP 694 nmol/L | 168
    PCT 9.51 µg/L | 168
    IL-6 32.5 U/L | 168
    LBP 25.3 U/L | 168
    HLA-DR 61.2% | 168
    catecholamines reduced | 168
    catecholamines discontinued | 168
    transferred to normal ward | 384
    prosthesis fitting | 384
    discharged to rehabilitation | 624
    discharged home | 1440
    <|eot_id|>
    