40 years old|0
    businessman|0
    admitted to intensive care unit (ICU)|0
    fever|-480
    chills|-480
    vomiting|-96
    seizures|-96
    decreased urine output|-96
    shock|0
    intubated|0
    mechanical ventilation|0
    icteric|0
    acute kidney injury|0
    dengue antigen non-structural (NS1) positive|0
    malaria negative|0
    enteric fever negative|0
    hematocrit 35.2%|0
    total leukocyte count 9600/mm³|0
    coagulopathy|0
    endotracheal bleed|0
    anuria|0
    progressively deteriorating liver function|0
    ongoing septic shock|0
    lung protective mechanical ventilation|0
    slow low efficiency daily dialysis|0
    vasopressors (noradrenaline)|0
    broad spectrum antibiotics (ceftriaxone)|0
    artesunate|0
    dengue IgM positive|0
    Leptospira IgM positive|0
    HEV IgM positive|0
    malaria negative|0
    enteric fever negative|0
    hepatitis A negative|0
    hepatitis B negative|0
    hepatitis C negative|0
    human immunodeficiency virus negative|0
    serum procalcitonin rising trends|0
    blood culture no growth|0
    endotracheal culture no growth|0
    urine culture no growth|0
    died|144
    no renal biopsy|0
    no liver biopsy|0
    fever persisted|0
    thrombocytopenia|0
    liver dysfunction|0
    renal dysfunction|0
    dengue antigen positivity|0
    hypovolemic shock|0
    septic shock|0
    endothelial dysfunction|0
    coagulopathy|0
    thrombocytopenia|0
    cerebral edema|0
    disseminated intravascular coagulation|0
    triple co-infection|0
    hemodynamically unstable|0
    