67 years old | 0
female | 0
admitted to the hospital | 0
past medical history of sternoclavicular septic arthritis | -672
recurrent bacteremia | -672
previous bacterial endocarditis | -672
end-stage renal disease | -672
on hemodialysis | -672
persistent cough | 0
dysphagia to solid foods | 0
chest radiograph | 0
computed tomography angiogram | 0
large true aneurysm of the proximal right subclavian artery | 0
cardiac clearance | 0
consent for open repair | 0
operative exposure | 12
partial median sternotomy | 12
right infraclavicular extension | 12
partial right claviculectomy | 12
clavicle reconstruction deferred | 12
dissection of aneurysm | 12
highly inflamed and fibrous mediastinal/periclavicular tissue | 12
right internal jugular vein ligated and divided | 12
multiple enlarged collateral veins ligated and divided | 12
excision of aneurysm | 12
right phrenic nerve identified and protected | 12
right vertebral artery identified | 12
innominate-to-right subclavian arterial bypass | 12
reimplantation of the right common carotid artery | 12
Rifampin-soaked Dacron graft used | 12
specimens sent for pathologic analysis | 12
postoperative moderate head and neck edema | 12
endotracheal ventilation | 12
head elevation | 12
extubated on postoperative day 7 | 168
transferred out of intensive care unit on postoperative day 9 | 216
discharged to rehabilitation facility on postoperative day 20 | 480
final pathology demonstrated chronic osteomyelitis of clavicular head | 480
right subclavian artery specimen revealed partial wall necrosis and organized thrombus | 480
microbiologic analysis confirmed methicillin-sensitive Staphylococcus aureus | 480
6-week course of intravenous cefazolin | 480
converted to cephalexin for life-long suppressive therapy | 480
free from recurrent bacteremia | 480
no residual head or neck edema | 480
minimal change in upper extremity functioning | 480
denies any vasculogenic symptoms | 480