39 years old | 0
African-American male | 0
admitted to the hospital | 0
weakness | -72
decreased appetite | -72
suspected sepsis | 0
vancomycin | 0
meropenem | 0
Candida glabrata in urine cultures | 0
chronic indwelling Foley catheter | -672
urinary retention | -672
transferred to general medical floor | 120
osteomyelitis | 240
Stage IV sacral decubitus ulcer | 240
exposed bone | 240
negative blood cultures | 240
Candida albicans in urine cultures | 672
failure to thrive | 48
body mass index 14.7 kg/m2 | 48
percutaneous endoscopic gastrostomy tube placement | 288
elevated alkaline phosphatase | 0
elevated aspartate aminotransferase | 0
elevated alanine aminotransferase | 0
brittle diabetes | 0
hypoglycemic episodes | 0
insulin glargine | 0
50% dextrose boluses | 0
NPH insulin | 1224
glycemic goals | 0
leukocytosis | 816
abdominal computed tomography scan | 864
right-sided pyelonephritis | 864
left-sided hydronephrosis | 864
left-sided hydroureter | 864
micafungin | 900
urology consultation | 888
repeat abdominal computed tomography scan | 912
pyelonephritis in both kidneys | 912
filling defects | 912
mild debris along the bladder base | 912
fungus balls/mycetomas | 912
urine cultures with C. glabrata and C. albicans | 960
blood cultures with C. glabrata | 960
switched to high-dose fluconazole | 960
nephrostomy tube placement | 1080
systemic antifungal therapy | 1080
renal ultrasound | 1296
fungal balls | 1296
renal impairment | 1296
estimated glomerular filtration rate 10-30 mL/min/1.73 m2 | 1296
intermittent hemodialysis | 1344
placement of right nephrostomy tube | 1416
discontinued fluconazole | 1416
initiated systemic AmBd | 1416
LFTs significantly worsened | 1488
Naranjo adverse drug reaction probability scale score of 5 | 1488
LFTs returned to near baseline | 1512
code status changed to do not resuscitate | 1512
stopped 5% dextrose infusion | 1584
expired | 1584