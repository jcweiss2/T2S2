70 years old | 0
female | 0
admitted to the hospital | 0
lower abdominal pain | -24
fever | -24
nausea | -24
vomiting | -24
diaphoresis | -24
right ovarian cyst | -24
acute appendicitis | -24
congestive heart failure | -8760
atrial fibrillation | -8760
hypertension | -8760
right coronary artery 90% stenosis | -8760
digoxin | -8760
dilatrend | -8760
nitrate | -8760
telmisartan | -8760
thiazide | -8760
electrocardiogram showed AF | 0
left ventricular hypertrophy | 0
cardiomegaly | 0
pleural effusion | 0
ejection fraction 55% | 0
left atrial enlargement | 0
right atrial enlargement | 0
eccentric hypertrophy | 0
decreased mobility of the inferior wall of the left ventricle | 0
moderate aortic valve insufficiency | 0
aortic valve sclerosis | 0
mild aortic stenosis | 0
severe posterior mitral valve leaflet calcification | 0
mitral valve width 1.92 cm2 | 0
chronic cerebral infarction | -8760
dysarthria | -8760
dehydration | 0
prerenal azotemia | 0
serum creatinine 1.7 mg/dl | 0
fluid therapy | 0
serum creatinine 1.3 mg/dl | 12
glycopyrrolate 0.2 mg IM | -0.5
premedicated | -0.5
blood pressure 130/50 mmHg | 0
ventricular response 90-100 times/min | 0
arterial oxygen saturation 97% | 0
right radial artery cannulation | 0
induction of anesthesia | 0
lidocaine 2% | 0
propofol | 0
remifentanil | 0
rocuronium 40 mg | 0
endotracheal intubation | 0
central venous catheterization | 0
ventilation with 100% O2 | 0
systolic BP 130-150 mmHg | 0
diastolic BP 40-60 mmHg | 0
ventricular response 100-110 times/min | 0
central venous pressure 8-9 mmHg | 0
effect site concentration 2.5-3.0 µg/ml propofol | 0
effect site concentration 2.0 ng/ml remifentanil | 0
lower abdomen laparotomy | 0
small bowel infarction | 0
transesophageal echocardiography | 0
thrombus in left atrial appendage | 0
segmental resection and intestinal anastomosis | 0
anticoagulation therapy | 72
low molecular weight heparin | 72
oral warfarin | 120
cardioversion | 672
normal sinus rhythm | 672
discharged | 720