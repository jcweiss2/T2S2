19 years old|0
male|0
presented to the Emergency Department|-120
fever|-120
arthralgia|-120
myalgia|-120
headache|-120
intermittent productive cough|-120
yellowish sputum|-120
chest heaviness|-120
dyspnea at rest|-120
diarrhea|-120
reduced oral intake|-120
denied history of travelling|0
denied recent jungle activities|0
stayed in the military base camp|0
no past medical illness|0
no previous hospitalization|0
never sought medical treatment|0
conscious|0
dehydrated|0
cold peripheries|0
febrile|0
temperature of 38.5 °C|0
hypotensive|0
blood pressure of 81/53 mmHg|0
tachycardic|0
heart rate of 146 beats per minute|0
tachypnoeic|0
respiratory rate of 30 breaths per minute|0
oxygen saturation of 75–80%|0
15L high flow mask|0
coarse crepitation over both lower zone of lungs|0
tenderness at epigastric region|0
palpable liver around 5 cm below costal margin|0
no cervical lymph nodes palpable|0
no inguinal lymph nodes palpable|0
no axillary lymph nodes palpable|0
hemoglobin of 11.3 g/dL|0
low white blood cell of 0.5 × 106/L|0
neutrophil predominance (86.1%)|0
platelet count of 80 × 106/L|0
C-reactive protein of 28.28 mg/dL|0
acute kidney injury|0
serum sodium 137 mmol/L|0
potassium 3.7 mmol/L|0
urea 14 mmol/L|0
creatinine of 206 μmol/L|0
liver function tests normal except serum albumin of 22 g/dL|0
creatinine kinase 351 IU/L|0
arterial blood gases: pH 7.378|0
pCO2 37 mmHg|0
pO2 52.7 mmHg|0
O2 saturation of 89%|0
HCO3 21.7 mmol/L|0
Dengue NS-1 Antigen negative|0
Dengue IgG antibody negative|0
Dengue IgM antibody negative|0
chest radiograph showed consolidation of right upper lobe and left lower lobes|0
diagnosis of severe community acquired pneumonia (CAP)|0
resuscitated with normal saline|0
non-invasive ventilation|0
blood pressure remained hypotensive|0
required inotropic support|0
commenced intravenous ceftriaxone|0
commenced azithromycin|0
condition deteriorated|0
intubation|0
mechanical ventilation in ICU|0
persistent type 2 respiratory failure|0
bronchoscopy done|48
copious amount of haemoserous secretion|48
greenish secretion|48
repeated chest radiograph showed worsening consolidation|48
early changes of abscess formation|48
antibiotics upgraded to intravenous meropenem|48
antibiotics upgraded to cloxacillin|48
antiviral oseltamivir added|48
required continuous venous-venous haemofiltration|48
severe metabolic acidosis|48
oliguric acute kidney injury|48
persistent spiking of temperature|72
worsening septic parameters|72
refractory hypotension|72
patient died|72
blood cultures negative|72
atypical bacterial serologies negative|72
Leptospiral serologies negative|72
Hepatitis B serology undetected|72
Hepatitis C serology undetected|72
HIV serology undetected|72
respiratory viruses screening negative|72
tracheal aspiration positive for MDR Acinetobacter baumannii|72
bronchoalveolar lavage positive for MDR Acinetobacter baumannii|72
MDR Acinetobacter baumannii susceptible only to polymyxin B|72
minimum inhibitory concentration (MIC) of 0.5 μg/ml|72
MDR Acinetobacter baumannii resistant to penicillin group|72
resistant to ampicillin/sulbactam|72
resistant to third generation cephalosporins|72
resistant to fluoroquinolone|72
resistant to carbapenem group|72
smoker|0
