25 years old | 0
primigravida | 0
male infant | 0
40 + 2 weeks’ gestation | 0
spontaneous onset of labor | 0
fetal distress | 0
ventouse-assisted delivery | 0
birth weight 3940 grams | 0
resuscitation with mask ventilation | 0
intubated | 0.13
transferred to NICU | 0
synchronized intermittent positive pressure ventilation (SIPPV) | 0
gentamicin 4 mg/kg 24-hourly | 0
benzyl penicillin 60 mg/kg 12-hourly | 0
neutropenia | 18
left shift | 18
elevated C-reactive protein (CRP; 60 mg/L) | 18
elevated procalcitonin (68.55 µg/L) | 18
lumbar puncture | 23
normal cell count | 23
negative for pathogens | 23
placental surface eSwab | 23
Gram-negative diplococci | 23
Neisseria meningitidis | 23
molecular testing | 23
blood cultures negative | 0.48
heel-prick blood in EDTA | 5.5
N. meningitidis genogroup W DNA | 5.5
benzylpenicillin dosage decreased | 13.5
cefotaxime 50 mg/kg 12-hourly | 13.5
maternal bloods taken | -2.5
elevated leucocyte count | -2.5
neutrophil count | -2.5
mother remained well | 0
baby improved | 13.5
discharged home | 192
contact tracing | 192
chemoprophylaxis with ciprofloxacin | 192
vaccination with quadrivalent conjugate meningococcal vaccine | 192
counseling | 192
funisitis | 0
chorioamnionitis | 0
maternal and fetal inflammatory response | 0
extubated | 13.5