45 years old | 0  
    male | 0  
    admitted to the hospital | 0  
    first symptoms: fever | -144  
    first symptoms: mild dyspnoea | -144  
    first symptoms: fatigue | -144  
    presented to the emergency department | -144  
    computed tomography of the thorax showed mild ground-glass opacities | -144  
    nasopharyngeal swab for SARS-CoV-2 tested negative | -144  
    transferred to the intensive care unit | -138  
    diagnosis of cardio-septic shock | -138  
    pyretic | -138  
    hypoxic (SpO2 85%) | -138  
    severe biventricular impairment | -138  
    metabolic acidosis (pH 7.26; lactate 9 mmol/L) | -138  
    non-invasive mechanical ventilation | -138  
    inotropic support with noradrenaline | -138  
    inotropic support with adrenaline | -138  
    empiric antibiotic therapy | -138  
    worsening hypotension | -134  
    persistent metabolic acidosis | -134  
    intra-aortic balloon pump (IABP) placed | -134  
    conditions remained critical but stable | -128  
    bronchoscopy performed | -128  
    bronchoalveolar lavage tested positive for SARS-CoV-2 | -128  
    clinical stabilization | -108  
    IABP removed | -108  
    complete weaning from inotropic support | -108  
    transferred to the Cardiology department | -102  
    decent clinical condition | -102  
    haemodynamically stable | -102  
    cardiac MRI: severe biventricular dysfunction | -102  
    augmented T1 mapping | -102  
    signs of acute myocarditis | -102  
    myocardial biopsy of the right ventricle | -90  
    histology revealed mild lymphohistiocytic infiltrate | -90  
    diffuse platelet clots | -90  
    Parvovirus B-19 DNA detected | -90  
    SARS-CoV-2 RNA not detected | -90  
    Levosimendan 0.5 μg/kg/min administered | -84  
    persistent severe ventricular impairment | -84  
    intense fatigue | -84  
    discussion with immuno-rheumatologist | -78  
    subcutaneous Anakinra 100 mg bid started | -78  
    clinical conditions ameliorated | 0  
    blood tests ameliorated | 0  
    echocardiography revealed significant improvement of biventricular function | 0  
    discharged | 168  
    first follow-up: good clinical conditions | 432  
    mild effort dyspnoea | 432  
    stable improvement of biventricular function at MRI | 432  
    LVEF 47% | 432  
    RVEF 48% | 432  
    normalization of T1 mapping | 432  
    second follow-up: good clinical conditions | 672  
    no more dyspnoea for mild effort | 672  
    cardiac MRI: normalization of biventricular function | 672  
    LVEF 55% | 672  
    RVEF 56% | 672  
    admitted to ICU | 0  
    shortness of breath | 0  
    confusion | 0  
    severe asthenia | 0  
    arterial blood pressure 75/50 mmHg | 0  
    heart rate 120 bpm | 0  
    peripheral oxygen saturation 85% | 0  
    diffuse bilateral reduction in vesicular breath sounds | 0  
    tachypnoea | 0  
    axillary temperature 37.8°C | 0  
    ECG showed sinus tachycardia | 0  
    diffuse repolarization abnormalities | 0  
    low peripheral voltages | 0  
    mild leukocytosis (WBC 11.1 ×10^9/L) | 0  
    thrombocytopenia (54 ×10^9/L) | 0  
    high sensitive troponin T increased (max 39 ng/dL) | 0  
    peak NT-proBNP 17,000 pg/mL | 0  
    C-reactive protein 285 mg/L | 0  
    chest X-ray: vascular congestion | 0  
    bilateral interstitial alterations | 0  
    transthoracic echocardiography: LVEF 25% | 0  
    TAPSE 12 mm | 0  
    diffuse wall hypokinesia | 0  
    mild biventricular dilatation | 0  
    no significant valvular disease | 0  
    thoracic CT: minute bilateral ground-glass opacities | 0  
    absence of coronary artery stenosis | 0  
    absence of aortic disease | 0  
    nasopharyngeal swab for SARS-CoV-2 RNA negative | 0  
    epidemiological investigation revealed contact with colleague from Lodi | 0  
    colleague’s parents had fever | 0  
    bronchoalveolar lavage detected SARS-CoV-2 RNA | 0  
    repeated nasopharyngeal swabs negative | 0  
    repeated blood cultures negative | 0  
    treated with non-invasive mechanical ventilation | 0  
    hydroxychloroquine 200 mg bid | 0  
    large-spectrum empirical antibiotic therapy | 0  
    needed mechanical circulatory support with IABP | 0  
    inotropes (noradrenaline 0.15 μg/kg/min) | 0  
    inotropes (adrenaline 0.15 μg/kg/min) | 0  
    worsening hypotension | 0  
    severe metabolic acidosis | 0  
    hyper-lactacidaemia | 0  
    pH 7.26 | 0  
    base excess −10 mmol/L | 0  
    lactates 9 mmol/L | 0  
    mechanical circulatory support attempted with IABP | 0  
    weaned from IABP and inotropes | 0  
    transferred to Clinical Cardiology department | 0  
    cardiac MRI confirmed severe biventricular dysfunction | 0  
    higher T1 and T2 mapping | 0  
    absence of late gadolinium enhancement | 0  
    myocardial biopsy: mild lymphohistiocytic inflammatory infiltrate | 0  
    no myocardial necrosis | 0  
    diffuse platelets clots | 0  
    Parvovirus B19 DNA detected | 0  
    SARS-CoV-2 RNA not detected in cardiac tissue | 0  
    levosimendan 0.05 μg/kg/min infusion | 0  
    collegial discussion with immunology consultant | 0  
    off-label therapy with Anakinra 100 mg b.i.d. | 0  
    echocardiography showed LVEF 40-45% | 0  
    TAPSE 18 mm | 0  
    no arrhythmias recorded | 0  
    discharged with optimal medical therapy | 0  
    Metoprolol 50 mg daily | 0  
    Ramipril 2.5 mg daily | 0  
    Spironolactone 37 mg daily | 0  
    Furosemide 25 mg daily | 0  
    6-month therapy with Anakinra | 0  
    clinical conditions improved | 168  
    blood tests improved | 168  
    echocardiography improvement | 168  
    cardiac MRI at follow-up: biventricular improvement | 432  
    absence of late gadolinium enhancement | 432  
    T1 and T2 mapping normalization | 432  
    complete recovery of biventricular function | 672  
    LVEF 55% | 672  
    RVEF 56% | 672  

