77 years old | 0
    male | 0
    admitted to the hospital | 0
    abdominal distension | -168
    increased abdominal girth | -168
    diarrhea | -168
    infrequent vomiting | -168
    weight loss | -168
    anorexia | -168
    no abdominal pain | 0
    mild metabolic alkalosis | 0
    slight elevation of C-reactive protein | 0
    contracted gallbladder | 0
    thick gallbladder | 0
    gallbladder stones | 0
    gas bubbles in gallbladder | 0
    cholecystocolonic fistula suspected | 0
    abdominal distension persisted | 0
    diarrhea persisted | 0
    HIDA scan showed no gallbladder filling | 24
    cystic duct occlusion | 24
    ERC performed | 24
    common bile duct free of stones | 24
    right hepatic duct free of stones | 24
    left hepatic duct free of stones | 24
    cystic duct occlusion confirmed | 24
    sphincterotomy performed | 24
    pancreatic stent placed | 24
    fever | 20
    hypotension | 20
    tachycardia | 20
    transferred to ICU | 20
    CT scan showed free intraabdominal fluid | 20
    normal serum amylase | 20
    normal serum lipase | 20
    biliary sepsis suspected | 20
    open abdominal exploration | 20
    hepatic flexure adherent to gallbladder | 20
    fistulous tract identified | 20
    stones retrieved from gallbladder | 20
    colonic mucosa biopsied | 20
    frozen section analysis | 20
    partial cholecystectomy | 20
    fulguration of remaining mucosa | 20
    acute cholecystitis | 20
    chronic cholecystitis | 20
    hepatic flexure resected | 20
    external drainage tube placed | 20
    hospitalized for two weeks | 336
    nocturnal desaturation | 336
    central sleep apnea | 336
    discharged | 336
    right upper quadrant abscess | 504
    antibiotics administered | 504
    percutaneous drainage | 504
    uneventful follow-up | 8760
    