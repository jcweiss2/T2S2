57 years old | 0
male | 0
admitted to the hospital | 0
diagnosed as Philadelphia-positive ALL | -168
remission-induction chemotherapy | -168
intra-thecal chemotherapy | -168
hospital day 1 | 0
initial vital signs stable | 0
blood pressure 110/60 mmHg | 0
pulse rate 80/min | 0
respiratory rate 20/min | 0
body temperature 36.4℃ | 0
pre-transplant conditioning chemotherapy | 96
fludarabine | 96
melphalan | 96
anti-thymocyte immunoglobulin | 96
ciprofloxacin | 96
itraconazole syrup | 96
acyclovir | 96
SCT | 288
neutropenia | 288
intermittent mild abdominal pain | 336
diarrhea | 336
C. difficile toxin assay | 96
C. difficile culture | 96
severe pain at the left chest wall | 432
severe pain at the left buttock | 432
severe pain at the left thigh | 432
localized swelling | 432
tissue edema | 432
empirical antibiotics | 432
piperacillin/tazobactam | 432
vancomycin | 432
complete blood cell count | 432
hemoglobin of 9.3 g/dL | 432
hematocrit of 25.2% | 432
white blood cells of 10/mm3 | 432
ANC 0/mm3 | 432
platelet 61,000/mm3 | 432
Ciprofloxacin stopped | 432
chest X-ray | 432
soft tissue swelling with air density | 432
blood pressure 92/60 mmHg | 432
heart rate 164/min | 432
oxygen saturation 83% | 432
normal saline | 432
oxygen via a simple facial mask | 432
vital signs stabilized | 432
chest and abdominal computed tomography | 432
multiple emphysematous soft tissue infection | 432
needle aspiration | 442
heart rate increased to 163/min | 442
blood pressure 98/63 mmHg | 442
planned to be transferred to intensive care unit | 442
cardiac arrest | 444
cardiopulmonary resuscitation | 444
died | 444
Clostridium perfringens isolated | 444
blood cultures | 444
culture of aspirated fluid | 444
chronic diarrhea | -720