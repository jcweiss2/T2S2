73 years old | 0
male | 0
admitted to the hospital | 0
lower back pain | 0
severe fatigue | 0
20-kg weight loss | 0
transitional cell bladder cancer | -48
invasion of the submucosa | -48
transurethral resection | -48
intravesical mitomycin | -48
recurrence of disease | -24
transurethral resection of a low-grade non-muscle-invasive tumor | -24
adjuvant therapy with intravesical BCG solution | -24
peripheral edema of the lower extremities | 0
pain on palpation cranial to the left iliac crest | 0
positron emission tomography scan | 0
pathologic activity of the abdominal aorta and left iliopsoas muscle | 0
thoracoabdominal computed tomography scan | 0
pseudoaneurysm of the abdominal aorta and surrounding infiltration | 0
mycotic aneurysm | 0
elective open aorta reconstructive surgery | 0
intravenous perioperative antibiotic prophylaxis with cephalosporin and metronidazole | 0
operation | 0
neoaortoiliac system bypass | 0
reconstructive repair with a bovine tube graft | 0
infected aneurysmal segment excised | 0
collection of softened, infected mushy tissue | 0
culture and biopsy specimens from the aorta and surrounding tissue | 0
resorbable sponge impregnated with gentamicin | 0
rifampicin applied to the cavity | 0
graft sutured | 0
greater omentum wrap plasty | 0
M. bovis in para-aortic tissue | 0
extensive granulomatous and necrotizing inflammation of the aorta | 0
histologic Ziehl-Neelsen staining | 0
DNA analyses | 0
M. bovis infection | 0
severe inflammatory response syndrome | 12
admitted to the intensive care unit | 12
acute-on-chronic renal insufficiency | 12
hemodialysis | 12
paralytic ileus | 12
chylous ascites | 12
paracentesis | 12
total parenteral nutrition | 12
administration of octreotide | 12
condition improved | 24
hemodialysis stopped | 24
production of chylous ascites diminished | 24
ileus resolved | 24
transferred to the general surgery ward | 24
transferred to a rehabilitation center | 144
antimicrobial treatment with rifampicin, ethambutol, and isoniazid | 144
fever | 216
generalized weakness | 216
malaise | 216
elevated C-reactive protein level | 216
leukocytosis | 216
fluid collection on the left dorsolateral side of the bovine aorta tube graft | 216
CT-guided drainage | 216
mycobacterium in the aspirated fluid | 216
treatment for active infection and paradoxical abscess formation | 216
antibiotic treatment regimen changed to rifampicin, ethambutol, and moxifloxacin | 216
paradoxical abscess formation treated with drainage and dexamethasone | 216
condition improved | 240
follow-up CT scan | 240
collection decreased | 240
discharged | 240