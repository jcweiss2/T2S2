26 years old | 0 | 0 
female | 0 | 0 
admitted to the hospital | 0 | 0 
rising levels of human chorionic gonadotropin | -336 | 0 
intermittent vaginal bleeding | -336 | 0 
vaginal ultrasound scan | -336 | 0 
intrauterine pregnancy | -336 | 0 
legal medical abortion | -336 | 0 
vaginal ultrasound | 0 | 0 
placental remnants in the uterus | 0 | 0 
surgical evacuation of the uterus | 0 | 0 
discharged | 12 | 12 
readmitted | 24 | 24 
temperature of 39.5°C | 24 | 24 
abdominal pain | 24 | 24 
severe endometritis | 24 | 24 
metronidazole | 24 | 48 
benzylpenicillin | 24 | 48 
gentamicin | 24 | 48 
deterioration | 48 | 48 
saturation fell to 90% | 48 | 48 
respiratory rate rose to around 40 breaths per minute | 48 | 48 
oxygen given by mask | 48 | 48 
temperature peaked at 40.7°C | 48 | 48 
C-reactive protein rose to around 300 mg/L | 48 | 48 
leukocytes to around 15 × 10^9/L | 48 | 48 
intubated | 48 | 48 
moved to the intensive care unit | 48 | 48 
CT scan | 48 | 48 
thrombophlebitis of the internal jugular vein | 48 | 48 
hepatomegaly | 48 | 48 
diagnosed with Lemierre's syndrome | 48 | 48 
benzylpenicillin discontinued | 48 | 48 
gentamicin discontinued | 48 | 48 
tazocin | 48 | 336 
clindamycin | 48 | 336 
metronidazole | 48 | 336 
heparin injections | 48 | 336 
recovered | 336 | 336 
discharged | 336 | 336 
infection with F. necrophorum | 0 | 336 
blood cultures | 48 | 48 
F. necrophorum cultivated from the patient's cervix | 48 | 48 
no symptoms from the oropharyngeal tract | 0 | 336 
respiratory support | 48 | 336 
antibiotics | 24 | 336 
anticoagulation | 48 | 336 
surgical drainage of abscesses | 48 | 336 
patient gave consent to the publication | 0 | 0 
no conflict of interest | 0 | 0