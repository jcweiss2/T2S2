33 years old | 0
male | 0
admitted to the emergency room | 0
severe abdominal pain | -720
vomiting | -720
abdominal pain continued after breakfast | 0
visited another hospital before admission | -720
pain did not diminish | -720
experienced minor mental deterioration | -720
transferred to the ER with suspected ileus | -720
vital signs upon arrival: BP 105/63 mmHg | 0
HR 69 beats/min | 0
SpO2 99% | 0
RR 20 rates/min | 0
body temperature 36.9℃ | 0
arterial blood gas analysis: pH 7.64 | 0
PaCO2 25.8 mmHg | 0
PaO2 111.1 mmHg |0
BE 8.3 mmol/L |0
chest radiograph |0
chest and abdominal CT |0
BP 83/66 mmHg |0
HR increased from 70 to 116 beats/min |0
administration of 100 ml crystalloid fluids |0
BP 124/88 mmHg |0
severe increase in stomach volume observed through CT |0
stricture in gastric pylorus and duodenum |0
attempted insertion of nasogastric tube unsuccessful |0
pneumomediastinum suggested |0
esophageal rupture suspected |0
right internal jugular vein catheterization |0
BP 84/44 mmHg |0
HR 113 beats/min |0
administration of 300 ml crystalloid solution |0
2 L/min oxygen via nasal cannula |0
SpO2 97% |0
esophageal rupture suspected 24 hours after vomiting |24
moved to operating room |24
fasting time 12 hours |24
preoperative blood tests: blood urea nitrogen 32 mg/dl |24
creatine 2.2 mg/dl |24
white blood cell 12,400/mm3 |24
clear consciousness |24
preoperative BP 80/50 mmHg |24
HR 125 beats/min |24
SpO2 94% on FIO2 0.21 |24
preoxygenation with 100% oxygen |24
SpO2 99% |24
general anesthesia induced |24
etomidate 15 mg |24
cisatracurium 20 mg |24
manual ventilation: TV 400-500 ml |24
RR 15 rates/min |24
PIP 15-25 cmH2O |24
ETCO2 30&ndash;40 mmHg |24
endotracheal intubation with DLT |24
breath sounds confirmed |24
tube position confirmed with bronchoscope |24
mechanical ventilation: PCV mode |24
PIP 20 cmH2O |24
PEEP 0 cmH2O |24
RR 12 rates/min |24
TV 500-600 ml |24
FIO2 1.0 |24
anesthesia maintained with desflurane 2 vol% |24
dopamine 5 µg/kg/min |24
systolic BP 90-110 mmHg |24
diastolic BP 50-70 mmHg |24
HR 110-120 beats/min |24
central venous pressure 14-16 cmH2O |24
ETCO2 30-35 mmHg |24
BIS 30-40 |24
right lateral position for left thoracotomy |24
single right lung ventilation |24
PCV mode: PIP 20 cmH2O |24
TV 300-400 ml |24
ABGA: pH 7.439 |24
PaCO2 36.5 mmHg |24
PaO2 154.3 mmHg |24
BE 1.3 mmol/L |24
SpO2 gradually decreased |24
manual ventilation performed |24
tube position confirmed |24
volatile anesthetics stopped |24
SpO2 80% |24
two-lung ventilation conducted |24
SpO2 not improved |24
breath sounds slightly decreased |24
consultation with thoracic surgeon |24
moved to supine position |24
SpO2 dropped to 70% |24
bilateral breath sounds low |24
DLT position confirmed |24
desaturation persisted |24
DLT replaced with single-lumen tube |24
manual ventilation maintained |24
ETCO2 25-35 mmHg |24
SpO2 dropped to 50% |24
ETCO2 10 mmHg |24
HR below 40 beats/min |24
systolic BP 50 mmHg |24
CPR performed |24
thoracic compressions |24
epinephrine 1 mg injected twice |24
bilateral breath sounds disappeared |24
bilateral tension pneumothorax suspected |24
20 gauge angiocatheter inserted left mid-clavicle |24
air leakage confirmed |24
right mid-clavicle angiocatheter inserted |24
air leakage with brown liquid |24
SpO2 increased to 90% |24
HR improved to 70-80 beats/min |24
systolic BP 100-120 mmHg |24
SpO2 94-95% |24
BIS score above 10 |24
CPR terminated |24
emergency chest radiograph |24
chest tube inserted right chest |24
chest tube inserted left chest |24
breath sounds recovered |24
SpO2 100% |24
stomach contents gushing out |24
air leaking from right chest tube |24
severe lung parenchymal damage suspected |24
changed to left-lung ventilation |24
DLT inserted again |24
right thoracotomy performed |24
suctioned 500 ml stomach contents |24
lung irrigation |24
chemical burn observed |24
esophageal rupture on left side |24
right thoracotomy |24
ruptures in epiphrenic esophagus and subphrenic stomach |24
distal esophagectomy |24
esophagogastrostomy |24
feeding jejunostomy |24
surgical time 11 hours |24
fluids administered: colloid 4500 ml |24
crystalloid 4050 ml |24
packed red blood cells 2 pints |24
estimated blood loss 1000 ml |24
urine output 1700 ml |24
ABGA: pH 7.429 |24
PaCO2 31.3 mmHg |24
PaO2 367.7 mmHg |24
BE -2.2 mmol/L |24
tube replaced with single-lumen |24
transferred to ICU |24
chest radiography: no pulmonary edema |24
mechanical ventilation: assisted control mode |24
pressure 14 cmH2O |24
RR 12 breaths/min |24
PEEP 6 cmH2O |24
FIO2 0.6 |24
fentanyl infusion 20-40 µg/h |24
ABGA 2 hours post-op: pH 7.43 |24
PaCO2 31 mmHg |24
PaO2 211 mmHg |24
BE -2 mmol/L |24
drowsy mental status |24
mechanical ventilation continued |24
FIO2 decreased to 0.4 |24
ABGA: pH 7.39 |24
PaCO2 35 mmHg |24
PaO2 169 mmHg |24
BE -2.0 mmol/L |24
vital signs stable |24
SpO2 99% on FIO2 0.4 |24
mechanical ventilation stopped |120
T-piece applied |120
extubated |168
moved to general ward |192
vital signs stable |192
mental status alert |192
SpO2 97% on 3 L/min oxygen |192
left chest tube removed |264
right chest tube removed |600
discharged |768
