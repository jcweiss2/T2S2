32 years old | 0
male | 0
smoker | 0
occasional drinker | 0
technician in a factory | 0
sudden onset severe abdominal pain | -24
syncope | -24
hypotension (systolic blood pressure 50+) | -24
no change in bowel habit | 0
no recent loss of appetite | 0
no recent loss of weight | 0
never experienced abdominal pain like this before | 0
severely tender abdomen | 0
tense abdomen | 0
bedside ultrasound demonstrated free fluid | 0
large 8x9cm AAA | 0
CT aortogram confirmed tortuous and aneurysmal dilatation of the abdominal aorta | 0
abdominal aorta measuring up to 10.8 × 10.8 cm in axial dimension | 0
abdominal aorta measuring 24.1 cm in cranio-caudal length | 0
extends into the left common iliac artery | 0
proximal aspect involving the origin of the bilateral renal arteries | 0
large retroperitoneal hematoma | 0
emergency open abdominal aortic aneurysm repair | 0
difficult access | 0
haemodynamic instability | 0
need for an expedited procedure | 0
aortic cross clamp applied beneath the right renal artery | 0
aortic cross clamp applied just proximal to left renal artery | 0
bifurcated aortic graft anastomosed proximally | 0
no need for renal artery implantation | 0
anastomosed distally to the bilateral common iliac arteries | 0
on table angiogram of the left lower limb | 0
pale left lower limb intraoperatively | 0
abrupt cut-off at the level of the left popliteal artery | 0
transverse arteriotomy over the left common femoral artery | 0
Fogarty balloon catheter used to trawl out multiple thrombi | 0
final angiogram demonstrated in-line flow to the foot via the anterior tibial artery | 0
foot pulses palpable | 0
strong foot pulses | 0
transferred to the intensive care unit (ICU) | 0
extubated on post-operative day (POD) 1 | 24
intensive chest physiotherapy | 24
incentive spirometry | 24
nasogastric feeding started on POD2 | 48
oral diet by POD 6 | 144
developed a fever on the 4th day of ICU stay | 96
fever secondary to basal atelectasis | 96
empirically started on piperacillin-tazobactam | 96
piperacillin-tazobactam stopped 4 days later | 192
negative septic work up | 192
down-trending inflammatory markers | 192
pro-calcitonin level within normal limits | 192
surgical sites healing well | 192
no hematoma at surgical sites | 192
no signs of infection at surgical sites | 192
acute kidney injury during ICU stay | 96
managed with proper hydration | 96
normalising of renal function | 192
transient liver enzyme rise | 96
transient liver enzyme rise resolved gradually | 192
preserved coagulation profile | 192
clinically stable by POD 12 | 288
independently mobile by POD 12 | 288
fit for discharge from hospital by POD 12 | 288
discharged from hospital | 288
histopathological examination revealed degenerative changes of the aortic wall | 0
aortic rupture | 0
no granulomas | 0
no giant cells | 0
no obliterative phlebitis | 0
no storiform fibrosis | 0
no malignancy | 0
not suggestive of tuberculosis | 0
no vasculitic changes | 0
no IgG4 sclerosing disease | 0
no evidence of infective process in the aortic wall | 0
etiology of AAA of interest | 0
large size AAA | 0
young age at presentation | 0
multiple investigations while in hospital | 0
returned to Vietnam after discharge | 288
lost to follow up | 288
genetic testing not arranged | 288
mother had significant bilateral hallux valgus | 0
youngest sibling has pectus carinatum | 0
no known cardiac disease in the family | 0
no known lung disease in the family | 0
no known rheumatological disease in the family | 0
taller than peers | 0
height 179 cm | 0
body mass index 24.2 kg/m2 | 0
average head width 19 cm | 0
average head length 22 cm | 0
normal arched palate | 0
triangular uvula centre | 0
mild pectus excavatum | 0
no obvious scoliosis | 0
no truncal striae | 0
unusually long and slender fingers | 0
unusually long and slender toes | 0
no deformities | 0
no positive thumb sign | 0
bilateral pes planus | 0
arachnodactyly | 0
keloid at midline laparotomy wound | 0
high C-reactive protein (241.6 mg/L) | 0
elevated CRP remained on discharge (71.6 mg/L) | 288
elevated erythrocyte sedimentation rate (35 mm/h) | 0
no evidence of atheroma on imaging | 0
normal serum cholesterol | 0
normal homocysteine level | 0
no tell-tale clinical features of rheumatological disorders | 0
no dry eyes | 0
no xerostomia | 0
no abnormal hair loss | 0
no rashes | 0
no concomitant aortic root involvement | 0
no cardiac involvement | 0
echocardiography not performed | 0
explained need for genetic testing | 288
offered free genetic testing | 288
