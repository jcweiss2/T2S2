43 years old | 0
    male | 0
    diagnosed with epileptic disorder | -240
    phenytoin 100 mg thrice daily | -240
    sudden onset of fluid-filled lesions | -48
    fluid-filled lesions increased in number | -48
    fluid-filled lesions increased in surface area | -48
    blisters started bursting out releasing watery fluid | -48
    developed fever | -48
    developed easy fatigability | -48
    developed breathlessness | -48
    symptoms progressively increased | -48
    symptoms worsened | -48
    admitted to the hospital | 0
    severe respiratory distress | 0
    gasping for breath | 0
    unconscious | 0
    not responding to deep stimuli | 0
    low saturation | 0
    blood pressure not recordable | 0
    intubated | 0
    mechanical ventilation | 0
    inotropes started | 0
    multiple ruptured bullae all over the body | 0
    erythematous skin | 0
    oral mucosa involved | 0
    conjunctival mucosa involved | 0
    provisional diagnosis of SJS | 0
    elevation in cardiac biomarkers | 0
    echocardiogram revealed global hypokinesia | 0
    prothrombin time 15 s | 0
    activated partial thromboplastin time 32 s | 0
    platelet count 143,000 L/mm3 | 0
    normal liver function tests | 0
    ICU care | 0
    inotropes continued | 0
    hydrocortisone 100 mg injection started | 0
    myocarditis managed conservatively | 0
    switched to sodium valproate 1000 mg twice a day | 0
    renal parameters deranged | 12
    blood pressure 80/60 mmHg | 12
    Glasgow coma scale score 4/15 | 12
    near-normal leukocyte count | 12
    no improvement in clinical parameters | 12
    no improvement in biochemical parameters | 12
    sudden cardiac arrest | 18
    revived | 18
    sustained another cardiac arrest | 19
    declared dead | 19
    <|eot_id|>

  43 years old | 0
male | 0
diagnosed with epileptic disorder | -240
phenytoin 100 mg thrice daily | -240
sudden onset of fluid-filled lesions | -48
fluid-filled lesions increased in number | -48
fluid-filled lesions increased in surface area | -48
blisters started bursting out releasing watery fluid | -48
developed fever | -48
developed easy fatigability | -48
developed breathlessness | -48
symptoms progressively increased | -48
symptoms worsened | -48
admitted to the hospital | 0
severe respiratory distress | 0
gasping for breath | 0
unconscious |8
not responding to deep stimuli |0
low saturation |0
blood pressure not recordable |0
intubated |0
mechanical ventilation |0
inotropes started |0
multiple ruptured bullae all over the body |0
erythematous skin |0
oral mucosa involved |0
conjunctival mucosa involved |0
provisional diagnosis of SJS |0
elevation in cardiac biomarkers |0
echocardiogram revealed global hypokinesia |0
prothrombin time 15 s |0
activated partial thromboplastin time 32 s |0
platelet count 143,000 L/mm3 |0
normal liver function tests |0
ICU care |0
inotropes continued |0
hydrocortisone 100 mg injection started |0
myocarditis managed conservatively |0
switched to sodium valproate 1000 mg twice a day |0
renal parameters deranged |12
blood pressure 80/60 mmHg |12
Glasgow coma scale score 4/15 |12
near-normal leukocyte count |12
no improvement in clinical parameters |12
no improvement in biochemical parameters |12
sudden cardiac arrest |18
revived |18
sustained another cardiac arrest |19
declared dead |19