80 years old | 0 | 0 
female | 0 | 0 
non-smoker | 0 | 0 
hypertension | 0 | 0 
admitted to the hospital | 0 | 0 
acute dyspnea | -24 | 0 
fecal incontinence | -6.67 | -6.67 
left hemiplegia | -6.67 | -6.67 
dextroversion | -6.67 | -6.67 
dysarthria | -6.67 | -6.67 
vomiting | -6.67 | -6.67 
impaired consciousness | -6.67 | 0 
Japan coma scale score of Ⅱ-10 | -6.67 | 0 
right thalamus and putamen bleeding | -6.67 | 0 
Glasgow coma scale score 12 | 0 | 0 
systolic blood pressure 91 mmHg | 0 | 0 
respiratory rate 24/min | 0 | 0 
oxygen saturation of arterial blood 86% | 0 | 0 
poor oral hygiene | 0 | 0 
diminished breath sounds on the left side | 0 | 0 
coarse crackles in the right lung | 0 | 0 
decrease in breath sounds in the front of the chest | 0 | 0 
respiratory condition deteriorated | 0 | 2 
endotracheal intubation | 2 | 2 
mechanical ventilation | 2 | 240 
bilateral infiltration | 2 | 2 
admitted to the intensive care unit | 2 | 2 
leukocyte count 1900/μL | 2 | 2 
C-reactive protein level 3.6 mg/dL | 2 | 2 
respiratory failure | 2 | 2 
partial pressure of oxygen in arterial blood 64 mmHg | 2 | 2 
hepatorenal function normal | 2 | 240 
extensive infiltration shadows | 2 | 2 
hematoma extending from the right basal ganglia and putamen to the thalamus | 2 | 2 
cerebral edema | 2 | 2 
consolidations admixture with ground-glass opacities | 2 | 2 
A-DROP score corresponded to patient age | 2 | 2 
increased blood urea nitrogen | 2 | 2 
decreased SpO2 | 2 | 2 
impaired consciousness | 2 | 2 
antigen test for coronavirus disease 2019 negative | 2 | 2 
Mendelson's syndrome | 2 | 240 
aspiration bacterial pneumonia | 2 | 240 
sputum culture showed Streptococcus agalactiae and Klebsiella oxytoca | 24 | 24 
leukocytopenia | 2 | 24 
low serum CRP level | 2 | 24 
elevated WBC | 24 | 240 
elevated serum CRP level | 24 | 240 
management in the ventilator mode | 24 | 240 
meropenem | 24 | 240 
levofloxacin | 24 | 240 
partial pressure of oxygen in arterial blood/fraction of inspired oxygen 128.75 | 24 | 24 
prednisolone | 24 | 240 
infiltration shadows improved | 240 | 240 
extubated | 240 | 240 
transferred to the Department of Neurosurgery | 528 | 528 
transferred to a rehabilitation hospital | 528 | 528