60 years old | 0
female | 0
admitted to the emergency unit | 0
pain | -48
paresthesia | -48
coolness of the right lower leg and foot | -48
cesarean section | -8760
cold toes | 0
capillary filling lasting more than 5 s | 0
absent distal pulses in both legs | 0
computed tomography angiography | 0
floating thrombus in the abdominal aorta | 0
thromboembolism of the entire right deep femoral artery | 0
thromboembolism of the distal part of the left deep femoral artery | 0
sustained flow in both superficial femoral arteries | 0
occlusion of the third segment of the right popliteal artery | 0
thromboembolus in the posterior tibial artery | 0
marginal recanalization | 0
surgical thromboembolectomy | 0
treated with LMWH | 0
treated with proton pump inhibitor | 0
treated with analgesic therapy | 0
treated with cefuroxime | 0
transfusions of deplasmatized red blood cells | 0
positive PCR test for SARS-CoV-2 | 0
treated with oral amoxicillin and clavulanic acid | 14
treated with intravenous PPI | 14
treated with subcutaneous LMWH | 14
homozygous MTHFR C677T gene mutation | 14
discharged | 336
nausea | 6720
jaundice | 6960
admitted to the intensive care unit | 6960
ALI of unknown etiology | 6960
liver damage | 6960
fulminant liver failure | 6960
acute hepatocellular injury | 6960
DILI | 6960
grade 3 hepatic encephalopathy | 6960
mechanical ventilation | 6960
tonic-clonic seizures | 6960
diffuse brain edema | 6960
brain edema progression | 6960
death | 6972
autopsy not performed | 6972
rivaroxaban 15 mg BID | 336
PPI QD | 336