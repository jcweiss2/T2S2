22 years old | 0
male | 0
admitted to the hospital | 0
fever | -360
escharotic and purpuric skin lesions | -360
self-administered ibuprofen | -168
self-administered diclofenac sodium | -168
cephalosporin antibiotics | -96
history of alcoholism | -8760
body temperature 39°C | 0
pulse 120 bpm | 0
blood pressure 154/108 mmHg | 0
height 166 cm | 0
weight 90 kg | 0
severe obesity | 0
black necrotic eschar | 0
subcutaneous nodules | 0
enlarged lymph nodes | 0
purpuric and necrotic crusted lesions | 0
thrombosis in the small saphenous vein | 0
thrombosis in the great saphenous vein | 0
thrombosis in the cephalic vein | 0
cerebral infarction | 0
intracranial infection | 0
lung infection | 0
pleurisy | 0
pericardial effusion | 0
pain in the skin lesions | 48
pain in the back | 48
headache | 48
vertigo | 48
sputum-free cough | 48
diarrhea | 48
stomach ache | 48
abdominal pain | 168
hematemesis | 168
blood in the stool | 168
occult blood tests positive | 168
gastrointestinal bleeding | 168
pulmonary embolisms | 168
liver damage | 168
multiple embolisms | 168
inflammatory | 168
difficulty breathing | 240
irritability | 240
progressive decline in blood oxygen saturation | 240
respiratory failure | 240
sedative drugs | 240
right subclavian vein puncture | 240
catheterization | 240
intravenous hypernutrition | 240
fiberoptic bronchoscopy | 240
liver function damage | 240
renal function damage | 240
hypokalemia | 240
hyperchloremia | 240
hypernatremia | 240
metabolic acidosis | 240
continuous coma | 240
continuous renal replacement therapy | 480
improved consciousness | 480
tar-like stools | 480
positive occult blood test | 480
increased PLT | 480
extubated | 480
oxygen administered by mask | 480
returned to the Dermatology Department | 528
blood chloride increased | 576
oxygen partial pressure 48% | 576
carbon dioxide partial pressure 23% | 576
HGB 48 g/L | 576
transferred to the ICU | 576
femoral artery puncture catheterization | 576
monitoring by PiCCO | 576
radial artery puncture catheterization | 576
invasive blood pressure monitoring | 576
peripheral puncture central venous catheterization | 576
active bloody stools | 720
bruise | 720
edema | 720
T 37°C–39°C | 864
HGB 80 g/L | 864
returned to the Dermatology Department | 900
red liquid drained from the gastric tube | 984
palpitations | 984
shortness of breath | 984
convulsions | 984
breathing difficulty symptoms worsened | 1056
mask given at 66–78% oxygen saturation | 1056
transferred to the ICU | 1056
thoracentesis catheter drainage | 1056
tracheal intubation | 1056
mechanical ventilation | 1056
condition gradually improved | 1248
T 37°C–37.8°C | 1248
PLT 355 × 10^9/L | 1248
coagulation function improved | 1248
stable condition | 1344
normal body T | 1344
returned to dermatology | 1356
gastroscopy | 1356
varicose veins in the fundus of the stomach | 1356
chronic non-atrophic gastritis | 1356
portal venous system CTA | 1584
splenic infarction | 1584
thrombosis of the portal vein | 1584
thrombosis of the hepatic arteriovenous | 1584
thrombosis of the inferior vena cava | 1584
skin lesion area significantly reduced | 1608
texture became soft | 1608
no tenderness | 1608
purpura-like skin lesions subsided | 1608
vital signs stable | 1608
laboratory indicators stable | 1608
weight dropped to 46 kg | 1608
discharged | 1608