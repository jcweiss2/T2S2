11 years old | 0
female | 0
admitted to the hospital | 0
high fever | -72
nausea | -72
severe weakness | -72
myalgia | -72
main body ache | -72
conscious | 0
pale | 0
ill | 0
body temperature 39.5°C | 0
pulse 120 bpm | 0
blood pressure 110/75 mmHg | 0
no rash | 0
no spontaneous bleeding | 0
no jaundice | 0
hemoglobin 14.8 g/dl | 0
hematocrit 40% | 0
platelet count 140000/mm3 | 0
Dengue IgM antibodies positive | 0
SARS-COV2 antigen nasopharynx test negative | 0
clinical diagnosis suspect of Dengue fever | 0
standard diet | 0
feverish | 24
looked ill | 24
short of breath | 24
nausea | 24
abdominal bloating | 24
platelet count 78000/mm3 | 24
platelet count decreased dramatically to 15000/mm3 | 72
blood pressure 110/90 mmHg | 72
pulse 90 bpm | 72
chest X-ray revealed remarkable pleura effusion | 72
pleural effusion index 38.13% | 72
managed in intensive care unit | 72
severe abdominal pain | 96
abdominal ultrasonography showed acalculous cholecystitis | 96
liver function test elevated AST 151 IU/L | 96
liver function test elevated ALT 59 IU/L | 96
C-reactive protein level increased 14.4 mg/L | 96
managed as DHF and AAC complications | 96
conservative treatment | 96
intravenous antibiotics | 168
no blood transfusion | 168
no hematoma | 168
abdominal pain | 96
abdominal bloating sensation | 96
condition improved gradually | 168
discharged | 168
liver function enzyme restored after treatment | 168
sharp acute abdominal pain | 72
abdominal pain lasted 3 days | 72
abdominal bloating sensation lasted 3 days | 72
platelet count decreased until 4th day | 96
thrombocytopenia | 96
liver dysfunction | 96
elevated transaminase enzymes | 96
no jaundice | 96
acute acalculous cholecystitis confirmed | 96
thickened gallbladder wall over 3.5 mm | 96
increased CRP marker | 96
abnormal liver function test | 96
gallbladder wall thickening | 96
pericholecystic fluid | 96
mucosal membrane sludge | 96
gallbladder distension | 96
improved with conservative therapy | 168
adequate intravenous fluid therapy | 168
analgesic | 168
antibiotics | 168
