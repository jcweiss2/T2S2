55 years old | 0
    male | 0
    common cold | -168
    myalgia | -168
    fatigue | -168
    headaches | -168
    pleuritic chest pain | -168
    breathlessness on exertion | -168
    mild asthma | 0
    Beclomethasone | 0
    salbutamol | 0
    ex-smoker | 0
    body mass index 24.6 kg/m² | 0
    blood pressure 130/80 mmHg | 0
    pulse 110 bpm | 0
    temperature 38.2°C | 0
    decreased air entry on the right lung | 0
    coarse crackles | 0
    normal heart sounds | 0
    no murmurs | 0
    sinus tachycardia 113 bpm | 0
    PR interval 124 ms | 0
    QRS duration 99 ms | 0
    corrected QT interval 382 ms | 0
    no ST-T wave abnormalities | 0
    serum creatinine 85 µmol/L | 0
    alanine aminotransferase 216 IU/L | 0
    potassium level 5.4 mmoL/mL | 0
    magnesium 1.2 | 0
    corrected calcium 2.26 | 0
    sodium 138 | 0
    C-reactive protein 184 mg/L | 0
    haemoglobin 86 g/L | 0
    normocytic normochromic | 0
    platelets 670 × 10^9/L | 0
    WBC 18 × 10^9/L | 0
    neutrophilia | 0
    international normalized ratio 1.4 | 0
    activated partial thromboplastin time 27.2 s | 0
    right sided consolidation | 0
    Pseudomonas aeruginosa | 0
    community acquired P. pneumonia | 0
    oxygen | 0
    intravenous fluids | 0
    antibiotics meropenem | 0
    clarithromycin | 0
    central chest pain | 96
    inferior ST elevation myocardial infarction | 96
    occlusion mid segment of left circumflex artery | 96
    drug-eluting stent | 96
    left anterior descending disease | 96
    atrial fibrillation | 96
    ventricular bigeminy | 96
    dual antiplatelet therapy aspirin | 96
    ticagrelor | 96
    rapid respiratory deterioration | 120
    intubation | 120
    ventilation | 120
    maximum oxygenation | 120
    bronchoscopy | 120
    diuresis | 120
    antibiotic escalation | 120
    type 1 respiratory failure | 120
    proning attempts | 120
    inhaled nitric oxide | 120
    COVID-19 negative | 120
    Murray score 2.5 | 120
    RESP score 5 | 120
    veno(venous ECMO | 144
    retrieval to tertiary centre | 144
    multiple segmental pulmonary emboli | 144
    sub-segmental pulmonary emboli | 144
    left lower lung lobe embolus | 144
    right lower lobe anterior sub-segmental embolus | 144
    no right heart strain | 144
    necrotizing pneumonia | 144
    pleural effusion | 144
    minimal basal consolidation | 144
    peripheral ground glass opacification | 144
    severely impaired left ventricular systolic function | 144
    mild dilatation right ventricle | 144
    moderate to severe impairment right ventricular systolic function | 144
    cardiac output 3.5 L/min | 144
    T-wave inversion inferior leads | 144
    QTc 515 ms | 144
    amiodarone loading dose 300 IV | 144
    amiodarone 900 mg IV | 144
    AF controlled | 144
    ventricular ectopy controlled | 144
    QT prolongation | 144
    antibiotic regimen amikacin | 144
    ceftazidime | 144
    linezolid | 144
    noradrenaline | 144
    potassium level 5.3 mmoL/mL | 144
    magnesium 1.6 | 144
    corrected calcium 2.49 | 144
    temperature 36.1°C | 144
    AF with ventricular rate 140-150 bpm | 168
    increased ventricular ectopy burden | 168
    ventricular bigeminy | 168
    self-terminating ventricular tachycardia | 168
    mean arterial pressure below 59 mmHg | 168
    noradrenaline requirement increased 0.06-0.18 µg/kg/min | 168
    electrolyte replenishment | 168
    renal replacement therapy | 168
    amiodarone reloading | 168
    metoprolol 25 mg TDS | 168
    esmolol 50 mcg/kg/min | 168
    bradycardia | 168
    hypotension | 168
    first degree AV block | 168
    QTc prolongation 550 ms | 168
    lidocaine infusion ineffective | 168
    worsening cardiogenic shock | 168
    AF | 168
    ventricular tachycardia | 168
    ventricular ectopy | 168
    severely impaired left ventricular systolic function | 168
    repeat coronary angiography | 192
    patent LCx stent | 192
    two drug-eluting stents LAD | 192
    arrhythmia burden not improved | 192
    short-acting beta-blockers restarted | 192
    amiodarone when QTc below 480 ms | 192
    QTc prolongation 550 ms | 288
    Torsade de pointes | 288
    ventricular fibrillation | 288
    CPR | 288
    direct current cardioversion | 288
    return of spontaneous circulation | 288
    AF with high VE burden | 288
    persistent VE | 312
    AF | 312
    bradycardic episodes | 312
    noradrenaline requirement increased | 312
    atrial pacemaker insertion | 336
    AAI 90 bpm | 336
    cessation of VE | 432
    AF cessation | 432
    noradrenaline requirement reduction | 432
    decannulated from ECMO | 648
    secondary-prevention implantable cardioverter defibrillator | 864
    repatriated to local ICU | 1080
    sepsis | 1080
    death | 1080

<|eot_id|>