74 years old | 0
white | 0
female | 0
admitted to the hospital | 0
low-grade fever | -48
dry cough | -48
shortness of breath | -48
elective right total knee replacement | -168
post-operative course | -168
pain | 0
redness | 0
swelling | 0
essential hypertension | 0
obesity | 0
myasthenia gravis | 0
osteoarthritis | 0
body temperature | 0
blood pressure | 0
pulse | 0
respiratory rate | 0
oxygen saturation | 0
bilateral rhonchi | 0
rales | 0
patchy air space opacity | 0
pneumonia | 0
rapid nucleic acid amplification test | 0
nasopharyngeal swab | 0
broad-spectrum antibiotics | 0
cefepime | 0
levofloxacin | 0
supportive care | 0
supplemental oxygen | 0
mild diarrhea | 72
generalized weakness | 72
fatigue | 72
intravenous immunoglobulin | 72
mild MG exacerbation | 72
arterial blood gases | 0
complete blood count | 0
basic metabolic profile | 0
mild absolute lymphopenia | 0
anemia | 0
pH | 0
pCO2 | 0
pO2 | 0
bicarbonate | 0
creatinine kinase | 144
lactic acid | 144
lactate dehydrogenase | 144
ferritin | 144
interleukin-6 | 144
progressively increasing SOB | 24
oxygen requirements | 24
nasopharyngeal swab results | 96
SARS-CoV-2 | 96
hydroxychloroquine | 96
azithromycin | 96
zinc sulfate | 96
oral vitamin C | 96
blood and sputum cultures | 96
broad-spectrum antibiotics discontinued | 96
SOB worsened | 144
oxygen requirements | 144
drowsy | 144
moderate distress | 144
unable to protect airways | 144
blood pressure | 144
heart rate | 144
temperature | 144
respiratory rate | 144
bilateral alveolar infiltrates | 144
interstitial edema | 144
ARDS | 144
intubated | 144
mechanical ventilation | 144
norepinephrine | 144
septic shock | 144
colchicine | 144
cytokine storm | 144
high-dose vitamin C | 168
clinical condition improved | 192
norepinephrine support stopped | 192
CXR | 240
improvement of pneumonia | 240
interstitial edema | 240
spontaneous breathing trial | 240
CPAP/PS | 240
ABGs | 240
pH | 240
pCO2 | 240
pO2 | 240
bicarbonate | 240
extubated | 240
oxygen saturation | 384
CXR | 384
infiltrates | 384
interstitial edema | 384
discharged | 384
hydroxychloroquine treatment | 480
azithromycin treatment | 480
colchicine treatment | 192
high-dose vitamin C infusion | 480
oral zinc sulfate | 480
inpatient physical rehabilitation | 384
occupational rehabilitation | 384
quarantine | 384