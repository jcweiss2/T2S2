hepatitis C-related cirrhosis | 0 | 0 | Factual
recurrent hepatic encephalopathies | 0 | 0 | Factual
chronic portal vein thrombosis | 0 | 0 | Factual
liver transplantation | 0 | 0 | Factual
end-to-side anastomosis of the donor portal vein to the superior mesenteric vein | 0 | 0 | Factual
end-to-end bile duct anastomosis | 0 | 0 | Factual
massive venous bleeding from local varices | 0 | 0 | Factual
iliac conduit construction | 0 | 0 | Factual
normal liver graft function | 0 | 0 | Factual
stenosis of the bile duct anastomosis | -6720 | -3360 | Factual
biliary leakage | -6720 | -3360 | Factual
elevated liver enzymes | -6720 | -3360 | Factual
pigtail treatment | -3360 | -3360 | Factual
FCSCEMS insertion | -3024 | -3024 | Factual
persisting leakage | -3024 | -1680 | Factual
stent extraction | -1680 | -1680 | Factual
hepatitis C reinfection | -1680 | 0 | Factual
recurrent stenosis of the biliary anastomosis | -1680 | 0 | Factual
ERCP | -1680 | 0 | Factual
balloon dilatations | -1680 | 0 | Factual
pigtail placements | -1680 | 0 | Factual
stent placements | -1680 | 0 | Factual
biopsy-proven significant fibrosis | -8760 | -8760 | Factual
treatment with pegylated interferon and ribavirin | -8760 | -6720 | Factual
elective ERCP | 0 | 0 | Factual
portobiliary fistula | 0 | 0 | Factual
hemobilia | 0 | 0 | Factual
FCSEMS placement | 0 | 0 | Factual
prophylactic antibiotic treatment with ciprofloxacin | 0 | 0 | Factual
septic shock | 48 | 48 | Factual
admission to the intensive care unit | 48 | 48 | Factual
hemodynamic support | 48 | 48 | Factual
empiric broad-spectrum antibiotic treatment | 48 | 48 | Factual
computed tomography | 48 | 48 | Factual
angiography | 48 | 48 | Factual
chronic obliteration of the iliac conduit | 48 | 48 | Factual
partial perfusion of the hepatic artery by gastroduodenal collaterals | 48 | 48 | Factual
anuric kidney failure | 48 | 48 | Factual
continuous venovenous hemofiltration | 48 | 192 | Factual
intermittent hemodialysis | 192 | 672 | Factual
evaluation for liver re-transplantation | 4032 | 4032 | Factual
FCSEMS replacement | 4032 | 4032 | Factual
no evidence of persisting leakage | 4032 | 4032 | Factual
no relevant stenosis | 4032 | 4032 | Factual
no recurrent stenosis or portobiliary fistula | 4032 | 12000 | Factual