73 years old | 0
female | 0
hypertension | 0
syphilis | 0
type 2 diabetes mellitus | 0
admitted to the hospital | 0
altered mental status | 0
mechanical fall | -720
pruritic scalp | -720
purulent drainage from sinuses on the scalp | -720
temperature of 97.9°F | 0
heart rate of 127 bpm | 0
respiratory rate of 22 breaths/min | 0
blood pressure of 144/80 mmHg | 0
oxygen saturation of 98% on room air | 0
oriented to person and place, but not to time | 0
face, scalp and right ear were erythematous and edematous | 0
large fluctuant mass with purulent drainage over the occipital and parietal portions of the scalp | 0
posterior auricular mass without signs of active drainage | 0
hyperglycemia to 700 | 0
anion gap metabolic acidosis with serum bicarbonate of 20 | 0
ketonuria | 0
non-contrast head computed tomography (CT) | 0
extensive multifocal scalp swelling along the right temporal, right posterior parietal and left frontal regions | 0
no acute intracranial abnormalities | 0
diabetic ketoacidosis | 0
cellulitis of the scalp | 0
concern for underlying abscesses | 0
continuous infusion of insulin | 0
broad-spectrum coverage with intravenous Vancomycin and Cefepime | 0
incision and drainage of scalp lesion | 48
10-cm subgaleal abscess with large amounts of purulence evacuated | 48
initial admission blood cultures grew MRSA | 72
continued on intravenous Vancomycin and Cefepime | 72
paranasal sinus CT with intravenous contrast | 72
no involvement | 72
transesophageal echocardiogram | 72
no evidence for endocarditis | 72
pulse irrigation of the wounds and sharp debridement | 96
involvement of plastic surgery | 96
serial bedside debridements | 96
scalp wound measured 20 cm in length, 10 cm in width and 2 cm depth | 96
right posterior auricular wound measured 7 × 7 × 2 cm | 96
wounds of the scalp and post-auricular region were definitively closed with split-thickness skin grafts | 120
split-thickness skin grafts harvested from the right thigh | 120
100% take of the grafts | 168
discharged on hospital day 32 | 768
intravenous Vancomycin to complete a full 7-week course | 768