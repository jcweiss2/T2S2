8 years old | 0
female | 0
admitted for severe bilateral optic neuritis | 0
admitted for longitudinally extensive transverse myelitis (LETM) | 0
March 2008 | 0
3 infusions of methylprednisolone | 0
oral tapering steroids | 0
fully recovered | 0
five months later | 360
another LETM occurred | 360
presence of AQP4-Ab in serum | 360
diagnosis of NMOSD | 360
following 9 years | 79200
intensive immunosuppression by immunoadsorptions | 79200
intensive immunosuppression by plasma exchanges | 79200
mycophenolate mofetil | 79200
RTX | 79200
9 severe relapses | 79200
permanent visual disability | 79200
right amblyopia | 79200
visual acuity OD=0.1 | 79200
visual acuity OS=0.8 | 79200
Expanded Disability Status Scale=3 | 79200
RTX pediatric protocol | 79200
2 infusions with interval of 2 weeks | 79200
375 mg/m2 for each infusion | 79200
initially at each relapse | 79200
then every 6 months since 2013 | 79200
September 2014 | 11520
RTX infusion-related reaction | 11520
July 2015 | 17424
hospitalization in intensive care unit for anaphylactic-like reaction related to RTX | 17424
following infusions performed in intensive care unit | 17424
persistence of clinical activity | 17424
B-cells still detected despite RTX | 17424
severe sepsis related to central catheter infection | 17424
introduction of subcutaneous OFA in August 2017 | 19848
one injection of 20 mg every week for 4 weeks | 19848
one injection of 20 mg every 4 weeks | 19848
2018 | 21768
detection of antibodies against RTX | 21768
therapeutic change | 21768
2 years of follow-up | 35040
30 injections of OFA | 35040
no further relapse | 35040
November 2019 | 43392
clinical examination normal except visual disability | 43392
Expanded Disability Status Scale=3 | 43392
January 2019 | 40032
MRI revealed no radiologic activity | 40032
atrophy of optic nerves | 40032
persistent spinal cord lesion from C2 to T5 | 40032
perfect tolerance | 40032
no anaphylactic-like event | 40032
no infectious event | 40032
complete B-cell depletion | 40032
no lymphopenia | 40032
no hypogammaglobulinemia | 40032
