55 years old | 0
female | 0
RA | -7200
treated with prednisolone | -7200
treated with methotrexate | -7200
treated with etanercept | -7200
fever | -72
progressive fatigue | -2160
malaise | -2160
anorexia | -2160
oral bleeding | -2160
weight loss | -2160
admitted to the hospital | 0
body temperature 37.5 | 0
blood pressure 120/80 mmHg | 0
pulse rate 104 beats per minute | 0
respiratory rate 18 breaths per minute | 0
pale conjunctiva | 0
oral ulcer | 0
advanced multiple symmetrical joint deformities | 0
fine rales on both lower lung fields | 0
hemoglobin 7.7 g/dL | 0
platelet count 40,000/mm3 | 0
white blood cell count 3,000/mm3 | 0
liver function tests abnormal | 0
rheumatoid factor 2,180 IU/mL | 0
antimycoplasma antibodies negative | 0
anti-HIV antibodies negative | 0
poorly-defined nodular opacities in both lower lung zones | 0
enlarged lymph nodes in the para-aortic area | 0
dyspnea | 96
oxygen saturation dropped below 80% | 96
intubated | 96
transferred to the intensive care unit | 96
pulmonary hemorrhage suspected | 96
diffuse bilateral pulmonary consolidation | 96
diffuse consolidation and ground-glass attenuation | 96
small bilateral pleural effusions | 96
enlarged lymph nodes with central attenuation | 96
minimal pericardial effusion | 96
diffuse hypokinesia | 96
left ventricular ejection fraction 36% | 96
hypocellular marrow | 96
mucosal injection and fold thickening | 96
intravenous immunoglobulin | 96
solucortef | 96
azithromycin | 96
ceftriaxone | 96
amikacin | 96
meropenem | 240
ciprofloxacin | 240
condition improved | 960
chest radiograph showed complete resolution | 960
normal LV systolic function | 960
ejection fraction 70% | 960
without hypokinesia | 960
adenovirus positive | 960
discharged | 960
maintained oral medication | 960
prednisolone | 960
celecoxib | 960
hydroxychloroquine sulfate | 960
methotrexate | 960
without complications | 960
without aggravating arthralgia | 960