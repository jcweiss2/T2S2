54 years old | 0
female | 0
rheumatoid arthritis | 0
uncontrolled diabetes mellitus type II | 0
neuropathy | 0
hypothyroidism | 0
transferred | 0
acute idiopathic necrotizing pancreatitis | 0
multiple prior episodes of pancreatitis | -4320
sepsis | -4320
infected pseudocyst | -4320
requiring pressor support | -4320
acute respiratory distress syndrome | -4320
acute kidney injury | -4320
deep vein thrombosis | -4320
pulmonary embolism | -4320
requiring anticoagulation | -4320
retroperitoneal drainage catheter placed | -48
enlarging abscess | -48
no subcapsular hepatic hematoma | -48
normal hepatic parenchymal enhancement | -48
admitted to surgical intensive care unit | 0
critical condition | 0
stable condition | 0
anticoagulation therapy continued | 0
progressive abdominal pain | 24
low drain output | 24
imaging demonstrated appropriate drain position | 24
persistent collection | 24
tissue-plasminogen activator injected | 48
fresh blood in drainage catheter | 72
hypotensive | 72
decreased hemoglobin | 72
anemic baseline of 7.6 gm/dL | 72
hemoglobin decreased to 6.2 gm/dL | 72
platelet count within normal limits | 72
coagulation panel within normal limits | 72
liver enzymes within normal limits | 72
resuscitation | 72
crystalloid solution | 72
blood transfusions | 72
pressors not initiated | 72
unenhanced CT demonstrating hemoperitoneum | 72
heterogeneously hyperdense subcapsular collections | 72
perihepatic collections | 72
contrast-enhanced CT confirmed active hemorrhage | 72
active hemorrhage in gallbladder fossa | 72
active hemorrhage into perihepatic hematoma | 72
percutaneous endovascular embolization | 72
gelatin foam | 72
detachable coil | 72
transfusion of 5 units packed red blood cells | 72
transfusion of 2 units fresh frozen plasma | 72
transfusion of 400 mL albumin | 72
blood pressure stabilized | 72
hemoglobin stabilized | 72
remained in critical condition | 72
bedbound | 72
anticoagulation not restarted | 72
serum transaminases increased | 120
alkaline phosphatase increased | 120
bilirubin increased | 120
hemoglobin decreased from 8.4 gm/dL to 6.8 gm/dL | 120
follow-up contrast-enhanced CT | 120
increased size of hepatic subcapsular hematoma | 120
marked mass effect on liver | 120
new ill-defined hypoattenuation of liver parenchyma | 120
hepatic ischemia | 120
multiple punctate areas of contrast extravasation | 120
continued active bleeding | 120
hepatic angiography | 120
punctate areas of contrast blush | 120
cystic artery remained occluded | 120
no embolization performed | 120
anticoagulation remained discontinued | 120
blood products administered | 120
crystalloid resuscitation administered | 120
laboratory indicators worsened | 120
concern for developing liver failure | 168
surgical evaluation | 168
laparoscopy demonstrated inflammatory adhesions | 168
large organized hematoma | 168
hematoma could not be suctioned | 168
hematoma could not be morcellated | 168
hand port utilized | 168
diffuse oozing from liver parenchyma | 168
right subcostal incision | 168
hepatic subcapsular hematoma evacuated | 168
packs placed for hemostasis | 168
subhepatic hematoma evacuated | 168
cholecystectomy performed | 168
retroperitoneal necrosectomy performed | 168
feeding jejunostomy tube placed | 168
primary closure | 168
repeat laboratories showed improvement | 168
alkaline phosphatase improvement | 168
ALT improvement | 168
AST improvement | 168
bilirubin improvement | 168
no further bleeding events | 168
liver enzymes remained stable | 168
follow-up imaging 32 days after evacuation | 768
persistent areas of infarction | 768
follow-up imaging 5 months later | 3600
persistent wedge-shaped nonenhancement | 768
peripheral hepatic infarcts | 768
right portal vein restored | 768
protracted admission due to pancreatitis severity | 168
t-PA administration | 48
anticoagulants administration | 0
thrombolytics administration | 48
continued expansion of hematoma | 120
discontinuation of anticoagulation | 72
mass effect upon liver | 120
ischemia | 120
infarction | 120
peripheral hepatic parenchyma infarction | 120
narrowing of right portal vein | 120
decreased vascular inflow | 120
Page kidney-like mechanism | 120
increased pressure within capsule | 120
reduced arterial inflow | 120
coagulative necrosis due to pancreatic enzymes | 120
wedge-shaped infarction | 120
off-target embolization considered | 120
embolic material insufficient | 120
serial labs | 72
fluid resuscitation | 72
blood transfusions if indicated | 72
strict bed rest | 72
selective transcatheter embolization | 72
surgical control of bleeding | 168
electrocauterization | 168
hemostatic devices | 168
packing | 168
laparoscopy | 168
laparotomy | 168
extravasation from cystic artery | 72
embolized cystic artery | 72
weakened Glisson's capsule | 0
irritated hepatic surface | 0
pericapsular small arteries irritation | 0
hematoma formation | 0
exacerbated by anticoagulants | 0
exacerbated by thrombolytics | 48
active bleeding into subcapsular hematoma | 72
peripheral location of bleeding | 72
embolization not safely performed | 120
persistent contrast blushes | 120
mass effect worsened | 120
hepatic failure | 120
nonoperative management | 72
operative management | 168
persistent peri-hepatic bleeding | 120
