72 years old | 0
    male | 0
    weakness | -336
    fatigue | -336
    virtual consultation with general practitioner | -336
    conservative management | -336
    apprehensive about attending hospital | -336
    progressive dyspnea on exertion | -96
    limitation of physical activity | -96
    no chest pain | -96
    no palpitations | -96
    no ankle edema | -96
    increased urinary frequency | -96
    dark urine | -96
    no dysuria | -96
    no dysphagia | -96
    no bleeding per rectum | -96
    no abdominal pain | -96
    no weight loss | -96
    no fever | -96
    no rigors | -96
    no recent travel | -96
    admission | 0
    spike in temperature to 39.1°C | 0
    tachycardia 133 bpm | 0
    past medical history of benign prostatic hyperplasia | 0
    medication Dutasteride/tamsulosin 0.5/0.4 mg | 0
    physical examination: tachycardic | 0
    vital signs within normal range | 0
    no peripheral stigmata of cardiovascular disease | 0
    non-displaced apex beat | 0
    pansystolic murmur loudest at apex radiating into axilla | 0
    jugular venous pressure not raised | 0
    no peripheral edema | 0
    unremarkable respiratory examination | 0
    unremarkable gastrointestinal examination | 0
    unremarkable neurological examination | 0
    C-reactive protein 101 mg/L | 0
    high-sensitivity troponin T 500 ng/L | 0
    NT-proBNP 4337 pg/mL | 0
    ferritin 1498 ng/mL | 0
    electrocardiogram: sinus tachycardia with diffuse non-territorial ischemic changes | 0
    chest radiograph: ill-defined perihilar air-space opacities | 0
    transthoracic echocardiogram: dilated left ventricle | 0
    left ventricular internal diastolic dimension 6.9 cm | 0
    left ventricular ejection fraction 47% | 0
    thinned and akinetic inferior and inferoseptal walls | 0
    elevated LV filling pressure | 0
    moderate mitral regurgitation | 0
    elevated right ventricular systolic pressure >60 mmHg | 0
    electrocardiogram showing right ventricular strain pattern and S1Q3T3 | 0
    computed tomography pulmonary angiography (CTPA) performed | 0
    CTPA negative for pulmonary embolism | 0
    pulmonary edema | 0
    moderate bilateral pleural effusions | 0
    ground glass change | 0
    interlobular septal thickening | 0
    trace pericardial fluid | 0
    pericardial thickening | 0
    initial impression: systemic inflammatory response syndrome due to infectious process | 0
    investigated for COVID-19 | 0
    three nasal-pharyngeal swabs negative | 0
    differential diagnosis: heart failure of ischemic etiology | 0
    audible murmur | 0
    abnormal electrocardiogram | 0
    abnormal echocardiogram | 0
    elevated NT-proBNP | 0
    considered pulmonary embolism | 0
    admitted under general medical physician | 0
    cardiology team consulted on day 4 | 96
    infectious process ruled out | 96
    diagnostic coronary angiogram performed | 144
    occlusion of right coronary artery (RCA) at mid-vessel | 144
    collateralization from left coronary system | 144
    left coronary system free of significant disease | 144
    improved on intravenous diuretic therapy | 144
    reviewed by HF specialist team | 144
    institution of disease-modifying agents | 144
    discharged home | 168
    discharge diagnosis: ischemic HF with LV involvement due to RCA occlusion | 168
    prescription: Dutasteride/tamsulosin 0.5/0.4 mg | 168
    prescription: Pantoprazole 40 mg | 168
    prescription: Aspirin 75 mg | 168
    prescription: Clopidogrel 75 mg | 168
    prescription: Furosemide 40 mg | 168
    prescription: Atorvastatin 80 mg | 168
    prescription: Ramipril 2.5 mg | 168
    prescription: Bisoprolol 1.25 mg | 168
    plan for intensive medical management | 168
    discussed at heart team meeting regarding revascularization | 168
    case discussed with hospital heart team | 168
    consensus decision to proceed to cardiac magnetic resonance imaging (CMR) | 168
    CMR to assess viability of right coronary territory | 168
    re-presentation with NYHA class III symptoms | 600
    fatigue | 600
    night sweats | 600
    palpitations | 600
    treated with intravenous diuresis | 600
    repeat transthoracic echocardiogram: severe MR | 600
    restricted motion of posterior mitral valve leaflet | 600
    large LV saccular outpouching in basal inferior wall | 600
    CMR viability study performed | 648
    dilated LV with focal posterior saccular outpouching | 648
    aneurysmal segment dyskinetic with transmural late gadolinium enhancement | 648
    endocardial low signal consistent with thrombus | 648
    intact pericardium | 648
    organizing thrombus at base | 648
    saccular outpouching narrow neck compared to base | 648
    sudden progression from normal myocardium to attenuated layer | 648
    diagnosis of LV pseudoaneurysm (LVP) | 648
    LV ejection fraction 37% | 648
    severe secondary MR | 648
    tethered chordae | 648
    restricted motion of posterior mitral leaflet | 648
    assigned to bed rest | 648
    close monitoring in coronary care unit | 648
    findings discussed with patient and family | 648
    decision for surgical replacement of mitral valve and repair of LVP | 648
    intraoperative findings: severe ischemic MR | 816
    LV aneurysm 5x4 cm adherent to diaphragmatic pericardium | 816
    Perimount Magna Ease mitral valve placed | 816
    cuff of pericardium dissected | 816
    repair of pseudoaneurysm by direct closure | 816
    difficult postoperative course | 816
    26 days in intensive care | 816
    complications: arrhythmia | 816
    complications: cardiogenic shock | 816
    complications: ischemic sigmoid colitis | 816
    complications: bowel perforation | 816
    complications: sepsis | 816
    recuperated well | 816
    intensive rehabilitation | 816
    discharged home | 2472
    prescription: Atorvastatin 80 mg | 2472
    prescription: Bisoprolol 7.5 mg | 2472
    prescription: Furosemide 40 mg | 2472
    prescription: Aspirin 75 mg | 2472
    prescription: Apixaban 5 mg twice daily | 2472
    prescription: Pantoprazole 40 mg | 2472
    prescription: Ramipril 7.5 mg | 2472
    repeat echocardiogram: LV ejection fraction 26% | 2472
    akinetic inferior and inferolateral walls | 2472
    well-functioning mitral valve prosthesis | 2472
    no significant transvalvular or paravalvular regurgitation | 2472

    