44 years old|0
African-American|0
woman|0
presented to the Hematology/Oncology clinic|0
weakness|0
fatigue|0
HTLV associated T-cell lymphoma/leukemia|0
allogenic bone marrow transplant|0
disease relapse|0
graft failure|0
blood transfusion dependence|0
disseminated aspergillosis|0
skin involvement|0
lung involvement|0
oral posaconazole|0
high dose micafungin|0
left tunneled internal jugular catheter|0
oral acyclovir|0
oral levofloxacin|0
monthly inhaled pentamidine|0
hypotensive (83/57 mmHg)|0
tachycardic (117 bpm)|0
afebrile|0
non-tender ulceration|0
right distal leg|0
urchin diameter 2 cm|0
no erythema|0
no discharge|0
no induration|0
left internal jugular tunneled catheter|0
catheter exit site no erythema|0
catheter exit site no drainage|0
admitted to the intensive care unit|0
sepsis|0
blood cultures obtained from central line|0
blood cultures obtained from periphery|0
empirical treatment with cefepime|0
empirical treatment with vancomycin|0
leukopenia (2.0 K/uL)|0
absolute neutrophil count 0.04 K/uL|0
low hemoglobin (10.2 g/dL)|0
thrombocytopenia (25 K/uL)|0
high creatinine (1.24 mg/dL)|0
elevated transaminases (AST 505 U/L)|0
elevated transaminases (ALT 477 U/L)|0
chest computed tomography bilateral perihilar nodules|0
chest computed tomography pulmonary nodules|0
unchanged from previous images one month ago|0
hypotension worsened|0
norepinephrine infusion|24
antibiotic therapy escalated from cefepime to meropenem|24
vancomycin continued|24
transaminitis|24
intravenous isavuconazole substituted for posaconazole|24
intravenous micafungin continued|24
gram-positive rods in blood cultures|48
Cellulosimicrobium sp. identified by MALDI-TOF|48
in vitro susceptibility testing|48
benzyl penicillin MIC 0.012 ug/mL|48
levofloxacin MIC >32 ug/mL|48
vancomycin MIC 0.38 ug/mL|48
catheter related bloodstream infection|48
tunneled catheter removed|48
catheter tip grew Cellulosimicrobium sp.|48
clinical improvement|48
resolution of hypotension|48
resolution of acute renal failure|48
resolution of transaminitis|48
meropenem discontinued|48
oral levofloxacin resumed|48
repeat blood cultures negative|72
discharged|168
pneumonia|216
death|216
