69 years old | 0
male | 0
admitted to the hospital | 0
generalized abdominal pain | -192
multiple episodes of bilious vomiting | -192
obstipation | -96
diabetic | 0
chronic alcoholic | 0
tachycardia | 0
abdominal distension | 0
generalized tenderness | 0
leucocytosis | 0
ultrasonography | 0
prominent fluid filled small bowel loops | 0
sluggish peristalsis | 0
CECT of abdomen and pelvis | 0
large hyperdense calculus | 0
dilated small bowel loops | 0
gall bladder partially dilated | 0
suspicious fistulous communication | 0
multiple air foci | 0
Rigler's triad | 0
diagnosis of GI | 0
exploratory laparotomy | 24
gallstone impacted in ileum | 24
enterotomy | 24
cholecystoduodenal fistula | 24
subtotal cholecystectomy | 24
primary closure of duodenal fistula | 24
chronic cholecystitis | 48
reactive lymphadenitis | 48
full diet | 120
suture line healthy | 120
left abdominal drain removed | 192
right abdominal drain removed | 216
respiratory infection | 288
shock | 288
acute kidney injury | 288
intubated and ventilated | 288
blood transfusions | 288
intravenous antibiotics | 288
inotropic support | 288
electrolyte corrections | 288
pneumonia | 504
sepsis | 504
death | 504