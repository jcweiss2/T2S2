42 years old | 0
female | 0
admitted to the hospital | 0
dyspnea | -96
enduring cough | -96
influenza A (H1N1) | -96
oseltamivir | -96
blood pressure 90/60 mm Hg | 0
pulse rate 100 beats per minute | 0
respiratory rate 22 breaths per minute | 0
body temperature 36.3 | 0
oxygen saturation 93.3% | 0
coarse breathing sounds | 0
peribronchial consolidations | 0
multifocal ground glass opacities | 0
hypoxemia | 0
hemoglobin 13.8 g/dL | 0
white blood cell count 4640 cells/mm3 | 0
neutrophils 77.4% | 0
platelet count 161000 cells/mm3 | 0
C-reactive protein 30.24 mg/dL | 0
serum albumin 3.7 g/dL | 0
aspartate aminotransferase 35 U/L | 0
alanine aminotransferase 27 U/L | 0
total bilirubin 0.9 mg/dL | 0
serum creatinine 1.8 mg/dL | 0
tracheobronchial wall thickening | 0
multifocal patchy consolidations | 0
nodular opacities with cavitations | 0
severe mucosal inflammation | 0
sloughing | 0
diffuse cobblestone-like multiple mucus swelling of exudates | 0
partial obstruction of airways | 0
pseudomembranous tracheobronchitis | 0
respiratory failure | 24
mechanical ventilation | 24
Methicillin-sensitive Staphylococcus aureus | 24
tube thoracotomy | 48
bilateral pneumothoraces | 48
infected pneumatoceles | 48
colistin | 72
improvement of dyspnea | 1200
improvement of radiologic findings | 1200
pigtail catheter removal | 1200
follow-up bronchoscopy | 1080
discharged | 1248