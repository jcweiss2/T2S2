46 years old | 0
female | 0
breast implants | 0
thyroidectomy | 0
admitted to the hospital | 0
headache | 0
vomiting | 0
neurological deterioration | 0
hyposthenia of the left hemisome | 0
cerebral CT scan | 0
intraparenchymal hemorrhage | 0
rupture of an internal carotid artery aneurysm | 0
emergency evacuation of the haematoma | 0
clipping of the aneurysm | 0
transferred to the intensive care unit | 0
fever | -144
Escherichia coli urinary tract infection | -144
treated with gentamicin | -144
neutrophilic leukocytosis | -96
thrombocytopenia | -96
procalcitonin value of 1.15 ng/mL | -96
blood cultures revealed R. mannitolilytica and R. pickettii | -96
R. mannitolilytica susceptible to ciprofloxacin and trimethoprim-sulfamethoxazole | -96
R. pickettii susceptible to ciprofloxacin and trimethoprim-sulfamethoxazole | -96
fever persisted | -96
treated with ciprofloxacin | -96
additional blood cultures performed | -72
Candida parapsilosis | -72
R. pickettii | -72
R. mannitolilytica | -72
cultures of the removed central venous catheter negative | -72
transthoracic echocardiogram showed no signs of cardiac vegetations | -72
funduscopic examinations negative | -72
MRI showed thrombosis of the internal carotid artery | -72
anticoagulant therapy with enoxaparin | -72
clearance of candidemia | -48
trimethoprim-sulfamethoxazole added to the antimicrobial regimen | -48
antibiotic treatment discontinued | 0
R. pickettii and R. mannitolilytica bacteraemia relapsed | 168
treated with trimethoprim-sulfamethoxazole and ciprofloxacin | 168
cranioplasty surgery | 216
fever | 320
R. pickettii grown from blood cultures | 320
ciprofloxacin administered | 320
progressive clinical improvement | 320
transferred to a rehabilitation centre | 320
completed an eight-week therapy course | 448
no further relapse of Ralstonia infection | 720