18-year-old male|0
autoimmune cirrhosis|0
admitted to the hospital|0
diagnosed with autoimmune cirrhosis|-8760
listed for liver transplantation|0
massive variceal hemorrhage|0
ostium secundum|-17520
percutaneous Amplatzer|-17520
propranolol|0
azathioprine|0
vitamin E|0
multivitamin supply|0
leukopenia|0
anemia|0
thrombocytopenia|0
alkaline phosphatase elevation|0
total serum bilirubin elevation|0
direct bilirubin elevation|0
indirect bilirubin elevation|0
CHILD A score|0
MELD score 11|0
variceal banding|0
normal chest X-rays|0
desaturation during surgery|0
right superior lobar atelectasis|0
right inferior lobar atelectasis|0
positive pressure therapy|0
purulent tracheal secretions|0
clinical sepsis|120
intensive care unit admission|120
increased cholestasis|120
endoscopic retrograde cholangiopancreatography|120
biliary stenting|120
transesophageal echocardiography|120
persistent tracheal secretions|720
sputum cultures|720
Aspergillus spp. identification|720
thoracic CT scan|720
multiple lung nodes|720
tree-in-bud opacities|720
pulmonary Aspergillus|720
posaconazole|720
caspofungin|720
amphotericin B|720
aciclovir|720
left hemiplegia|720
severe headache|720
mental status changes|720
brain MRI|720
right frontal lesions|720
right parietal lesions|720
perilesional edema|720
brain biopsy|720
multiple organ failure|1152
death|1152
copper deposits in liver|0
aldehyde fuchsin study|0
periodic acid-Schiff study|0
periseptal copper deposits|0
focal intracanalicular cholestasis|0
Wilson's disease|0
Trucut liver biopsy|96
hepatocanalicular cholestasis|96
apoptotic hepatocytes|96
Kupffer cells with pigment|96
sinusoidal congestion|96
mild acute cellular rejection|96
Banff score 4/9|96
portal swelling|96
ductulitis|96
endotheliitis|96
cytomegalovirus negative|96
cerebral collection|1152
H&E staining|1152
PAS-D staining|1152
Ziehl-Neelsen staining|1152
Gram staining|1152
Gomori staining|1152
brain parenchyma edema|1152
necrosis|1152
neutrophil infiltration|1152
apoptotic cells|1152
Aspergillus hyphae|1152
necrotizing encephalitis|1152
measles|432
tachycardia|432
fever|432
altered state of consciousness|432
rapid neurological deterioration|1152
