85 years old | 0
    woman | 0
    arrived at the emergency room | 0
    cardiac arrest | 0
    cardiopulmonary resuscitation | 0
    spontaneous circulation | 0
    urinary tract infection | -720
    left pleuritic pain | -72
    cough | -72
    dementia | 0
    arterial hypertension | 0
    diabetes mellitus type II | 0
    depression | 0
    sedation effects | 0
    no brain reflexes | 0
    mydriatic pupils | 0
    leukocytosis | 0
    neutrophilia | 0
    type II myocardial infarction | 0
    right basal consolidation | 0
    septic shock of pulmonary origin | 0
    myocardial infarction | 0
    admitted to the intensive care unit | 0
    antibiotics | 0
    piperacillin 4.5 gr QID | 0
    clarithromycin 500 mg BID | 0
    vasopressor | 0
    norepinephrine | 0
    mechanical ventilator support | 0
    brain CT scan | 0
    diffuse brain edema | 0
    subfalcine herniation | 0
    transtentorial herniation | 0
    sedation withdrawal | 48
    Glasgow Coma Scale score of 3/15 | 48
    absence of brainstem reflexes | 48
    complete brain MRI scan | 72
    BOLD signal | 72
    DTI acquisitions | 72
    second cardiac arrest | 72
    unsuccessful cardiopulmonary resuscitation | 72
    deceased | 72
    DTT | 72
    disruption of ventral tegmental tracts | 72
    disruption of dorsal tegmental tracts | 72
    reduction in FA values | 72
    hyperconnected FC | 72
    anticorrelated brain regions | 72
    correlated brain regions | 72
    