64 years old | 0
    male | 0
    admitted to the hospital | 0
    general malaise | -72
    fever | -72
    chills | -72
    pronounced nuchal swelling on the left side | -72
    pronounced facial swelling on the left side | -72
    left-sided microtia | 0
    complete absence of meatus acusticus | 0
    diabetes mellitus type 2 | 0
    arterial hypertension | 0
    valsartan 160 mg/d | 0
    left-sided head-and-neck edema | 0
    herpetiform-grouped vesicles around the left ear | 0
    herpetiform-grouped vesicles on the nose | 0
    yellowish crusts | 0
    formation of bullae in the perioral region | 0
    leukocytosis | 0
    white blood cell count of 25.7 | 0
    thrombocytopenia of 64 Gpt/L | 0
    lowered hematocrit of 0.245 L/L | 0
    hemoglobin of 5.1 mmol/L | 0
    erythrocyte count of 2.5 Tpt/L | 0
    neutrophilia of 13.8 Gpt/L | 0
    lymphopenia of 11% | 0
    increased number of large unstained cells with 2 Gpt/L | 0
    C-reactive protein (CRP) of 333 mg/L | 0
    HIV tests negative | 0
    antibiotic treatment with sultamicillin | -24
    facial swelling worsened | 24
    diagnostic ultrasound | 24
    thoracic computerized tomography (CT) | 24
    diagnosis of impetiginized herpes zoster | 24
    antibiotic treatment changed to clindamycin | 24
    aciclovir 3 × 500 mg/d | 24
    pain management using metamizole sodium | 24
    minor clinical improvement | 48
    11% blasts in peripheral blood | 48
    bone marrow biopsy suggested | 48
    malodorous oozing | 72
    formation of bullae | 72
    increasing edema | 72
    firm infiltrates on left chin | 72
    firm infiltrates on left submandibular region | 72
    skin biopsies taken | 72
    histopathology nonspecific | 72
    putrid inflammation | 72
    vesicles dissemination suggesting zoster generalisatus | 72
    increased dosage of aciclovir to 10 mg/kg | 72
    pain sensations become worse | 72
    pregabalin started | 72
    certoparin sodium 3000 I.E. anti-Xa/d | 72
    CRP increased to >400 mg/L | 96
    leukocytosis of 28.4 Gpt/L | 96
    procalcitonin increased to 3.65 ng/mL | 96
    suspicion of septicemia | 96
    transferred to intensive care unit | 96
    central venous access by subclavian catheter | 96
    treatment with piperacillin | 96
    levofloxacin | 96
    acyclovir every 8 hours | 96
    prednisolone | 96
    developed doughy stool | 120
    antibiosis changed to vancomycin | 120
    stool samples for Clostridium difficile negative | 120
    reduction of vesiculation | 120
    reduction of edema | 120
    CT performed | 168
    bone marrow biopsy performed | 168
    atypical myelopoiesis | 168
    reduced atypical erythropoiesis | 168
    micromegakaryocytic megakaryopoiesis | 168
    10% of bone marrow blasts | 168
    myelodysplastic syndrome (MDS) | 168
    refractory anemia | 168
    blast excess II (RAEB II) | 168
    karyotype 46/XY | 168
    translocations t(2;12)(p13; q13) | 168
    translocations t(6;9)(p22;q34) | 168
    erythrocyte concentrates required | 168
    pain in right arm | 336
    erythematous skin surrounding subclavian catheter | 336
    catheter removed | 336
    microbial cultures of the tip negative | 336
    vena subclavia thrombosis | 336
    soft tissue hematoma | 336
    oozing of the scalp | 360
    oozing of the ear helix | 360
    Pseudomonas aeruginosa identified | 360
    intensified diuresis | 360
    progressive edema | 360
    cytoreductive treatment with azacitidine | 360
    anemia | 360
    thrombocytopenia | 360
    erythrocyte concentrates | 360
    thrombocyte concentrates | 360
    herpes zoster persisted | 360
    intravenous infusion of varicella immunoglobulin | 408
    anaphylactic shock | 408
    managed by intensive care | 408
    septic shock | 408
    died | 432