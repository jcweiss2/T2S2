76 years old | 0
male | 0
admitted to the hospital | 0
pancreatic adenocarcinoma | -672
metastasis to the liver | -672
diastolic heart failure | -672
atrial fibrillation | -672
coronary artery disease | -672
severe hyponatremia | 0
sodium level of 116 mmol/L | 0
x-ray findings consistent with pneumonia | 0
broad-spectrum antibiotics | 0
fluid for hyponatremia | 0
transferred to the intensive care unit | 0
jugular vein distention | 0
lower extremity pitting edema | 0
transthoracic echocardiogram | 0
normal left ventricular cavity size | 0
mildly reduced systolic function | 0
septal flattening | 0
left atrial enlargement | 0
suspected MV vegetation | 0
severe mitral regurgitation | 0
tricuspid regurgitation | 0
elevated RV systolic pressure | 0
type 2 and type 3 pulmonary arterial hypertension | 0
ill-defined thickening in the TV leaflets | 0
afebrile | 0
leukocytosis | 0
recent urethral instrumentation | -24
blood cultures | 0
infectious disease specialist | 0
transesophageal echocardiogram | 24
normal left ventricular size and function | 24
ejection fraction of 60%-65% | 24
normal RV size and function | 24
hypermobile interatrial septum | 24
no left atrial or left atrial appendage thrombus | 24
vegetations on the atrial aspect of MV leaflets | 24
severe mitral regurgitation | 24
systolic flow reversal in the pulmonary vein | 24
vegetation on the TV leaflet | 24
tricuspid regurgitation | 24
RVSP 47 mm Hg | 24
negative blood cultures | 96
polymerase chain reaction testing negative | 96
workup for antiphospholipid syndrome unremarkable | 96
discontinued apixaban | -672
recommended low molecular weight heparin or unfractionated heparin | 0
computed tomography imaging of the head | 0
discontinued broad-spectrum antibiotics | 0
started on enoxaparin | 48
expired | 168