29 years old | 0
male | 0
unresponsive | -120
out-of-hospital cardiac arrest | -120
cardiac pulmonary resuscitation | -120
admitted to the hospital | 0
VF | -120
defibrillator-delivered electrical shocks | -120
intubated | 0
ventilation/oxygenation | 0
return of spontaneous circulation | 0
sinus tachycardia | 0
no chest pain | 0
no palpitations | 0
no syncope | 0
no SCD prior to admission | 0
blood pressure 122/70 mmHg | 0
temperature 38.5 °C | 0
pulse 102 bpm | 0
respiratory 22 bpm | 0
moist rales | 0
normal physical examinations | 0
no history of previous disease | 0
no family history of SCD | 0
type 1 Brugada ECG pattern | 0
coved-type ST-segment elevations | 0
negative T-wave | 0
brother with type 2 Brugada ECG pattern | -672
amaurosis | -672
ECG changes | 0
induced-hypothermia protocol | 0
sedation | 0
analgesia | 0
continuous renal replacement therapy | 0
Linezolid injection | 0
Sulperazon injection | 0
Mycamine injection | 0
correcting water-electrolyte and acid-base balance | 0
nutritional support | 0
protecting hepatorenal function | 0
tracheotomy | 480
no further episodes of VT/VF | 480
various ECG changes | 480
refused ICD | 480
brother received Reveal LINQ Insertable Cardiac Monitor | 480
recommended genetic testing | 480
no arrhythmia episodes after discharge | 2592
good physical condition | 2592
normal sinus rhythm | 2592
remote monitoring | 2592
no ventricular arrhythmia | 2592
pulmonary infection | 0
sepsis | 0
multiple organ dysfunction syndrome | 0
hypoxic ischemic encephalopathy | 0
elevated creatine kinase | 0
elevated CK-MB | 0
elevated urea | 0
elevated creatinine | 0
elevated serum alanine transaminase | 0
elevated aspartate aminotransferase | 0
elevated total bilirubin | 0
elevated direct bilirubin | 0
elevated procalcitonin | 0
elevated D-dimer | 0
elevated fibrinogen degradation products | 0
elevated activated partial thromboplastin time | 0
elevated brain natriuretic peptides | 0
normal electrolytes | 0
echocardiography revealed no structural disease | 0
chest radiography revealed pulmonary infection | 0
head computed tomography did not reveal infarction or hemorrhage | 0
fever | -120
treated with antipyretics | 0
education and lifestyle measures | 0
CPR | -120