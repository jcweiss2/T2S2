developed pancytopenia | -504
received broad anti-infective treatment | -504
developed tachycardia | -72
developed hypotension | -72
developed lactic acidosis | -72
admitted to pediatric intensive care unit | 0
transthoracic echocardiography revealed severely impaired left ventricular ejection fraction | 0
electrocardiogram showed sinus tachycardia with incomplete right bundle branch block | 0
NT-proBNP was 19 384 pg/ml | 0
high-sensitive troponin T was 53.7 pg/ml | 0
fluid therapy was started | 0
noradrenaline was started | 0
dobutamine was started | 0
milrinone was started | 0
deep sedation was initiated | 0
mechanical ventilation was initiated | 0
lactate acidosis worsened | 12
va-ECMO was initiated | 12
va-ECMO blood flow was 3.3 l/min | 12
mean arterial pressure was 45 torr | 12
noradrenaline was administered at 80 µg/min | 12
vasopressin was administered at 2 units/h | 12
levosimendan was administered at 0.5 mg/h | 12
hydrocortisone was administered at 200 mg/d | 12
CVVHDF was started | 12
anti-infective therapy was continued | 12
linezolid was replaced by vancomycin | 12
PCT was 2.37 ng/ml | 12
CRP was 2.98 mg/dl | 24
mean arterial blood pressure declined to 40 torr | 24
LVEF further decreased below 10% | 24
levosimendan infusion was stopped | 24
acute ischemic injury of non-cannulated leg developed | 24
right femoral artery was dissected | 24
Dacron conduit was sewed on right femoral artery | 24
second arterial cannula was introduced | 24
ECBF was enhanced to 4-5 l/min | 24
MAP was maintained at 40-50 torr | 24
PCT levels rose to 42.5 ng/ml | 48
Hickman catheter was explanted | 48
broad-complex tachycardia occurred | 48
esmolol was administered | 48
metoprolol was administered | 48
left ventricular function further decreased | 48
aortic valve ceased to open | 48
second venous cannula was placed into left atrium | 48
ECBF reached 5-6 l/min | 48
lactate levels peaked at 29 mmol/l | 48
lactate levels fell | 72
MAP rose from 30 torr | 72
cerebral oximetry showed sufficient regional oxygen saturation | 72
left ventricle was unloaded | 72
therapeutic anticoagulation was ensured | 72
PCT peaked with 80.4 ng/ml | 72
CRP peaked with 7.23 mg/dl | 72
leukocytes remained low at 300/µl | 72
high-sensitive troponin T increased to 343 pg/ml | 72
creatine kinase MB increased to 178 U/l | 72
all microbial specimens collected remained negative | 72
viral myocarditis was excluded | 72
cardiac systolic function gradually recovered | 120
ECMO cannulas in left femoral vessels were removed | 120
ECMO was completely removed | 168
LVEF had recovered to approximately 30% | 168
mean arterial pressures were 60-70 torr | 168
CVVHDF could be stopped | 168
leucocyte count recovered to 1000/µl | 312
normal values were reached spontaneously | 720
respirator weaning was reached | 792
allogenic stem cell transplantation was performed | 1008
patient was discharged to rehabilitation facility | 1344
LVEF recovered to approximately 40% | 1344