45 years old| 0
male | 0
admitted to the emergency department | -216
cough | -216
sore throat | -216
oxygen saturation 88% | -216
heart rate 104 beats per minute | -216
blood pressure 105/75 mmHg | -216
temperature 38.5 °C | -216
SARS-CoV-2 infection positive | -216
COVID-19 pneumonia | -216
antiviral (favipiravir) | -216
dexamethasone | -216
LMWH (enoxaparin) | -216
oxygen support 3/L | -216
d-dimer level 660 μg/L | -216
oxygen support decreased | -216
antiviral treatment completed | -216
discharged | -168
left upper quadrant pain | 0
left flank pain | 0
mild tenderness in left upper quadrant | 0
no peritonitis findings | 0
leukocytosis 17.2 × 10∧3/μL | 0
d-dimer 310 μg/L | 0
troponin 0.001 | 0
splenic hypodense area on abdominal CT | 0
thoracic CT ground-glass opacities | 0
oral intake stopped | 0
intravenous hydration | 0
nonopioid analgesics | 0
enoxaparin dose increased | 0
sudden onset chest pain | 24
ST segment elevation | 24
acute inferior MI | 24
consultation with cardiologists | 24
no cardiac thrombus | 24
emergency coronary angiography | 24
RCA stent placement | 24
coronary intensive care unit admission | 24
haemodynamically stable | 24
transferred to general surgery clinic | 24
regressive abdominal pain | 48
insignificant analgesics | 48
oral intake increased | 48
epigastric tenderness regressed | 48
left hypochondrial tenderness regressed | 48
discharged | 48
acetylsalicylic acid | 48
ticagrelor | 48
lupus anticoagulant negative | 48
antiphospholipid syndrome negative | 48
normal spleen on ultrasonography | 216
no intra-abdominal fluid | 216
no abscess collection | 216
meningococcal vaccine not needed | 216
Haemophilus influenza vaccine not needed | 216
follow-up imaging not indicated | 216
