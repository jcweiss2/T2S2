46 years old | 0
male | 0
ulcerative colitis | 0
malaise | -72
fever | -72
loss of appetite | -72
admission | 0
blood pressure 124/46 mmHg | 0
heart rate 122 beats per min | 0
SpO2 98% | 0
respiratory rate 16/min | 0
body temperature 40.2°C | 0
alert | 0
chills | 0
nausea | 0
cardiac arrest | 0
chest compression | 0
tracheal intubation | 0
ventricular fibrillation | 0
defibrillation | 0
adrenaline | 0
Brugada syndrome | 0
coved-type ST elevation in V1 and V2 | 0
fever subsided | 0
acetaminophen | 0
hypercalcemia | 0
hypotension | 12
septic shock | 12
ulcerative colitis exacerbation | 12
tazobactam-piperacillin | 12
vasopressors | 12
extubation | 48
fever reoccurred | 120
liver abscess | 120
meropenem | 120
vancomycin | 120
puncture drainage | 120
infection controlled | 720
pilsicainide test | 720
implantable cardioverter defibrillator | 720
discharged | 720
sudden death | -8760
high parathyroid hormone levels | 720
abnormal uptake in the anterior mediastinum | 720
tumor resection | 720
ectopic parathyroid adenoma | 720
nonfunctional pituitary adenomas | 720
nonfunctional adrenal tumors | 720
multiple endocrine neoplasia type 1 | 720