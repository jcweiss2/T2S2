35 years old | 0
male | 0
common variable immune deficiency (CVID) | -6720
monthly maintenance intravenous immunoglobulin (IVIG) infusions | -6720
fever | -744
headache | -744
shortness of breath | -744
asthma | -10080
hypertension | -10080
depression | -10080
swam in the Tennessee River | -1008
smoked 1.5 packs of cigarettes per day | -10080
consumed alcohol | -10080
smoked marijuana | -10080
son had CVID | -10080
construction worker | -10080
disabled | -10080
admitted to the hospital | 0
febrile | 0
tachycardic | 0
left maxillary sinus tenderness | 0
White blood cell (WBC) count 1.0 × 10−3/μL | 0
neutrophils 36% | 0
lymphocytes 50% | 0
monocytes 14% | 0
hemoglobin (Hb) 9.4 g/dL | 0
platelets 53 × 10−3/μL | 0
serum electrolytes normal | 0
renal function tests normal | 0
liver function tests normal | 0
Chest X-ray chronic blunting of right costo-phrenic angle | 0
Chest X-ray clear lung fields | 0
Chest X-ray normal cardiac silhouette | 0
Computed tomography (CT) of the paranasal sinuses pan sinus mucosal thickening | 0
intravenous vancomycin | 0
ceftazidime | 0
levofloxacin | 0
blood cultures negative | 0
urinalysis normal | 0
tick-borne panel negative | 0
Cytomegalovirus polymerase chain reaction (CMV-PCR) negative | 0
monospot negative | 0
bone marrow biopsy pancytopenia | 0
bone marrow biopsy no blasts | 0
bone marrow biopsy no organisms | 0
micafungin | 120
transferred to our facility | 120
dyspneic | 120
temperature 39.4 °C | 120
heart rate 118/min | 120
oxygen saturation (SpO2) 93% | 120
nasal oxygen at 11 L/min | 120
massive splenomegaly | 120
bilateral crackles in lower lung fields | 120
no rash | 120
no lymphadenopathy | 120
no meningeal signs | 120
no focal neurologic deficits | 120
WBC 1.94 × 10−3/μL | 120
neutrophils 48% | 120
lymphocytes 36.6% | 120
monocytes 14.4% | 120
basophils 0.5% | 120
Hb 9.8 g/dL | 120
platelets 51 × 10−3/μL | 120
prothrombin time 18.4 s | 120
serum electrolytes normal | 120
renal function tests normal | 120
serum aspartate aminotransferase (AST) 60 U/L | 120
total protein 5.0 g/dL | 120
albumin 2.5 g/dL | 120
liver function tests normal | 120
C-reactive protein elevated | 120
plasma procalcitonin elevated | 120
lactate dehydrogenase (LDH) 476 U/L | 120
serum ferritin 3016 ng/mL | 120
blood smear atypical lymphocytes | 120
blood smear pancytopenia | 120
blood smear toxic granulation of neutrophils | 120
Chest x-ray linear reticular opacities | 120
Chest x-ray opacities extending from hila to periphery | 120
CT chest extensive bilateral confluent alveolar opacities | 120
CT chest sub pleural sparing | 120
CT chest moderate left pleural effusion | 120
CT chest small right pleural effusion | 120
CT chest multiple pre- and para-tracheal lymph nodes | 120
CT chest massive splenomegaly | 120
blood cultures (bacterial, acid fast bacilli and fungal) sent | 120
Human Immunodeficiency Virus (HIV) 1,2 antigen-antibody negative | 120
urine Legionella antigen negative | 120
urinalysis normal | 120
serum beta-d-glucan sent | 120
cryptococcal antigen sent | 120
serum and urine for Histoplasma and Blastomyces antigens sent | 120
intravenous vancomycin | 120
piperacillin-tazobactam | 120
doxycycline | 120
transfer to intensive care unit | 144
empiric liposomal amphotericin B | 144
lumbar puncture | 144
cerebrospinal fluid analysis normal | 144
nasal endoscopic exam | 144
no invasive fungal disease | 144
serum beta-D glucan elevated | 168
Histoplasma antigen in serum positive | 168
Histoplasma antigen in urine positive | 168
afebrile | 192
hypoxemia improved | 192
switched to oral itraconazole | 288
discharged home | 288
fungal blood cultures grew Histoplasma capsulatum | 456
clinically improved | 1440
blood cell counts improved | 1440
itraconazole levels adequate | 1440
splenomegaly resolved | 2160
gained weight | 2880
symptom free | 2880
urine Histoplasma antigen negative | 4320
itraconazole stopped | 4320