22 years old | 0
female | 0
headache | -48
neck pain | -48
vomiting | -48
diarrhea | -48
abdominal pain | -48
photophobia | -48
malaise | -48
Pfizer vaccine second dose | -48
no history of COVID-19 infection | 0
tachycardic | 0
pyrexial | 0
normal blood pressure | 0
suspected meningitis | 0
ceftriaxone | 0
acyclovir | 0
CSF sampling unremarkable | 0
persistent fever over 40°C | 72
tachycardia | 72
severe hypoxia | 72
lactatemia | 72
hypotension | 72
unresponsive to IV fluids | 72
admitted to ITU | 72
high-flow nasal oxygen | 72
vasopressors | 72
fatigued | 72
intubated | 72
ventilated | 72
hypotension (cardiovascular) | 90
hypoxia (respiratory) | 90
azotemia | 90
oliguria | 90
nonabsorption of feeds | 90
diarrhea (GI) | 90
focused intensive care echocardiogram showed well filled but poorly contracting right and left ventricles | 90
commenced on dobutamine | 90
renal dysfunction | 90
severe metabolic acidosis | 90
progressive severe hyperpyrexia | 90
commenced on hemofiltration | 90
CT chest/abdomen | 90
multiple enlarged mesenteric lymph nodes | 90
moribund | 90
diagnostic laparoscopy | 90
multiple mesenteric lymph node enlargement | 90
minimal ascites | 90
small left ovarian cyst | 90
lymph node biopsy | 90
ascitic sampling | 90
no source of sepsis | 90
all microbiological sampling negative | 90
ciprofloxacin | 90
vancomycin | 90
meropenem | 90
no clinical improvement | 90
diagnosis of MIS-A | 90
IV immunoglobulin | 90
methylprednisolone daily for 5 days | 90
resolution of hyperpyrexia | 126
resolution of cardiovascular instability | 126
decreasing oxygen requirements | 126
extubated | 168
repeat echo showed normal ventricular function | 168
full recovery | 312
discharged home | 312
raised white cell count | 0
CRP 349 mg/L | 0
CSF clear appearance | 0
no cells detected | 0
Gram stain negative | 0
no organisms in culture | 0
chest X-ray no acute findings | 0
CT head no acute pathology | 0
CT abdomen and pelvis Day 3 postadmission showed significant mesenteric lymphadenopathy | 72
all body fluid and blood cultures negative | 0
CMV and EBV IgG and IgM positive | 0
vasculitis and autoimmune screen negative | 0
transthoracic echocardiogram no evidence of vegetation | 0
biventricular dysfunction | 0
lymph node biopsy suggestive of marked suppurative inflammation | 0
acute vasculitic changes | 0
three negative SARS-CoV-2 PCR tests | 0
COVID-19 antibodies positive | 0
macrophage activation syndrome considered | 0
mildly elevated ferritin | 0
no hypofibrinogenemia | 0
no cytopenias in more than two lineages | 0
