newborn female | 0
born at 24 weeks + 3 days | 0
breech presentation | 0
cord prolapse | 0
birth weight of 645 g | 0
HIV negative mother | 0
Apgar score of 4 | 0
Apgar score of 8 | 5
mechanical ventilation | 0
central umbilical catheters | 0
total parenteral nutrition | 0
empiric antibiotics | 0
skin sensors | 0
late-onset sepsis | 216
Escherichia coli bacteremia | 216
antimicrobial therapy with cefepime | 216
adhesive patch removal | 480
skin abrasion | 480
erythema | 480
induration | 480
plaque with necrotic center | 480
ulcer | 528
subcutaneous cell tissue | 528
necrotic area | 528
intensive treatment by wound care team | 480
healings | 480
hydrating dermal wound dressings | 480
sodium alginate | 480
carboxymethylcellulose | 480
hydrocolloids | 480
thermic instability | 528
metabolic acidosis | 528
hyperglycemia | 528
hypotension | 528
clinical deterioration | 528
cutaneous mucormicosis | 528
skin biopsy | 528
empiric antifungal treatment | 528
liposomal amphotericin B | 528
fungal biomarkers | 528
serum galactomannan | 528
1,3 beta-D-glucan | 528
refractory shock | 552
renal failure | 552
death | 564
fungal cultures | 528
Rhizopus spp. | 528
histopathology | 528
broad aseptate hyphae | 528
right angle branching | 528
Mucorales | 528
mass spectroscopy | 528
MALDI-TOF MS | 528
polymerase chain reaction | 528
PCR | 528
Rhizopus arrhizus | 528
fungal blood cultures | 528 
R. arrhizus | 528 
R. oryzae | 528 
Mucor | 528 
Lichtheimia | 528 
Absidia | 528 
R. microsporus | 528 
Lichtheimia corymbifera | 528 
Absidia corymbifera | 528 
necrotizing cellulitis | 528 
cutaneous aspergillosis | 528 
hyalohyphomycosis | 528 
Fusarium | 528 
necrotizing fasciitis | 528 
clostridial gas gangrene | 528 
sepsis-associated purpura fulminans | 528 
bacterial cellulitis | 528 
pyoderma gangrenosum | 528 
surgical debridement | 528 
anti-fungal treatment | 528 
L-AmB | 528 
ischemic necrosis | 528 
leukocytes | 528 
anti-fungal agents | 528 
tissue necrosis | 528 
cellulitis | 528 
ulcer | 528 
necrotic eschar | 528 
skin abscesses | 528 
gangrenous form | 528 
superficial infection | 528 
vesicle | 528 
pustule | 528 
erythematous plaque | 528 
necrotic plaque | 528 
papule | 528 
infection control | 528 
aggressive approach | 528 
diagnostic methods | 528 
microbiology | 528 
histopathology | 528 
mass spectrometry | 528 
molecular studies | 528 
etiological diagnosis | 528 
informed consent | 0 
Institutional Ethics Committee | 0 
Clínica Universitaria Bolivariana | 0 
Universidad Pontificia Bolivariana | 0 
Álvaro Hoyos | 0 
María Adelaida Mejía | 0 
Verónica Herrera | 0 
Andrés Soto | 0 
Clara Rico | 0 
Alejandro Díaz-Díaz | 0