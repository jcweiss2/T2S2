18 years old | 0
male | 0
admitted to the hospital | 0
ulcerative colitis | -9
infliximab | -9
infliximab | -22
acute respiratory deterioration | 0
septic shock | 0
moderate acute respiratory distress syndrome | 0
acute kidney failure | 0
invasive ventilation | 0
renal replacement therapy | 0
septic cardiomyopathy | 0
reduced systolic left ventricular function | 0
reduced systolic right ventricular function | 0
left ventricular ejection fraction <15% | 0
venoarterial extracorporeal membrane oxygenation | 24
percutaneous approach | 24
multistage cannula | 24
arterial cannula | 24
distal limb perfusion | 24
microaxial left ventricular assist device | 48
ejection fraction improved | 72
progressive colitis | 72
pancolitis | 72
gastrointestinal bleeding | 72
subtotal colectomy | 96
revision surgeries | 168
packing | 168
depacking | 168
recurrent intra-abdominal bleeding | 168
heart function recovered | 264
perfusion recovered | 264
transaminase levels decreased | 264
ECMELLA support removed | 264
transferred to general ward | 936
discharged | 1464
topical corticosteroids | 1464
improved general condition | 1824