4 years old | 0
male | 0
admitted to the hospital | 0
headaches | -48
vomiting | -48
tonic-clonic seizure | -48
subacute hydrocephalus | 0
COVID-19 positive | 0
asymptomatic | 0
external ventricular drain (EVD) placed | 0
noncontrast computed tomography (CT) of the brain | 0
satisfactory catheter placement | 0
interval reduction in ventriculomegaly | 0
magnetic resonance imaging (MRI) of the brain | 0
membrane obstructing the right foramen of Monro | 0
congenital malformation | 0
hydrocephalus | 0
magnetic resonance venography | 24
cervical spine MRI | 24
new left-sided hemiparesis | 72
repeat MRI | 72
magnetic resonance angiography (MRA) | 72
new diffusion restriction indicative of infarctions | 72
vasculitis or vasospasm | 72
stroke workup initiated | 72
echocardiography | 72
coagulopathy workup | 72
D-dimer levels | 72
protein S level | 72
homozygous 4G/4G for the plasminogen activator inhibitor type 1 (PAI-1) gene | 72
cerebrospinal fluid (CSF) infectious studies | 72
empirical treatment with exogenous steroids | 72
intracranial pressure monitoring | 72
ventricular endoscopy | 120
membranous obstruction at the right foramen of Monro | 120
septum pellucidotomy | 120
external CSF drainage continued | 120
surveillance MRI/MRA | 168
interval resolution of vascular findings | 168
discharged | 240