41 years old|0
male|0
chronic hepatitis C infection|-8760
IV drug use|-8760
smoking 15 cigarettes per day for the past 10 years|-8760
no current illicit drug abuse|-8760
altered mental status|0
fever|0
diffuse myalgia|0
flu-like symptoms|-120
fever|-120
muscle pain|-120
severe fatigue|-120
presyncopal event|0
intubated|0
mechanical ventilation|0
no nausea|-8760
no vomiting|-8760
no diarrhea|-8760
no skin rashes|-8760
blood pressure 144/95 mmHg|0
heart rate 130 beats/minute|0
oral temperature 101.9°F|0
respiratory rate 18 breaths/minute|0
oxygen saturation 97% on room air|0
AMS|0
toxic appearance|0
moderate distress|0
normocephalic head|0
atraumatic head|0
no palpable masses|0
no visible masses|0
poor dentition|0
no lymphadenopathy|0
no jugular venous distention|0
no carotid bruits|0
tachycardia|0
normal S1|0
normal S2|0
no murmurs|0
no thrills|0
clear breath sounds|0
symmetric breath sounds|0
no crackles|0
no wheezes|0
no rhonchi|0
soft abdomen|0
non-distended abdomen|0
non-tender abdomen|0
normal bowel sounds|0
no organomegaly|0
good skin turgor|0
mild cyanosis|0
no rashes|0
no lesions|0
no lower-extremity edema|0
radial pulses 3+|0
posterior tibial pulses 3+|0
dorsalis pedis pulses 3+|0
Glasgow coma score 8|0
sinus tachycardia|0
ventricular rate 115|0
normal axis|0
PR duration 138 milliseconds|0
no ST abnormalities|0
no T wave abnormalities|0
no acute chest X-ray abnormalities|0
normal CT head scan|0
white blood cell count 18 600/mm³|0
hemoglobin 14.1 g/dL|0
platelet count 50 000/mm³|0
CRP 24.3 MG/DL|0
lactic acid 3.1 mmol/L|0
normal chemistry panel|0
normal renal function|0
normal liver function|0
normal electrolytes|0
blood cultures sent|0
intravenous ceftriaxone|0
intravenous vancomycin|0
initial diagnosis meningitis|0
lumbar puncture not done|0
admitted to intensive care unit|0
extubated|24
encephalopathy improved|24
mechanical ventilation weaning trials|24
blood cultures grew MSSA|24
no skin wounds|24
no lacerations|24
no oral lesions|24
TTE performed|24
normal ejection fraction|24
no valvular heart disease|24
no vegetations|24
repeat blood cultures|168
blood cultures continued to grow MSSA|168
CT chest bilateral diffuse alveolar disease|168
septic emboli|168
bilateral pleural effusions|168
worsening respiratory distress|168
repeat TTE performed|168
no vegetations|168
no valvular heart disease|168
TEE performed|216
moderate mitral regurgitation|216
30×30 mm vegetation|216
consultation with cardiothoracic surgery|216
mitral valve replacement|504
intraoperative findings|504
resection of abscess|504
blood cultures no growth after 7 days|168
mental status improved|504
clinical status improved|504
discharged|600
