69 years old | 0
male | 0
ischaemic heart disease | 0
chronic liver disease | 0
adrenal incidentaloma | 0
arterial hypertension | 0
diabetes mellitus type 2 | 0
hyperuricaemia | 0
dyslipidaemia | 0
bacteraemia | -720
ESBL-producing Escherichia coli | -720
Klebsiella pneumoniae | -720
fever | 0
dyspnoea | 0
dizziness | 0
diffuse abdominal pain | 0
elevated plasma C-reactive protein | 0
elevated plasma procalcitonin | 0
negative blood culture | 0
heterogeneous liver | 0
cholelithiasis | 0
laparoscopic cholecystectomy | 24
hepatic lesions | 24
calcified biliary hamartomas | 24
K. pneumoniae in sample | 24
discharged | 168
bacteraemia | 720
ESBL-producing K. pneumoniae | 720
abdominal contrast-enhanced CT scan | 720
liver with increased dimensions | 720
heterogeneous texture | 720
multiple calcified lesions | 720
granulomas | 720
hypodense area | 720
MRI | 744
nodular lesions | 744
probable calcifications | 744
morphological alteration of liver | 744
hypertrophy | 744
chronic hepatopathy | 744
hepatobiliary scintigraphy | 744
normal appearance of bile ducts | 744
no obstruction | 744
multidisciplinary meeting | 744
hypothesis of liver transplant | 744
ruled out | 744
meropenem | 768
amikacin | 768
piperacillin and tazobactam | 768
ceftriaxone | 768
favourable clinical evolution | 896
discharged | 1344
sepsis | 2016
bacteriaemia | 2016
ESBL-producing K. pneumoniae | 2016
extended cycle of antibiotic therapy | 2016
meropenem | 2016
discharged | 2176
prophylactic antibiotics | 2176
ciprofloxacin | 2176
annual MRI | 2176
no relapse | 8760
no symptoms | 8760
prophylactic antibiotic | 8760
ciprofloxacin | 8760
annual MRI | 8760