57 years old | 0
male | 0
admitted to the hospital | 0
fever | -168
cough | -168
ischaemic stroke | -1820
patent foramen ovale | -1820
percutaneous closure | -1820
febrile | 0
cough | 0
dyspnoea | 0
mild oxygen desaturation | 0
sinus tachycardia | 0
bilateral lung crackles | 0
no murmur | 0
no sign of heart failure | 0
nasopharyngeal swab tested positive for SARS-CoV-2 | 0
hydroxychloroquine therapy | 0
antiviral agents therapy | 0
worsening hypoxaemia | 72
ARDS | 72
mechanical ventilation | 72
paroxysmal atrial fibrillation | 240
low molecular weight heparin therapy | 240
new onset of worsening fever | 336
haemoculture tested positive for MRSA | 336
TTE performed | 336
mild mitral regurgitation | 336
mild impairment of left ventricular systolic function | 336
TOE performed | 480
endocarditis vegetation on the aortic valve | 480
mild eccentric aortic valve regurgitation | 480
ventilator-associated pneumonia | 480
Klebsiella pneumoniae infection | 480
teicoplanin therapy | 480
ceftazidime/avibactam therapy | 480
linezolid therapy | 504
fosfomycin therapy | 528
improvement of clinical status | 528
reduction of inflammatory markers | 528
discharged from ICU | 720
transferred to Sub-ICU | 720
transferred to rehabilitation hospital | 888
TTE performed | 1104
smaller vegetation | 1104
no sign of significant regurgitation | 1104
new TTE scheduled | 1440