44 years old | 0
female | 0
Kuwaiti | 0
HER-2/Neu + score of +3 | 0
infiltrating ductal carcinoma of the right breast | 0
admitted to the hospital | 0
hyporesponsive | 0
tachycardic | 0
hypotensive | 0
temperature of 101.8°F | 0
mechanically ventilated | 0
multiple rounds of chemotherapy | -720
radiation | -720
craniotomy for resection of a tumor | -720
increased intracranial pressure (ICP) | -48
aspiration pneumonia | -48
intubation | -48
meropenem | 0
presumed pneumonia | 0
possible meningitis | 0
septic shock | 0
magnetic resonance imaging of the brain | 0
mild hydrocephalus | 0
large enhancing cavitary lesion in the right hemisphere | 0
craniotomy | 72
ventricular drain | 72
elevated ICP | 72
Epidural and intracavitary swabs | 72
CSF cultures | 72
heavy growth of Enterococcus faecalis | 72
vancomycin | 72
nonresponsive | 72
no use of analgesics or sedatives | 72
ampicillin plus gentamicin | 120
all subsequent CSF cultures remained positive | 120
tried to open her eyes | 240
regain her strength on the right side | 240
extubated | 288
verbally communicate | 288
intraventricular vancomycin | 432
vancomycin administered intraventricularly via the ventriculostomy drain | 432
normal-sized ventricles | 432
CSF drainage frequently remained less than 50 mL/d | 432
vancomycin of 10 mg administered intraventricularly every 3 days | 432
intraventricular vancomycin administered on August 27 | 432
intraventricular vancomycin administered on August 30 | 456
intraventricular vancomycin administered on September 3 | 480
first CSF culture returned negative | 504
subsequent cultures remained negative | 504
restart chemotherapy | 720
infection free | 4320
physical therapy | 4320
positive improvements | 4320