47 years old | 0
    female | 0
    referred to hospital for postoperative bleeding | 0
    postoperative bleeding following vaginal hysterectomy | -72
    vaginal hysterectomy | -96
    third-degree uterovaginal prolapse | -96
    conscious | 0
    drowsy | 0
    tachypneic | 0
    heart rate 120 beats per minute | 0
    blood pressure 90/60 mm Hg | 0
    peripheries cold | 0
    peripheries clammy | 0
    low hemoglobin 6.2 g/dl | 0
    emergency laparotomy | 0
    re-exploration | 0
    low blood pressure | 0
    inotropic support | 0
    triple lumen central venous access secured | 0
    fluid resuscitation | 0
    colloid 1 liter | 0
    packed red blood cells 2 units | 0
    general anesthesia | 0
    left radial artery cannulated | 0
    invasive hemodynamic monitoring | 0
    ligation of bilateral internal iliac arteries | 0
    continuous ooze | 0
    fresh frozen plasma 4 units | 0
    packed red blood cells 3 units | 0
    dopamine 10-15 μg/kg/min | 0
    mean BP 65 mm Hg | 0
    admitted to ICU | 0
    elective ventilation | 0
    disseminated intravascular coagulopathy on second day | 24
    managed with blood products | 24
    managed with cryoprecipitate | 24
    dopamine up to 20 μg/kg/min | 72
    acute respiratory distress syndrome | 72
    increasing ventilatory support | 72
    tracheostomy on seventh day | 168
    ventilatory support continued for 15 days | 168
    dusky discoloration of digits both hands | 72
    extremities cold | 72
    unstable hemodynamic status | 72
    deferred decannulation | 120
    left thumb, index, middle finger worsening discoloration | 120
    left radial artery cannula removed | 120
    vascular surgery opinion sought | 120
    Doppler ultrasound partial thrombosis | 120
    arterial pulsation well felt | 120
    enoxaparin started | 120
    IV dextran started | 120
    stellate ganglion block attempted | 120
    nitroglycerine ointment applied | 120
    right hand discoloration improved | 144
    left hand digits not improved | 144
    digits turning dark | 144
    digits became blackish | 168
    clear line of demarcation | 168
    dry gangrene | 168
    pulmonary rehabilitation | 672
    psychiatric rehabilitation | 672
    amputation of gangrenous digits | 672
    brachial plexus block | 672
    