13 years old | 0
male | 0
atopic dermatitis | 0
not fully vaccinated | 0
presented to the emergency department | 0
progressive fatigue | -96
hypoactivity | -96
slurred speech | -96
lower extremity weakness | -120
progressive | -120
hypoactivity associated with lower extremity weakness | -120
slurred speech | -72
multiple episodes of choking | -72
urinary incontinence | -72
fecal incontinence | -72
difficulty breathing | -24
drooling of saliva | -24
ascending weakness | -24
inability to bear weight | -24
septic shock | 0
IV fluid boluses | 0
systolic blood pressure 100 | 0
hypoxemia | 0
metabolic acidosis | 0
right upper lobe collapse | 0
pneumonia | 0
diffuse infiltrates | 0
early ARDS | 0
non-invasive ventilation | 0
clinical deterioration | 0
decreasing level of consciousness | 0
CT scan of brain | 0
no bleeding | 0
no mass | 0
intubation | 0
mechanical ventilation | 0
MRI Brain normal | 0
broad spectrum antibacterial | 0
transferred to pediatric intensive care unit | 0
WBC 6000 | 0
elevated CRP | 0
elevated ESR | 0
disseminated intravascular coagulopathy | 0
platelets 57000 | 0
INR 1.4 | 0
fibrinogen 456 | 0
D-dimer 0.36 | 0
history of inability to bear weight | -24
choking | -72
absent deep tendon reflexes | 0
negative Babinski reflex | 0
Guillain-Barre syndrome | 0
IVIG treatment | 0
lumbar puncture not done | 0
blood cultures positive for Streptococcus pneumoniae | 48
Mycoplasma pneumoniae serology negative | 0
nasal wash for influenza negative | 0
severe ARDS | 96
hypoxia | 96
respiratory acidosis | 96
continued deterioration | 96
died | 96
