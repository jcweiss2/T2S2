63 years old | 0
male | 0
history of smoking | -8760
hypertension | -8760
vascular disease | -8760
diagnosis of adenocarcinoma | -120
clinically T3 | -120
N3 | -120
M0 | -120
poorly differentiated | -120
stadium IIIB | -120
concurrent chemoradiation therapy | -120
carboplatin/etoposide chemotherapy | -120
radiation therapy | -120
4-dimensional volumetric-modulated arc therapy | -120
target volume for irradiation | -120
mean lung dose | -120
mean heart dose | -120
maximal dose to mediastinal structures | -120
dysphagia grade 3 | -48
weight loss | -48
gastroscopy | -48
radiation esophagitis | -48
stenosis | -48
nasogastric tube | -48
tube feeding | -48
sepsis | 0
acute dyspnea | 0
right sided thoracic pain | 0
reduced right sided airflow | 0
tachycardia | 0
hypotension | 0
saturation of 85% | 0
C-reactive protein of 348 mg/L | 0
leukocytosis of 24.8 × 10^9/L | 0
atelectasis | 0
right sided pleural effusion | 0
mediastinal air configuration | 0
pneumonia | 0
empyema | 0
admitted to intensive care unit | 0
noninvasive ventilation | 0
intravenous broad-spectrum antibiotics | 0
fluid resuscitation | 0
bronchoscopy | 0
bronchopleural fistula | 0
chest tube | 0
drainage of empyema | 0
repeated CT scan | 10
decrease of empyema | 10
consolidations | 10
mediastinal air configuration remained unchanged | 10
no signs of cancer recurrence | 10
multidisciplinary consultation | 14
optimize patient’s condition | 14
enteral feeding | 14
antibiotics | 14
surgical coverage of fistula | 14
pedicled latissimus dorsi flap | 14
surgery | 21
harvesting of latissimus dorsi muscle flap | 21
thoracotomy | 21
defect reached | 21
salvage pneumonectomy considered | 21
pedicled latissimus dorsi flap draped and fixated | 21
ventilator showed insignificant air leak | 21
bronchoscopy showed full coverage of defect | 21
intrathoracic chest tube | 21
lung reinsufflated | 21
wound closed | 21
recovered well | 27
transferred to surgical ward | 27
limited air leakage | 29
drain removed | 31
dismissed to rehabilitation center | 36
readmitted | 630
hemoptysis | 630
pneumonia | 630
anemia | 630
bronchoscopy | 630
large defect of intermediate bronchus | 630
palliative care started | 630
died | 882