38 years old | 0
female | 0
flank pain | -120
fever | -120
raised total leukocyte counts | -120
normal creatinine | -120
pyuria | -120
urine culture grew Escherichia coli | -120
noncontrast computerized tomography of kidney, ureter, and bladder | -120
obstructive calculus in the left lower ureter | -120
ureteroscopy | 0
spinal anesthesia | 0
antibiotics | 0
thick pus drained from the left pelvicalyceal system | 0
ureteric catheter placement | 0
calculus fragmentation with Lithoclast | 0
double-J stent placement | 0
high-grade fever | 6
hypotension | 6
acute respiratory distress syndrome | 6
vasopressors | 6
ventilator support | 6
Gram-negative septicemia | 6
blood parameters repeated | 6
urine and blood culture samples taken | 6
antibiotics stepped up | 6
fluid resuscitation | 6
dopamine | 6
norepinephrine | 6
ventilator support in prone position | 6
acrocyanosis of all four limbs | 6
coagulation panel within normal limits | 6
cardiac evaluation | 6
vasopressors needed for 5 days | 6
acrocyanosis progressed to all four-limb peripheral gangrene | 72
multispecialty management started | 72
conservative local debridement | 72
secondary skin grafting | 72
sympathetic blockade | 72
left below-elbow amputation | 120
right below-knee amputation | 120
loss of all fingers and toes of the other two limbs | 120
discharged | 600