38 years old | 0
female | 0
Caucasian | 0
admitted to the Emergency Department | 0
complaint of malaise | -96
fever | -96
coughing | -96
diarrhea | -96
scleroderma | -6720
treated with chloroquine | -6720
hypotensive | 0
tachycardic | 0
prolonged capillary refill time | 0
administered 3 L of crystalloid fluid | 0
transferred to the Intensive Care Unit | 0
arterial hypotension | 20
norepinephrine infusion | 20
lactate level peaked | 20
norepinephrine infusion reached 0.4 mcg/kg/min | 20
left ventricular impairment | 20
pericardial effusion | 20
dobutamine infusion | 20
intubated | 20
sedated | 20
large spectrum antibiotic | 20
cardiac arrest | 20
cardiopulmonary resuscitation | 20
cardiac tamponade | 20
pericardiocentesis | 20
peripheral venoarterial non-heparin-coated extracorporeal membrane oxygenation | 20
heparin infusion | 20
continuous renal replacement therapy | 20
intra-aortic balloon pump | 48
improvement of hemodynamic condition | 48
lactate levels dropped | 48
requirement of vasopressor agents lessened | 48
improvement of peripheral tissue perfusion | 48
diagnostic hypothesis of viral myocarditis | 48
reversion of organ failures | 48
recovery of left ventricular function | 48
pulseless acute left lower limb ischemia | 48
IABP removal | 48
weaned off ECMO | 120
extubated | 120
vasopressor administration discontinued | 240
left femoral artery thrombectomy | 240
angioplasty | 240
irreversible limb ischemia | 240
deep venous thrombosis | 240
ultrasound scan | 240
platelet count 179,000/mm³ | 240
hypoxemic respiratory failure | 288
septic shock | 288
ventilator-associated pneumonia | 288
reintubation | 288
continuous sedation | 288
broad-spectrum antibiotics | 288
high-dose vasopressors | 288
CRRT maintained | 288
platelet count fallen | 288
nadir of 20,000/mm³ | 312
heparin-induced thrombocytopenia suspected | 312
4 Ts score applied | 312
anti-platelet factor 4/heparin enzyme-linked immunosorbent assay positive | 312
heparin infusion ceased | 312
fondaparinux administration | 312
anti-factor Xa chromogenic assays | 312
platelet count improvement | 336
tracheostomy | 360
debridement of necrotic areas | 360
transtibial amputation | 360
fondaparinux ceased | 360
clinically relevant non major bleeding | 360
blood products transfusion | 360
reoperation for hemostasis | 360
CRRT transitioned to intermittent hemodialysis | 384
renal function recovery | 384
last hemodialysis session | 552
left sided pleural effusion | 720
diagnostic thoracentesis | 720
hemothorax | 720
RBC transfusion | 720
chest tube placement | 720
pleural empyema | 720
pulmonary abscess | 720
lung decortication | 720
antimicrobial therapy | 720
anticoagulant therapy transitioned to oral apixaban | 720
discharged home | 2160