78 years old | 0
man | 0
admitted to Intensive Care Unit | 0
urgent surgical repair of stent-grafting endoleak | -120
urgent surgical repair of aortobronchial fistula | -120
thoracic endovascular repair of descending thoracic aorta aneurysm | -43800
acute renal failure | 96
elevated inflammatory markers | 96
bacteremia | 96
refractory shock | 96
therapy with broad-spectrum antibiotics | 96
no evidence of bleeding | 96
CT-scan revealed thickened esophageal wall | 96
CT-scan revealed small gas bubbles near aortic stent graft | 96
referred to department for upper endoscopy | 96
fistula on posterior surface of middle third of esophagus | 96
aortic stent observed | 96
diagnosis of aortoesophageal fistula | 96
esophageal stenting with covered self-expanding esophageal stent | 96
medical treatment optimized with intravenous proton pump inhibitors | 96
medical treatment optimized with parenteral nutrition | 96
maintaining broad-spectrum antibiotics | 96
no signs of hemorrhage | 672
no signs of infection | 672
recovered from shock | 672
subsequent suspension of amines | 672
subsequent suspension of ventilator support | 672
clinical improvement | 672
patient died unexpectedly | 672
rupture of aortic arch | 672
aortoesophageal fistula secondary to previous thoracic endovascular repair technique | 96
upper gastrointestinal bleeding absent | 96
new-onset fever | 96
esophageal stenting improved septic shock | 672
esophageal stenting prevented bleeding | 672
autopsy identified rupture of aortic arch | 672
