87 years old | 0
    man | 0
    referred to the oncologic center | -1200
    abnormal prostate-specific antigen (PSA) determination | -1200
    physical examination | -1200
    abnormal digital rectal examination | -1200
    firm prostate gland | -1200
    prostate cancer | -1200
    prostatic biopsy | -1200
    Gleason score 7 (3 + 4) adenocarcinoma | -1200
    radionuclide bone scan | -1200
    abnormal uptake in several ribs | -1200
    bone metastasis | -1200
    hypertension | -1200
    chronic kidney disease | -1200
    estimated creatinine clearance of 20 mL/min | -1200
    amlodipine | -1200
    hydrochlorothiazide | -1200
    no anticoagulants | -1200
    no non-steroidal anti-inflammatory drugs | -1200
    no personal history of abnormal bleeding | -1200
    no familial history of abnormal bleeding | -1200
    no altered blood clotting test at diagnosis | -1200
    surgical castration | -960
    significant decrease of the PSA determinations | -960
    nadir of 9 ng/dL | -960
    castration-resistant disease | -768
    PSA levels rose again | -768
    peripheral anti-androgen blockade with bicalutamide | -768
    decline in transient PSA determinations | -768
    rising PSA within 12 months | -576
    second-line therapy with prednisone 5 mg twice daily | -576
    stabilization of the PSA levels at around 20.0 ng/dL | -576
    gross hematuria | 0
    back pain | 0
    spontaneous skin hematomas | 0
    admitted to the emergency department | 0
    severe anemia | 0
    hemoglobin determination of 4.8 g/dL | 0
    red-blood-cell transfusion | 0
    prothrombin time (PT) of 14.7 seconds | 0
    83% of activity | 0
    active partial thromboplastin time (aPTT) of 97.7 seconds | 0
    fibrinogen level of 406 mg/dL | 0
    active partial thromboplastin time not corrected after mixing study | 0
    no lupus anticoagulants identified | 0
    normal liver function tests | 0
    abnormal bleeding | 0
    laboratory abnormalities | 0
    presence of an inhibitor of the coagulation factor | 0
    diagnosis of AHA confirmed | 0
    FVIII < 1% | 0
    FVIII inhibitor quantified as 864 Bethesda Units (BU) | 0
    PSA level stable | 0
    computerized tomography (CT) scan | 0
    no signs of new metastasis | 0
    no evidence of cancer progression | 0
    iliopsoas hematoma | 0
    treatment initiated with prednisone 1 mg/kg per day | 0
    no improvement during the first 48 hours | 48
    daily dose of 100 mg of azathioprine added | 48
    hematuria ceased | 48
    hemoglobin level remained stable | 48
    no signs of new skin hematomas | 48
    no homeostatic agents necessary | 0
    CT study showed no further enlargement of the iliopsoas hematoma | 144
    hematoma-associated back pain improved | 144
    asymptomatic | 144
    discharged after 17 days of hospitalization | 408
    progressive fall of the inhibitor titles | 408
    lowest quantification of 7.6 UBTH | 408
    increase of the coagulation FVIII levels (28%) | 408
    no other hemorrhage phenomenon | 408
    admitted to the Intensive Care Unit | 1872
    diagnosis of pneumonia | 1872
    died due to septic shock | 1872

  