36 years old|0
male|0
diabetic|0
admitted to the hospital|0
high-grade fever|-2160
multiple swellings around joints|-2160
weight loss of 10 kg|-2160
no cough|0
no dyspnoea|0
no abdominal pain|0
episode of septic shock|-2160
fever persisted|-2160
swellings did not respond|-2160
antibiotics (cefaperazone/sulbactum, amikacin, levofloxacin)|-2160
blood cultures were sterile|0
significant proteinuria|0
chest CT showing patchy infiltrates in lungs without cavity, nodules or lymphadenopathy|0
Granulomatosis with polyangiitis considered as differential diagnosis|0
anti-neutrophil cytoplasmic antibody negative|0
anti-proteinase 3 negative|0
anti-myeloperoxidase negative|0
Rheumatoid factor negative|0
anti-nuclear antibody negative|0
HIV negative|0
empirical steroids|0
worsening of symptoms|0
enlargement of swellings|0
no past history of tuberculosis|0
no recurrent infections|0
no alcoholism|0
no intravenous drug abuse|0
no exposure to dust|0
no bird droppings exposure|0
no animal handling exposure|0
no agriculture work exposure|0
cachectic|0
bilateral knee joint contractures|0
diffuse, multiple, tender and firm nodules deep in muscle plane|0
hepatosplenomegaly|0
multiple bilateral lung nodules|0
musculoskeletal ultrasound showing multiple intramuscular densities|0
fine needle aspiration from lesions inconclusive|0
gram stains negative|0
acid fast stains negative|0
polymyositis considered unlikely|0
undifferentiated arthritis considered unlikely|0
aseptic systemic abscess considered unlikely|0
other connective tissue disease considered unlikely|0
high dose of insulin (86 IU/day)|0
continued febrile|0
nodules developed into abscesses|0
vancomycin|168
pus drained from abscesses|168
drank untreated water from a waterfall|-720
melioidosis suspected|0
blood culture isolated Burkholderia pseudomallei|0
diagnosis of melioidosis confirmed|0
administered intravenous ceftazidime|0
fever subsided|672
pyomyositis resolved|672
lung nodules subsided|672
underwent eradication phase with oral cotrimoxazole|672
repeat contrast CT scan showing clearance of lung nodules|4032
managed diabetes with metformin|672
underwent physical therapy|672
complete resolution of symptoms|4032
return to baseline function|4032
