15 years old | 0
male | 0
mild asthma | 0
involved in road traffic accident | -120
not wearing helmet | -120
collided with car | -120
Glasgow Coma Scale 6 | -120
Oxygen saturation 75% | -120
intubated | -120
respiratory failure | -120
airway protection | -120
Chest xray shows massive right haemothorax | -120
segmented fracture of 6th posterior rib | -120
Ipsilateral chest tube inserted | -120
300 ml of blood drained | -120
transferred to Hospital University Sains Malaysia | -120
CT of brain reveals subarachnoid haemorrhage | -120
punctate intracerebral haemorrhage | -120
burr hole | -120
intracranial pressure monitoring | -120
transferred to Intensive Care Unit | -96
ventilator support | -96
inotropic support | -96
Noradrenaline 0.1-0.2 mcg/kg/min | -96
extubated | -72
reintubated | -64
febrile | -64
temperature 38-40°C | -64
Bronchoscopy | -64
purulent secretions | -64
blood cultures grew Burkholderia pseudomallei | -64
tracheal secretions cultures grew Burkholderia pseudomallei | -64
bronchoalveolar lavage fluid cultures grew Burkholderia pseudomallei | -64
Gram stain showed gram negative bacilli | -64
safety-pin appearance | -64
sensitive to amoxicillin-clavulanate | -64
sensitive to ceftazidime | -64
sensitive to doxycycline | -64
sensitive to imipenem | -64
sensitive to trimethoprim-sulfamethoxazole | -64
Hepatitis B screening negative | -64
Hepatitis C screening negative | -64
HIV screening negative | -64
syphilis screening negative | -64
CXR shows right hemithorax consolidations | -64
low to moderate ventilator setting | -64
minimal inotropic support | -64
extubated | 168
discharged to general ward | 504
IV Meropenem 1g 8-hourly | -56
deescalated to IV Ceftazidime 2g 8-hourly | 0
oral trimethoprim/sulfamethoxazole | 168
eradication phase | 168