79 years old | 0
female | 0
surgery on the medial collateral ligament | -7200
TKA | -8760
fell from a height of about 50 cm | -1
overstretched the right knee | -1
right knee pain | -1
admitted to the hospital | 0
periprosthetic tibial fracture | 0
popliteal artery injury | 0
right dorsalis pedis artery was not palpable | 0
transferred to emergency and critical care medicine center | 0
computed tomography angiography | 0
emergency surgery for revascularization | 0
semicircular partial rupture of the popliteal artery | 0
anastomosis between the popliteal and posterior tibial arteries | 0
damage to the popliteal vein | 0
excision of the injured area | 0
end-to-end anastomosis | 0
external fixation across the knee | 0
internal fixation | 264
Felix classification IIB | 264
anatomical locking plates | 264
screws inserted forwards and backwards of the keel of the tibial implant | 264
antibiotic treatment | 312
surgical-site sepsis | 312
debridement | 336
exposed plate covered using the gastrocnemius muscle flap | 504
infection resolved | 1200
partial weight-bearing | 2160
bone union confirmed | 3600