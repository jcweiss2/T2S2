23 years old | 0
    pregnant | 0
    female | 0
    presented to the emergency room | 0
    high-grade fever | 0
    high-grade fever for one week | 0
    abnormal movements of her eyes | -120
    abnormal movements of her limbs | -120
    no history of drug intake | 0
    no history of toxin intake | 0
    restless | 0
    appeared sick | 0
    blood pressure 90/50 mm Hg | 0
    pulse rate 120 beats/minute | 0
    respiratory rate 32 breaths/minute | 0
    oxygen saturation 96% on room air | 0
    bilateral basal crepitations | 0
    typical ‘cigarette burn’ eschar | 0
    conscious | 0
    oriented to time | 0
    oriented to place | 0
    oriented to person | 0
    opsoclonus | 0
    myoclonic jerks involving all four limbs | 0
    normal tone | 0
    normal power | 0
    normal deep tendon reflexes | 0
    no features of parkinsonism | 0
    no bradykinesia | 0
    no rigidity | 0
    no features of cerebellar dysfunction | 0
    normal finger-nose test | 0
    normal heel-knee-shin test | 0
    normal tandem gait test | 0
    elevated leukocyte count | 0
    thrombocytopenia | 0
    deranged renal function | 0
    deranged hepatic function | 0
    elevated total bilirubin | 0
    elevated aspartate aminotransferase | 0
    elevated alanine transaminase | 0
    multiorgan dysfunction | 0
    normal serum sodium | 0
    normal serum potassium | 0
    normal serum magnesium | 0
    normal serum calcium | 0
    emergency cesarean section | 0
    intensive care admission | 0
    treated with injectable azithromycin | 0
    supportive management | 0
    diagnosis of scrub typhus confirmed by IgM ELISA | 0
    negative vasculitis markers | 0
    negative autoimmune antibody profile | 0
    negative paraneoplastic antibody profile | 0
    negative HIV serology | 0
    negative hepatitis B serology | 0
    negative hepatitis C serology | 0
    negative VDRL test | 0
    normal brain MRI with contrast | 0
    normal cerebrospinal fluid examination | 0
    normal electroencephalography | 0
    normal PET-CT | 0
    OMS gradually resolved over the next two weeks | 168
    