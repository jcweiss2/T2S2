64 years old | 0
male | 0
hypertension | 0
hiatal hernia | 0
osteoarthritis | 0
acute worsening of chronic lower back pain | -336
progressive weakness in lower extremities | -336
use of cane | -336
use of walker | -336
non-ambulant | -336
subjective fevers | -336
temperature of 100.1°F | 0
blood pressure normal | 0
respiratory rate normal | 0
heart rate normal | 0
no distress | 0
cachectic | 0
disheveled | 0
poor dentition | 0
regular heart rate | 0
regular rhythm | 0
normal S1 | 0
normal S2 | 0
no murmurs | 0
clear lungs | 0
bilateral air entry | 0
crepitus in both knees | 0
limping gait | 0
Kernig’s sign obscured | 0
Brudzinski’s sign obscured | 0
chronic bilateral knee pain | 0
congenital deformation of right knee | 0
smoker | 0
40 pack-years | 0
occasional alcohol use | 0
occasional marijuana use | 0
denies intravenous drugs | 0
toxicology positive for oxycodone | 0
leukocytosis of 25,500 | 0
89% neutrophils | 0
no bands | 0
sedimentation rate of 44 | 0
lactic acid 1.6 | 0
anion gap 18 | 0
thoracic spine CT | 0
lumbar spine CT | 0
multilevel central canal compromise | 0
bilateral neural foraminal compromise | 0
no evidence of abscess | 0
cavitary lesion in left lower lobe | 0
circumferential thick wall | 0
left inferior renal pole abnormalities | 0
blood cultures grew S. aureus | 0
started on vancomycin | 0
TTE performed | 0
ejection fraction 65% | 0
normal valves | 0
no vegetations | 0
clinical picture worsened | 24
altered mental status | 24
nuchal rigidity | 24
lumbar puncture | 24
meningitis | 24
cerebrospinal fluid leukocytosis of 1157 | 24
culture positive for S. aureus | 24
HIV negative | 24
HSV negative | 24
PPD negative | 24
spine MRI | 24
osteomyelitis at T12-L1 | 24
renal infarcts | 24
continued febrile | 24
vancomycin MIC <2 mg/mL | 24
trough previous to 4th dose 11 | 24
repeat trough 18.4 | 24
repeat blood cultures at 48 hours | 48
repeat blood cultures at 96 hours | 96
clinical deterioration | 144
tachypnea | 144
hypoxia | 144
new systolic 2/6 murmur | 144
louder over cardiac apex area | 144
bilateral respiratory crackles | 144
new right hemiparesis | 144
upgoing Babinski reflex | 144
switched to nafcillin | 72
blood culture confirmed methicillin susceptibility | 72
head MRI | 144
multiple infarcts | 144
non-vascular pattern | 144
TEE | 144
severe mitral regurgitation | 144
severe tricuspid regurgitation | 144
1.5 cm vegetation on mitral valve | 144
transferred to ICU | 144
MSSA bacteremia | 144
IE | 144
osteomyelitis | 144
meningitis | 144
ischemic stroke | 144
renal infarcts | 144
pulmonary infarcts | 144
continued nafcillin | 144
resolution of leukocytosis | 144
resolution of fever | 144
mental status improvement | 144
indications for mitral valve replacement | 144
not feasible due to embolic stroke | 144
follow up TTE | 672
worsening mitral valve involvement | 672
worsening tricuspid valve involvement | 672
mitral valve replacement | 672
tricuspid valve replacement | 672
completed 8 weeks of nafcillin | 1344
discharged | 1344
dual-chamber pacemaker | 1344
persistent 3rd degree AV block | 1344
