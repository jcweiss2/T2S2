33 years old | 0
female | 0
chronic hypersensitivity pneumonitis | -672
dyspnea | -672
high-dose glucocorticoids | -672
azathioprine | -672
admitted to the hospital | 0
mechanical ventilation | -672
 FiO2 0.21 | -672
brain dead donor | -24
traumatic brain injury | -24
donor lungs explantation | 0
secretions in main bronchi | 0
swabs sent for bacterial culture | 0
thoracic cavity accessed | 0
clamshell incision | 0
lung transplantation | 0
induction immunosuppression | 0
intravenous basiliximab | 0
intravenous methylprednisolone | 0
surgery completed | 10
shifted to Intensive Care Unit | 10
immunosuppression | 10
intravenous methylprednisolone | 10
oral tacrolimus | 10
histopathological examination | 10
airway-centric fibrosis | 10
FiO2 0.4 | 0
bilateral diffuse alveolar opacities | 24
echocardiography | 24
normal ejection fraction | 24
primary graft dysfunction | 24
antibody-mediated rejection | 24
hospital-acquired infection | 24
direct crossmatch | 0
negative results | 0
intravenous colistin | 24
intravenous vancomycin | 24
extubated | 48
preemptive noninvasive ventilation | 48
culture from bronchial swabs | 24
MDR Klebsiella pneumoniae | 24
blood culture | 24
bronchoalveolar lavage fluid | 24
intravenous tigecycline | 72
vancomycin stopped | 72
tacrolimus withheld | 72
basiliximab withheld | 72
oral prednisolone | 72
fever | 24
respiratory failure | 24
bilateral empyema | 120
intravenous fosfomycin | 120
intrapleural irrigation | 120
partial clearing of lung opacities | 168
weaned off NIV | 168
high-flow nasal cannula | 168
nasal prongs | 168
acute onset hypotension | 288
fresh blood in chest drains | 288
surgical re-exploration | 288
anterior wall of right ventricle punctured | 288
sternal wire | 288
repaired | 288
refractory septic shock | 336
hospital-acquired pneumonia | 336
death | 336
biopsy of transplanted lung | 288
no evidence of graft rejection | 288