56 years old | 0
female | 0
morbidly obese | 0
no history of cardiac disease | 0
feeling poorly | -72
cough | -72
fatigue | -72
found on bedroom floor | -1
nonresponsive | -1
without palpable pulse | -1
chest compressions initiated | -1
automated external defibrillator used | -1
automated rhythm analysis | -1
shock advised | -1
shock delivered | -1
patient awakened | 0
admitted to medical intensive care unit | 0
diagnosed with Klebsiella pneumonia | 0
treated over 2-week course | 0
echocardiogram demonstrated normal heart | 24
no arrhythmias during hospital course | 24
cardiac electrophysiologist consulted | 24
implantable cardioverter-defibrillator considered | 24
rhythm strip from AED obtained | 48
review of rhythm strip revealed incorrect interpretation | 48
sinus tachycardia misinterpreted as ventricular arrhythmia | 48
shock presumably awakened patient | -1
discharged from hospital | 336