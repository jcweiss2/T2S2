29 years old | 0
female | 0
Crohn’s disease for 10 years | -87600
left colon involvement | -87600
perianal fistula | -87600
Infliximab monotherapy | -87600
peri-anal abscess drainage 1 year ago | -8760
failed Certolizumab Pegol | -8760
pregnancy (35th week) | 0
mild peri-anal pain | 0
discharged following reassuring clinical examination | 0
worsening pain | 120
admitted for fetal monitoring and colorectal evaluation | 120
anal stricture | 120
white blood cell count 13500 | 120
C-reactive protein 115 mg/L | 120
perineal ultrasound showing 9-ml fluid collection | 120
intravenous ceftriaxone | 120
intravenous metronidazole | 120
emergency cesarean section due to fetal distress | 132
tachycardia (HR 124 bpm) | 144
hypotension (MAP 62 mmHg) | 144
perianal pain progressed | 144
diffuse hyperemia | 144
swelling of the vulva | 144
purple discoloration of the skin | 144
Fournier’s gangrene | 144
wide drainage | 144
debridement | 144
necrosis of the ischiorectal fat | 144
foul-smelling purulent discharge | 144
visualization of healthy tissue | 144
rectal ulcers | 144
fistulous opening with purulent discharge | 144
anal sphincter spared from necrosis | 144
laparoscopic loop ileostomy | 144
intraoperative colonic lavage | 144
vacuum-assisted therapy | 144
hydrocolloid paste | 144
polymicrobial infection | 144
Eschericia Coli | 144
Citrobacter freundii complex | 144
Candida albicans | 144
antibiotics adjusted | 144
discharged from Intensive Care Unit after 3 days | 144
postoperative day 14 | 336
4 debridements | 336
vacuum-therapy exchanges | 336
perineal defect closed with unilateral medial thigh advancement flap | 336
draining seton placed in suprasphincteric fistula | 336
discharged after 28 days of hospitalization | 672
medial thigh flap completely healed | 2160
no signs of infection | 2160
seton kept in place | 2160
Infliximab monotherapy resumed | 2160
ileostomy reversal planned | 2160
baby recovered well | 144
fetal distress | 132
oligohydramnios | 132
negative HIV serology | 0
no other clinical comorbidities | 0
unremarkable prenatal care | 0
