18 years old | 0
male | 0
admitted to hospital | 0
fever | -72
shortness of breath | -72
weight loss | -216
lethargy | -216
swallowing difficulties | -216
bilateral interstitial infiltrates | 0
empirical therapy for community-acquired pneumonia | 0
intubated | 0
hypoxic respiratory failure | 0
widespread nodular infiltrates | 0
mediastinal abscess | 0
septic | 0
high-dose vasopressors | 0
hemodynamic instability | 0
lung-protective mechanical ventilation | 0
prone positioning | 0
negative cultures from bronchoalveolar lavage | 0
negative viral PCR assays | 0
Ziehl-Neelsen staining negative | 0
indeterminable IGRA for tuberculosis | 0
antibiotic therapy | 0
empirical corticosteroids | 0
immunoglobulins | 0
transbronchial biopsies | 18
bilateral tension pneumothoraces | 18
pneumopericardium | 18
subcutant emphysema | 18
veno-venous ECMO therapy | 18
microscopy of transbronchial biopsies revealed acid-fast bacilli | 18
tuberculosis treatment initiated | 18
rifampicin | 18
isoniazide | 18
ethambutol | 18
pyrazinamide | 18
growth of Mycobacterium tuberculosis detected | 26
granulomas in bone marrow aspirate | 26
granulomas in liver biopsies | 26
granulomas in lung biopsies | 26
dysphagia | 0
mediastinal abscess | 0
multiple bullae | 336
persistent pneumothoraces | 336
subtherapeutic levels of isoniazid | 336
subtherapeutic levels of rifampicin | 336
multi-resistant Pseudomonas aeruginosa | 336
Stenotrophomonas maltophilia | 336
inhaled colistin | 336
tobramycin | 336
intravenous amikacin | 336
meropenem | 336
ceftazidime/avibactam | 336
low serum levels of amikacin | 336
signs of recovery | 45
increasing lung compliance | 45
re-expansion of lungs | 45
weaned from ECMO | 50
thrombocytopenia | 50
minor bleedings from puncture sites | 50
sensory symptoms in lower limbs | 50
discharged from ICU | 76
resumed previous activities | 120