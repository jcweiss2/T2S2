47 years old | 0
man | 0
presented to hospital | 0
symptoms typical of COVID-19 infection | -48
fever | -48
sweats | -48
cough | -48
shortness of breath | -48
COVID-19 diagnosis (nasopharyngeal swab) | 0
right basal atelectasis (CXR) | 0
inpatient duration | 0
ventilatory support (2 days) | 72
continuous positive airway pressure | 72
cardiovascular inotropic support not required | 0
dexamethasone treatment | 0
discharged | 504
represented with chest pain | 336
shortness of breath (recurrence) | 336
COVID-19 negative tests | 336
large left hydropneumothorax (CTPA) | 336
air fluid levels in left lower pleural cavity | 336
unclear differential between parenchymal abscess, necrotic lung, empyema | 336
right lung patchy basal consolidation | 336
small air fluid collection (COVID-19 infection) | 336
empirical antimicrobial therapy (clarithromycin, piperacillin/tazobactam) | 336
antibiotics escalation to meropenem | 336
intercostal drain insertion | 336
pleural fluid pH 7.1 | 336
microbiology cultures negative | 336
failed drainage of pleural cavity | 336
left uniportal video-assisted thoracoscopy | 1008
left pleural washout and decortication intent | 1008
intraparenchymal pathology | 1008
dark-colored, friable, necrotic lower lobe | 1008
left lower lobectomy | 1008
antibiotics continued post-surgery | 1008
fall in white cell count | 1008
fall in C reactive protein | 1008
sinus tachycardia (2 weeks) | 1008
resolved sinus tachycardia at discharge | 1008
no further surgical intervention required | 1008
antibiotics discontinued at discharge | 1008
mobile and independent in activities | 1008
no subsequent readmission | 1008
clear pleural spaces (CXR at discharge) | 1008
loss of left hemithorax volume (post lobectomy) | 1008
macroscopic inspection findings | 1008
microscopic evaluation findings | 1008
lytic therapy not considered | 336
