46 years old | 0
male | 0
admitted to the hospital | 0
ulcerative colitis | -672
malaise | -72
fever | -72
loss of appetite | -72
chills | -72
nausea | -72
blood pressure 124/46 mmHg | 0
heart rate 122 beats per min | 0
SpO2 98% | 0
respiratory rate 16/min | 0
body temperature 40.2°C | 0
cardiac arrest | 0
chest compression | 0
tracheal intubation | 0
ventricular fibrillation | 0
defibrillation | 0
adrenaline administered | 0
coved-type ST elevation in V1 and V2 | 0
Brugada syndrome | 0
hypercalcemia | 0
hypotension | 2
septic shock | 2
tazobactam-piperacillin administered | 2
vasopressors administered | 2
extubation | 48
fever reoccurred | 120
liver abscess | 120
meropenem administered | 120
vancomycin administered | 120
puncture drainage | 120
infection controlled | 720
pilsicainide test positive | 720
implantable cardioverter defibrillator implanted | 720
discharged | 720
sudden death in family history | -100000
ectopic parathyroid adenoma | 720
high parathyroid hormone levels | 720
abnormal uptake in the anterior mediastinum | 720
tumor resection | 720
nonfunctional pituitary adenoma | 720
nonfunctional adrenal tumor | 720
multiple endocrine neoplasia type 1 | 720
electrocardiogram taken on October 4, 2021 | -100000
electrocardiogram taken on June 28, 2021 | -100000
electrocardiogram taken on March 24, 2021 | 0
electrocardiogram taken on September 25, 2017 | -100000
J point elevation | -100000
early repolarization | -100000
inferolateral early repolarization | -100000