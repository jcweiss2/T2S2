78 years old | 0
man | 0
high-grade T1 urothelial carcinoma | 0
status post-transurethral resection of bladder tumor | 0
intravesical BCG instillation | -1344
fever | 0
rigors | 0
altered mental status | 0
shortness of breath | 0
denies cough | 0
denies chest pain | 0
no urinary symptoms | 0
no gastrointestinal symptoms | 0
BCG instillation done day before presentation | -24
temperature of 102.8 F | 0
pulse rate of 92/min | 0
respiratory rate of 40/min | 0
blood pressure 78/45 mmHg | 0
oxygen saturation of 93% on ambient air | 0
appears toxic | 0
dehydrated | 0
in respiratory distress | 0
asymmetric chest expansion | 0
dullness to percussion | 0
decreased tactile fremitus on the left side | 0
reduced air entry on auscultation | 0
unremarkable cardiovascular examination | 0
marked leukocytosis | 0
white cell count of 27,200/microliter | 0
hemoglobin of 11.5 g/dL | 0
lactate was markedly elevated at 7.8 meq/L | 0
high anion gap metabolic acidosis | 0
creatinine of 2.31 mg/dL | 0
blood urea nitrogen of 28 mg/dL | 0
sputum culture with gram stain showed normal oral flora | 0
urinary streptococcal antigen negative | 0
urinary legionella antigen negative | 0
chest X-ray revealed left basilar pneumonia | 0
chest X-ray revealed small left pleural effusion | 0
CT head showed no acute intracranial abnormalities | 0
preliminary blood culture negative | 0
intubated | 0
placed on ventilation | 0
commenced on vasopressors | 0
intravenous Vancomycin | 0
intravenous Piperacillin-Tazobactam | 0
septic shock | 0
community-acquired pneumonia | 0
possible urinary tract infection | 0
completion of several courses of broad-spectrum antibiotics | 0
continued low-grade pyrexia | 0
failed to improve clinically | 0
suspicion for systemic BCG dissemination | 0
blood cultures for acid-fast bacilli returned positive | 0
Mycobacteria bovis confirmed | 0
broad-spectrum antibiotics discontinued | 0
commenced on Isoniazid | 0
commenced on Ethambutol | 0
commenced on Rifampicin | 0
improved clinically | 0
discharged | 120
completed 2 months of triple therapy | 0
maintenance therapy with Rifampicin and Isoniazid | 0
return for follow up with infectious disease team | 0
