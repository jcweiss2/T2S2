39 years old | 0
Spanish | 0
male | 0
malnutrition | 0
alcohol abuse | 0
drug abuse | 0
smoking | 0
pulmonary tuberculosis | 0
cured pulmonary tuberculosis | 0
admitted to the Emergency Department | 0
temperature of 38°C | 0
abdominal pain | 0
7-day diarrhea | 0
no recent travel history | 0
never traveled outside of Europe | 0
no reported oral-anal sexual contact | 0
no history of receiving corticosteroids | 0
no history of immunosuppressant medication | 0
tachycardia | 0
tachypnea | 0
leucocytosis of 14×10^9/l | 0
raised serum transaminases | 0
inflammatory markers | 0
C-reactive protein level of 308 mg/l | 0
procalcitonin level of 39 ng/l | 0
abdominal CT scan | 0
multiple liver abscesses in the right liver lobe | 0
liver segments I and III | 0
empirical antibiotic treatment with i.v. meropenem | 0
acute clinical deterioration | -120
transferred to surgical Intensive Care Unit | 0
endotracheally intubated | 0
mechanical ventilation started | 0
vasopressor support | 0
septic shock | 0
percutaneous CT-guide drainage of the liver abscesses | 0
micro-biological samples obtained | 0
on the 5th day of admission in ICU | 120
liver aspirate revealed structures compatible with E. histolytica trophozoites | 120
genomic DNA isolated | 120
detection of Entamoeba histolytica DNA by real-time PCR | 120
RT-PCR positive in liver aspirate | 120
stool samples positive for E. histolytica | 120
bacterial cultures negative | 120
diagnosis of intestinal and extraintestinal amebiasis | 0
i.v. metronidazole added | 0
oral paromomycin | 0
respiratory deterioration | 168
thoracoabdominal CT scan | 168
bilateral pleural effusion | 168
abscess in the right lower pulmonary lobe | 168
small disseminated intraabdominal abscesses | 168
on the 10th day of admission | 240
amebic skin lesions appeared on the chest and face | 240
bronchial aspirate | 240
pleural drainage | 240
blood | 240
skin biopsy | 240
RT-PCR positive in all samples | 240
HIV serology negative | 240
PCR negative for Acanthamoeba spp | 240
PCR negative for Balamuthia mandrillaris | 240
PCR negative for Naegleria fowleri | 240
on the 15th day of ICU stay | 360
neurological symptoms with aphasia | 360
right-sided hemiplegia | 360
cranial CT scan | 360
multiple brain abscesses in left basal ganglia | 360
right temporal lobe | 360
right lenticular nucleus | 360
conservative management | 360
no brain samples obtained | 360
i.v. metronidazole therapy | 360
neurological symptoms improved | 360
full recovery of language | 360
slight paresis in the right arm | 360
end-of-treatment CT scans | 1680
residual liver abscesses | 1680
residual brain abscesses | 1680
co-infection of liver abscesses by Staphylococcus epidermidis | 0
Clostridium difficile pseudomembranous colitis | 0
discharged after 16-week stay | 2688
currently stable | 2688
rehabilitating | 2688
