18 years old | 0
male | 0
admitted to the hospital | 0
orthotopic heart transplant | 0
familial hypertrophic cardiomyopathy | -672
immunosuppressant regimen | 0
prednisone | 0
mycophenolate mofetil | 0
tacrolimus | 0
extubated | -48
shortness of breath | -72
hypoxic respiratory failure | -72
endotracheal intubation | -72
mechanical ventilation | -72
hemodynamically unstable | -72
vasopressor support | -72
increased white blood cell count | -72
neutrophils | -72
bands | -72
lymphocytes | -72
monocytes | -72
renal function tests | -72
liver function tests | -72
blood cultures | -72
broad-spectrum antibiotics | -72
vancomycin | -72
cefepime | -72
azithromycin | -72
computed tomography of the chest | -72
bilateral pulmonary consolidations | -72
air bronchograms | -72
bilateral pneumothoraces | -72
bronchoscopy | -96
bronchial washings | -96
bronchoalveolar lavage | -96
Candida albicans | -96
blood cultures | -120
no microbial growth | -120
repeat CT chest | -120
worsening diffuse pulmonary consolidations | -120
bronchoscopy | -216
BAL cultures | -216
mycobacteria | -216
Mycoplasma pneumoniae | -216
Legionella | -216
BAL viral cultures | -216
adenovirus | -216
Cytomegalovirus | -216
influenza | -216
parainfluenza | -216
respiratory syncytial virus | -216
blood CMV viral load | -216
HIV serology | -216
serum cryptococcal antigen | -216
serum Aspergillus galactomannan assay | -216
serum (1→3)-β-D-glucan assay | -216
urine for Histoplasma antigen | -216
BAL cytology | -216
acute inflammatory cells | -216
Gomori's methenamine silver stain | -216
cystic forms of Pneumocystis jirovecii | -216
Aspergillus species | -216
voriconazole | -216
micafungin | -216
combination therapy | -216
dramatic response | -192
vasopressor support discontinued | -192
therapeutic voriconazole trough levels | -192
micafungin discontinued | -192
intravenous voriconazole transitioned to oral route | -192
maintenance therapy | -192
review of day 4 posttransplant BAL fungal cultures | -192
Aspergillus species | -192
Candida colonies | -192
gardening | -192
spreading mulch | -192
donor-derived infection | -192
nosocomial environmental source | -192
Aspergillus contamination | -192
other organ recipients | -192
hospital construction | -192
renovation | -192
Infection Prevention team | -192
air sampling cultures | -192
patient's room | -192
adjacent rooms | -192
mold spore concentrations | -192
basidiospore variety | -192
Aspergillus spore | -192
immunosuppression decreased | -192
bilateral chest tubes | -192
persistent air leak | -192
antifungal therapy | -192
discharged | 1008
voriconazole maintenance monotherapy | 1008
repeat serum Aspergillus galactomannan assay | 1008
voriconazole therapy | 1008
pulmonary recovery | 1008
clinical signs of relapse | 1008
Aspergillus infection | 1008