42 years old | 0
    female | 0
    admitted to the hospital | 0
    fever | -168
    diffuse abdominal pain | -168
    discomfort during intercourse | -168
    complete blood count revealed no abnormalities | 0
    blood cultures negative for bacteria and fungi | 0
    urine cultures negative for bacteria and fungi | 0
    colposcopy | 0
    abnormal area in the cervix | 0
    Papanicolaou test showed abnormal cells | 0
    cervical colposcopic biopsies | 0
    endocervical curettage | 0
    cone biopsy | 0
    cervical intraepithelial neoplasia (CIN) grade 3 | 0
    squamous cell carcinoma | 0
    chemotherapy | 0
    radiotherapy | 0
    full clinical recovery | 0
    discharged home | 0
    hospitalized with diabetes mellitus | 8760
    abdominal distension | 8760
    appetite loss | 8760
    hypoalbuminemia | 8760
    intestinal sub occlusion | 8760
    actinic stenosis | 8760
    bowel resection | 8760
    jejunostomy | 8760
    parenteral nutrition | 8760
    antibiotic therapy | 8760
    adhesions between bowel loops | 8760
    mucous fistula | 8760
    corrective enterectomy | 8760
    fecal content | 8760
    intestinal evisceration | 8760
    aponeurotic dehiscence | 8760
    surgical wound infection | 8760
    Pseudomonas aeruginosa infection | 8760
    Citrobacter sp. infection | 8760
    Acinetobacter sp. infection | 8760
    sepsis | 8760
    generally worsening clinical condition | 8760
    intravenous vancomycin | 8760
    imipenem | 8760
    metronidazole | 8760
    readmitted to the intensive care unit | 8760
    fever episodes | 8760
    severe abdominal pain | 8760
    weakness | 8760
    respiratory distress | 8760
    elevated urea | 8760
    elevated creatinine | 8760
    leukopenia | 8760
    low hemoglobin | 8760
    low platelets | 8760
    venous blood samples collected | 8760
    blood cultures processed for mycological diagnosis | 8760
    direct examination with India ink | 8760
    culture on Sabouraud Dextrose Agar medium | 8760
    budding capsulated yeast cells | 8760
    blood cultures positive after five days of growth | 8760
    colonies grew | 8760
    contrasted budding encapsulated yeast cells | 8760
    nonfermentative colonies | 8760
    absence of KNO3 utilization | 8760
    caffeic acid negative | 8760
    urease positive | 8760
    utilization of lactose | 8760
    d-glucuronate | 8760
    d-gluconate | 8760
    melibiose | 8760
    Cryptococcus laurentii bloodstream infection | 8760
    bronchoalveolar lavage | 8760
    cerebrospinal fluid analysis | 8760
    cryptococcal latex agglutination | 8760
    no fungi detected | 8760
    minimal inhibitory concentrations determined | 8760
    sensitive to amphotericin B | 8760
    sensitive to fluconazole | 8760
    persistent elevated urea | 8760
    persistent elevated creatinine | 8760
    fluconazole treatment | 8760
    intravenous fluconazole | 8760
    central venous catheter removal | 8760
    significant improvement | 8760
    discharged home | 8760
    immunosuppressed due to radio and chemotherapy | 0
    diabetic status | 0
    multiple catheters and invasive medical devices | 0
    possible source of fungaemia | 0
    catheter tip removed during antifungal treatment | 8760
    nosocomial infection | 0
    susceptible patient | 0
    immunosuppressive therapies | 0
    contact with Cryptococcus laurentii | 0
    developed nosocomial infection | 0
    expand beyond environmental niche | 0
    recognized human pathogen | 0