52 years old | 0
Indian | 0
woman | 0
presented to hospital | 0
one-week history of right-sided retro#orbital pain | -168
right-sided retro-orbital pain | -168
facial swelling | -168
no other significant past medical history | 0
apyrexial | 0
pulse rate of 100 min–1 | 0
confused | 0
right-sided periorbital cellulitis | 0
decreased visual acuity in the right eye | 0
full range of extraocular muscle movements | 0
ipsilateral mild facial nerve weakness (House-Brackmann classification grade II) | 0
neutrophilic leukocytosis (31.6 x 109/L) | 0
C-reactive protein of 456 mg/L | 0
random blood glucose of 56.1 mmol/L | 0
urine dipstick analysis identified the presence of ketones | 0
blood gas analysis confirmed a metabolic acidosis | 0
clinical diagnosis of diabetic ketoacidosis | 0
treated with intravenous fluid replacement | 0
intravenous antibiotics (co-amoxiclav and metronidazole) | 0
insulin sliding scale | 0
CT of the head including both orbits confirmed right periorbital cellulitis | 0
stranding of the extraconal adipose tissue consistent with Chandler classification grade II | 0
no evidence of intra-orbital collection | 0
no intracranial extension | 0
complete opacification of the right nasal cavity | 0
complete opacification of the maxillary sinuses | 0
complete opacification of the frontal sinuses | 0
presumed source of sepsis | 0
endoscopic exploration under general anaesthesia | 0
large necrotic mass in the right nasal cavity | 0
biopsies sent for histopathology | 0
biopsies sent for microscopy | 0
biopsies sent for sensitivity | 0
histopathological assessment revealed fungal invasion | 0
fungal hyphae broad and distorted | 0
fungal hyphae branching at right angles | 0
surrounded by extensive necrotic debris | 0
no septae | 0
right nasal cavity exenterated | 0
paranasal sinuses exenterated | 0
irrigated | 0
parenteral amphotericin B added to treatment regime | 0
initial transient improvement in temperature | 0
initial transient improvement in conscious level | 0
cranial neuropathies persisted | 0
deteriorated becoming more confused | 0
losing vision completely from the right eye | 0
MRI scan of the head revealed right frontal cerebritis | 0
early abscess formation | 0
direct extension from nasal cavity into frontal lobes | 0
through cribiform plate | 0
re-accumulation of fluid | 0
thickening of the mucosa in the paranasal sinuses | 0
disease affecting sphenoid sinuses | 0
disease affecting ethmoid sinuses | 0
right maxillectomy performed via lateral rhinotomy approach | 0
orbital exenteration | 0
right eye necrotic | 0
frontal sinus opened | 0
mass extending into dura | 0
dura opened | 0
necrotic cerebral parenchyma removed | 0
repeated irrigation | 0
transferred to Intensive Care Unit | 0
failed to recover | 0
died | 144
generalized seizure | 144
