7 years old | 0
male | 0
Hispanic | 0
admitted to the hospital | 0
non-productive cough | -720
history of asthma | -720
albuterol inhaler | -720
non-bloody, non-bilious emesis | -720
fever | -720
temperature 104 | -720
decreased appetite | -720
4 pound weight loss | -720
denies pets in the home | 0
denies recent travel | 0
denies sick contacts | 0
denies foreign or new foods | 0
denies animal or insect bites | 0
denies fevers | 0
denies diarrhea | 0
denies constipation | 0
denies chills | 0
asthma well controlled | 0
fully immunized | 0
no allergies to medications | 0
unremarkable family history | 0
previous normal growth and development | 0
no surgical history | 0
non-tender, palpable, mobile lymphadenopathy | 0
lungs clear to auscultation | 0
para-tracheal mass | 0
CT scan | 0
paratracheal mass with supraclavicular lymph nodes | 0
teratoma | 0
thymoma | 0
lymphoma | 0
thyroid related tumor | 0
granulomatous type process | 0
Ceftriaxone | 0
white blood cell count 6.8 × 10^3/mL | 0
hemoglobin 11.5 g/dL | 0
platelets 307 × 10^3/mL | 0
neutrophil 23% | 0
lymphocytes 46% | 0
monocytes 12% | 0
eosinophils 18% | 0
ESR 30 mm/hr | 0
CRP < 0.012 mg/dL | 0
LDH 197 U/L | 0
uric acid 2.7 mg/dL | 0
comprehensive metabolic panel normal | 0
glucose normal | 0
bilirubin normal | 0
urinalysis normal | 0
TSH/T4 normal | 0
HIV negative | 0
PPD negative | 0
homovanillic acid normal | 0
vanillylmandelic acid normal | 0
angiotensin converting enzyme normal | 0
ANCA negative | 0
MRI of the brain normal | 0
blood cultures negative | 0
stool cultures negative | 0
serum cryptococcal antigen positive | 0
repeat serum cryptococcal antigen negative | 72
histoplasmosis H band negative | 0
M band antibody positive | 0
thoracotomy | 0
purulent fluid from the mass | 0
biopsies from the mediastinal lymph nodes | 0
biopsies from the right upper lung lobe | 0
biopsies from the mediastinal nodule | 0
biopsies from the mediastinal mass | 0
post-op pneumothorax | 24
right-sided chest tube | 24
spinal tap | 48
cerebral spinal fluid analysis normal | 48
necrotizing granulomatous inflammation with calcification | 0
itraconazole | 0
12 week course of itraconazole | 0
Hydrocodone/Acetaminophen | 0
Ketorolac | 0
incentive spirometry | 0
serial chest x-rays | 0
progressive improvement of post-op pneumothorax | 0
chest tube removed | 168
intermittent fevers | 0
cultures returning negative | 0
afebrile >24 h prior to discharge | 240
discharged | 288
repeat serum cryptococcal antigen test negative | 336
compliant to the 12 week course of itraconazole | 0
levels of itraconazole adjusted | 336
asymptomatic at each follow up | 0
finished course of itraconazole | 1008
reported no return of symptoms | 1008