33 years old | 0
female | 0
admitted to the hospital | 0
papillary thyroid carcinoma | -672
epilepsy | -672
medication for epilepsy | -672
laparoscopic distal gastrectomy | -672
stomach cancer | -672
left hemithyroidectomy | 0
left central compartment neck node dissection | 0
preoperative laboratory findings unremarkable | 0
preoperative ultrasonogram revealed hypoechoic nodule | 0
surgical history of laparoscopic distal gastrectomy | -672
fever | 12
pain at the surgical site | 12
intravenous antipyretics | 12
nausea | 24
tachycardia | 24
high fever | 24
hypotension | 24
septic shock | 24
admitted to the surgical intensive care unit | 24
empirical antibiotics | 24
carbapenem | 24
vancomycin | 24
massive hydration | 24
vasopressors | 24
neck computed tomography scan | 24
chest computed tomography scan | 24
abdomen computed tomography scan | 24
deep neck emphysema | 24
focal pneumomediastinum | 24
infiltration in the anterior neck and mediastinum | 24
abscess formation | 24
exploration of the infected site | 24
edematous changes | 24
massive irrigation | 24
closed-suction drains | 24
bedside thoracostomy | 24
blood cultures | 24
wound cultures | 24
no bacterial growth | 24
general condition stabilized | 168
vital signs stabilized | 168
transferred to the general ward | 168
interval reduction in fluid collection | 168
multidisciplinary approach | 168
video-assisted thoracic surgery | 168
esophagogram | 168
no leakage of the contrast | 168
bronchospasm | 192
retransferred to the surgical ICU | 192
extubated | 216
transferred to the general ward | 216
discharged | 504
infection status acceptable | 8760
follow-up CT scans | 8760
no sign of fluid collection | 8760