abdominal pain | -130
nausea | -130
vomiting | -130
elevated liver enzyme alanine aminotransferase | -130
positive autoimmune antibody | -130
elevated immunoglobulin G | -130
coarse liver surface | -130
liver biopsy | -130
overlap syndrome predominantly with features of an autoimmune hepatitis | -130
high dose of ursodeoxycholic acid | -130
prednisolone 40 mg daily | -130
reduction of prednisolone | -14
azathioprine 50 mg | -6
mild heartburn | -48
abdominal pain worsened | -24
nausea | -24
vomiting | -24
diarrhea | -24
admission to emergency room | 0
abdominal tenderness | 0
mild fever | 0
tachycardia | 0
tachypnea | 0
reduced white blood cells | 0
reduced platelets | 0
decreased neutrophil level | 0
elevated C-reactive protein level | 0
elevated liver enzymes | 0
prothrombin time international normalized ratio | 0
huge stomach with layered wall thickening | 0
air in the stomach wall | 0
decrease of mucosal enhancement | 0
necrotizing gastritis | 0
septic shock | 0
intravenous hydration | 0.5
antibiotic treatment | 0.5
transfer to intensive care unit | 0.5
hypotension | 0.5
inotropics | 1
fluid treatment | 1
increased blood pressure | 2
heart rate slowing | 3
stress-induced cardiomyopathy | 3
ejection fraction of less than 10% | 3
extracorporeal membrane oxygenation | 3
cardiac arrest | 3
pulseless electrical activity | 3
cardiopulmonary resuscitation | 3
death | 3