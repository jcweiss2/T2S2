25 years old | 0
female | 0
presented to the emergency department | -48
returning from Ghana | -48
no prophylactics taken | -48
febrile | -48
diarrhea | -48
hypotension | -48
blood smear positive for malaria | -48
suspected Plasmodium falciparum | -48
normal hemoglobin (15.3 g/dL) | -48
high lactate dehydrogenase (275 IU/L) | -48
discharged with doxycycline | -48
returned to the emergency department | 72
worsening symptoms | 72
inability to tolerate oral medications | 72
chills | 72
nausea | 72
vomiting | 72
dizziness | 72
generalized malaise | 72
admitted to the intensive care unit | 72
diagnosed with septic malaria | 72
diagnosed with influenza | 72
acute kidney injury | 72
creatinine of 2.5 | 72
BUN of 58 | 72
lactate 3.2 | 72
unable to transfer to hospitals with artesunate | 72
hospital acquired intravenous artesunate from CDC | 72
hemoglobin 13.6 g/dL | 72
thrombocytopenic (platelets 12,000) | 72
anemic (Hgb 7.9 g/dL) | 72
received several units of blood | 72
lab tests consistent with hemolytic anemia (reticulocyte count 6.2%, LDH 512 U/L, hematocrit 29.1%) | 96
discharged | 96
followed up with weekly labs for 4 weeks | 240
elevated reticulocyte count | 240
elevated hemoglobin | 240
decreased haptoglobin | 240
decreased lactate dehydrogenase | 240
delayed hemolytic anemia | 240
