68 years old | 0
female | 0
para 3 | 0
postmenopausal bleeding | -672
transvaginal ultrasound scan | -672
endometrial thickness of 5 mm | -672
outpatient hysteroscopy | 0
endometrial biopsy not possible | 0
abdominal pain | 15
nausea | 15
vomiting | 15
fever | 15
sweats | 15
rigors | 15
tachycardic | 15
hypotensive | 15
oxygen saturation of 92% | 15
high vaginal swab sent | 15
bloods in A and E were normal | 15
computed tomography scan of the abdomen and pelvis | 15
desaturation | 16
temperature spiked to 38.1°C | 16
blood pressure falling to 84/48 mm Hg | 16
arterial blood gases done | 16
normal pH | 16
lactate of 3.6 | 16
admitted to the Intensive Treatment Unit | 16
septic shock | 16
inotropic support | 16
started on augmentin | 16
started on metronidazole | 16
stat dose of gentamicin | 16
procalcitonin more than 10.0 μg/L | 16
metronidazole replaced with gentamicin | 24
fever started coming down | 24
lactate levels started decreasing | 24
maximum lactate of 4.25 | 24
stable enough to be stepped down to high dependency unit | 72
augmentin replaced by 1.2 g benzylpenicillin QDS | 72
clindamycin added | 72
inotropes stopped | 72
transferred to the gynecology ward | 72
afebrile | 120
vitals stable | 120
antibiotics switched to oral formulations | 120
discharged home | 192
normal CT scan | 15
no perforation | 15
no pelvic collection | 15
HVS revealed a growth of beta-hemolytic Group A Streptococci | 24
blood cultures revealed a growth of beta-hemolytic Group A Streptococci | 24
diagnosis of septic shock following GAS | 24