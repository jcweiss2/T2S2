65 years old | 0
male | 0
presented to tertiary hospital emergency department | 0
diarrhea | -48
hypotensive | 0
blood pressure 70/40 mmHg | 0
febrile | 0
temperature 38.4 °C | 0
vomited 5 times | -48
brown stools | -48
green stools | -48
denied blood in stool | 0
denied mucous in stool | 0
denied pain | 0
granddaughter with diarrheal illness | -72
contact with granddaughter 1-2 days prior | -72
no significant past medical history | 0
no medication | 0
unvaccinated for rotavirus | 0
distended abdomen | 0
non-tender abdomen | 0
resonant to percussion | 0
bowel sounds audible | 0
clear chest | 0
equal air entry to both lungs | 0
peripheral limb pulses not palpable | 0
cool peripheries | 0
hemoglobin 160 g/L | 0
white cell count 18.1×10⁹/L | 0
platelet count 128×10⁹/L | 0
hypokalemia | 0
potassium 2.7 mmol/L | 0
C-reactive protein 144 mg/L | 0
procalcitonin 235 µg/L | 0
ferritin 2708 µg/L | 0
creatinine 286 µmol/L | 0
raised from baseline creatinine 83 µmol/L | -48
lactate 6.9 mmol/L | 0
sterile blood cultures | 0
sterile urine cultures | 0
negative respiratory swabs | 0
rotavirus detected in feces | 0
negative for norovirus | 0
negative for sapovirus | 0
negative for astrovirus | 0
negative for adenovirus | 0
negative for ova, cysts, parasites | 0
negative for Clostridium difficile | 0
negative cerebrospinal fluid tuberculosis | 0
negative cerebrospinal fluid cryptococcal antigen | 0
negative cerebrospinal fluid cultures | 0
high sensitivity troponin 834 ng/L | 0
serial troponin 1062 ng/L | 24
type-2 acute myocardial infarction | 0
electrocardiogram anteroinferior T-wave inversion | 0
echocardiogram no ventricular dysfunction | 0
echocardiogram no valvular dysfunction | 0
alanine transaminase 1124 U/L | 0
aspartate transaminase 1101 U/L | 0
ischemic liver injury | 0
negative hepatitis screen | 0
negative hepatitis A serology | 0
negative hepatitis B serology | 0
negative hepatitis C serology | 0
negative HIV serology | 0
urinary albumin/creatinine ratio 112.7 mg/mmol | 0
concerns for glomerulonephritis | 0
negative glomerulonephritis screen | 0
acute tubular necrosis | 0
atypical ANCA pattern | 0
negative myeloperoxidase immunofluorescence | 0
negative proteinase-3 immunofluorescence |
