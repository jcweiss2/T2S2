57 years old | 0
    female | 0
    intractable low back pain | 0
    severely impaired mobility | 0
    lumbar laminectomy | -8760
    fusion with posterior spinal instrumentation between L2 and S1 | -8760
    motor strength 4/5 in lower limbs | 0
    decreased sensation in bilateral dermatomes from L1 to S1 | 0
    adjacent segment disease | -8760
    revision surgery of posterior laminectomies (T11-L1) | 0
    posterior spinal fusion with bilateral transpedicular instrumentation from T10 to S1 | 0
    hemovac drain placed into epidural space | 0
    severe headache | 48
    somnolence | 48
    left hemiparesia | 48
    intraprenchymal hemorrhage in right parietal lobe | 48
    subarachnoid hemorrhage | 48
    bilateral symmetrical cerebellar hemorrhages | 48
    pneumocephalus | 48
    hemovac drain removed | 48
    drain exit site closed with single suture | 48
    admitted to Intensive Care Unit | 48
    antiedema treatment (dexamethasone) | 48
    antiepileptic treatment (levatiracetam) | 48
    in-patient rehabilitation | 48
    cognitive impairment | 48
    residual dysphagia | 48
    neurogenic bladder | 48
    referred to nursery clinic for ongoing rehabilitation | 48
    died of aspiration pneumonia | 2160
    sepsis | 2160
    