74 years old | 0
    male | 0
    presented unconscious | 0
    florid shock | 0
    intubation | 0
    initial hemodynamic stabilization | 0
    transferred to cardiac intensive care unit | 0
    presumed devastating cardiac event | 0
    extremis | 0
    initial objective presentation | 0
    usual state of health until two weeks prior | -336
    reactive airway disease began to worsen | -336
    progression of winter | -336
    taking Karo syrup with ephedrine (Forcalide syrup) | -61320
    reactive airway disease | 0
    accidental ingestion of gasoline | -672
    pharmacist prepared Karol-Ephedrine syrup | -61320
    symptoms worsened two weeks prior to admission | -336
    doubled daily intake of Karol-Ephedrine syrup | -336
    respiratory system improved | -336
    returned to usual daily activities | -336
    second week | -168
    dull epigastric pain | -168
    progressed to periodic bouts of extreme pain | -168
    fever | -168
    anorexia | -168
    continued consumption of double dose of Karol-Ephedrine syrup | -168
    disoriented | 0
    febrile | 0
    experiencing constant extreme abdominal pain | 0
    diagnosis of septic shock | 0
    suspicion of abdominal source | 0
    intubated | 0
    sedated | 0
    not chemically paralyzed | 0
    abdomen rigid | 0
    abdomen markedly distended | 0
    progression of severe episodes of epigastric pain | 0
    STAT portable chest radiograph demonstrated massively dilated stomach | 0
    STAT abdominal radiograph demonstrated massively dilated stomach | 0
    decompressed loops of small bowel | 0
    nasogastric tube placed | 0
    rush of air released | 0
    200 ml of blood-stained bilious fluid released | 0
    emergently taken to operating room | 0
    exploratory laparotomy | 0
    more than 3 liters of transudative ascites evacuated | 0
    sepsis | 0
    acute abdomen | 0
    stomach decompressed due to nasogastric tube | 0
    extensive necrosis along greater curvature | 0
    dependent portion of the body of the stomach necrosis | 0
    multiple microperforations along greater curvature | 0
    palpable pulses present in vessels supplying greater curvature | 0
    no evidence of visceral vascular occlusive disease | 0
    subtotal gastrectomy | 0
    Roux-en-Y cardiojejunostomy | 0
    tolerated procedure well | 0
    discharged from hospital | 0
    discontinued use of Karol-Ephedrine syrup | 0
    no complications associated with gastrointestinal ischemia | 0
    chronic gastritis | 0
    microvascular thrombosis | 0
    full thickness necrosis | 0
    multiple gastric perforations | 0
    presence of ephedrine in Karol-Ephedrine syrup | 0
    presence of ephedrine in serum | 0
    hematoxylin and eosin staining demonstrated chronic gastritis | 0
    hematoxylin and eosin staining demonstrated microvascular thrombosis | 0
    hematoxylin and eosin staining demonstrated full thickness necrosis | 0
    hematoxylin and eosin staining demonstrated multiple gastric perforations | 0
    diagnosis of isolated gastric ischemia | 0
    discontinuation of Forcalide syrup | 0
    physicians discontinued prescribing Forcalide syrup | 0
    pharmacy discontinued dispensing Forcalide syrup | 0
    <|eot_id|>
    
  74 years old | 0
male | 0
presented unconscious | 0
florid shock | 0
intubation | 0
initial hemodynamic stabilization | 0
transferred to cardiac intensive care unit | 0
presumed devastating cardiac event | 0
extremis | 0
initial objective presentation | 0
usual state of health until two weeks prior | -336
reactive airway disease began to worsen | -336
progression of winter | -336
taking Karo syrup with ephedrine (Forcalide syrup) | -61320
reactive airway disease | 0
accidental ingestion of gasoline | -672
pharmacist prepared Karol-Ephedrine syrup | -61320
symptoms worsened two weeks prior to admission | -336
doubled daily intake of Karol-Ephedrine syrup | -336
respiratory system improved | -336
returned to usual daily activities | -336
second week | -168
dull epigastric pain | -168
progressed to periodic bouts of extreme pain | -168
fever | -168
anorexia | -168
continued consumption of double dose of Karol-Ephedrine syrup | -168
disoriented | 0
febrile |)