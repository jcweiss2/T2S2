47 years old | 0
male | 0
admitted to the hospital | 0
fever | -72
sore throat | -72
left-sided neck swelling | -72
generalized fatigue | -72
myalgia | -72
blood pressure 100/65 mmHg | 0
heart rate 115 beats/min | 0
temperature 38.9 °C | 0
respiratory rate 20 breath/min | 0
oxygen saturation 100 % | 0
congested throat | 0
left-sided mild posterior lymphadenopathy | 0
high C-reactive protein | 0
slight rise in serum creatinine | 0
high international normalized ratio (INR) | 0
SARS-CoV-2 infection | 0
hydroxychloroquine | 0
azithromycin | 0
cefuroxime | 0
transferred to a quarantine facility | 0
diarrhea | 48
vomiting | 48
mild diffuse abdominal pain | 48
severe abdominal pain | 48
right lower quadrant abdominal pain | 48
low blood pressure | 48
high inflammatory markers | 48
procalcitonin elevation | 48
acute kidney injury | 48
transaminitis | 48
bilateral reticular infiltrates | 48
diffuse abdominal tenderness | 48
guarding | 48
meropenem | 48
resuscitated with crystalloid fluids | 48
transferred to the intensive care unit (ICU) | 48
CT scan of the abdomen | 48
no evidence of bowel perforation | 48
no appendiceal inflammation | 48
diffuse paracolic gutters fat stranding | 48
mild free fluid | 48
bilateral mild pleural effusion | 48
consolidations | 48
filling defect at superior mesentery vein | 48
CT angiogram of the abdomen | 72
no acute thrombosis | 72
major abdominal arterial system patent | 72
high serum lipase | 72
high serum amylase | 72
sepsis workup | 72
blood cultures | 72
urine cultures | 72
sputum cultures | 72
conservative treatment | 72
pain settled | 120
kidney and liver injury improved | 120
inflammatory markers trending down | 120
discharged | 168
follow-up phone call | 168
asymptomatic | 168