79 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
hypertension | 0 | 0 | Factual
ischemic heart disease | 0 | 0 | Factual
severe symptomatic aortic stenosis | 0 | 0 | Factual
coronary artery bypass graft surgery | -7920 | -7920 | Factual
mitral valve repair | -7920 | -7920 | Factual
preprocedural transthoracic echocardiography | -1 | 0 | Factual
severe aortic stenosis | -1 | 0 | Factual
aortic valve area 0.6 cm2 | -1 | 0 | Factual
transvalvular maximal and mean gradients 61 and 33 mm Hg | -1 | 0 | Factual
left ventricular ejection fraction of 45% | -1 | 0 | Factual
right transcarotid approach | 0 | 0 | Factual
fluoroscopic and transesophageal echocardiographic guidance | 0 | 0 | Factual
TEE probe | 0 | 1 | Factual
SAPIEN 3 valve | 0 | 1 | Factual
prosthesis in good position | 1 | 1 | Factual
no visible paravalvular leak | 1 | 1 | Factual
gastric aspiration | 1 | 1 | Factual
blood-tinged secretions | 1 | 1 | Factual
extubated | 1 | 1 | Factual
transferred to the intensive care unit | 1 | 1 | Factual
progressive chest pain | 2 | 2 | Factual
shivering | 2 | 2 | Factual
computed tomography | 2 | 2 | Factual
pneumomediastinum | 2 | 2 | Factual
right hydropneumothorax | 2 | 2 | Factual
esophageal perforation | 2 | 2 | Factual
right thoracic drain | 2 | 2 | Factual
serosanguinous liquid | 2 | 2 | Factual
esophagogastroscopy | 2 | 2 | Factual
4-cm vertical perforation | 2 | 2 | Factual
right thoracotomy | 7 | 7 | Factual
repair of esophageal perforation | 7 | 7 | Factual
primary closure of the esophageal wall | 7 | 7 | Factual
intercostal muscular flap | 7 | 7 | Factual
thoracic drains | 7 | 7 | Factual
pneumonia | 7 | 720 | Factual
severe delirium | 7 | 720 | Factual
congestive heart failure | 7 | 720 | Factual
pulmonary edema | 7 | 720 | Factual
died | 720 | 720 | Factual
vertebral osteophytes | -672 | 0 | Factual
anterior vertebral osteophytes | -672 | 0 | Factual
diffuse idiopathic skeletal hyperostosis | -672 | 0 | Factual
esophageal stricture | 0 | 0 | Negated
Zenker's diverticulum | 0 | 0 | Negated
fibrosis from prior chest radiation | 0 | 0 | Negated
ulceration caused by medication | 0 | 0 | Negated
severe cardiomegaly | 0 | 0 | Negated
large calcified lymph nodes | 0 | 0 | Negated
dysphagia | 0 | 0 | Negated
odynophagia | 0 | 0 | Negated
aspiration | 0 | 0 | Negated
cervical osteophytes | -672 | 0 | Factual
thoracic osteophytes | -672 | 0 | Factual
esophageal compression | -672 | 0 | Possible
esophageal laceration | 0 | 1 | Factual
transesophageal probe | 0 | 1 | Factual
general anesthesia | 0 | 1 | Factual
MitraClip implantation | 0 | 0 | Hypothetical
left atrial appendage occlusion | 0 | 0 | Hypothetical