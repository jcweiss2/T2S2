26 years old | 0
woman | 0
referred to the department | 0
rising levels of human chorionic gonadotropin | 0
intermittent vaginal bleeding | 0
legal medical abortion | -1008
vaginal ultrasound scan confirmed intrauterine pregnancy | -1008
new vaginal ultrasound revealed placental remnants in the uterus | -0
surgical evacuation of the uterus | 0
operation without complications | 0
discharged | 6
readmitted | 24
temperature of 39.5°C | 24
abdominal pain | 24
suspecting severe endometritis | 24
metronidazole administered intravenously | 24
benzylpenicillin administered intravenously | 24
gentamicin administered intravenously | 24
deteriorated within 24 hours | 48
saturation fell to 90% | 48
respiratory rate rose to around 40 breaths per minute | 48
oxygen given by mask | 48
temperature peaked at 40.7°C | 48
C-reactive protein rose to around 300 mg/L | 48
leukocytes rose to around 15 × 10^9/L | 48
moved to the intensive care unit | 48
intubated | 48
rapid deterioration of respiratory function | 48
CT scan performed | 48
thrombophlebitis of the internal jugular vein | 48
hepatomegaly | 48
diagnosed with Lemierre's syndrome | 48
benzylpenicillin discontinued | 48
gentamicin discontinued | 48
tazocin administered | 48
clindamycin administered | 48
metronidazole administered | 48
treated with heparin injections | 48
respiratory support | 672
antibiotics at the intensive care unit | 672
week in standard hospital ward | 1344
recovered | 1680
discharged | 1680
no symptoms from the oropharyngeal tract | 48
blood cultures showed infection with F. necrophorum | 48
F. necrophorum cultivated from the cervix | 48
infection originated from the cervix | 48
Infection following surgical evacuation | 0
common occurrence | 0
common infective agents include Neisseria gonorrhoeae | 0
Chlamydia trachomatis | 0
Gardnerella vaginalis | 0
anaerobic bacteria | 0
infections treated with oral antibiotics | 0
Fusobacterium necrophorum common in urogenital tract | 0
normally not pathogenic | 0
hematogenous spread supported | 48
no symptoms from oropharyngeal tract | 48
F. necrophorum cultivated from cervix | 48
infection reached internal jugular vein | 48
spread hematogenously | 48
pulmonary embolisms | 48
arthritis | 48
abscesses | 48
early diagnosis crucial | 48
correct treatment crucial | 48
CT of neck and lungs diagnostic | 48
antibiotic treatment with metronidazole and beta-lactamase inhibitor | 48
anticoagulation considered | 48
respiratory support necessary | 48
surgical drainage of abscesses necessary | 48
patient consent to publication | 0
no conflict of interest | 0
