70 years old | 0
female | 0
admitted to the hospital | 0
symptom onset of weakness | -48
polyuria | -48
elevated blood glucose | -48
syncope | 0
negative RT-PCR swab for COVID-19 | 0
prophylactic anticoagulation started | 0
transthoracic echocardiogram | 24
dilated right ventricle | 24
computed tomography pulmonary angiogram | 48
pulmonary embolism | 48
clot in transit | 48
therapeutic anticoagulation started | 48
repeat RT-PCR swab for COVID-19 returns positive | 48
transferred for percutaneous aspiration thrombectomy with AngioVac | 48
patient died during the procedure | 72
hypertension | 0
hyperlipidaemia | 0
diabetes | 0
supraventricular tachycardia | 0
denies fever | 0
denies chills | 0
denies sore throat | 0
denies cough | 0
denies chest pain | 0
denies dyspnoea | 0
initial blood pressure 84/55 mmHg | 0
pulse 72 b.p.m. | 0
oxygen saturation 88% on room air | 0
respiratory rate 16/min | 0
temperature 36.6°C | 0
no jugular venous distension | 0
normal heart and lung sounds | 0
no peripheral oedema | 0
blood pressure and oxygenation improved | 24
hydration | 24
insulin | 24
antibiotics | 24
prophylactic dose anticoagulation | 24
droplet precautions | 24
contact isolation | 24
differential diagnosis included hypovolaemia | 24
differential diagnosis included sepsis | 24
syncope and hypoxaemia | 24
suspicion for acute PE | 24
myocardial infarction | 24
arrhythmia | 24
heart failure | 24
underlying COVID-19 suspected | 24
chest X-ray unremarkable | 24
head computed tomography unremarkable | 24
electrocardiogram showed sinus rhythm | 24
S1, Q3, T3 pattern | 24
prolonged QTc | 24
T-wave inversions | 24
hyperglycaemia | 24
elevated anion gap | 24
serum creatinine | 24
lactate | 24
D-dimer | 24
C-reactive protein | 24
pro-BNP | 24
INR | 24
serial troponin T-tests negative | 24
urine positive for ketones | 24
urine positive for white cells | 24
initial nasopharyngeal swab for COVID-19 negative | 0
bedside echocardiogram | 24
moderately dilated right ventricle | 24
mild hypokinesis | 24
elevated right ventricular systolic pressure | 24
patient remained comfortable | 24
haemodynamically stable | 24
saturation 98% on 3 L of oxygen | 24
dyspnoea | 48
desaturation | 48
pulse 80 b.p.m. | 48
blood pressure 132/78 mmHg | 48
computed tomography pulmonary angiogram | 48
saddle PE | 48
bilateral filling defects | 48
thrombus in the right atrium | 48
repeat echo | 48
highly mobile clot in transit | 48
repeat nasopharyngeal swab for COVID-19 positive | 48
therapeutic dose anticoagulation | 48
intravenous heparin | 48
transferred to intensive care unit | 48
evaluated by multidisciplinary institutional Pulmonary Embolism Response Team | 48
percutaneous aspiration thrombectomy with adjunctive intra-pulmonary and catheter-directed thrombolysis | 48
AngioVac device | 72
patient decompensated | 72
rescue thrombectomy | 72
Inari FlowTriever device | 72
intra-pulmonary and systemic thrombolysis | 72
patient arrested | 72
patient died | 72