8-year-old boy | 0
admitted to the hospital (regional) | 0
flame burn injury | 0
intubated | 0
ventilated | 0
burns debridement | 0
Total Body Surface Area affected by burns (61%) | 0
retrieved to tertiary PICU (LCCH) | -24
donor sites harvested | 72
burns debrided | 72
significant blood loss | 72
no grafting completed | 72
Split Skin Graft (SSG) on day 6 | 144
SSG posterior torso | 144
SSG buttocks | 144
SSG posterior upper thighs | 144
SSG right lower leg | 144
SSG bilateral upper arms | 144
post-operative orders requiring ventilation | 144
post-operative orders requiring deep sedation | 144
post-operative prone positioning | 144
minimal movement allowed | 144
avoidance of shear forces over graft sites | 144
sepsis on day 6 | 144
systemic inflammatory response | 144
respiratory deterioration | 144
difficult ventilation | 144
chest x-ray showing multifocal atelectasis | 144
no spontaneous cough | 144
increasing ventilator requirements | 144
raised peak inspiratory pressures | 144
retained secretions | 144
systemic unwellness | 144
hemodynamic instability | 144
episodes of hypotension | 144
requiring fluid resuscitation | 144
requiring inotropes | 144
conventional physiotherapy techniques limited | 144
repositioning using bed tilt | 144
manual hyperinflation | 144
saline lavage | 144
suction | 144
passive joint mobility | 144
limited effectiveness | 144
secretions remaining difficult to access | 144
palpable secretions post intervention | 144
MetaNeb® implementation | 144
consultation with LCCH PICU Medical Consultants | 144
consultation with USA centers | 144
MetaNeb® attached to oxygen source | 144
open-ended bagging circuit (FiO2 1.0) | 144
Continuous High Frequency Oscillation mode (230 bpm) | 144
10-minute treatments | 144
occlusion ring placement | 144
inline nebuliser with normal saline | 144
pressure maintained (10-20 cmH2O) | 144
variable volume breaths | 144
secretion mobilization evaluated | 144
reconnection to bagging circuit | 144
manual hyperinflation with expiratory flow bias | 144
suction via ETT | 144
treatment cycle repeated | 144
secretions no longer palpable | 144
ETT mucus clearance minimal | 144
outcome measures: sputum volume | 144
outcome measures: sputum quality | 144
outcome measures: CXR | 144
outcome measures: PIP values | 144
vital signs monitoring | 144
transient blood pressure decrease (MAP <10 mmHg) | 144
recovery without intervention | 144
4 days of treatment (twice daily) | 168
resolution of focal CXR changes | 168
reduction in secretions | 168
reduction in PIP (25%) | 168
extubation without incident | 168
MetaNeb® via mouthpiece trialled post-extubation | 168
poorly tolerated | 168
discontinued due to behavioral issues | 168
lip pain | 168
lip swelling | 168
inhibited lip seal | 168
skin grafting on day 17 | 408
required intubation | 408
required ventilation | 408
required immobility | 408
MetaNeb® utilized during second phase | 408
optimized secretion clearance | 408
decreased risk of retained secretions | 408
decreased risk of lung infection | 408
no respiratory deterioration | 408
successful extubation | 408
conflict of interest (Hill-Rom funding) | 0
