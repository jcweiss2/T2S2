30 years old | 0
African American | 0
female | 0
admitted to the hospital | 0
shortness of breath on exertion | 0
chest pain with deep inspiration | 0
no recent infections | 0
physical examination did not yield any abnormalities | 0
VQ scan indicated high probability for pulmonary emboli | 0
pulmonary emboli in her right lobe | 0
chest x ray showed possible development of small bilateral pleural effusions | 0
multiple nodular opacities scattered throughout the lungs | 0
CT scan of the abdomen showed moderate alveolar consolidation | 0
pulmonary infarct or pneumonia | 0
EKG was normal | 0
2D echocardiograms were normal | 0
no indication of endocarditis | 0
Heparin drip was initiated | 0
high fevers during her hospital stay | 24
tachycardia | 24
blood cultures were positive | 24
Gram positive cocci in pairs and clusters | 24
Staphylococcus species | 24
S. caprae | 24
vancomycin was started | 24
S. aureus was ruled out | 48
antibiotics were changed to Kefzol | 48
fever resolved | 72
significant clinical improvement | 72
urinalysis indicated the presence of E. coli | 72
E. coli was sensitive to all 17 antimicrobial agents | 72
Ciprofloxacin was administered | 72
treated the urinary tract infection | 96
echocardiogram did not reveal any evidence of endocarditis | 96
no indication that the patient recently visited a farm | 0
no contact with goats | 0
no transplants | 0
no internal fixation for orthopedic prosthesis | 0
no foreign subject implants | 0
discharged | 120