31 years old | 0
female | 0
SLE | -8760
stage IV lupus nephritis | -8760
prior stroke | -8760
intravenous drug use | -8760
cardiogenic shock | 0
mental status changes | 0
elevated jugular venous pressure | 0
prominent v wave | 0
body temperature 36.3°C | 0
blood pressure 95/66 mm Hg | 0
heart rate 94 beats/min | 0
hemoglobin 10.3 g/dL | 0
white blood cell count 18.9 × 10^9/L | 0
platelet count 64 × 10^9/L | 0
international normalized ratio 3.6 | 0
creatinine level 1.7 mg/dL | 0
drug studies positive for narcotics | 0
drug studies positive for cannabis | 0
antiphospholipid serology normal | 0
blood cultures negative | 0
infectious endocarditis considered | 0
broad-spectrum intravenous antibiotics | 0
mitral valve replacements | -720
NBTE | -720
aggressive immunosuppression | -720
anticoagulation | -720
dehisced mitral valve prosthesis | 0
severe mitral regurgitation | 0
perivalvular regurgitation | 0
annular pseudoaneurysm | 0
fourth sternotomy | 24
mitral valve annulus reconstruction | 24
bioprosthesis integration | 24
left atrial dome reconstruction | 24
interatrial septal incision reconstruction | 24
postbypass TEE | 24
extracorporeal membrane oxygenation | 24
left ventricular ejection fraction 25% | 24
sluggish flow in left atrium | 24
multiple blood product transfusions | 24
layered thrombus in left atrium | 120
surgical clot removal | 120
thrombus reaccumulation | 120
extracorporeal membrane oxygenation withdrawn | 120
death | 120
autopsy declined | 120