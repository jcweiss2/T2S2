19 years old | 0
    male | 0
    mild asthma | 0
    scratched by a cat | 0
    fever | 0
    deep venous thrombosis in left leg | 0
    fondaparinux | -168
    apixaban | -168
    macroscopic hematuria | -48
    leg edema | -48
    asthenia | -48
    persistent fever | -48
    lethargic | 0
    Glasgow Coma Scale 15/15 | 0
    blood pressure 100/66 mm Hg | 0
    sinus tachycardia 120 beats per minute | 0
    mitral murmur | 0
    hemocultures taken | 0
    piperacillin started | 0
    ceftriaxone/gentamicin | 24
    Haemophilusparainfluenzae | 24
    hemoglobin 6.3 g/dL | 0
    red blood cells transfused | 0
    anterograde amnesia | 0
    cerebral computed tomography | 0
    nuclear magnetic resonance scan | 0
    large hematoma in left occipitoparietal region | 0
    multiple bilateral microhemorrhage | 0
    hematoma next to right cerebellum | 0
    hematoma in right occipital region | 0
    multiple ischemic microlesions | 0
    left cerebellar ischemic stroke | 0
    intracerebral mycotic aneurysm of left posterior cerebral artery | 0
    embolization | 0
    transthoracic echocardiography | 0
    large vegetation 20 mm | 0
    mobile echo dense masses >15 mm on mitral valve | 0
    significant mitral valve prolapse | 0
    septic shock | 0
    intubated | 0
    sedated | 0
    norepinephrine started | 0
    dobutamine started | 0
    wake-up test | 0
    obeying commands | 0
    no neurological deficits | 0
    emergency surgery | 48
    minimal cardiopulmonary bypass (MCBP) | 48
    right radial arterial line | 48
    left internal jugular central venous line | 48
    intubated | 48
    ventilated | 48
    sedated with propofol | 48
    sedated with sufentanil | 48
    hemodynamically supported with norepinephrine | 48
    tranexamic acid 1 g intravenously | 48
    tranexamic acid infusion 10 mg/kg/h | 48
    MCPB primed with lactated Ringer’s solution | 48
    retrograde priming technique | 48
    Hb dropped to 7.8 | 48
    hematocrit 23% | 48
    red blood cells transfused | 48
    Hb 8.5–8.8 g/dL | 48
    hematocrit 25%–26% | 48
    mean arterial blood pressure above 70 mm Hg | 48
    norepinephrine peak infusion rate 1 mg/h | 48
    anterograde cold cardioplegia | 48
    retrograde cold cardioplegia | 48
    central body temperature cooled to 33°C | 48
    temperature increased to 36.8°C | 48
    transesophageal echocardiography | 48
    large vegetations | 48
    damage of mitral annulus | 48
    biological mitral valve replacement | 48
    cerebral oximetry above 60 | 48
    right hemisphere oxygen saturation 53 | 48
    activated clotting time 133 seconds | 48
    heparin 10,000 units | 48
    ACT peak 401 seconds | 48
    ACT 283 seconds | 48
    ACT 289 seconds | 48
    protamine 100 mg | 48
    ACT normalized 126 seconds | 48
    MCBP time 74 minutes | 48
    aortic clamping time 56 minutes | 48
    MCBP weaning 18 minutes | 48
    atrioventricular pacemaker stimulation | 48
    fresh frozen plasma transfused | 48
    platelets transfused | 48
    transferred to intensive care unit | 48
    norepinephrine 0.032 mg/h | 48
    reoperation to remove thromboemboli from left popliteal artery | 432
    ventilation-acquired pneumonia | 432
    tracheostomy | 432
    percutaneous gastric feeding | 432
    rehabilitation medicine | 672
    good neurological recovery | 672
    no loss in memory capacity | 672
    no neurological deficits | 672
    discharged home | 672
    bilateral emboli into legs | 672
    residual bilateral claudication | 672
    control nuclear magnetic resonance | 672
    resorption of occipital hematoma | 672
    resorption of left cerebellar hematoma | 672
    