54 years old | 0
male | 0
presented to the hospital | 0
pre-syncope | 0
syncope lasting <5 min | 0
sudden onset | 0
left-sided chest tightness | 0
chest tightness self-resolved after 2 min | 0
under review by general practitioner | -2928
generalized fatigue | -2928
weight loss | -2928
physical examination | 0
weight of 41 kg | 0
blood pressure of 96/60 mm Hg |; 0
unremarkable cardiac examination | 0
unremarkable respiratory examination | 0
diffuse erythematous rash in left lower limb | 0
electrocardiography demonstrated normal sinus rhythm | 0
raised troponin concentration of 1,268 ng/l | 0
eosinophil count of 7.6 × 109/l | 0
referred to cardiology | 0
review at cardiac center | 0
myocarditis diagnosis | 0
CMR imaging showed eosinophilic myocarditis | 0
coronary angiography revealed no coronary artery disease | 0
working diagnosis of EM | 0
secondary causes sought | 0
decision to perform skin biopsy | 0
cardiac biopsy considered | 0
improved clinically | 0
discharged | 0
prescriptions for edoxaban | 0
prescriptions for prednisolone | 0
scheduled follow-up in rheumatology clinic in 2 weeks | 0
missed follow-up appointment | 432
presented to cardiology clinic 2 months later | 432
neck swelling | 432
urgently admitted to hospital | 432
eosinophil count rise to 19.7 × 109 cells/l | 432
decision to increase prednisolone dose | 432
CT neck demonstrated lymphadenopathy | 432
lymphadenopathy confirmed as T-cell lymphoma on biopsy | 432
decision for chemotherapy with cyclophosphamide | 432
deteriorated from sepsis secondary to cholecystitis | 432
new onset seizures | 432
reduction in consciousness with GCS 9/15 | 432
head CT demonstrated multiple bilateral acute infarctions | 432
infarct areas not amenable to thrombectomy | 432
GCS score continued to deteriorate | 432
transferred to intensive care unit | 432
investigations for bilateral cerebral infarcts | 432
medical history: hepatitis B | 0
medical history: asthma | 0
medical history: intravenous drug use | 0
medical history: excessive alcohol use | 0
differential diagnosis: ischemic stroke secondary to EM | 432
differential diagnosis: reduced GCS score | 432
differential diagnosis: seizures | 432
differential diagnosis: intracranial bleeding | 432
differential diagnosis: malignancy | 432
differential diagnosis: intracerebral infection | 432
CMR demonstrated subendocardial late gadolinium enhancement | 432
CMR showed increased signal on STIR images | 432
mild LV systolic impairment (EF 50%) | 432
skin biopsy revealed eczematous changes | 432
bone marrow biopsy revealed no increase in eosinophils | 432
axillary lymph node biopsy confirmed T-cell lymphoma | 432
head CT revealed frontal infarcts | 432
head CT revealed parietal infarcts | 432
head CT revealed left temporo-occipital infarcts | 432
critical care echocardiography demonstrated apical tear | 432
preserved apical architecture suggestive of intramural tear | 432
small apical cavity in continuity with LV cavity | 432
small mobile structures attached to dissected myocardium | 432
color flow Doppler revealed diastolic flow in apical cavity | 432
pulse wave Doppler demonstrated diastolic flow into apical cavity | 432
pulse wave Doppler demonstrated systolic flow out of apical cavity | 432
cyclophosphamide therapy begun | 432
partial response to cyclophosphamide | 432
eosinophil count reduction to 20-30 × 109 cells/l | 432
multidisciplinary team decision for palliation | 432
poor prognosis | 432
