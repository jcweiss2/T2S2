49 years old | 0
male | 0
admitted to the hospital | 0
bronchiectasis | -672
fibrosis of the middle lobe | -672
dyspnea | -72
recurrent hemoptysis | -72
nonproductive cough | -72
conservative management | -72
progressive decrease in physical endurance | -72
deterioration of the quality of life | -72
CT scan of the chest | -24
fibroatelectasis of the right middle lobe | -24
echocardiography | -24
large atrial septal defect | -24
biventricular enlargement | -24
severe mitral and tricuspid regurgitation | -24
mitral prolapse | -24
moderate pulmonary artery hypertension | -24
multidisciplinary evaluation | -12
simultaneous procedure proposed | -12
thoracoscopic uniportal cardiac intervention | -12
lobectomy | -12
written informed consent | -12
single 4 cm thoracoport placed | 0
femoral artery and vein cannulation | 0
CPB | 0
position of the venous cannula confirmed | 0
cross-clamping of the aorta | 0
antegrade cardioplegia | 0
approach to the right atrium and interatrial septum | 0
mitral valve ring annuloplasty | 0
De Vega annuloplasty of the tricuspid valve | 0
closure of the interatrial septal defect | 0
heparin reversal | 0
middle lobe vein isolated | 0
middle lobe vein tied | 0
middle lobe vein clipped | 0
middle lobe vein transected | 0
middle lobe bronchus and artery divided | 0
parenchymal bridge between the middle and upper lobes divided | 0
surgery completed | 332
extubated | 3
transferred from the intensive care unit | 24
chest tube removed | 96
discharged home | 192
follow-up | 7200
exercise tolerance improved | 7200
hemoptysis resolved | 7200
normalization of the cardiac chamber dimensions | 7200
absence of regurgitation | 7200