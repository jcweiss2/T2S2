41 years old | 0
female | 0
admitted to the hospital | 0
ischemic stroke | -72
right hemiplegia | -72
Broca’s aphasia | -72
dizziness | 48
vomiting | 48
Kussmaul breathing | 48
lowered response to verbal commands | 48
hyperglycemia | 48
metabolic acidosis | 48
DKA | 48
arterial blood gas analysis | 48
urine analysis | 48
ketone 3+ | 48
aggressive hydration | 48
insulin pump | 48
bicarbonate infusion | 48
electrolyte correction | 48
transferred to the intensive care unit | 48
serum ketone body | 72
metabolic acidosis with respiratory compensation | 72
comatose | 120
hemodynamic instability | 120
brain MRI | 120
acute infarction lesions | 120
brain swelling of infarction lesions | 120
midline shift | 120
occlusion of bilateral ICA | 120
glycerol | 120
endotracheal intubation | 120
echocardiograms | 120
normal left ventricle contractility | 120
no evidence of thrombus or vegetation formation | 120
mechanical ventilation | 120
coma | 120
respiratory failure | 120
severe hyperglycemia | 120
compassionate extubation | 696
expired | 696
T1DM | -7440
hypertension | -2190
hyperlipidemia | -1752
hyperthyroidism | -1092
methimazole | -1092
aspirin | -1092
atorvastatin | -1092
regular subcutaneous insulin injections | -1092
medical control | -1092
right central facial palsy | 0
right hemiplegia | 0
Brunnstrom stage | 0
functional status | 0
ambulate with use of a quad cane | 0
feed herself | 0
Broca’s aphasia | 0
body temperature | 0
pulse | 0
blood pressure | 0
breathing | 0
neurological examinations | 0
glycohemoglobin level | 48
hyperglycemia | 48
normal thyroid function | 48
urine analysis | 48
ketonuria | 48
pyuria | 48
blood examinations | 48
arterial blood gas analyses | 48
thyroid function | 48
stroke survey | 120
bilateral MCA and bilateral ACA territory infarction | 120
BICAO | 120
T1DM with DKA | 120
aggressive hydration | 48
insulin pumping | 48
electrolyte correction | 48
vasopressors | 120
glycerol | 120
mechanical ventilation | 120
coma | 120
respiratory failure | 120
severe hyperglycemia | 120
poor prognosis | 696
compassionate extubation | 696
expired | 696
bilateral internal carotid artery occlusion | -72
ischemic stroke | -72
left corona radiata | -72
bilateral frontal lobe | -72
parietal lobe | -72
inpatient rehabilitation programs | -72
no major accidents | -72
recurrent stroke | -72
urinary tract infection | -72
pneumonia | -72
transferred to our ward | 0
further rehabilitation | 0
significant right hemiplegia | 0
ambulate with use of a quad cane | 0
alert | 0
Broca’s aphasia | 0
dizziness | 48
vomiting | 48
Kussmaul breathing | 48
lowered response to verbal commands | 48
hyperglycemia | 48
persisted | 48
arterial blood gas analysis | 48
metabolic acidosis | 48
pH | 48
PCO2 | 48
HCO3- | 48
base excess | 48
urine analysis | 48
ketone 3+ | 48
DKA | 48
suspected | 48
transferred to the intensive care unit | 48
aggressive hydration | 48
insulin pump | 48
bicarbonate infusion | 48
electrolyte correction | 48
serum ketone body | 72
metabolic acidosis with respiratory compensation | 72
comatose | 120
hemodynamic instability | 120
brain MRI | 120
acute infarction lesions | 120
brain swelling of infarction lesions | 120
midline shift | 120
occlusion of bilateral ICA | 120
glycerol | 120
endotracheal intubation | 120
echocardiograms | 120
normal left ventricle contractility | 120
no evidence of thrombus or vegetation formation | 120
mechanical ventilation | 120
coma | 120
respiratory failure | 120
severe hyperglycemia | 120
compassionate extubation | 696
expired | 696