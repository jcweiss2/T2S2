48 years old | 0
woman | 0
G6P2042 | 0
presented to the emergency department | 0
fever | -360
chills | -360
diffuse abdominal pain | -360
uterine artery embolization | -360
uterine fibroids | -360
abnormal uterine bleeding | -360
dysmenorrhea | -360
hypertension | 0
obesity class III | 0
cholecystectomy |>
thyroidectomy | 0
left knee meniscal repair | 0
temperature of 101.5F | 0
heart rate of 110 beats per minute | 0
respiratory rate of 24–37 breaths per minute | 0
distended abdomen | 0
diffusely tender abdomen | 0
scant blond‑tinged vaginal discharge | 0
white blood cell count of 26,300 | 0
91% neutrophils | 0
computed tomography of abdomen and pelvis | 0
distended uterus | 0
intra-cavitary uterine masses | 0
gas in uterus | 0
air–fluid level | 0
sepsis | 0
pyomyoma | 0
broad-spectrum intravenous antibiotics | 0
Cefepime | 0
flagyl | 0
amikacin | 0
fluid resuscitation | 0
lactated ringers | 0
exploratory laparotomy | 0
hysterectomy | 0
bilateral salpingectomy | 0
small bowel resection | 0
primary end-to-end anastomosis | 0
frozen section of uterus | 0
negative for malignancy | 0
ovaries spared | 0
post-operative transfer to surgical intensive care unit | 0
prolonged course of antibiotics | 0
discharged from hospital | 504
incidental finding of poorly differentiated serous carcinoma of the fallopian tube | 504
staging procedure | 720
stage 1a fallopian tube carcinoma | 720
following up with oncology service | 720
