24 years old | 0
female | 0
26 weeks pregnant | 0
admitted to the emergency department | 0
abdominal pain | -120
abdominal distension | -120
constipation | -120
increasing severity of abdominal pain | -120
no significant past medical or surgical history | 0
uneventful menstrual and antenatal history | 0
dehydrated | 0
hypotension | 0
tachycardia | 0
tachypnea | 0
asymmetrically distended abdomen | 0
tenderness all over the abdomen | 0
empty rectum on digital examination | 0
vaginal examination not suggestive of threatened preterm labour | 0
elevated white cell count | 0
clear urine analysis | 0
distended bowel loop on ultrasound scan | 0
moderate amount of free fluid in the peritoneal cavity | 0
single viable fetus | 0
dilated large bowel on abdominal X-ray | 0
abnormal gas pattern on abdominal X-ray | 0
coffee bean appearance on abdominal X-ray | 0
sigmoid volvulus on abdominal X-ray | 0
sigmoidoscopy | 0
twisted sigmoid colon on sigmoidoscopy | 0
failure to negotiate the obstruction on sigmoidoscopy | 0
foetal distress | 0
deceleration in heart rate | 0
decision to perform caesarean section | 0
decision to explore the abdomen for IO | 0
initial resuscitation | 0
taken to the emergency theatre for laparotomy | 0
midline laparotomy | 0
enormously distended sigmoid loop | 0
ischemic and gangrenous changes | 0
no signs of perforation | 0
necrosis due to twisted sigmoid mesocolon | 0
gangrenous colon displaced posteriorly by the pregnant uterus | 0
lower segment caesarean section | 0
delivery of a male preterm infant | 0
preterm infant weighing 750 g | 0
admitted to the neonatal ICU | 0
mechanical ventilation due to lung immaturity | 0
resection of the gangrenous sigmoid colon | 0
Hartmann’s procedure | 0
end colostomy | 0
closure of the rectal stump | 0
uneventful post-operative course | 0
discharged home on the 9th post-operative day | 216
child discharged home after 10 weeks in the neonatal ICU | 720
reversal of Hartmann’s procedure | 4320
bowel continuity restored through colo-rectal anastomosis | 4320