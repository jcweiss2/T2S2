20 years old | 0
female | 0
exposure to upper tract respiratory infection | -168
cough | -72
yellow sputum | -72
intermittent fever | -72
night sweats | -72
dyspnea | -24
admitted to urgent care | 0
community acquired pneumonia | 0
antibiotics initiated | 0
admitted to ICU | 0
denies GI symptoms | 0
denies rash | 0
denies arthralgia | 0
denies thromboembolic disease | 0
denies chest pain | 0
denies leg pain | 0
denies leg swelling | 0
oral contraceptive | 0
intubation | 72
non-invasive positive pressure ventilation failed | 72
severe hypoxemia | 0
arterial blood gas testing | 0
chest X-ray revealed diffuse bilateral opacities | 0
enterovirus/rhinovirus detected | 0
high PEEP | 0
low tidal volume ventilation | 0
hypoxemia | 0
hypercapnia | 0
ECMO initiated | 72
vancomycin | 0
piperacillin-tazobactam | 0
levofloxacin | 0
high-dose intravenous vitamin C initiated | 72
AP chest X-ray imaging | 120
improvement in bilateral lung opacities | 120
bronchoscopy | 168
negative for bacterial or fungal respiratory pathogens | 168
histoplasma antigen negative | 168
blastomyces antigen negative | 168
aspergillus antigen negative | 168
legionella antigen negative | 168
furosemide | 168
daily negative fluid balance | 168
lung gas exchange improved | 168
ECMO decannulation | 168
extubation | 168
vitamin C dosing reduced | 168
discharged home | 288
follow-up exam | 720
completely recovered | 720
follow-up chest X-ray film | 720