32 years old | 0
female | 0
admitted to the hospital | 0
fever | -840
rash | -720
cough | -840
treated with cefalexin | -840
cefalexin stopped | -785
itchy rash appeared | -720
fever returned | -720
hospitalized | 0
diagnosed with erythema multiforme | 0
weight-loss capsule | -720
antiallergic treatment | 0
prednisone | 0
levofloxacin | 0
cefuroxime | 0
yellowish watery diarrhea | 6
infectious diarrhea | 6
treated with Bifidobacterium | 6
diarrhea got worse | 12
transferred to ICU | 12
signs of MOF | 12
FMT treatment plan | 12
high-dose intravenous methylprednisolone | 12
intravenous immune globulin | 12
anti-EBV and CMV treatment | 12
ganciclovir | 12
FMT | 12
first FMT | 12
second FMT | 18
body temperature dropped | 18
MODS symptoms recurred | 18
blood cultures remained sterile | 18
third FMT | 24
stool output declined | 24
stools became well-formed | 24
fourth FMT | 30
frequency and volume of stools returned to normal | 30
inflammatory markers reduced | 18
CRP reduced | 18
PCT reduced | 18
ESR reduced | 18
IL-6 reduced | 18
aspartate aminotransferase decreased | 30
alanine aminotransferase decreased | 30
level of consciousness improved | 30
EBV and CMV DNA levels returned to normal | 30
discharged | 1440
abdominal CT scan | 0
thickening of the walls of the small intestine | 0
hepatosplenomegaly | 0
normal-sized abdominal lymph nodes | 0
intestinal flora examination | 0
decreased levels of beneficial bacteria | 0
Bifidobacterium | 0
Lactobacillus | 0
Clostridium | 0
antibiotic treatment stopped | 12
FMT procedures | 12
donor feces infusion | 12
total of 4 FMT | 12
FMT frequency | 12
once every 6 days | 12
serum inflammatory markers analysis | 12
IL-6 examined | 12
PCT analyzed | 12
CRP analyzed | 12
ESR analyzed | 12
statistical analysis | 30
linear regression analysis | 30
Pearson test | 30
OTU analysis | 30
PC analysis | 30
CANOCO software | 30
P value | 30
intestinal microflora analysis | 30
16S rRNA gene-based sequencing | 30
genomic DNA isolated | 30
DNA samples examined | 30
NanoDrop spectrophotometer | 30
agarose gel electrophoresis | 30
V3V4 regions amplified | 30
PCR products purified | 30
sequencing library prepared | 30
TruSeq DNA Kit | 30
Illumina MiSeq sequencer | 30
QIIME pipeline | 30
raw sequences processed | 30
tags clustered | 30
OTUs assigned | 30
Greengenes database | 30
bacterial composition analyzed | 30
phyla | 30
classes | 30
orders | 30
families | 30
genera | 30
principal component analysis | 30
bacterial genera | 30
clustering tree | 30
Firmicutes phylum increased | 36
Bacteroidetes phylum increased | 39
Proteobacteria phylum decreased | 39
Lachnospiraceae family enriched | 39
Ruminococcaceae family enriched | 39
Veillonellaceae family enriched | 39
Roseburia increased | 39
Dialister increased | 39
Prevotella increased | 39
Bacteroides increased | 39
Oscillospira increased | 39
Faecalibacterium increased | 39
intestinal failure | 0
DIHS | 0
MODS | 12
MOF | 12
severe diarrhea | 6
FMT effective | 30
intestinal microflora restored | 30
microecological balance restored | 30
intestinal barrier function restored | 30
mucosal barrier function restored | 30
Bifidobacteria increased | 30
Lactobacillus increased | 30
Bacteroides increased | 30
Escherichia coli decreased | 30
B/E ratio restored | 30
anaerobic to aerobic bacteria ratio restored | 30
intestinal microflora analysis | 30
16S rRNA gene-based sequencing | 30
genomic DNA isolated | 30
DNA samples examined | 30
NanoDrop spectrophotometer | 30
agarose gel electrophoresis | 30
V3V4 regions amplified | 30
PCR products purified | 30
sequencing library prepared | 30
TruSeq DNA Kit | 30
Illumina MiSeq sequencer | 30
QIIME pipeline | 30
raw sequences processed | 30
tags clustered | 30
OTUs assigned | 30
Greengenes database | 30
bacterial composition analyzed | 30
phyla | 30
classes | 30
orders | 30
families | 30
genera | 30
principal component analysis | 30
bacterial genera | 30
clustering tree | 30
FMT treatment | 12
FMT effective | 30
intestinal microflora restored | 30
microecological balance restored | 30
intestinal barrier function restored | 30
mucosal barrier function restored | 30
Bifidobacteria increased | 30
Lactobacillus increased | 30
Bacteroides increased | 30
Escherichia coli decreased | 30
B/E ratio restored | 30
anaerobic to aerobic bacteria ratio restored | 30
DIHS diagnosed | 0
DIHS treatment | 12
FMT effective | 30
intestinal microflora restored | 30
microecological balance restored | 30
intestinal barrier function restored | 30
mucosal barrier function restored | 30
Bifidobacteria increased | 30
Lactobacillus increased | 30
Bacteroides increased | 30
Escherichia coli decreased | 30
B/E ratio restored | 30
anaerobic to aerobic bacteria ratio restored | 30
MODS treated | 12
MOF treated | 12
severe diarrhea treated | 12
FMT effective | 30
intestinal microflora restored | 30
microecological balance restored | 30
intestinal barrier function restored | 30
mucosal barrier function restored | 30
Bifidobacteria increased | 30
Lactobacillus increased | 30
Bacteroides increased | 30
Escherichia coli decreased | 30
B/E ratio restored | 30
anaerobic to aerobic bacteria ratio restored | 30