30 years old | 0
female | 0
anorexia nervosa | -8760
body mass index 11 kg/m2 | 0
nausea | -72
vomiting | -72
diarrhea | -72
abdominal pain | -72
previous hospitalisations | -720
severe weakness | -720
electrolyte disbalance | -720
anemia | -720
emaciated | 0
dehydrated | 0
distended abdomen | 0
generalized peritonitis | 0
hypovolemic shock | 0
heart rate 92/min | 0
blood pressure 70/30 mmHg | 0
hypothermic 34.3 °C | 0
tachypneic up to 30/min | 0
oxygen saturation 98% | 0
metabolic acidosis | 0
electrolyte derangement | 0
sodium 116 mmol/L | 0
potassium 3.9 mmol/L | 0
chloride 85 mmol/L | 0
bicarbonate 10 mmol/L | 0
blood urea nitrogen 94 mg/dL | 0
anion gap 21 mmol/L | 0
creatinine 3.01 mg/dL | 0
microcytic anemia | 0
white blood cell count 14,200/mm3 | 0
hemoglobin 10.7 g/dL | 0
hematocrit 31% | 0
mean corpuscular volume 73 fL | 0
platelets 546,000 /mm3 | 0
abdominal X-ray | 0
computer tomography scan | 0
extensive portal venous gas | 0
bowel wall pneumatosis | 0
aggressive resuscitation | 0
intravenous crystalloids | 0
infusion of sodium bicarbonate | 0
nasogastric tube | 0
broad spectrum systemic antibiotics | 0
admission to the intensive care unit | 0
hemodynamic status unstable | 3
addition of vasoactive agents | 3
exploratory laparotomy | 6
bowel resection | 6
control of sepsis source | 6
necrosis of the entire small bowel | 6
necrosis of the right hemicolon | 6
death | 6