62 years old | 0
female | 0
total abdominal hysterectomy | -672
bilateral salpingo-oophorectomy | -672
uterine fibroid | -672
endometrial polyp | -672
ovarian cyst | -672
incisional hernia | -672
laparoscopic dual mesh repair | -504
severe abdominal pain | 0
abdominal wall tenderness | 0
erythema | 0
urgent contrast Computed Tomography | 0
urinary bladder perforation | 0
surgical emphysema | 0
necrotizing fasciitis | 0
emergency debridement | 0
intra-operation cystoscopy | 0
mesh erosion into urinary bladder | 0
vesico-cutaneous fistula | 0
urethral catheter insertion | 0
septic shock | 0
inotropic support | 0
mechanical ventilation | 0
antibiotics | 0
repeated debridement | 24
removal of mesh | 168
repair of urinary bladder defect | 168
abdominoplasty | 336
condition stabilized | 336
cystogram | 336
no leakage from urinary bladder | 336
transferred to general ward | 336
transferred to rehabilitation bed | 336
wound healing | 504
satisfactory condition | 504