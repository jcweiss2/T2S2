73 years old | 0
female | 0
fever | -168
asthenia | -168
odynophagia | -168
daily episodes of a small volume of epistaxis through the left nasal cavity | -168
denied expelling any foreign body through the oral or nasal cavity | -168
treated in the Emergency Unit | -24
referred to the otorhinolaryngology service of a tertiary hospital | 0
cacosmia | -26208
foul-smelling nasal crusts | -26208
diabetes | 0
hypertension | 0
afebrile | 0
oriented | 0
cooperative | 0
crackles in the lung bases | 0
mucopurulent secretion in the left external auditory canal | 0
peritonsillar bulging | 0
hyperemia | 0
extended to the soft palate | 0
initial suspicion of peritonsillar abscess | 0
puncture of the oral bulge | 0
no secretion drained | 0
hospitalized | 0
intravenous antibiotic therapy with ceftriaxone | 0
intravenous antibiotic therapy with clindamycin | 0
second puncture | 24
no drainage | 24
evidence of larvae coming out through the mouth | 24
evidence of larvae coming out through the left nostril | 24
developed septicemia | 24
transferred to the intensive care unit | 24
decreased level of consciousness | 24
blood desaturation | 24
requiring intubation | 24
mechanical ventilation | 24
Iodoform applied to the oral cavity | 24
Iodoform applied to the nasal passages | 24
ivermectin administered through the nasogastric tube | 24
wide-spectrum antibiotics with piperacillin/tazobactam | 24
wide-spectrum antibiotics with vancomycin | 24
otorhinolaryngological examination performed daily | 24
removal of larvae | 24
approximately 150 larvae removed after 72 h | 96
computed tomography of the nose | 24
computed tomography of paranasal sinuses | 24
computed tomography of temporal bones | 24
computed tomography of skull | 24
computed tomography of lung | 24
complete removal of the larvae in the oral cavity | 96
complete removal of the larvae in the nasal cavity | 96
died due to respiratory failure secondary to pneumonia | 720
