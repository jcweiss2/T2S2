39 years old | 0
female | 0
virgo intacta | 0
admitted to the hospital | 0
history of heavy menstrual bleeding | -672
submucous leiomyoma | -672
hysteroscopy | -24
GnRH agonists | -24
difficult entry into the uterine cavity | -24
leiomyoma incompatible with resection | -24
discharged home | -24
mild pelvic pain | 24
vomiting | 24
no fever | 24
no bleeding | 24
ultrasound | 24
no free pelvic fluid | 24
no leukocytosis | 24
normal C-reactive protein | 24
paracetamol | 24
discharged | 24
intermittent fever | 96
abdominal pain | 96
distension | 96
multiple episodes of vomiting | 96
normotensive | 120
normal heartrate | 120
tympanic temperature | 120
facial flushing | 120
distal hypoperfusion | 120
cold extremities | 120
mottled skin | 120
IV fluid infusion | 120
large-spectrum antibiotics | 120
blood samples | 120
urine samples | 120
vaginal ultrasound | 120
normal-sized uterus | 120
leiomyoma | 120
no signs of perforation | 120
virtual uterine cavity | 120
retro-uterine position | 120
limited mobility | 120
endometriosis | 120
fluid-filled cystic mass | 120
dilated right fallopian tube | 120
transferred to intermediate care unit | 120
leukocytosis | 120
neutrophilia | 120
elevated C-reactive protein | 120
anuric status | 120
acute renal lesion | 120
blood creatinine | 120
primary metabolic alkalosis | 120
arterial blood gasometry | 120
abdominal X-ray | 120
distension of stomach | 120
distension of small bowel | 120
no pneumoperitoneum | 120
CT scan | 120
marked distension of gastric chamber | 120
proximal small bowel | 120
fluid collection in pelvis | 120
emergency exploratory laparotomy | 144
ruptured right fallopian tube | 144
hemoperitoneum | 144
generalized pelvic infection | 144
ampicillin-sensitive E. coli | 144
sub-total hysterectomy | 144
bilateral adnexectomy | 144
transferred to intensive care unit | 144
stage 4 multiple organ failure | 144
mechanical ventilation | 144
vasopressors | 144
hypoperfusion acute kidney injury | 144
fluid resuscitation | 144
aminergic support | 144
full recovery of kidney function | 240
discharged home | 288
oral antibiotics | 288
histological findings | 288
acute salpingitis | 288
peritonitis | 288
endometriotic cysts | 288
uterine leiomyomas | 288
no uterine perforation | 288
hormone replacement therapy | 288