Here is the table of events and timestamps:

48 years old | 0
male | 0
admitted to the Emergency Service | 0
toothache | -96
dyspnea | -96
chest pain | -96
sweating | -96
tachyarrhythmia | -96
sore throat | -96
fever | -96
treated at home with ceftriaxone-steroids-based | -96
gross swelling of the lower right cheek | -96
submandibular and mental regions were erythematous and warm on palpation | -96
difficulties in opening the jaw | -96
inflammatory changes in the mucous membrane of his oral cavity | -96
WBC count increased | -48
neutrophils increased | -48
C-reactive protein increased | -48
urgently orotracheal intubation | -48
left pleural effusion | -48
mediastinitis | -48
right parapharyngeal abscess | -48
odontogenic infection | -48
drainage of the right neck | -48
left chest drain | -48
intravenous antibiotic therapy | -48
clinical condition worsened | -46
transferred to an Intensive Care Unit | -46
chest and neck CT scan | -44
air collection in the right submandibular, in the left carotid, in the retroesophageal and pretracheal spaces | -44
collections characterized by air and fluids in the upper, anterior, and posterior mediastinum | -44
cervical necrotizing fasciitis with DNM derived | -44
bilateral pleural effusions | -44
additive pleural drain | -44
chest and neck CT angiography | -42
abscesses in the cervical spaces, an extensive mediastinal empyema, a left pleural effusion and right hydropneumothorax | -42
aggressive mediastinal debridement and VATS | -42
mediastinal empyema | -42
anterior and posterior mediastinum spaces | -42
1100 mL of yellow-brown secretion | -42
incision and drainage of the neck abscesses | -42
oral tooth extraction | -42
purulent fluid in the cavity below was drained and packed | -42
microscopy and culture of aspirated fluids and abscesses | -42
growth of Streptococcus anginosus, Gemella morbillorum, and Staphylococcus lagdunensis | -42
antibiotic therapy initiated | -42
Amoxicillin 1000 mg intravenously | -42
Metronidazole 500 mg intravenously | -42
dismissed in better health conditions | -7