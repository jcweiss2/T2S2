 \n\n

\boxed{
46 years old | 0  
male | 0  
Asian-Indian | 0  
no history of alcohol consumption | 0  
diagnosed with tropical chronic pancreatitis | -157680  
oral pancreatic enzyme therapy | -157680  
non-insulin-dependent diabetes mellitus | -157680 + 25920  
glucotrol (glipizide) 5 mg daily | -157680 + 25920  
steady midepigastric pain | -6  
dull pain | -6  
radiating pain through back | -6  
exacerbated by food intake | -6  
recurrent pain | -6  
lasted between 1 and 3 days | -6  
completely well in interval phase | -6  
hospitalized for pain control with narcotics | -6  
discharged | -6  
returning with continuing epigastric pain | -48  
increasing intensity of pain | -48  
nausea | -48  
vomiting | -48  
no documented fever | -48  
CT scan | -48  
fatty atrophy of both the pancreatic head and uncinate process | -48  
large calcifications in the pancreatic duct | -48  
possible obstruction at the level of the neck | -48  
marked upstream ductal dilatation of 1.5 cm | -48  
admitted for management of pain secondary to chronic pancreatitis | 0  
similar pain and fever | -1488  
CT scan in India | -1488  
chronic atrophic calcific pancreatitis | -1488  
dilated pancreatic duct (7 mm) | -1488  
intraductal calculi | -1488  
ERCP in India | -1488  
confirmed findings on pancreatography | -1488  
medically managed and discharged | -1488  
fever | 48  
chills and rigors | 48  
severe sepsis | 48  
septic shock | 48  
transferred to the medical intensive care unit | 48  
intubated for hypoxemic respiratory failure | 48  
acute respiratory distress syndrome | 48  
multiorgan failure | 48  
administration of broad-spectrum antibiotics | 48  
vasopressor support | 48  
activated recombinant human protein C | 48  
ultrasound of the abdomen | 48  
markedly dilated pancreatic duct (1.9 cm) | 48  
8.7 × 7.6 mm calculus within the duct | 48  
diffusely echogenic pancreas | 48  
prominent common bile duct | 48  
no obvious obstructing calculi | 48  
emergency ERCP | 48  
major papilla of Vater expelling frank pus | 48  
no evidence of papillitis, tumor, or previous sphincterotomy | 48  
evacuation of more than 5 ml of yellow pus | 48  
normal biliary tree without stones | 48  
marked dilatation of the main pancreatic duct | 48  
single distal calculus | 48  
evacuation of approximately 20 ml of pus | 48  
placement of 5-cm-long 5 F stent | 48  
no more pus draining | 48  
assumed ASPD | 48  
contrast enhanced CT scan | 72  
inflammatory changes within the fat surrounding the body and tail of the pancreas | 72  
edema | 72  
diminished dilatation of the pancreatic duct | 72  
distal migration of calculus towards the sphincter of Oddi | 72  
no evidence of pancreatic necrosis or fluid collection | 72  
bilateral moderate pleural effusions | 72  
clinical improvement | 96  
stabilization of hemodynamic parameters | 96  
blood cultures grew Klebsiella ornithinolytica | 96  
extubated | 96  
transferred from the intensive care unit | 96  
completed antibiotic course | 264  
discharged home | 264  
follow-up examination at 1 month | 744  
follow-up examination at 3 months | 2208  
no further complications | 2208  
} \n
Note: The timestamps for events that occurred in the past relative to the current admission (e.g., diagnosis of tropical chronic pancreatitis, development of diabetes mellitus) are approximated based on the provided timeline. The exact number of hours is calculated assuming 3 years and 2 months (1104 days) for the interval between the initial diagnosis and the current admission. \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
} \n
}