60 years old | 0
Malay lady | 0
admitted to the hospital | 0
right otalgia | 0
purulent otorrhea | 0
diagnosed with right malignant otitis externa | 0
started on intravenous Augmentin | 0
bony destruction of external auditory canal | -120
bony destruction of mastoid | -120
bony destruction of right mandibular fossa | -120
osteomyelitis of the right temporal bone | -120
Infectious disease consult | 120
started on intravenous linezolid | 120
started on intravenous piperacillin/tazobactam | 120
severe sepsis | 192
metabolic acidosis | 192
acute renal failure | 192
intubated | 192
managed in the surgical intensive care unit | 192
cultures performed on pus | 192
grew multi-resistant staphylococcus aureus | 192
grew pseudomonas aeruginosa | 192
urine culture grew Candida albicans | 192
antibiotic regime changed to intravenous meropenem | 192
antibiotic regime changed to intravenous vancomycin | 192
started on intravenous caspofungin | 192
anuric | 240
started on dialysis | 240
started on sustained low efficiency dialysis | 240
converted to continuous veno-venous hemodialysis | 288
abdominal distension | 288
abdominal X-ray performed | 288
mottled lucencies over the gastric lumen | 288
computed tomography scan of the abdomen and pelvis | 288
extensive gastric intramural gas | 288
exploratory laparotomy | 336
intra-operative findings revealed an infarcted stomach | 336
total gastrectomy | 336
vasculature of the coeliac axis had good palpable pulsations | 336
vasculature of the superior mesenteric artery had good palpable pulsations | 336
persistent hypotension | 408
bradycardia | 408
maximal inotropic support | 408
passed away | 432
total gastric infarction | 432
widely disseminated fungal organisms | 432
infarction of the entire gastric wall | 432
fungal organisms disseminated through the entire gastric wall | 432
fungal organisms within the vascular channels | 432
spores and hyphae of variable irregular sizes | 432
branching at right angles | 432
poorly controlled type 2 diabetes mellitus | -10000
bone marrow transplant for acute myeloid leukemia | -10000 
right malignant otitis externa | 0 
refractory to antibiotic treatment | 120 
follow up computed tomography scan | 120 
bony destruction | 120 
osteomyelitis | 120 
sepsis | 192 
metabolic acidosis | 192 
acute renal failure | 192 
intubated and managed in the surgical intensive care unit | 192 
multi-resistant staphylococcus aureus | 192 
pseudomonas aeruginosa | 192 
Candida albicans | 192 
intravenous meropenem | 192 
intravenous vancomycin | 192 
intravenous caspofungin | 192 
anuric | 240 
dialysis | 240 
sustained low efficiency dialysis | 240 
continuous veno-venous hemodialysis | 288 
abdominal distension | 288 
abdominal X-ray | 288 
mottled lucencies over the gastric lumen | 288 
computed tomography scan of the abdomen and pelvis | 288 
extensive gastric intramural gas | 288 
exploratory laparotomy | 336 
intra-operative findings revealed an infarcted stomach | 336 
total gastrectomy | 336 
persistent hypotension | 408 
bradycardia | 408 
maximal inotropic support | 408 
passed away | 432 
total gastric infarction | 432 
widely disseminated fungal organisms | 432 
infarction of the entire gastric wall | 432 
fungal organisms disseminated through the entire gastric wall | 432 
fungal organisms within the vascular channels | 432 
spores and hyphae of variable irregular sizes | 432 
branching at right angles | 432 
mucormycosis | 432 
invasive mycormycosis | -10000 
immunocompromised states | -10000 
diabetes | -10000 
Acquired Immunodeficiency Syndrome (AIDS) | -10000 
malnutrition | -10000 
defects in host phagocytes | -10000 
corticosteroid use | -10000 
organ or stem cell transplantation | -10000 
gastrointestinal mucormycosis | 432 
infection of the alimentary tract | 432 
ingestion of the spores | 432 
stomach | 432 
colon | 432 
ileum | 432 
duodenum | 432 
jejunum | 432 
arterial invasion | 432 
arterial thrombosis | 432 
tissue infarction | 432 
necrosis | 432 
venous invasion | 432 
hemorrhage | 432 
aseptate, wide, ribbon-like hyphae | 432 
branching at right angles | 432 
anti-fungal treatment | 432 
surgery | 432 
debulking the fungal infection | 432 
resection of all the infected necrotic tissue | 432 
liposomal or lipid complex amphotericin B | 432 
surgical debridement | 432 
reversal of the predisposing condition | 432 
controlling hyperglycaemia | 432 
limiting the use of glucocorticosteroids | 432 
reducing the dosage in immunosuppressed patients | 432 
ischemic gut | 432 
immunocompromised patients | 432 
extended surgical intensive care unit stay | 432 
mucormycosis/fungal infections of the gut | 432 
early consult by the infectious disease specialty | 432 
appropriate anti-fungal treatment | 432 
timely implementation of subsequent surgical management | 432 
better recognition of mucormycosis | 432 
prompt management | 432 
better outcomes | 432