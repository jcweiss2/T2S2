57 years old | 0
female | 0
non-smoker | 0
non-drinker | 0
good past health | 0
sore throat | -168
runny nose | -168
productive cough | -168
high fever | 0
sinus tachycardia | 0
skin erythema | 0
crepitus | 0
oxygen saturation maintained | 0
retropharyngeal gas | 0
consolidative changes at the right lower zone | 0
metabolic acidosis | 0
multiple gas locules in bilateral deep cervical spaces | 0
loculated right pleural effusion | 0
right chest wall subcutaneous emphysema | 0
deep neck space infection | 0
descending mediastinitis | 0
empyema thoracis | 0
emergency surgical debridement | 0
drainage | 0
necrotic fascia and muscle debrided | 0
turbid fluid drained | 0
neck wound laid open | 0
gauze packed | 0
multiple right lower posterior teeth extracted | 0
severe periodontitis | 0
chest drains inserted | 0
high dose inotropes | 0
intubated | 0
daily wound examination | 0
daily dressing | 0
second look wound exploration | 72
debridement | 72
residual collection drained | 72
tracheostomised | 72
feeding tube inserted | 72
inotropic support | 0
ventilatory support | 0
primary closure of neck wound | 432
tracheostomy decanalised | 432
swallowing rehabilitation | 432
discharged | 1440
necrotizing inflammation | 0
C. parapsilosis | 0
Peptostreptococcus micros | 0
Bacteroides pyogenes | 0
Prevotella buccae | 0
intravenous anidulafungin | 0
broad-spectrum antibiotics | 0