2 years old | 0
    male | 0
    admitted to the local hospital | 0
    collapse | 0
    unresponsive | 0
    crying | 0
    persistently altered level of consciousness | 0
    normal vital signs | 0
    dual heart sounds | 0
    clear chest | 0
    soft abdomen | 0
    nontender abdomen | 0
    generalized poor tone | 0
    no neurological deficits | 0
    no significant medical history | 0
    no antenatal history | 0
    no regular medications | 0
    intravenous ceftriaxone | 0
    aciclovir | 0
    mild neutrophilia | 0
    hypokalaemia | 0
    metabolic acidosis | 0
    improved level of consciousness | 24
    transferred to tertiary center | 24
    sepsis | 24
    meningitis | 24
    atypical seizures | 24
    marked dysmetria | 48
    dysphagia | 48
    deranged coagulation profile | 48
    international normalized ratio 1.7 | 48
    activated partial thromboplastin time 62 | 48
    fibrinogen level 0.9 | 48
    blood cultures | 48
    infectious serology | 48
    autoimmune screen | 48
    vasculitic screen | 48
    lumbar puncture | 48
    possible bite mark on lip | 48
    snake venom-specific enzyme immunoassay | 48
    acute respiratory distress | 72
    transferred to pediatric intensive care unit | 72
    encephalopathy | 72
    intubation | 72
    ventilation | 72
    cryoprecipitate | 72
    methylprednisolone | 72
    normal echocardiogram | 72
    MRI with contrast | 96
    multiple acute ischemic infarctions | 96
    no hemorrhage | 96
    antibiotics ceased | 120
    antivirals ceased | 120
    corticosteroids ceased | 120
    extubated | 120
    positive Eastern Brown snake venom | 120
    resolved dysmetria | 144
    resolved dysphagia | 144
    discharged | 192
    ongoing rehabilitation | 192
    physical therapy | 192
    occupational therapy | 192
    good recovery | 192
    meeting developmental milestones | 192
    