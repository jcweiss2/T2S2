60 years old | 0
male | 0
admitted to the emergency department | 0
acute anaemia | 0
fever | 0
poorly controlled diabetes mellitus | -720
laparoscopic radical cystectomy | -720
bilateral pelvic lymph node dissection | -720
urinary diversion | -720
discharged | -720
septic shock | 0
haemorrhagic shock | 0
diffuse extravasation of the contrast medium | 0
right external iliac artery disruption | 0
broad-spectrum antibiotics | 0
imipenem | 0
open exploratory operation | 0
extensive adhesion formation | 0
inflammation | 0
vessel split of the right external iliac artery | 0
vascular stent insertion | 0
transferred to the intensive care unit | 0
Klebsiella pneumoniae subsp. Pneumoniae isolated | 72
blood culture | 72
standard drug susceptibility test | 72
tigecycline | 72
imipenem | 72
vital signs became normal | 504
blood tests became normal | 504
repeat enhanced CT | 744
no effusion of the contrast medium | 744
discharged | 816
follow-up | 8760
no relapse | 10512