47 years old | 0
    man | 0
    admitted to the hospital | 0
    persistent severe headache | -1080
    chronic smoker | 0
    nonalcoholic | 0
    subarachnoid hemorrhage | -1080
    hydrocephalus | 0
    external ventricular drain | 0
    aneurysm clipping | 0
    ventriculoperitoneal shunt | 0
    elective ventilation | 0
    extubation | 24
    fever | 72
    hypotension | 72
    deterioration in sensorium | 72
    sepsis suspected | 72
    fluid resuscitation | 72
    antibiotics | 72
    noradrenaline infusion | 72
    vasospasm suspected | 72
    repeat digital subtraction angiography | 72
    complete aneurysm clipping confirmed | 72
    no vasospasm | 72
    sepsis source not identified | 72
    abdominal distension | 120
    persisting fever | 120
    ascites | 120
    bilateral pleural effusion | 120
    severe hypoalbuminemia | 120
    intravenous albumin administered | 120
    respiratory effort interference | 120
    failed ventilator weaning | 120
    elevated lipase | 120
    CT abdomen ordered | 120
    edematous pancreas | 120
    peripancreatic fat stranding | 120
    acute pancreatitis | 120
    antibiotics continued | 120
    antipyretics | 120
    total parental nutrition | 120
    sensorium fluctuations | 168
    VP shunt externalization | 168
    neurologic status improved | 168
    ascitic fluid testing | 168
    no infection | 168
    abdominal distension subsiding | 336
    tracheostomy | 336
    ventilator weaning | 336
    GCS improvement | 336
    enteral feedings initiated | 336
    lipase normalization | 336
    shifted to ward | 336
    fever recurrence | 504
    altered sensorium | 504
    shunt tube infection signs | 504
    Klebsiella identified | 504
    antibiotics adjusted | 504
    septic shock | 504
    death | 672
    
    
    47 years old | 0
    man | 0
    admitted to the hospital | 0
    persistent severe headache | -1080
    chronic smoker | 0
    nonalcoholic | 0
    subarachnoid hemorrhage | -1080
    hydrocephalus | 0
    external ventricular drain | 0
    aneurysm clipping |0
    ventriculoperitoneal shunt |0
    elective ventilation |0
    extubation |24
    fever |72
    hypotension |72
    deterioration in sensorium |72
    sepsis suspected |72
    fluid resuscitation |72
    antibiotics |72
    noradrenaline infusion |72
    vasospasm suspected |72
    repeat digital subtraction angiography |72
    complete aneurysm clipping confirmed |72
    no vasospasm |72
    sepsis source not identified |72
    abdominal distension |120
    persisting fever |120
    ascites |120
    bilateral pleural effusion |120
    severe hypoalbuminemia |120
    intravenous albumin administered |120
    respiratory effort interference |120
    failed ventilator weaning |120
    elevated lipase |120
    CT abdomen ordered |120
    edematous pancreas |120
    peripancreatic fat stranding |120
    acute pancreatitis |120
    antibiotics continued |120
    antipyretics |120
    total parental nutrition |120
    sensorium fluctuations |168
    VP shunt externalization |168
    neurologic status improved |168
    ascitic fluid testing |168
    no infection |168
    abdominal distension subsiding |336
    tracheostomy |336
    ventilator weaning |336
    GCS improvement |336
    enteral feedings initiated |336
    lipase normalization |336
    shifted to ward |336
    fever recurrence |504
    altered sensorium |504
    shunt tube infection signs |504
    Klebsiella identified |504
    antibiotics adjusted |504
    septic shock |504
    death |672
    

    
    <|eot_id|>
    
  