44 years old | 0
    male | 0
    heart transplant | - (assumed prior to admission, exact time unclear; assigned 0)
    tacrolimus | - (prior to admission, exact time unclear; assigned 0)
    End-Stage Renal Disease (ESRD) | - (prior to admission, exact time unclear; assigned 0)
    hemodialysis | - (prior to admission, exact time unclear; assigned 0)
    recently treated CMV viremia | - (prior to admission, exact time unclear; assigned 0)
    necrotizing pancreatitis | - (prior to admission, exact time unclear; assigned 0)
    chills | -96
    decreased appetite | -96
    worsening non-bloody emesis | -96
    dull left upper quadrant abdominal pain | -96
    radiation to the back | -96
    no shortness of breath | -96
    no fever | -96
    no diarrhea | -96
    no blood in the stool | -96
    blood pressure 90/61 mmHg | 0
    heart rate 110 beats per minute | 0
    temperature 98.1 °F | 0
    respiratory rate 18 per minute | 0
    scleral icterus | 0
    decreased bibasilar breath sounds | 0
    moderate abdominal tenderness | 0
    left flank | 0
    left upper abdominal quadrant | 0
    no palpable mass | 0
    1+ bilateral pedal edema | 0
    sinus tachycardia | 0
    no ischemic changes | 0
    mild pulmonary edema | 0
    WBC 8.3 k/uL | 0
    hemoglobin 10.2 g/dL | 0
    platelet count 90 k/uL | 0
    BUN/creatinine 45/5.8 | 0
    elevated high sensitivity troponin 2479 pg/mL | 0
    BNP 600 | 0
    AST 2645 U/L | 0
    ALT 2935 U/L | 0
    ALP 106 U/L | 0
    lipase 61 U/L | 0
    total bilirubin 3.5 mg/dL | 0
    conjugated bilirubin 2.1 mg/dL | 0
    reduced left ventricular size | 0
    hyperdynamic systolic function |)