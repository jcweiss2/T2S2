60 years old | 0
male | 0
hypertension | 0
admitted to the hospital | 0
left eye swelling | -168
pain | -168
erythema | -168
circulatory shock | 0
sepsis | 0
broad-spectrum intravenous antibiotics | 0
Vancomycin | 0
Gentamycin | 0
Meropenem | 0
Clindamycin | 0
aggressive fluid resuscitation | 0
oxygen supplementation | 0
diffuse left orbital cellulitis | 0
no intraorbital collection | 0
no intracerebral vascular thrombosis | 0
inflammatory picture | 0
CRP 560 | 0
WBC 19.80 | 0
Neutrophils 18.60 | 0
Lymphocytes 0.70 | 0
Hb 154 | 0
Creatinine 792 | 0
K+ 3.7 | 0
Blood glucose 7.1 | 0
respiratory compromise | 2
haemodynamic instability | 2
intubation | 2
ventilatory support | 2
vasopressor treatment | 2
IVIg | 4
emergency transfer | 4
surgical intervention | 4
left periorbital swelling | 4
necrosis of the upper eyelid | 4
abscess of the lower eyelid | 4
debridement | 4
septic shock | 4
multiorgan failure | 4
Meropenem | 4
Clindamycin | 4
Ceftriaxone | 4
Linezolid | 4
Beta-haemolytic Group A Streptococcus | 4
Staphylococcus Aureus | 4
penicillin | 4
erythromycin | 4
trimethoprim | 4
gentamycin | 4
flucloxacillin | 4
condition stabilization | 28
repeat CT orbit | 28
persistent soft tissue swelling | 28
no orbital breach | 28
no collections | 28
discharge from hospital | 456
wound healing | 2196
no visual deficit | 2196
reconstructive surgery | 2196