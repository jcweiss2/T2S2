34 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
primary refractory acute myeloblastic leukemia | -8760 | -8760 | Factual
multiple relapses | -8760 | 0 | Factual
allogeneic bone marrow transplant | -648 | -648 | Factual
delayed engraftment | -648 | 0 | Factual
prolonged severe neutropenia | -648 | 0 | Factual
vancomycin-resistant Enterococcus | -648 | 0 | Factual
Streptococcus viridans | -648 | 0 | Factual
Streptococcus mitis | -648 | 0 | Factual
bacteremia | -648 | 0 | Factual
tedizolid | -648 | 0 | Factual
cefepime | -648 | 0 | Factual
Flagyl | -648 | 0 | Factual
daptomycin | -648 | 0 | Factual
acute abdominal pain | 0 | 0 | Factual
filgrastim | 0 | 0 | Factual
acyclovir | 0 | 0 | Factual
Bactrim | 0 | 0 | Factual
caspofungin | 0 | 0 | Factual
fever | 0 | 0 | Factual
tachycardia | 0 | 0 | Factual
hypotension | 0 | 0 | Factual
tachypnea | 0 | 0 | Factual
ill appearing | 0 | 0 | Factual
distended abdomen | 0 | 0 | Factual
localized peritonitis | 0 | 0 | Factual
white cell count 0.2 x 10^9 /L | 0 | 0 | Factual
absolute neutrophil count (ANC) of zero | 0 | 0 | Factual
anemic | 0 | 0 | Factual
hemoglobin of 7 g/L | 0 | 0 | Factual
thrombocytopenic | 0 | 0 | Factual
platelet count of 10 x 10^9 /L | 0 | 0 | Factual
lactic acid of 3.1 mmol/L | 0 | 0 | Factual
CT scan | 0 | 0 | Factual
segmental ischemia of the small bowel | 0 | 0 | Factual
exploratory laparotomy | 0 | 24 | Factual
ischemic bowel segment | 0 | 24 | Factual
small bowel resection | 0 | 24 | Factual
primary anastomosis | 0 | 24 | Factual
norepinephrine | 0 | 24 | Factual
vasopressin | 0 | 24 | Factual
transesophageal echo | 0 | 24 | Factual
intensive care unit | 24 | 48 | Factual
pressors weaned | 24 | 48 | Factual
extubated | 24 | 48 | Factual
transferred to the floor | 48 | 48 | Factual
diet advanced | 72 | 72 | Factual
passed flatus | 72 | 72 | Factual
new fevers | 96 | 96 | Factual
increased abdominal pain | 96 | 96 | Factual
lactic acidosis | 96 | 96 | Factual
respiratory decompensation | 96 | 96 | Factual
neutropenic | 96 | 96 | Factual
white cell count of 0.1x 10^9 /L | 96 | 96 | Factual
ANC 0 | 96 | 96 | Factual
lactic acid 3.7 mmol/L | 96 | 96 | Factual
amphotericin B | 96 | 96 | Factual
repeat CT scan | 96 | 96 | Factual
necrotic small bowel | 96 | 96 | Factual
expedited pathology report | 96 | 96 | Factual
invasive fungal forms | 96 | 96 | Factual
mucormycosis | 96 | 96 | Factual
hematologic dissemination | 96 | 96 | Factual
septic emboli | 96 | 96 | Factual
comfort measures | 120 | 120 | Factual
died | 120 | 120 | Factual