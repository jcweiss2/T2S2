21 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
obese | 0 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
cough | -72 | 0 | Factual
fever | -72 | 0 | Factual
shortness of breath | -72 | 0 | Factual
pleuritic chest pain | -72 | 0 | Factual
light-headedness | -24 | 0 | Factual
near syncope | -24 | 0 | Factual
dyspnoea | -24 | 0 | Factual
COVID-19 | 0 | 0 | Factual
sub-massive pulmonary embolism | 0 | 0 | Factual
unfractionated heparin | 0 | 12 | Factual
hypotensive | 12 | 12 | Factual
massive pulmonary embolism | 12 | 12 | Factual
catheter-directed thrombolysis | 12 | 18 | Factual
improved clinically | 18 | 24 | Factual
plans made for discharge | 24 | 24 | Factual
acute respiratory failure | 72 | 72 | Factual
hypotension | 72 | 72 | Factual
intubated | 72 | 72 | Factual
cardiac arrest | 72 | 72 | Factual
return of spontaneous circulation | 72 | 72 | Factual
vasopressors | 72 | 120 | Factual
veno-arterial extracorporeal membrane oxygenation | 72 | 240 | Factual
recurrent massive pulmonary embolism | 72 | 72 | Factual
repeat catheter-directed thrombolysis | 72 | 78 | Factual
ventilation parameters improved | 120 | 120 | Factual
vasopressors discontinued | 120 | 120 | Factual
weaning of ECMO began | 120 | 240 | Factual
deep venous thrombus | 120 | 120 | Factual
inferior vena cava filter | 120 | 120 | Factual
low-molecular-weight heparin | 120 | 0 | Factual
septic shock | 240 | 240 | Factual
right thigh haematoma | 336 | 336 | Factual
compartment syndrome | 336 | 336 | Factual
surgical debridement | 336 | 336 | Factual
rivaroxaban | 336 | 0 | Factual
discharged | 1248 | 1248 | Factual
home | 1608 | 1608 | Factual
anticoagulated | 1608 | 0 | Factual
no major adverse events | 1936 | 1936 | Factual