42 years old | 0
female | 0
admitted to the hospital | 0
stag horn calculus | 0
hyperparathyroidism | 0
morbid obesity | 0
BMI of 75 | 0
limited exercise tolerance | 0
obstructive sleep apnea | 0
BiPAP | 0
hypertension | 0
diabetes | 0
acid reflux disease | 0
hepatitis C | 0
smoker | 0
postoperative nausea and vomiting | 0
no known drug allergies | 0
insulin | 0
lisinopril | 0
hydrochlorothiazide | 0
atorvastatin | 0
aspirin | 0
venlafaxine | 0
trazodone | 0
rosuvastatin | 0
heart rate 77/min | 0
BP 93/53 mmHg | 0
respiration 16/min | 0
SpO2 93% on room air | 0
decreased thyromental distance | 0
interincisor distance 4 cm | 0
elevated parathyroid hormone | 0
elevated calcium | 0
premedicated with 30 ml of 0.3 molar sodium citrate | 0
IV ranitidine 50 mg | 0
20 G intravenous cannula placed on right foot | 0
arterial line in right radial artery | 0
invasive blood pressure monitoring | 0
arterial line for frequent blood sampling | 0
transferred to operating room | 0
placed on RAMP | 0
standard ASA monitoring | 0
preoxygenated for 3 minutes | 0
rapid sequence induction | 0
propofol 300 mg | 0
suxamethonium 160 mg | 0
trachea intubated with size 7.5 endotracheal tube | 0
MAC 4 blade with grade I view | 0
anesthesia maintained with oxygen/air | 0
sevoflurane | 0
intermittent doses of rocuronium | 0
neck explored | 0
multiple frozen sections sent for identification | 0
fat tissue identified | 0
surgery duration four-and-a-half hours | 0
resection of left inferior parathyroid adenoma | 0
parathyroid hormone levels normalized in 15 minutes | 0
extensive neck dissection | 0
resultant edema | 0
planned to keep intubated in ICU | 0
extubate on following day | 0
transferred to ICU intubated and ventilated | 0
propofol infusion started at 20 μg/kg/min | 0
not tolerating endotracheal tube | 0
propofol escalated to 80 μg/kg/min | 0
propofol dose 4 mg/kg/h | 0
failed spontaneous breathing test | 0
oxygen requirements increasing | 0
respiratory failure secondary to basal atelectasis | 0
ventilator-associated pneumonia | 0
postoperative day 3 | 72
creatinine kinase 66900 IU/l | 72
myoglobin 19470 ng/ml | 72
rhabdomyolysis diagnosed | 72
urine output declining | 72
creatinine 3.1 mg/dl | 72
BUN 41 mg/dl | 72
acute renal failure | 72
septic shock secondary to urinary tract infection | 72
ventilator-associated pneumonia | 72
inotropic support with norepinephrine | 72
metabolic acidosis | 72
base deficit more than 10 mmol/l | 72
PRIS suspected | 72
propofol infusion stopped | 72
lorazepam and fentanyl for sedation | 72
dialyzed for acute renal failure | 72
postoperative day 10 | 240
rhabdomyolysis resolved | 240
renal failure resolved | 240
multiple extubation attempts failed | 240
tracheostomy on postoperative day 16 | 384
large decubitus ulcer | 384
frequent debridement | 384
awaiting palliative care | 384
died on postoperative day 65 | 1560
fall from bed | 1560
tracheostomy occlusion in prone position | 1560
propofol infusion syndrome | 72
acute event recovery | 240
death from other causes | 1560
hyperparathyroidism |+0
