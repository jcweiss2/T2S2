69 years old | 0
    female | 0
    referred to tertiary referral center | 0
    recurrent UTIs | 0
    problems during monthly iBC change | 0
    surgery for spondylolisthesis | -1440
    stress urinary incontinence | -1056
    treated with increasing number of pads | -1056
    addressed to iBC | -1056
    iBC changed monthly | -1056
    abdominal ultrasound | 0
    computed tomography | 0
    bladder stone | 0
    videourodynamic study | 0
    defunctionalized bladder | 0
    addressed to uterus-sparing simple cystectomy | 0
    uretero?ileal?cutaneous diversion according to Bricker | 0
    operative time 215 minutes | 0
    antibiotic prophylaxis with Cefazolin | 0
    active chronic cystitis with follicular and eosinophilic features | 0
    mucosa ulcers | 0
    septic on third POD | 72
    severe lumbar pain | 72
    Escherichia coli colonization | 72
    Pseudomonas aeruginosa colonization | 72
    Candida glabrata colonization | 72
    pancreatic edema | 72
    conservative approach attempted | 72
    septic shock on 18th POD | 432
    Enterococcus faecium positive | 432
    Pseudomonas aeruginosa positive | 432
    Acinetobacter spp positive | 432
    urgent exploratory laparotomy | 432
    acute necrotizing hemorrhagic pancreatitis | 432
    medical therapy continued | 432
    abdominopelvic washing surgeries | 432
    other septic episodes | 432
    stay in intensive care for 95 days | 432
    discharged after 141 days | 3384
    IV grade Clavien-Dindo complications | 3384
    well-functioning urinary diversion at follow-up | 3384
    no significant urinary tract conditions at follow-up | 3384
  