54 years old | 0
man | 0
presented with acutely discharging sinus | 0
abscess to right proximal tibia | 0
complex orthopaedic history | 0
infected non-union | 0
elective right tibial osteotomy | 0
past medical history included well-controlled asthma | 0
obstructive sleep apnoea | 0
hypertension | 0
deep vein thrombosis | 0
pericarditis | 0
generally unwell | 0
swinging fever | 0
Staphylococcus aureus bacteraemia | 0
started on flucloxacillin intravenously | 0
echocardiogram requested | 0
right knee radiographs showed non-union of the proximal tibia | 0
evidence of sequestrum | 0
CT scan confirmed | 0
right tibial exploration | 0
debridement conducted | 0
tissue sampling | 0
instillation of CERAMENT G | 0
application of spanning external fixator | 0
six tissue samples grew methicillin-sensitive S. aureus | 0
Proteus mirabilis | 0
Enterobacter | 0
oral rifampicin added | 0
transthoracic echo showed echogenic mobile structure behind mitral valve leaflet | 0
queried as endocarditis vegetation | 0
flucloxacillin increased to six times per day | 0
postoperative complications included significant pain | 0
acute kidney injury stage III | 0
hypovolaemia | 0
improved following intravenous fluid administration | 0
episodes of fever resolved | 0
postoperative day 5 | 120
difficult night with pain | 120
commenced 75 mg pregabalin two times per day | 120
commenced 100 mg tapentadol modified release every 12 hours | 120
pregabalin increased to 150 mg two times per day | 120
already taking 25 mg amitriptyline one time per day | 0
already taking 150 mg sertraline one time per day | 0
already taking 20 mg ketamine up to four times per day as required | 0
patient deteriorated | 144
impression of sepsis secondary to tibial infection | 144
impression of infective endocarditis | 144
possibility of serotonin syndrome raised | 144
commenced on tapentadol one dose | 144
commenced on pregabalin | 144
already taking sertraline and amitriptyline | 144
hyperthermia (41°C at highest) | 144
tachycardia | 144
tachypnoea | 144
tremor | 144
hyperreflexia | 144
agitation | 144
bilateral inducible ankle clonus | 144
diagnosis of serotonin syndrome | 144
serotoninergic medications suspended | 144
critical care involvement requested | 144
admitted to critical care unit | 144
blood cultures taken at initial temperature rise | 144
grew Proteus mirabilis | 144
meropenem added | 144
flucloxacillin increased to every four hours | 144
creatine kinase rose to 6490 U/L | 144
tenderness to mid anterior thigh | 144
urgent MRI ruled out myositis | 144
vital signs settled after cessation of medications | 144
last significant temperature rise of 39.5°C | 216
day 7 | 168
CK dropped to 205 U/L | 168
stepped down to the ward | 168
avoided requiring level 2 or 3 interventions | 168
transoesophageal echo conducted | 168
no criteria for infective endocarditis | 168
previously reported abnormality not significant | 168
discharged from intensive care unit | 168
CRP 276 mg/L | 144
CRP rose to 354 mg/L | 144
WCC 7.8×10^9/L | 144
neutrophils 6.7×10^9/L | 144
lymphocytes 0.6×10^9/L | 144
creatinine 138 µmol/L | 144
alkaline phosphatase 138 U/L | 144
discharged on 6-week course of antibiotics | 432
further orthopaedic procedure on right knee | 432
currently has circular fixator in place | 432
pin site infections | 432
ongoing issues with pain | 432
episode of deep vein thrombosis in right leg | 432
walking fully weight bearing | 432
help of crutches | 432
listed for removal of external fixator | 432
application of cast | 432
blood culture grew P. mirabilis | 144
positive blood culture for P. mirabilis | 144
raised CRP | 144
no raise in WCC | 144
no raise in neutrophils | 144
initial fever developed following initiation of pregabalin | 144
significant deterioration overnight following single dose of tapentadol | 144
administration of tapentadol at 00:30 a.m. | 144
clinical deterioration started around 04:44 a.m. | 144
hallucinations | 144
feeling irritable | 144
restless | 144
extreme hot sweats | 144
high temperatures | 144
verbal abuse | 144
anxiety | 144
irritation | 144
serotonin syndrome diagnosis | 144
