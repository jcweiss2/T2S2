43 years old | 0
    male | 0
    admitted to the hospital | 0
    left facial swelling | -336
    left hemifacial swelling | -336
    left hemifacial pain | -336
    fever | -240
    diabetes mellitus | -672
    insulin treatment | -672
    left cheek trismus | 0
    left cheek skin thinning | 0
    left cheek crepitation | 0
    elevated HbA1C (17.1) | 0
    high WBC count (15170/μL) | 0
    low hemoglobin (10.5 g/dL) | 0
    elevated hs-CRP (212.94 mg/L) | 0
    high glucose level (242 mg/dL) | 0
    low sodium (134 mmol/L) | 0
    low albumin (2.3 g/dL) | 0
    facial CT showing multiple abscesses with air bubbles | 0
    facial CT showing pleomorphic wall-enhancing lesions | 0
    LRINEC score 10 | 0
    surgical decompression | 0
    tachycardia | 24
    hypotension | 24
    septic shock | 24
    elevated procalcitonin (1.140 ng/mL) | 72
    K. pneumoniae in blood cultures | 72
    chest X-ray showing multiple nodules | 0
    chest CT showing septic emboli | 48
    chest CT showing pneumonia | 48
    abdominopelvic CT showing renal abscesses | 72
    intravenous meropenem | 24
    intravenous levofloxacin | 24
    antibiotic change to cefotaxime | 72
    seizures due to metabolic encephalopathy | 72
    addition of metronidazole | 144
    renal PCD insertion | 168
    improvement in hs-CRP | 168
    improvement in WBC | 168
    albumin recovery (≥3 g/dL) | 168
    facial CT showing decreased abscesses | 600
    APCT showing resolved renal abscesses | 1080
    HbA1C decrease to 4.9 | 1080
    resolved trismus | 4320
    discharge | 672