92 years old | 0
male | 0
admitted to the hospital | 0
general deterioration | 0
diabetes mellitus | 0
systemic hypertension | 0
stroke | 0
temperature of 34°C | 0
blood pressure of 70/30 mmHg | 0
pulse rate of 115 per minute | 0
respiratory rate of 22 per minute | 0
Glasgow Coma Scale of 8 out of 15 | 0
urinary tract infection | 0
septic shock | 0
transferred to the intensive care unit | 0
intravenous fluids | 0
vasopressors | 0
mechanical ventilation | 0
imipenem-cilastatin | 0
ciprofloxacin | 0
extended-spectrum beta-lactamase (ESBL)-producing Escherichia coli | 0
resistant to ciprofloxacin | 0
susceptible to imipenem | 0
susceptible to gentamicin | 0
ciprofloxacin replaced with gentamicin | 24
clinical conditions improved | 168
gentamicin discontinued | 240
imipenem-cilastatin discontinued | 336
fever up to 38.6°C | 576
hypotension | 576
peripheral blood leukocytosis | 576
white blood cell count 18×109/L | 576
80% neutrophils | 576
dull percussion sound | 576
reduced breath sounds in the left lung | 576
chest x-ray showed left lung consolidation | 576
chest x-ray showed large pleural effusion | 576
pigtail catheter inserted | 576
drain pleural effusion | 576
fluid analysis revealed protein at 52.0 g/L | 576
fluid analysis revealed lactate dehydrogenase at 1477 IU/L | 576
fluid analysis revealed pH at 7.0 | 576
fluid analysis revealed white blood cells at 8450 | 576
96% neutrophils | 576
ventilator-associated pneumonia | 576
pleurisy | 576
colistin methanesulfonate started | 576
imipenem-cilastatin 500 mg four times daily | 576
pneumothorax | 672
pigtail catheter replaced with intercostal chest drain | 672
pleural fluid showed ESBL-producing E. coli | 672
pleural fluid showed carbapenem-resistant Acinetobacter baumannii | 672
febrile | 672
continued to require high dose vasopressor infusions | 672
lack of clinical improvement | 672
intra-pleural colistin methanesulfonate added | 672
drain clamped for 2 hours | 672
drain resumed | 672
improvement in patient’s condition | 792
peripheral white blood cell count dropped to 8.8×109/L | 792
reduced need for ventilation | 792
discontinuation of vasopressor support | 792
pleural fluid sample taken | 816
Proteus mirabilis | 816
successful microbiological clearance | 816
imipenem switched to meropenem | 816
intra-pleural colistin methanesulfonate discontinued | 816
intravenous colistin methanesulfonate discontinued | 816
meropenem continued | 816
pleural fluid culture negative for A. baumannii and E. coli | 888
intercostal drain removed | 1008
resolution of infection signs | 1008
resolution of effusion | 1008
clinically stable | 1008
no further episodes of sepsis | 1008
attempts to wean off mechanical ventilation unsuccessful | 1008
acute myocardial ischemia | 1608
passed away | 1608
