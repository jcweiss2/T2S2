69 years old | 0
male | 0
admitted to the hospital | 0
severe sepsis | 0
Pulseless electrical activity (PEA) cardiac arrest | 0
cardiopulmonary resuscitation (CPR) | 0
return of spontaneous circulation | 0
hypotensive | 0
tachycardic | 0
fluid boluses | 0
metaraminol boluses | 0
tracheal intubation | 0
mechanical ventilation | 0
arterial blood gas analysis | 0
severe metabolic acidosis | 0
treatment initiated | 0
central venous catheter (CVC) inserted | 0
norepinephrine infusion | 0
sustained oliguria | 0
systemic acidosis | 0
CVVH initiated | 0
double lumen hemofiltration catheter inserted | 0
chest radiograph | 0
CVC and hemofiltration catheter tips adjacent | 0
precipitous hypotension | 0
PEA arrest | 0
spontaneous circulation restored | 0
CVVH recommenced | 24
fluid boluses | 24
epinephrine boluses | 24
norepinephrine infusion rate increased | 24
massive fluctuations in blood pressure | 24
CVVH stopped | 39
norepinephrine requirement reduced | 39
hemodynamic stability restored | 39
hemofiltration catheter withdrawn | 39
repeat chest radiograph | 39
CVVH resumed | 45
little hemodynamic instability | 45
no significant increase in vasopressor infusion rate | 45