67 years old | 0
male |9
neck pain | -2160
ground-level fall | -2160
no signs or symptoms of radiculopathy | 0
no signs or symptoms of myelopathy | 0
physical examination | 0
5/5 strength on manual motor testing | 0
decreased sensation to light touch involving right ear, face, and neck | 0
normal upper and lower extremity reflexes | 0
negative Hoffman’s sign | 0
negative Babinski reflex | 0
negative Romberg sign | 0
normal tandem gait | 0
radiographs of cervical spine | 0
persistent neck pain refractory to over-the-counter pain medications | 0
advanced imaging | 0
CT scan of cervical spine | 0
destructive lesion with peripheral sclerosis | 0
MRI scan of cervical spine | 0
T2 hyperintense enhancing mass | 0
extradural extension displacing spinal cord | 0
no evidence of myelomalacia | 0
mass extension into odontoid, anterior arch, right lateral mass of C1, right C2–3 neural foramen, right transverse process of C3, complete encasement of right vertebral artery | 0
CT-guided needle biopsy | 0
pathology consistent with chordoma | 0
CT scan of chest, abdomen, pelvis | 0
no evidence of metastatic disease | 0
temporary balloon occlusion of right vertebral artery | 0
embolization of right vertebral artery | 0
harvesting corticocancellous struts and cancellous autograft | 0
exposure of spine from occiput to C7 | 0
ligation of right vertebral artery | 0
laminectomy at C1 | 0
partial laminectomies at C2 and C3 | 0
osteotomies through lateral mass of C2 and vertebral body of C3 | 0
transection of right C2 and C3 nerve roots | 0
posterior instrumentation from occiput to C7 | 0
placement of rib allograft and fibular allograft struts | 0
placement of cancellous iliac crest autograft | 0
tracheostomy | 0
mandibulotomy and transmandibular approach | 0
exposure of anterior cervical spine | 0
ligation of right vertebral artery at C4 | 0
discectomy at C3–4 | 0
excision of posterior longitudinal ligament | 0
mobilization of tumor specimen | 0
intraoperative pathologist review demonstrating negative margins | 0
free vascularized fibular graft (FVFG) | 0
dural tear at clivus | 0
anastomosis of vasculature to facial artery and vein | 0
repair of mandibulotomy | 0
placement into halo vest | 0
disorientation postoperatively | 24
CT scan of head demonstrating cerebellar hemorrhage | 24
progressive recovery of neurological function | 24
febrile with leukocytosis | 120
decline in strength and mentation | 120
CT scan of neck with contrast | 120
fluid collections in operative bed | 120
aspiration of fluid collections | 120
placement of drains | 120
beta-2 transferrin positive | 120
Serratia marcescens infection | 120
initiation of meropenem and vancomycin | 120
improvement in strength and mentation | 168
severe dysphagia | 0
nasogastric tube feeds | 0
percutaneous endoscopic gastrostomy (PEG) tube placement | 600
tracheostomy decannulation | 600
discharge home | 768
CT scan at 3 months postoperatively | 2160
early osseous bridging | 2160
lifelong suppressive antibiotics | 2160
intact strength in extremities | 2160
CT scan at 5 months postoperatively | 3600
complete fusion of FVFG | 3600
removal of halo vest | 3600
initiation of isometric neck exercises | 3600
proton beam radiation | 4320
annual follow-up | 57600
no tumor recurrence | 57600
solid circumferential arthrodesis | 57600
endoscopic swallow evaluation at 3.5 years | 30240
thinning of posterior pharyngeal wall | 30240
plate removal | 30240
improvement in posterior pharyngeal wall | 34560
Neck Disability Index improvement | 57600
death from unrelated condition | 97680
