18 years old | 0
male | 0
type II diabetes | -1080
intravenous medications | -168
intravenous medications for a week | -168
intermittent high-grade fever | -168
generalized dull-aching abdominal pain | -168
turbid urine | -168
decrease in urine output | -168
swelling of both feet | -168
admitted to the hospital | 0
conscious | 0
afebrile | 0
tachycardic | 0
renal angle tenderness bilaterally | 0
high total leukocyte counts with left shift | 0
elevated urea and creatinine levels | 0
pyuria with leukocyte esterase positivity | 0
activated partial thromboplastin time was prolonged | 0
sepsis-induced coagulopathy | 0
ultrasound of the kidneys revealed enlarged kidneys with bilateral renal abscesses | 0
emergency ultrasound-guided drainage of renal abscesses | 0
pus drained was sent for bacterial, fungal, and mycobacterial smear and culture | 0
GenExpert polymerase chain reaction test for Mycobacterium tuberculosis was negative | 0
X-ray chest and electrocardiogram were normal | 0
intravenous meropenem | 0
renal impairment | 0
intravenous voriconazole | 0
intravenous amphotericin B | 0
cultures from both renal abscesses revealed growth of Aspergillus fumigatus | 0
worsening renal function | 0
acute pulmonary edema | 0
hyperkalemia | 0
metabolic acidosis | 0
hemodialysis | 0
noninvasive ventilation | 0
sudden cardiac arrest | 24
aspiration | 24
succumbed to his illness | 24