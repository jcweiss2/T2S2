73 years old | 0
female | 0
abdominal pain | -72
dizziness | -72
decompensated cirrhosis | 0
abdominal infection | 0
spontaneous peritonitis | 0
hypoproteinemia | 0
ARDS | 0
septic shock | 0
noninvasive ventilation | 0
perioral herpes infection | 48
perioral wound | 48
local bleeding | 0
crusting of blood | 0
Prothrombin time 15.9 sec | 0
partial thromboplastin time 34.5 sec | 0
albumin 27.9 g/L | 0
alanine aminotransferase 56 U/L | 0
total bilirubin 129.4 μmol/L |"0
neutrophils 79.2% | 0
hemoglobin 87 g/L | 0
platelet count 48 × 109/L | 0
high sensitivity C-reactive protein 77 mg/L | 0
oral antiviral drugs | 0
topical penciclovir | 0
mupirocin | 0
wet application of topical nitrocilin | 0
antiviral treatment | 0
furacilin | 0
local epinephrine injection | 0
topical thrombin lyophilized powder | 0
wet wound healing approach | 0
discharged | 0
