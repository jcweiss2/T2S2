44 years old | 0
male | 0
pulmonary sarcoidosis | -336
endobronchial ultrasound (EBUS) bronchoscopy | -336
pleuritic chest pain | 0
fever | 0
chills | 0
night sweats | 0
chest pain | 0
chest pain (continuous) | 0
chest pain (sharp) | 0
chest pain (relieved with leaning forward) | 0
tachycardia (110 beats/min) | 0
oxygen saturation (92% on room air) | 0
mild distress | 0
distant heart sounds | 0
no pericardial rubs | 0
oral temperature (97.9°F/36.6°C) | 0
blood pressure (110/71 mm Hg) | 0
no pulsus paradoxus |# 第4章 网络层
