77 years old | 0
female | 0
menopause | -9360
adenocarcinoma | -72
endometrial cytology | -72
magnetic resonance imaging (MRI) | -72
primary malignant tumor | -72
cervical cancer | -72
fluid accumulation in uterine cavity | -72
cervical biopsy | -72
Stage IIB cervical cancer | -72
concurrent chemoradiotherapy (CCRT) | 0
cisplatin | 0
whole-pelvis irradiation | 0
brachytherapy | 0
fever | 72
malaise | 72
COVID-19 negative | 72
discharged from outpatient clinic | 72
decreased consciousness | 96
worsening general condition | 96
Glasgow Coma Scale (GCS) score of 13 | 96
white blood cell count (WBC) | 96
neutrophils | 96
lymphocytes | 96
C-reactive protein (CRP) | 96
computed tomography (CT) imaging | 96
extensive pyometra | 96
small inflammation of small intestine | 96
transcervical drainage | 120
intrauterine purulent material | 120
sepsis | 120
intravenous meropenem | 120
tracheal intubation | 120
anti-epileptic medication | 120
levetiracetam | 120
L. monocytogenes detected in pyometra material | 144
L. monocytogenes detected in blood culture | 144
ampicillin | 144
gentamicin | 144
lumbar puncture (LP) | 144
cerebral spinal fluid (CSF) pressure | 144
CSF examination | 144
FilmArray meningitis/encephalitis panel assay | 144
L. monocytogenes meningitis | 144
ganciclovir | 144
vital signs improved | 576
blood test results improved | 576
moved from intensive care unit | 576
able to open eyes spontaneously | 4032
state of consciousness stable | 4032
Glasgow Coma Scale (GCS) score of 8 | 4032