31 years old|0
male|0
alcohol use disorder|0
generalized fatigue|-72
weakness|-72
myalgias|-72
throat pain|-672
GAS pharyngitis|-672
positive throat culture|-672
completed azithromycin|-672
severe penicillin allergy|-672
fever|-168
chills|-168
nausea|-168
vomiting|-168
arthralgias|-168
myalgias|-168
fatigue|-168
weakness|-168
admitted to hospital|0
febrile|0
tachycardic|0
ill appearing|0
unremarkable cardiac exam|0
unremarkable pulmonary exam|0
unremarkable abdominal exam|0
neutrophilic leukocytosis|0
thrombocytopenia|0
hyponatremia|0
abnormal liver enzymes|0
elevated Nt-ProBNP|0
negative HIV|0
elevated troponin T|0
negative COVID-19 test|0
hepatic steatosis|0
negative acute viral hepatitis panel|0
bilateral striated nephrograms|0
perinephric fat stranding|0
bilateral pyelonephritis|0
mild hepatosplenomegaly|0
continued high fevers|168
worsening myalgias|168
worsening nausea|168
worsening vomiting|168
worsening leukocytosis|168
worsening thrombocytopenia|168
acute hypoxic respiratory failure|168
desaturation|168
chest x-ray|168
CT chest|168
diffuse interstitial markings|168
alveolar markings|168
ground-glass airspace consolidations|168
GAS bacteremia|168
erythromycin resistance|168
clindamycin resistance|168
started vancomycin|168
started cefepime|168
started doxycycline|168
high fevers|168
increasing oxygen requirements|168
non-invasive positive pressure ventilation|168
transferred to higher care|168
transthoracic echocardiogram|168
left ventricular ejection fraction 55–60%|168
thickened aortic valve|168
possible bicuspid aortic valve|168
severe aortic regurgitation|168
possible vegetation|168
Janeway lesions|168
splinter hemorrhages|168
conjunctival hemorrhages|168
desquamative rash|168
hemodynamic instability|168
worsening vital signs|168
worsening heart failure|168
worsening respiratory distress|168
urgent valve surgery|168
aortic root abscess|168
left ventricle involvement|168
partial aortic valve annuloplasty reconstruction|168
incision and drainage of root abscess|168
partial root repair|168
gram positive cocci in culture|168
recovered well|168
sterile blood cultures|168
discharged home|168
completed ceftriaxone|168
