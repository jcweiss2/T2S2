21 years old|0
male|0
blunt abdominal trauma|-?
high-speed collision|-?
major liver laceration|-?
admitted to secondary care hospital|-?
liver packing|-?
received 20 units of packed red blood cells|-?
received fresh frozen plasma|-?
transferred to Armed Forces Hospital|-?
required more blood|-?
required more FFP|-?
continued bleeding from liver laceration|-?
emergency right hepatectomy|-?
intubated|0
mechanical ventilation|0
intensive care unit admission|0
prolonged ICU course|0
pneumothorax|360
sepsis|360
bed sores|360
renal failure|360
coagulopathy|360
cardiac arrest on day 15|360
deranged liver enzymes|0
abnormal liver function|0
abdominal distension|0
bile drainage from abdominal drain|0
endoscopic retrograde cholangiopancreatography (ERCP)|?
confirmed major bile leak from left main bile duct|?
inserted 10 Fr 5 cm plastic stent|?
no sphincterotomy due to coagulopathy|?
improvement in abdominal distension|168
improvement in bile drainage|168
improvement in liver function|168
abdominal distension recurrence|?
deranged liver chemistry|?
high bilirubin|?
high alkaline phosphate|?
anticipated blocked or migrated stent|?
second ERCP|?
stent in place|?
good drainage|?
contrast injection into biliary tree|?
major leak from right hepatic duct stump|?
considered high risk for further surgery|?
plastic stent removed|?
leaking bile branch selectively cannulated|?
0.035 mm Boston Scientific guide wire used|?
metallic endovascular coil deployed|?
3/30 mm coil|?
injection of 1.5 ml NBCA and lipidol mixture|?
marked improvement in liver enzymes|?
marked improvement in bile drainage|?
general condition improved|?
discharged home|?
CT abdomen three months postintervention|2160
endovascular coil in place|2160
six months postdischarge|4320
abdominal pain|4320
low grade fever|4320
mild elevation in liver enzymes|4320
preserved liver function|4320
CT abdomen revealed dilated CBD|4320
radio-opaque object (migrated coil)|4320
treated with antibiotics|4320
ERCP three days after presentation|4320
CBD patent|4320
passed endovascular coil|4320
conflict of interest|0
funding|0
ethical approval|0
author contributions|0
blunt abdominal trauma|0
high-speed collision|0
major liver laceration|0
admitted to secondary care hospital|0
liver packing|0
received 20 units of packed red blood cells|0
received fresh frozen plasma|0
transferred to Armed Forces Hospital|0
required more blood|0
required more FFP|0
continued bleeding from liver laceration|0
emergency right hepatectomy|0
endoscopic retrograde cholangiopancreatography (ERCP)|0
confirmed major bile leak from left main bile duct|0
inserted 10 Fr 5 cm plastic stent|0
no sphincterotomy due to coagulopathy|0
abdominal distension recurrence|168
deranged liver chemistry|168
high bilirubin|168
high alkaline phosphate|168
anticipated blocked or migrated stent|168
second ERCP|168
stent in place|168
good drainage|168
contrast injection into biliary tree|168
major leak from right hepatic duct stump|168
considered high risk for further surgery|168
plastic stent removed|168
leaking bile branch selectively cannulated|168
0.035 mm Boston Scientific guide wire used|168
metallic endovascular coil deployed|168
3/30 mm coil|168
injection of 1.5 ml NBCA and lipidol mixture|168
marked improvement in liver enzymes|168
marked improvement in bile drainage|168
general condition improved|168
discharged home|216
