44 years old | 0
male | 0
admitted to the hospital | 0
fever over 39°C | -216
productive cough | -216
chest pain | -216
treatment with amoxicillin–clavulanate | -216
treatment with paracetamol | -216
anal fissure | -72000
COVID-19 diagnosed | 0
reverse transcriptase-PCR (RT-PCR) testing for SARS-CoV-2 | 0
nasopharyngeal swab | 0
plain film of the chest | 0
right infrahilar opacity | 0
bilateral peripheral reticular pattern | 0
C-reactive protein (CRP) 16.64 mg/dL | 0
procalcitonin (PCT) 0.29 ng/mL | 0
ferritin 1966 ng/mL | 0
D-dimer 1248 ng/mL | 0
international normalized ratio (INR) 1.53 | 0
lactate dehydrogenase (LDH) 380 U/L | 0
minimal neutrophilia | 0
interleukin-6 levels (<3.0 pg/mL) | 0
AST (38 UI/L) | 0
alanine aminotransferase (ALT) (28 UI/L) | 0
bilirubin (1.20 mg/dL) | 0
hepatitis serological tests | 0
hepatitis B virus vaccination | 0
blood and urine cultures | 0
Legionella pneumophila and Streptococcus pneumoniae urinary antigens | 0
Lopinavir/ritonavir 400/100 mg | 0
hydroxychloroquine 200 mg | 0
teicoplanin 400 mg | 48
piperacillin–tazobactam 4.5 g | 48
enoxaparin 4000 UI | 0
improvement of general conditions | 144
resolution of fever | 144
remission of cough | 144
low flow oxygen support | 144
CRP decreased | 144
D-dimer decreased | 144
AST increased | 144
ALT increased | 144
hyperammonaemia | 144
cholinesterase normal | 144
bilirubin normal | 144
alkaline phosphatase normal | 144
gamma-glutamyl transferase slightly increased | 144
treatment with lopinavir/ritonavir and hydroxychloroquine interrupted | 144
acetylcysteine administered | 144
lactulose administered | 144
ultrasound (US) examination of the abdomen | 144
lung high-resolution CT | 144
bi-basal dorsal consolidations | 144
traction bronchiectasis | 144
right inferior lobe | 144
COVID-19 pneumonia | 144
abdominal non-CE-CT | 144
no particular abdominal finding | 144
lung US examination | 144
progressive resolution of subpleural consolidations | 216
complete recovery | 216
no other symptom | 216
CRP normalised | 216
PCT normalised | 216
AST normalised | 216
ALT still increased | 216
D-dimer increased | 216
Echo-color-Doppler examination | 216
inferior vena cava and iliac–femoral–popliteal–infrapopliteal venous axis | 216
no deep thrombosis | 216
lung contrast-enhanced CT (CE-CT) | 216
reduction of consolidations | 216
residual ground glass opacity | 216
intraperitoneal free bubbles | 216
abdominal CE-CT | 216
pneumatosis intestinalis (PI) | 216
caecum and right colon | 216
no filling defects in abdominal aorta and its branches | 216
no portal venous air | 216
no free fluid collection | 216
ciprofloxacin 500 mg | 336
metronidazole 500 mg | 336
enoxaparin 4000 UI | 336
discharged | 432
asymptomatic | 576
abdominal non-CE-CT | 576
complete resolution of PI | 576
laboratory examinations normal | 576
D-dimer slightly increased | 576
ferritin slightly increased | 576
ALT slightly increased | 576
RT-PCR for SARS-CoV-2 negative | 576