29 years old | 0
pregnant | 0
female | 0
admitted to the hospital | 0
fever | -96
cough | -96
second pregnancy | 0
previous pregnancy | -7300
full-term caesarean delivery | -7300
regular antenatal visits | -672
body mass index 35 kg/m2 | 0
anomaly scan at 20 weeks | -672
glucose tolerance test at 24 weeks | -336
last routine antenatal visit | -336
X-ray showed patchy infiltrates | 0
nasopharyngeal swab confirmed COVID-19 | 0
prophylactic medication | 0
shifted to ICU | 72
antibiotic changed to intravenous piperacillin–tazobactam | 72
therapeutic dose of enoxaparin | 72
continuous positive airway pressure | 72
intubated and given mechanical ventilation | 96
midazolam | 144
fentanyl | 144
cisatracurium | 144
effective anticoagulation by heparin infusion | 144
ECMO insertion | 144
VV-ECMO circuit initiated | 144
transferred to Dubai Hospital | 144
fetal heart monitored | 144
repeat COVID-19 swab | 216
COVID-19 swab negative | 216
weaned off ECMO | 240
postdecannulation | 240
haemodynamic stability | 240
discharged from ICU | 336
monitored in general antenatal ward | 336
regular chest physiotherapy sessions | 336
fetal growth parameters normal | 336
Doppler Studies normal | 336
white blood cell count | 0
platelet count | 0
arterial blood gas analysis | 0
coagulation markers | 0
D-dimer | 0
septic markers | 0
blood sugar levels | 0
liver function tests | 0
renal function tests | 0
cardiac markers | 0
ferritin levels | 0
chest X-ray findings | 0
APTT levels | 144
discharged home | 552
outpatient antenatal visit | 672
fetal growth parameters normal | 672
scheduled for regular antenatal follow-ups | 672
transthoracic echocardiography | 672
taper prednisolone | 552
enoxaparin | 552
ambulating | 432
maintaining saturation | 432
haemodynamically stable | 432