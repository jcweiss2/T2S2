fever | -48
abdominal pain | -48
edema of the scrotum | -48
edema of the penis | -48
edema of the perineum | -48
edema of the right gluteal region | -48
hypertension | 0
osteoporosis | 0
hemorrhoids | 0
blood pressure 103/62 mmHg | 0
heart rate 135/min | 0
oxygen saturation 88% | 0
white blood cell count 13.11/μL | 0
C-reactive protein level 61.4 mg/dL | 0
serum creatinine 4.3 mg/dL | 0
blood urea 157 mg/dL | 0
blood sugar 142 mg/dL | 0
procalcitonin 8.53 ng/mL | 0
RT-PCR test for SARS-CoV-2 negative | 0
CT of the abdomen and the pelvis | 0
inflammatory infiltration of the subcutaneous tissues | 0
liquefaction and presence of gas in the subcutaneous tissues | 0
diagnosis of Fournier's gangrene | 0
antibiotic therapy started | 0
meropenem 1 g thrice daily | 0
metronidazole 500 mg thrice daily | 0
linezolid 600 mg twice daily | 0
resection of the necrotic tissues | 12
bilateral orchiectomy | 12
excision of the penile and scrotal skin | 12
transfer to ICU | 12
mechanical ventilation | 12
broad-spectrum antibiotics | 12
supportive and nutritional therapies | 12
colostomy | 24
wound debridement | 24
negative pressure wound therapy | 24
sedation discontinued | 48
recovery of consciousness | 48
extubation | 48
breathing on own with oxygen | 48
hemodynamically stable | 48
diuresis stimulated | 48
inflammatory markers decreased | 48
culture of pus material | 48
Escherichia coli | 48
Pseudomonas aeruginosa | 48
antibiotic therapy modified | 48
cephazolin 1g twice daily | 48
NPWT discontinued | 72
transfer to Department of Plastic Surgery | 72
free-skin grafts applied | 96
discharge | 1104
testosterone supplementation | 1104
physiotherapy | 1104
follow-up | 1104
colostomy reversal | 1104 
free-skin graft care | 1104
regular dressing changes | 1104