57 years old | 0
man | 0
visited emergency department | 0
dyspnea | -48
cough | -48
sputum | -48
left shoulder pain | -48
diaphoresis | -48
myalgia | -48
fever | -48
chilled sensation | -48
diabetes mellitus | -26208
well-controlled diabetes mellitus | -26208
linagliptin | -26208
metformin | -26208
30-pack year smoker | 0
alcohol consumption | 0
marble dust exposure | 0
industrial mask use | 0
raw gizzards consumption | -168
blood pressure 206/109 | 0
heart rate 123 beats/minute | 0
sinus tachycardia | 0
body temperature 38.2°C | 0
left hydropneumothorax | 0
pleural adhesion | 0
multiloculated left pleural effusion | 0
passive atelectasis | 0
pleural enhancement | 0
leukocytosis | 0
white blood cell count 24,300 cells/mm3 | 0
neutrophils 93% | 0
erythrocyte sedimentation rate 121 mm/hr | 0
C-reactive protein 45.8 mg/dL |9 0
arterial partial pressure of oxygen 50.9 mmHg | 0
oxygen applied | 0
hemoglobin A1c 6.9% | 0
aspartate aminotransferase 21 IU/L | 0
alanine aminotransferase 26 IU/L | 0
total bilirubin 0.5 mg/dL | 0
prothrombin time 1.18 INR | 0
albumin 3.0 g/dL | 0
turbid pleural fluid | 0
thick pleural fluid | 0
brownish-yellow pleural fluid | 0
foul odor pleural fluid | 0
exudative pleural fluid | 0
pleural fluid lactate dehydrogenase/serum lactate dehydrogenase 1.08 | 0
pleural fluid glucose 0 mg/dL | 0
pleural fluid white blood cell count 2,976 cells/mm3 | 0
pleural fluid pH 6.34 | 0
ceftriaxone | 24
levofloxacin | 24
clindamycin | 24
chest tube insertion | 24
admitted to intensive care unit | 24
esophago-gastro-duodenoscopy | 48
no esophageal injury | 48
K. kristinae identified | 144
piperacillin-tazobactam | 192
escalated levofloxacin | 192
relapsed fever | 264
discharged | 552
amoxicillin-clavulanic acid | 552
follow-up blood culture negative | 240
improved chest radiographic findings | 552
