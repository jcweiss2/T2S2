64 years old | 0
    male | 0
    obesity | 0
    recurrent olfactory groove meningioma | 0
    left-sided optic neuropathy | 0
    bifrontal craniotomy | -24
    endoscopic resection | -24
    empiric antibiotics | -24
    steroids | -24
    postoperative changes | 0
    pneumocephalus | 0
    new palpable collection below the scalp | 120
    worsening pneumocephalus | 120
    new large scalp collection | 120
    remained at preoperative neurologic baseline | 120
    disorientation | 168
    unsteady gait | 168
    worsening intracranial air | 168
    worsening extracranial air | 168
    mental status decline | 168
    respiratory status decline | 168
    bradycardia | 168
    tachypnea | 168
    hypoxia | 168
    disorientation | 168
    restlessness | 168
    minimal verbal output | 168
    hypoxic respiratory failure | 168
    endotracheal intubation | 168
    emergent bedside needle decompression | 168
    endoscopic exploration | 168
    repair of anterior cranial fossa defect | 168
    profound hypotension | 168
    vasopressors | 168
    diffuse pulmonary edema | 168
    unremarkable transthoracic echocardiogram | 168
    white blood cell count of 44 | 168
    erythrocyte sedimentation rate of 49 mm/h | 168
    C-reactive protein of 11.7 mg/dL | 168
    procalcitonin of 1.17 ng/mL | 168
    platelet count of 521 | 168
    lactate of 2.25 mmol/L | 168
    creatinine of 2.3 mg/dL | 168
    broad-spectrum antibiotics | 168
    negative cultures | 168
    improved pneumocephalus | 216
    laboratory parameters normalized | 264
    kidney function improved | 264
    vasopressors weaned off | 264
    extubated | 264
    CSF white blood cell count of 25 | 408
    CSF glucose of 111 mg/dL | 408
    CSF protein of 194 mg/dL | 408
    CSF lactic acid of 4.1 mmol/L | 408
    negative CSF cultures | 408
    improved to preoperative neurologic baseline | 264
    near-complete resolution of pneumocephalus | 1296
    