85 years old | 0
male | 0
farmer | 0
active lifestyle | 0
admitted to the hospital | 0
transferred to rehabilitation unit | 0
tetanus sequelae | 0
past medical history of atrial fibrillation | -720
past medical history of benign prostatic hypertrophy | -720
injured leg | -720
trismus | -720
hypertonia | -720
C. tetani infection | -720
treatment with immunoglobulins | -720
tetanus vaccination | -720
metronidazole | -720
transferred to ICU | -672
tracheostomy | -672
mechanical ventilation | -672
vasoactive support | -672
respiratory failure | -672
seizures | -672
baclofen | -672
midazolam | -672
diazepam | -672
electroencephalography | -672
slow cerebral activity | -672
opacity on chest radiography | -672
peripheral leukocytosis | -672
possible ventilator-associated pneumonia | -672
blood cultures | -672
tracheal secretion samples | -672
Klebsiella pneumoniae | -672
methicillin-sensitive Staphylococcus aureus | -672
piperacillin-tazobactam | -672
transferred to geriatric unit | -576
coma | -576
breathed spontaneously | -576
supplemental oxygen | -576
antibiotic therapy switched to linezolid | -504
VAP exacerbation | -504
meropenem | -504
septic shock | -504
cholestasis | -432
acute edematous pancreatitis | -432
endoscopic treatment postponed | -432
urinary tract infection | -360
multidrug-resistant organisms | -360
K. pneumoniae | -360
Acinetobacter baumannii | -360
Enterococcus faecalis | -360
colistin | -360
amoxicillin-clavulanate | -360
clinical condition improved | -288
eligible for rehabilitation | -288
MDRO isolation | 0
tracheal supplemental oxygen | 0
bladder catheter | 0
pressure ulcers | 0
sarcopenic | 0
low handgrip strength | 0
appendicular skeletal mass | 0
rehabilitative evaluations | 0
rehabilitation with good compliance | 24
Clostridioides difficile infection | 24
oral vancomycin | 24
atrial fibrillation | 72
third-degree atrioventricular block | 72
heart rate 30 beats/min | 72
single-chamber pacemaker implantation | 96
hyperkinetic delirium | 96
Pseudomonas aeruginosa bloodstream infection | 120
ceftazidime-avibactam | 120
amikacin | 120
SARS-CoV-2 | 120
remdesivir | 120
droplet isolation | 120
second recurrence of C. difficile | 168
fidaxomicin | 168
bloodstream infection | 216
Candida parapsilosis | 216
MSSA | 216
Candida tropicalis | 216
caspofungin | 216
cefazolin | 216
intravenous catheter | 216
piperacillin-tazobactam | 264
aztreonam | 264
ceftazidime-avibactam | 264
antibiotic resistance | 264
cefepime | 312
tracheostomy closure | 360
ENT specialist | 360
pulmonologist | 360
nutritional supplementation | 360
malnutrition | 360
sarcopenia | 360
motor point of view | 360
intensive rehabilitation | 360
infectious complications | 360
non-infectious complications | 360
postural transition | 432
assistance | 432
motor reconditioning | 432
respiratory reconditioning | 432
discharge | 480
posture transition training | 480
aided transfers | 480
axial stability | 480
balance improvement exercises | 480
standing position | 480
breath-movement coordination exercises | 480
thoracic expansion | 480
girdle opening exercises | 480
inhalation-exhalation exercises | 480
wheelchairs | 480
walkers | 480
mobility deficit | 480
safe postural transitions | 480
rehabilitation follow-up | 480
ENT follow-up | 480
geriatric follow-up | 480