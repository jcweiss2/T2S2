26 years old | 0
female | 0
G1P1 | 0
no known prior history of febrile urinary tract infection | 0
no known prior history of flank pain | 0
no known prior history of urolithiasis | 0
normal vaginal delivery | 0
no complications during delivery | 0
uneventful prenatal care | 0
two screening urine analyses and cultures done at 10 and 29 weeks of gestation | -672 and -504
no evidence of infection in urine analyses and cultures | -672 and -504
denies any signs of fever | -672 and -504
denies any lower urinary tract symptoms | -672 and -504
sinus tachycardia | 0
maximal heart rate of 142 beats per minute | 0
tachypnea | 0
dyspnea | 0
respiratory rate ranging between 20 and 24 breaths per minute | 0
hypotension | 0
maximal drop in systolic blood pressure by 30 mmHg | 0
refractory to fluid boluses | 0
no fever | 0
normally contracted uterus | 0
no abnormalities noted in physical exam | 0
elevated white count of 32,500/ml | 0
CT angiography of the chest | 0
huge lesion occupying the right kidney topography | 0
dedicated abdominal and pelvic MRI with Gadolinium | 0
large multi-loculated multi-septated cystic mass | 0
mass arising from the upper pole of the right kidney | 0
measuring 19.0 × 15.5 × 16.5 cm | 0
mass abutting the right hepatic lobe | 0
no definite infiltration | 0
mass effect on the aorta, celiac axis, portal confluence, gallbladder, and pancreas | 0
deviated to the left side | 0
no evidence of any filling defect or obstructing stone | 0
differential diagnosis included multilocular cystic nephroma, cystic renal carcinoma, or hydatid disease | 0
transferred to the Intensive Care Unit | 0
broad-spectrum antibiotic coverage with meropenem and vancomycin | 0
fever developed | 2
Tmax of 39.1 °C | 2
worsening of hemodynamics | 2
lowest mean arterial pressure reached 59 mmHg | 2
decision to proceed with surgical exploration | 2
extended Chevron incision | 4
huge right kidney identified | 4
ascending colon and duodenum medially retracted | 4
perinephric tissue easily dissected anteriorly and caudally | 4
extremely adherent posteriorly and superomedially | 4
attempts to elevate the kidney from the psoas fascia resulted in eruption of a large posterior cyst | 4
massive amount of purulent foul-smelling grey-brown fluid spilled over the field | 4
nephrectomy completed | 4
further cleaning of surrounding suspicious-looking fat tissues | 4
postoperative period uneventful | 4
hemodynamics improved significantly after resection | 4
discharged 4 days postoperatively | 96
heart rate and blood pressure completely normalized | 96
afebrile at the time of discharge | 96
urine and pus culture grew multi-sensitive Escherichia coli | 96
gross specimen weighted 1.26 kg | 96
consisting of a 17 × 16 × 10 cm kidney | 96
mass arising from the upper pole, tan yellow and soft with cystic areas and areas of necrosis | 96
histopathological examination revealed sheets of lipid-laden macrophages, histiocytes, and multinucleated giant cells | 96
involving the renal parenchyma and extending into the perinephric fat and adrenal gland | 96
no evidence of hydatid cyst disease | 96
GMS, PAS, and AFB stains were all negative for microorganisms | 96
diagnosis of xanthogranulomatous pyelonephritis (XGP) | 96
seen 2 weeks after discharge | 336
vital signs within normal range | 336
wound clean with no evidence of infection | 336