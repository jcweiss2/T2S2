55 years old | 0
female | 0
presented to the Emergency Department | 0
fever | -168
malaise | -168
fatigue | -168
decreased appetite | -168
productive cough | -168
abdominal pain | -168
watery diarrhea | -168
mental status changes | -168
nonresponsive to her name | -168
visual hallucinations | -168
denied headache | 0
denied loss of consciousness | 0
denied neck rigidity | 0
denied seizure | 0
denied focal neurological symptoms | 0
denied chest pain | 0
denied hemoptysis | 0
denied difficulty breathing | 0
allergy to penicillin | 0
returned from Ghana | -432
traveled to California | -168
denied malaria prophylaxis | 0
denied vaccination against yellow fever | 0
denied vaccination against hepatitis A virus | 0
developed symptoms in California | -168
discharged following unremarkable examination | -168
normal laboratory results | -168
became lethargic | 0
respiratory distress | 0
oral temperature 38.6°C | 0
heart rate 121 beats/min | 0
respiratory rate 45 breaths/min | 0
SpO2 93% on room air | 0
dry mucous membranes | 0
decreased bilateral breath sounds | 0
tenderness to palpation of left lower quadrant abdomen | 0
no jaundice | 0
no enlarged lymph nodes | 0
no splenomegaly | 0
lethargic | 0
confused | 0
Glasgow coma scale score 14 | 0
pupils equal, round, reactive to light | 0
no cranial nerve deficit | 0
no sensory deficit | 0
supple neck | 0
negative Brudzinski’s sign | 0
negative Kernig’s sign | 0
leukocytosis | 0
white cell count 19,800/µL | 0
neutrophils 44% | 0
lymphocytes 22% | 0
eosinophil 1% | 0
platelets 51,000/µL | 0
hemoglobin 11.8 g/dL | 0
hematocrit 35.3% | 0
red blood cell distribution width 16.9% | 0
lactate dehydrogenase 2714 U/L | 0
haptoglobin <8 mg/dL | 0
prothrombin time/international normalized ratio 14.9/1.4 | 0
troponin 0.161 ng/mL | 0
blood glucose 26 mg/dL | 0
blood urea nitrogen 157 mg/dL | 0
creatinine 7.52 mg/dL | 0
estimated glomerular filtration rate 6 mL/min | 0
bicarbonate 5 mmol/L | 0
anion gap 36 | 0
lactic acid 16.2 mmol/L | 0
sodium 131 mmol/L | 0
potassium 5.5 mmol/L | 0
chloride 91 mmol/L | 0
alanine transaminase 542 U/L | 0
aspartate transaminase 1328 U/L | 0
total bilirubin 14.5 mg/dL | 0
albumin 2.2 g/dL | 0
malaria smear positive | 0
parasitemia 25% | 0
ring forms/trophozoites | 0
developing gametocytes | 0
arterial blood gas pH 7.03 | 0
pCO2 20 | 0
HCO3 0 | 0
mental status deteriorated | 3
Glasgow coma scale score 10/15 | 3
intubated | 3
mechanically ventilated | 3
acute hypoxemic respiratory failure | 3
transferred to ICU | 3
severe malaria diagnosed | 0
Plasmodium falciparum malaria | 0
multi-organ failure | 0
respiratory failure | 0
renal failure | 0
hepatic failure | 0
septic shock | 0
disseminated intravascular coagulation | 0
acute toxic-metabolic encephalopathy | 0
cerebral malaria | 0
acute respiratory distress syndrome | 0
vasopressors started | 0
steroids started | 0
infectious disease consultation | 0
IV quinidine infusion | 0
IV doxycycline | 0
QTc monitoring | 0
blood glucose monitoring | 0
parasitemia monitoring | 0
CDC contacted | 0
artesunate requested | 0
empiric antibiotics started | 0
IV meropenem | 0
IV vancomycin | 0
exchange transfusion considered | 0
QTc prolongation | 24
quinidine switched to IV artesunate | 24
parasitemia improved | 24
acidosis improved | 24
decreased positive end-expiratory pressure | 24
decreased FiO2 requirements | 24
computed tomography of brain unremarkable | 24
lumbar puncture | 24
3 white blood cells per high-power field | 24
neutrophils 12% | 24
lymphocytes 48% | 24
monocytes 38% | 24
no organisms on gram stain | 24
vancomycin discontinued | 24
meropenem discontinued | 24
parasitemia decreased to 0.3% | 72
parasitemia negative | 144
multi-organ failure treated | 0
septic shock treated | 0
renal replacement therapy | 0
platelet transfusions | 0
clinically improving | 72
5-day course of IV artesunate | 0
5-day course of doxycycline | 0
additional 7-day course of oral doxycycline | 144
discharged to rehabilitation facility | 144
favorable outcome | 144
recuperation | 144
