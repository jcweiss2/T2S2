49 years old | 0
male | 0
history of alcohol abuse | 0
presented | 0
concern for esophageal rupture | 0
heavy alcohol consumption | -48
vomiting | -48
severe retrosternal chest pain | -48
severe dyspnea | -48
arrival at the hospital | 0
chest radiograph showed small left pneumothorax | 0
respiratory distress | 0
intubated | 0
admitted to medical intensive care unit | 0
interval chest radiograph showed enlarging left pneumothorax | 24
subcutaneous emphysema | 24
chest tube placed | 24
need for higher level of care | 24
concern for Boerhaave syndrome | 24
life-flighted to tertiary care medical center | -40
arrival at tertiary care center | 0
hypotensive | 0
requiring vasopressor support | 0
concerning for septic shock | 0
CT of chest with oral contrast | 0
diagnosis of esophageal perforation | 0
EGD identified 3-cm linear perforation in distal esophagus | 0
presentation >24 hours since initial event | 0
unstable clinical status | 0
decision to proceed with EndoVAC therapy | 0
EndoVAC procedure repeated every 3-4 days | 24
total of 6 EndoVAC sessions | 168
fed through Dobhoff tube | 0
fed through PEG-J | 168
granulation tissue noticed during fourth EndoVAC | 96
follow-up EGDs | 168
chest CT | 168
barium swallow | 168
confirmed complete healing of esophageal perforation | 168
nothing by mouth | 0
discharge home | N/A
percutaneous feeding tolerated | 168
healed esophageal perforation | 168
no leakage of contrast material | 168
healthy granulation tissue | 96
