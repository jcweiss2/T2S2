61 years old | 0
male | 0
bipolar disorder | -43800
admitted to the Emergency Unit | 0
decreased consciousness level | -120
lithium carbonate medication | -43800
sleepiness | -48
prostration | -48
mental confusion | -48
rigidity of the lower extremities | -48
insulin therapy | -43800
metformin | -43800
thyroxine (T4) | -43800
enalapril | -43800
atenolol | -43800
non-pale | 0
anicteric | 0
acyanotic | 0
rales in pulmonary base | 0
respiratory rate of 29 bpm | 0
irregular cardiac rhythm | 0
heart rate of 130 bpm | 0
blood pressure of 80 × 40 mmHg | 0
abdomen examination was normal | 0
hemoglobin = 12.5 g/dL | 0
hematocrit = 36% | 0
white blood cells (WBC) = 9500/mm³ | 0
platelets 207,000/mm3 | 0
multiple blood cultures negative | 0
chest X-radiography was normal | 0
lithium poisoning | 0
transferred to the intensive care unit (ICU) | 0
hemodialysis | 0
initial lithium serum level was 2.9 mmol/L | 0
creatinine: 2.3 mg/dL | 0
urea: 114 mg/dL | 0
potassium: 3.1 mEq/L | 0
sodium: 145mEq/L | 0
mechanical ventilation | 24
administration of dopamine | 24
brain tomography was normal | 24
electroencephalogram showed metabolic encephalopathy | 24
echocardiogram | 24
mildly dilated left atrium | 24
hypertrophy of the left ventricle | 24
left ventricular systolic function was normal | 24
creatine kinase-MB fraction CKMB level was 132 U/L | 24
cardiac troponin I was 20.92 μg/L | 24
cardiac catheterization | 24
atrial fibrillation | 0
ST segment elevation of 1 mm | 0
T-wave inversion | 0
left ventricular overload | 0
new event of atrial fibrillation | 24
low-ventricular response | 24
bradycardia (HR: 45 bpm) | 24
tachycardia (HR: 174b pm) | 24
electrical cardioversion | 24
ventricular tachycardia | 72
bradyarrhythmia | 72
implantation of temporary intravenous pacemaker | 72
pacemaker turned off | 120
serum lithium levels had decreased to 0.6 mmol/L | 120
control ECG showed sinus rhythm | 120
absence of arrhythmias | 120
tracheostomy | 120
hemorrhagic complications | 144
cardiorespiratory arrest | 144
pulseless electrical activity | 144
resuscitation manoeuvres were unsuccessful | 144
patient died | 144