62 years old | 0
female | 0
history of Ph + ALL | -2160
bone marrow biopsy | -2160
flow cytometry showing predominant immature B-cell population | -2160
expression of CD34 | -2160
expression of CD19 | -2160
expression of CD10 | -2160
expression of cytoplasmic CD79a | -2160
expression of TdT | -2160
induction chemotherapy with hyper-CVAD | -2160
intrathecal methotrexate for two cycles | -2160
nonoliguric acute kidney injury | -2160
hyper-CVAD therapy discontinued | -2160
switched to oral dasatinib | -2160
continued intrathecal methotrexate | -2160
sudden 10 out of 10 headaches | -48
neck pain | -48
back pain | -48
low-grade fever | -48
worsening generalized weakness | -48
increased difficulty with ambulation | -48
confusion | -24
last dose of intrathecal methotrexate | -96
febrile with temperature up to 101.5 degrees Fahrenheit | 0
tachycardic | 0
normotensive | 0
able to describe history | 0
progressively diaphoretic | 0
progressively lethargic | 0
neck stiffness | 0
hemoglobin 6.9 g/dL | 0
transfused with one unit of packed red blood cells | 0
white blood cell count 6.8 K/uL | 0
computed tomography imaging of head | 0
no acute process on head CT | 0
implanted spinal stimulator | 0
contraindication for MRI | 0
neurology consultation | 0
empiric antimicrobial therapy | 0
started on cefepime | 0
started on vancomycin | 0
started on ampicillin | 0
prophylactic fluconazole | 0
prophylactic acyclovir | 0
escalated to treatment-related dosing for acyclovir | 0
diagnostic lumbar puncture attempted | 24
unable to cooperate with procedure | 24
clinically deteriorate | 24
transferred to ICU | 24
agitated | 24
no longer followed commands | 24
rapid sequence intubation | 24
mechanical ventilation | 24
lumbar puncture performed | 24
cerebrospinal fluid cultures showed no growth | 24
negative PCR for herpes simplex virus | 24
negative PCR for varicella-zoster virus | 24
negative PCR for Lyme disease | 24
negative PCR for West Nile virus antibodies | 24
negative upper respiratory panel | 24
negative influenza testing | 24
negative SARS-CoV-2 PCR | 24
gradually improved | 24
hemodynamically stable | 24
extubation | 24
antimicrobial therapy discontinued | 24
prophylactic acyclovir continued | 24
not responding to commands | 24
no spontaneous eye opening | 24
no purposeful movement | 24
transitioned to general ward | 216
encephalopathic | 216
mentation rapidly improved | 240
limited conversations | 240
profound physical weakness | 240
strength began to improve | 240
nasogastric tube removed | 240
began to tolerate oral diet | 240
continued with physical and occupational therapy | 240
able to stand up with assistance | 264
no confusion | 288
no agitation | 288
back to baseline mentation | 288
fever resolved | 288
leukocytosis resolved | 288
recommended rehabilitation therapy | 288
declined extended care facility | 288
provided with home health care | 288
cessation of intrathecal methotrexate | 288
maintained on dasatinib | 288
started on blinatumomab | 288
no further episodes of encephalopathy | 288
