65 years old | 0
female | 0
admitted to the hospital | 0
complaining of worsening respiratory distress | 0
complaining of low back pain | 0
transferred to the intensive care unit | 0
took a drug containing bisphosphonate | -24
for the treatment of osteoporosis | -24
blood pressure was 132/85 mmHg | 0
pulse rate was 145/min | 0
hematocrit of 39% | 0
white-cell count of 10,300/mm3 | 0
serum urea nitrogen of 58 mg/dl | 0
creatinine 1.85 mg/dl | 0
serum sodium 128 mEq/L | 0
potassium 5 mEq/L | 0
chloride 101 mEq/L | 0
lactate dehydrogenase (LDH) was 345 | 0
serum glutamic oxaloacetic transaminase was (SGOT) 90 U/L | 0
creatine kinase (CK) was 422 U/L | 0
bilirubin was 3.07 mg/dl | 0
abnormal coagulation profile | 0
compatible with disseminated intravascular coagulation (DIC) | 0
contrast-enhanced computed tomography (CT) of the abdomen | 0
hypodense zone of the renal cortex | 0
hyperdense medulla | 0
no excretion of contrast media into the collecting system | 0
hemodialysis | 0
anticoagulation | 0
other supportive measures | 0
condition deteriorated | 0
died | 168
renal cortical necrosis | 0
bilateral renal cortical necrosis | 0
renal impairment | 0
acute renal failure | 0 
diffuse acute bilateral RCN | 0 
cortical necrosis | 0 
sepsis | -24 
septic shock | -24 
toxins | -24 
burns | -24 
trauma | -24 
hemorrhagic pancreatitis | -24 
abruptio placentae | -24 
vasoactive substances | -24 
cytotoxic substances | -24 
renal parenchymal damage | -24 
afferent arterioles | -24 
interlobular arteries | -24 
vasospasm | -24 
thrombosis | -24 
renal biopsy | 0 
percutaneous renal biopsy | 0 
CT scan | 0 
intensive care | 0 
dialysis | 0 
renal arteries are patent | 0 
renal cortical enhancement | 0 
subcapsular areas | 0 
juxtamedullary areas | 0 
medulla | 0 
renal tubular necrosis | 0 
renal arterial occlusion | 0 
renal arterial thromboembolism | 0 
striated nephrogram | 0 
wedge-shaped defects | 0 
nephrographic defects | 0 
high-density striations | 0 
renal cortex was not enhanced | 0 
renal medulla was well enhanced | 0 
parenchymal phase | 0 
arterial phase | 0 
CT scan shows | 0 
characteristic finding | 0 
lack of renal cortical enhancement | 0 
thin rim of viable tissue | 0 
dialysis and intensive care | 0 
high mortality and morbidity | 0 
second and third decade | 0 
predominantly female | 0 
pregnancy-related cases | 0 
hypotension | 0 
advanced age | 0 
high mortality | 0 
high morbidity | 0 
rare | 0 
renal cortical necrosis diagnosed | 0 
bilateral renal cortical necrosis diagnosed | 0 
acute renal failure diagnosed | 0 
renal impairment diagnosed | 0 
diffuse acute bilateral RCN diagnosed | 0 
cortical necrosis diagnosed | 0 
sepsis diagnosed | -24 
septic shock diagnosed | -24 
toxins diagnosed | -24 
burns diagnosed | -24 
trauma diagnosed | -24 
hemorrhagic pancreatitis diagnosed | -24 
abruptio placentae diagnosed | -24 
vasoactive substances diagnosed | -24 
cytotoxic substances diagnosed | -24 
renal parenchymal damage diagnosed | -24 
afferent arterioles diagnosed | -24 
interlobular arteries diagnosed | -24 
vasospasm diagnosed | -24 
thrombosis diagnosed | -24 
renal biopsy performed | 0 
percutaneous renal biopsy performed | 0 
CT scan performed | 0 
intensive care provided | 0 
dialysis provided | 0 
renal arteries patent confirmed | 0 
renal cortical enhancement confirmed | 0 
subcapsular areas confirmed | 0 
juxtamedullary areas confirmed | 0 
medulla confirmed | 0 
renal tubular necrosis diagnosed | 0 
renal arterial occlusion diagnosed | 0 
renal arterial thromboembolism diagnosed | 0 
striated nephrogram diagnosed | 0 
wedge-shaped defects diagnosed | 0 
nephrographic defects diagnosed | 0 
high-density striations diagnosed | 0 
renal cortex not enhanced confirmed | 0 
renal medulla well enhanced confirmed | 0 
parenchymal phase confirmed | 0 
arterial phase confirmed | 0 
CT scan shows confirmed | 0 
characteristic finding confirmed | 0 
lack of renal cortical enhancement confirmed | 0 
thin rim of viable tissue confirmed | 0 
dialysis and intensive care provided | 0 
high mortality and morbidity confirmed | 0 
second and third decade confirmed | 0 
predominantly female confirmed | 0 
pregnancy-related cases confirmed | 0 
hypotension confirmed | 0 
advanced age confirmed | 0 
high mortality confirmed | 0 
high morbidity confirmed | 0 
rare confirmed | 0 
renal cortical necrosis confirmed | 0 
bilateral renal cortical necrosis confirmed | 0 
acute renal failure confirmed | 0 
renal impairment confirmed | 0 
diffuse acute bilateral RCN confirmed | 0 
cortical necrosis confirmed | 0 
sepsis confirmed | -24 
septic shock confirmed | -24 
toxins confirmed | -24 
burns confirmed | -24 
trauma confirmed | -24 
hemorrhagic pancreatitis confirmed | -24 
abruptio placentae confirmed | -24 
vasoactive substances confirmed | -24 
cytotoxic substances confirmed | -24 
renal parenchymal damage confirmed | -24 
afferent arterioles confirmed | -24 
interlobular arteries confirmed | -24 
vasospasm confirmed | -24 
thrombosis confirmed | -24 
renal biopsy confirmed | 0 
percutaneous renal biopsy confirmed | 0 
CT scan confirmed | 0 
intensive care confirmed | 0 
dialysis confirmed | 0 
renal arteries patent confirmed | 0 
renal cortical enhancement confirmed | 0 
subcapsular areas confirmed | 0 
juxtamedullary areas confirmed | 0 
medulla confirmed | 0 
renal tubular necrosis confirmed | 0 
renal arterial occlusion confirmed | 0 
renal arterial thromboembolism confirmed | 0 
striated nephrogram confirmed | 0 
wedge-shaped defects confirmed | 0 
nephrographic defects confirmed | 0 
high-density striations confirmed | 0 
renal cortex not enhanced confirmed | 0 
renal medulla well enhanced confirmed | 0 
parenchymal phase confirmed | 0 
arterial phase confirmed | 0 
CT scan shows confirmed | 0 
characteristic finding confirmed | 0 
lack of renal cortical enhancement confirmed | 0 
thin rim of viable tissue confirmed | 0 
dialysis and intensive care confirmed | 0 
high mortality and morbidity confirmed | 0 
second and third decade confirmed | 0 
predominantly female confirmed | 0 
pregnancy-related cases confirmed | 0 
hypotension confirmed | 0 
advanced age confirmed | 0 
high mortality confirmed | 0 
high morbidity confirmed | 0 
rare confirmed | 0 
renal cortical necrosis confirmed | 0 
bilateral renal cortical necrosis confirmed | 0 
acute renal failure confirmed | 0 
renal impairment confirmed | 0 
diffuse acute bilateral RCN confirmed | 0 
cortical necrosis confirmed | 0 
sepsis confirmed | -24 
septic shock confirmed | -24 
toxins confirmed | -24 
burns confirmed | -24 
trauma confirmed | -24 
hemorrhagic pancreatitis confirmed | -24 
abruptio placentae confirmed | -24 
vasoactive substances confirmed | -24 
cytotoxic substances confirmed | -24 
renal parenchymal damage confirmed | -24 
afferent arterioles confirmed | -24 
interlobular arteries confirmed | -24 
vasospasm confirmed | -24 
thrombosis confirmed | -24 
renal biopsy confirmed | 0 
percutaneous renal biopsy confirmed | 0 
CT scan confirmed | 0 
intensive care confirmed | 0 
dialysis confirmed | 0 
renal arteries patent confirmed | 0 
renal cortical enhancement confirmed | 0 
subcapsular areas confirmed | 0 
juxtamedullary areas confirmed | 0 
medulla confirmed | 0 
renal tubular necrosis confirmed | 0 
renal arterial occlusion confirmed | 0 
renal arterial thromboembolism confirmed | 0 
striated nephrogram confirmed | 0 
wedge-shaped defects confirmed | 0 
nephrographic defects confirmed | 0 
high-density striations confirmed | 0 
renal cortex not enhanced confirmed | 0 
renal medulla well enhanced confirmed | 0 
parenchymal phase confirmed | 0 
arterial phase confirmed | 0 
CT scan shows confirmed | 0 
characteristic finding confirmed | 0 
lack of renal cortical enhancement confirmed | 0 
thin rim of viable tissue confirmed | 0 
dialysis and intensive care confirmed | 0 
high mortality and morbidity confirmed | 0 
second and third decade confirmed | 0 
predominantly female confirmed | 0 
pregnancy-related cases confirmed | 0 
hypotension confirmed | 0 
advanced age confirmed | 0 
high mortality confirmed | 0 
high morbidity confirmed | 0 
rare confirmed | 0 
renal cortical necrosis confirmed | 0 
bilateral renal cortical necrosis confirmed | 0 
acute renal failure confirmed | 0 
renal impairment confirmed | 0 
diffuse acute bilateral RCN confirmed | 0 
cortical necrosis confirmed | 0 
sepsis confirmed | -24 
septic shock confirmed | -24 
toxins confirmed | -24 
burns confirmed | -24 
trauma confirmed | -24 
hemorrhagic pancreatitis confirmed | -24 
abruptio placentae confirmed | -24 
vasoactive substances confirmed | -24 
cytotoxic substances confirmed | -24 
renal parenchymal damage confirmed | -24 
afferent arterioles confirmed | -24 
interlobular arteries confirmed | -24 
vasospasm confirmed | -24 
thrombosis confirmed | -24 
renal biopsy confirmed | 0 
percutaneous renal biopsy confirmed | 0 
CT scan confirmed | 0 
intensive care confirmed | 0 
dialysis confirmed | 0 
renal arteries patent confirmed | 0 
renal cortical enhancement confirmed | 0 
subcapsular areas confirmed | 0 
juxtamedullary areas confirmed | 0 
medulla confirmed | 0 
renal tubular necrosis confirmed | 0 
renal arterial occlusion confirmed | 0 
renal arterial thromboembolism confirmed | 0 
striated nephrogram confirmed | 0 
wedge-shaped defects confirmed | 0 
nephrographic defects confirmed | 0 
high-density striations confirmed | 0 
renal cortex not enhanced confirmed | 0 
renal medulla well enhanced confirmed | 0 
parenchymal phase confirmed | 0 
arterial phase confirmed | 0 
CT scan shows confirmed | 0 
characteristic finding confirmed | 0 
lack of renal cortical enhancement confirmed | 0 
thin rim of viable tissue confirmed | 0 
dialysis and intensive care confirmed | 0 
high mortality and morbidity confirmed | 0 
second and third decade confirmed | 0 
predominantly female confirmed | 0 
pregnancy-related cases confirmed | 0 
hypotension confirmed | 0 
advanced age confirmed | 0 
high mortality confirmed | 0 
high morbidity confirmed | 0 
rare confirmed | 0 
renal cortical necrosis confirmed | 0 
bilateral renal cortical necrosis confirmed | 0 
acute renal failure confirmed | 0 
renal impairment confirmed | 0 
diffuse acute bilateral RCN confirmed | 0 
cortical necrosis confirmed | 0 
sepsis confirmed | -24 
septic shock confirmed | -24 
toxins confirmed | -24 
burns confirmed | -24 
trauma confirmed | -24 
hemorrhagic pancreatitis confirmed | -24 
abruptio placentae confirmed | -24 
vasoactive substances confirmed | -24 
cytotoxic substances confirmed | -24 
renal parenchymal damage confirmed | -24 
afferent arterioles confirmed | -24 
interlobular arteries confirmed | -24 
vasospasm confirmed | -24 
thrombosis confirmed | -24 
renal biopsy confirmed | 0 
percutaneous renal biopsy confirmed | 0 
CT scan confirmed | 0 
intensive care confirmed | 0 
dialysis confirmed | 0 
renal arteries patent confirmed | 0 
renal cortical enhancement confirmed | 0 
subcapsular areas confirmed | 0 
juxtamedullary areas confirmed | 0 
medulla confirmed | 0 
renal tubular necrosis confirmed | 0 
renal arterial occlusion confirmed | 0 
renal arterial thromboembolism confirmed | 0 
striated nephrogram confirmed | 0 
wedge-shaped defects confirmed | 0 
nephrographic defects confirmed | 0 
high-density striations confirmed | 0 
renal cortex not enhanced confirmed | 0 
renal medulla well enhanced confirmed | 0 
parenchymal phase confirmed | 0 
arterial phase confirmed | 0 
CT scan shows confirmed | 0 
characteristic finding confirmed | 0 
lack of renal cortical enhancement confirmed | 0 
thin rim of viable tissue confirmed | 0 
dialysis and intensive care confirmed | 0 
high mortality and morbidity confirmed | 0 
second and third decade confirmed | 0 
predominantly female confirmed | 0 
pregnancy-related cases confirmed | 0 
hypotension confirmed | 0 
advanced age confirmed | 0 
high mortality confirmed | 0 
high morbidity confirmed | 0 
rare confirmed | 0 
renal cortical necrosis confirmed | 0 
bilateral renal cortical necrosis confirmed | 0 
acute renal failure confirmed | 0 
renal impairment confirmed | 0 
diffuse acute bilateral RCN confirmed | 0 
cortical necrosis confirmed | 0 
sepsis confirmed | -24 
septic shock confirmed | -24 
toxins confirmed | -24 
burns confirmed | -24 
trauma confirmed | -24 
hemorrhagic pancreatitis confirmed | -24 
abruptio placentae confirmed | -24 
vasoactive substances confirmed | -24 
cytotoxic substances confirmed | -24 
renal parenchymal damage confirmed | -24 
afferent arterioles confirmed | -24 
interlobular arteries confirmed | -24 
vasospasm confirmed | -24 
thrombosis confirmed | -24 
renal biopsy confirmed | 0 
percutaneous renal biopsy confirmed | 0 
CT scan confirmed | 0 
intensive care confirmed | 0 
dialysis confirmed | 0 
renal arteries patent confirmed | 0 
renal cortical enhancement confirmed | 0 
subcapsular areas confirmed | 0 
juxtamedullary areas confirmed | 0 
medulla confirmed | 0 
renal tubular necrosis confirmed | 0 
renal arterial occlusion confirmed | 0 
renal arterial thromboembolism confirmed | 0 
striated nephrogram confirmed | 0 
wedge-shaped defects confirmed | 0 
nephrographic defects confirmed | 0 
high-density striations confirmed | 0 
renal cortex not enhanced confirmed | 0 
renal medulla well enhanced confirmed | 0 
parenchymal phase confirmed | 0 
arterial phase confirmed | 0 
CT scan shows confirmed | 0 
characteristic finding confirmed | 0 
lack of renal cortical enhancement confirmed | 0 
thin rim of viable tissue confirmed | 0 
dialysis and intensive care confirmed | 0 
high mortality and morbidity confirmed | 0 
second and third decade confirmed | 0 
predominantly female confirmed | 0 
pregnancy-related cases confirmed | 0 
hypotension confirmed | 0 
advanced age confirmed | 0 
high mortality confirmed | 0 
high morbidity confirmed | 0 
rare confirmed | 0 
renal cortical necrosis confirmed | 0 
bilateral renal cortical necrosis confirmed | 0 
acute renal failure confirmed | 0 
renal impairment confirmed | 0 
diffuse acute bilateral RCN confirmed | 0 
cortical necrosis confirmed | 0 
sepsis confirmed | -24 
septic shock confirmed | -24 
toxins confirmed | -24 
burns confirmed | -24 
trauma confirmed | -24 
hemorrhagic pancreatitis confirmed | -24 
abruptio placentae confirmed | -24 
vasoactive substances confirmed | -24 
cytotoxic substances confirmed | -24 
renal parenchymal damage confirmed | -24 
afferent arterioles confirmed | -24 
interlobular arteries confirmed | -24 
vasospasm confirmed | -24 
thrombosis confirmed | -24 
renal biopsy confirmed | 0 
percutaneous renal biopsy confirmed | 0 
CT scan confirmed | 0 
intensive care confirmed | 0 
dialysis confirmed | 0 
renal arteries patent confirmed | 0 
renal cortical enhancement confirmed | 0 
subcapsular areas confirmed | 0 
juxtamedullary areas confirmed | 0 
medulla confirmed | 0 
renal tubular necrosis confirmed | 0 
renal arterial occlusion confirmed | 0 
renal arterial thromboembolism confirmed | 0 
striated nephrogram confirmed | 0 
wedge-shaped defects confirmed | 0 
nephrographic defects confirmed | 0 
high-density striations confirmed | 0 
renal cortex not enhanced confirmed | 0 
renal medulla well enhanced confirmed | 0 
parenchymal phase confirmed | 0 
arterial phase confirmed | 0 
CT scan shows confirmed | 0 
characteristic finding confirmed | 0 
lack of renal cortical enhancement confirmed | 0 
thin rim of viable tissue confirmed | 0 
dialysis and intensive care confirmed | 0 
high mortality and morbidity confirmed | 0 
second and third decade confirmed | 0 
predominantly female confirmed | 0 
pregnancy-related cases confirmed | 0 
hypotension confirmed | 0 
advanced age confirmed | 0 
high mortality confirmed | 0 
high morbidity confirmed | 0 
rare confirmed | 0 
renal cortical necrosis confirmed | 0 
bilateral renal cortical necrosis confirmed | 0 
acute renal failure confirmed | 0 
renal impairment confirmed | 0 
diffuse acute bilateral RCN confirmed | 0 
cortical necrosis confirmed | 0 
sepsis confirmed | -24 
septic shock confirmed | -24 
toxins confirmed | -24 
burns confirmed | -24 
trauma confirmed | -24 
hemorrhagic pancreatitis confirmed | -24 
abruptio placentae confirmed | -24 
vasoactive substances confirmed | -24 
cytotoxic substances confirmed | -24 
renal parenchymal damage confirmed | -24 
afferent arterioles confirmed | -24 
interlobular arteries confirmed | -24 
vasospasm confirmed | -24 
thrombosis confirmed | -24 
renal biopsy confirmed | 0 
percutaneous renal biopsy confirmed | 0 
CT scan confirmed | 0 
intensive care confirmed | 0 
dialysis confirmed | 0 
renal arteries patent confirmed | 0 
renal cortical enhancement confirmed | 0 
subcapsular areas confirmed | 0 
juxtamedullary areas confirmed | 0 
medulla confirmed | 0 
renal tubular necrosis confirmed | 0 
renal arterial occlusion confirmed | 0 
renal arterial thromboembolism confirmed | 0 
striated nephrogram confirmed | 0 
wedge-shaped defects confirmed | 0 
nephrographic defects confirmed | 0 
high-density striations confirmed | 0 
renal cortex not enhanced confirmed | 0 
renal medulla well enhanced confirmed | 0 
parenchymal phase confirmed | 0 
arterial phase confirmed | 0 
CT scan shows confirmed | 0 
characteristic finding confirmed | 0 
lack of renal cortical enhancement confirmed | 0 
thin rim of viable tissue confirmed | 0 
dialysis and intensive care confirmed | 0 
high mortality and morbidity confirmed | 0 
second and third decade confirmed | 0 
predominantly female confirmed | 0 
pregnancy-related cases confirmed | 0 
hypotension confirmed | 0 
advanced age confirmed | 0 
high mortality confirmed | 0 
high morbidity confirmed | 0 
rare confirmed | 0 
renal cortical necrosis confirmed | 0 
bilateral renal cortical necrosis confirmed | 0 
acute renal failure confirmed | 0 
renal impairment confirmed | 0 
diffuse acute bilateral RCN confirmed | 0 
cortical necrosis confirmed | 0 
sepsis confirmed | -24 
septic shock confirmed | -24 
toxins confirmed | -24 
burns confirmed | -24 
trauma confirmed | -24 
hemorrhagic pancreatitis confirmed | -24 
abruptio placentae confirmed | -24 
vasoactive substances confirmed | -24 
cytotoxic substances confirmed | -24 
renal parenchymal damage confirmed | -24 
afferent arterioles confirmed | -24 
interlobular arteries confirmed | -24 
vasospasm confirmed | -24 
thrombosis confirmed | -24 
renal biopsy confirmed | 0 
percutaneous renal biopsy confirmed | 0 
CT scan confirmed | 0 
intensive care confirmed | 0 
dialysis confirmed | 0 
renal arteries patent confirmed | 0 
renal cortical enhancement confirmed | 0 
subcapsular areas confirmed | 0 
juxtamedullary areas confirmed | 0 
medulla confirmed | 0 
renal tubular necrosis confirmed | 0 
renal arterial occlusion confirmed | 0 
renal arterial thromboembolism confirmed | 0 
striated nephrogram confirmed | 0 
wedge-shaped defects confirmed | 0 
nephrographic defects confirmed | 0 
high-density striations confirmed | 0 
renal cortex not enhanced confirmed | 0 
renal medulla well enhanced confirmed | 0 
parenchymal phase confirmed | 0 
arterial phase confirmed | 0 
CT scan shows confirmed | 0 
characteristic finding confirmed | 0 
lack of renal cortical enhancement confirmed | 0 
thin rim of viable tissue confirmed | 0 
dialysis and intensive care confirmed | 0 
high mortality and morbidity confirmed | 0 
second and third decade confirmed | 0 
predominantly female confirmed | 0 
pregnancy-related cases confirmed | 0 
hypotension confirmed | 0 
advanced age confirmed | 0 
high mortality confirmed | 0 
high morbidity confirmed | 0 
rare confirmed | 0 
renal cortical necrosis confirmed | 0 
bilateral renal cortical necrosis confirmed | 0 
acute renal failure confirmed | 0 
renal impairment confirmed | 0 
diffuse acute bilateral RCN confirmed | 0 
cortical necrosis confirmed | 0 
sepsis confirmed | -24 
septic shock confirmed | -24 
toxins confirmed | -24 
burns confirmed | -24 
trauma confirmed | -24 
hemorrhagic pancreatitis confirmed | -24 
abruptio placentae confirmed | -24 
vasoactive substances confirmed | -24 
cytotoxic substances confirmed | -24 
renal parenchymal damage confirmed | -24 
afferent arterioles confirmed | -24 
interlobular arteries confirmed | -24 
vasospasm confirmed | -24 
thrombosis confirmed | -24 
renal biopsy confirmed | 0 
percutaneous renal biopsy confirmed | 0 
CT scan confirmed | 0 
intensive care confirmed | 0 
dialysis confirmed | 0 
renal arteries patent confirmed | 0 
renal cortical enhancement confirmed | 0 
subcapsular areas confirmed | 0 
juxtamedullary areas confirmed | 0 
medulla confirmed | 0 
renal tubular necrosis confirmed | 0 
renal arterial occlusion confirmed | 0 
renal arterial thromboembolism confirmed | 0 
striated nephrogram confirmed | 0 
wedge-shaped defects confirmed | 0 
nephrographic defects confirmed | 0 
high-density striations confirmed | 0 
renal cortex not enhanced confirmed | 0 
renal medulla well enhanced confirmed | 0 
parenchymal phase confirmed | 0 
arterial phase confirmed | 0 
CT scan shows confirmed | 0 
characteristic finding confirmed | 0 
lack of renal cortical enhancement confirmed | 0 
thin rim of viable tissue confirmed | 0 
dialysis and intensive care confirmed | 0 
high mortality and morbidity confirmed | 0 
second and third decade confirmed | 0 
predominantly female confirmed | 0 
pregnancy-related cases confirmed | 0 
hypotension confirmed | 0 
advanced age confirmed | 0 
high mortality confirmed | 0 
high morbidity confirmed | 0 
rare confirmed | 0 
renal cortical necrosis confirmed | 0 
bilateral renal cortical necrosis confirmed | 0 
acute renal failure confirmed | 0 
renal impairment confirmed | 0 
diffuse acute bilateral RCN confirmed | 0 
cortical necrosis confirmed | 0 
sepsis confirmed | -24 
septic shock confirmed | -24 
toxins confirmed | -24 
burns confirmed | -24 
trauma confirmed | -24 
hemorrhagic pancreatitis confirmed | -24 
abruptio placentae confirmed | -24 
vasoactive substances confirmed | -24 
cytotoxic substances confirmed | -24 
renal parenchymal damage confirmed | -24 
afferent arterioles confirmed | -24 
interlobular arteries confirmed | -24 
vasospasm confirmed | -24 
thrombosis confirmed | -24 
renal biopsy confirmed | 0 
percutaneous renal biopsy confirmed | 0 
CT scan confirmed | 0 
intensive care confirmed | 0 
dialysis confirmed | 0 
renal arteries patent confirmed | 0 
renal cortical enhancement confirmed | 0 
subcapsular areas confirmed | 0 
juxtamedullary areas confirmed | 0 
medulla confirmed | 0 
renal tubular necrosis confirmed | 0 
renal arterial occlusion confirmed | 0 
renal arterial thromboembolism confirmed | 0 
striated nephrogram confirmed | 0 
wedge-shaped defects confirmed | 0 
nephrographic defects confirmed | 0 
high-density striations confirmed | 0 
renal cortex not enhanced confirmed | 0 
renal medulla well enhanced confirmed | 0 
parenchymal phase confirmed | 0 
arterial phase confirmed | 0 
CT scan shows confirmed | 0 
characteristic finding confirmed | 0 
lack of renal cortical enhancement confirmed | 0 
thin rim of viable tissue confirmed | 0 
dialysis and intensive care confirmed | 0 
high mortality and morbidity confirmed | 0 
second and third decade confirmed | 0 
predominantly female confirmed | 0 
pregnancy-related cases confirmed | 0 
hypotension confirmed | 0 
advanced age confirmed | 0 
high mortality confirmed | 0 
high morbidity confirmed | 0 
rare confirmed | 0 
renal cortical necrosis confirmed | 0 
bilateral renal cortical necrosis confirmed | 0 
acute renal failure confirmed | 0 
renal impairment confirmed | 0 
diffuse acute bilateral RCN confirmed | 0 
cortical necrosis confirmed | 0 
sepsis confirmed | -24 
septic shock confirmed | -24 
toxins confirmed | -24 
burns confirmed | -24 
trauma confirmed | -24 
hemorrhagic pancreatitis confirmed | -24 
abruptio placentae confirmed | -24 
vasoactive substances confirmed | -24 
cytotoxic substances confirmed | -24 
renal parenchymal damage confirmed | -24 
afferent arterioles confirmed | -24 
interlobular arteries confirmed | -24 
vasospasm confirmed | -24 
thrombosis confirmed | -24 
renal biopsy confirmed | 0 
percutaneous renal biopsy confirmed | 0 
CT scan confirmed | 0 
intensive care confirmed | 0 
dialysis confirmed | 0 
renal arteries patent confirmed | 0 
renal cortical enhancement confirmed | 0 
subcapsular areas confirmed | 0 
juxtamedullary areas confirmed | 0 
medulla confirmed | 0 
renal tubular necrosis confirmed | 0 
renal arterial occlusion confirmed | 0 
renal arterial thromboembolism confirmed | 0 
striated nephrogram confirmed | 0 
wedge-shaped defects confirmed | 0 
nephrographic defects confirmed | 0 
high-density striations confirmed | 0 
renal cortex not enhanced confirmed | 0 
renal medulla well enhanced confirmed | 0 
parenchymal phase confirmed | 0 
arterial phase confirmed | 0 
CT scan shows confirmed | 0 
characteristic finding confirmed | 0 
lack of renal cortical enhancement confirmed | 0 
thin rim of viable tissue confirmed | 0 
dialysis and intensive care confirmed | 0 
high mortality and morbidity confirmed | 0 
second and third decade confirmed | 0 
predominantly female confirmed | 0 
pregnancy-related cases confirmed | 0 
hypotension confirmed | 0 
advanced age confirmed | 0 
high mortality confirmed | 0 
high morbidity confirmed | 0 
rare confirmed | 0 
renal cortical necrosis confirmed | 0 
bilateral renal cortical necrosis confirmed | 0 
acute renal failure confirmed | 0 
renal impairment confirmed | 0 
diffuse acute bilateral RCN confirmed | 0 
cortical necrosis confirmed | 0 
sepsis confirmed | -24 
septic shock confirmed | -24 
toxins confirmed | -24 
burns confirmed | -24 
trauma confirmed | -24 
hemorrhagic pancreatitis confirmed | -24 
abruptio placentae confirmed | -24 
vasoactive substances confirmed | -24 
cytotoxic substances confirmed | -24 
renal parenchymal damage confirmed | -24 
afferent arterioles confirmed | -24 
interlobular arteries confirmed | -24 
vasospasm confirmed | -24 
thrombosis confirmed | -24 
renal biopsy confirmed | 0 
percutaneous renal biopsy confirmed | 0 
CT scan confirmed | 0 
intensive care confirmed | 0 
dialysis confirmed | 0 
renal arteries patent confirmed | 0 
renal cortical enhancement confirmed | 0 
subcapsular areas confirmed | 0 
juxtamedullary areas confirmed | 0 
medulla confirmed | 0 
renal tubular necrosis confirmed | 0 
renal arterial occlusion confirmed | 0 
renal arterial thromboembolism confirmed | 0 
striated nephrogram confirmed | 0 
wedge-shaped defects confirmed | 0 
nephrographic defects confirmed | 0 
high-density striations confirmed | 0 
renal cortex not enhanced confirmed | 0 
renal medulla well enhanced confirmed | 0 
parenchymal phase confirmed | 0 
arterial phase confirmed | 0 
CT scan shows confirmed | 0 
characteristic finding confirmed | 0 
lack of renal cortical enhancement confirmed | 0 
thin rim of viable tissue confirmed | 0 
dialysis and intensive care confirmed | 0 
high mortality and morbidity confirmed | 0 
second and third decade confirmed | 0 
predominantly female confirmed | 0 
pregnancy-related cases confirmed | 0 
hypotension confirmed | 0 
advanced age confirmed | 0 
high mortality confirmed | 0 
high morbidity confirmed | 0 
rare confirmed | 0 
renal cortical necrosis confirmed | 0 
bilateral renal cortical necrosis confirmed | 0 
acute renal failure confirmed | 0 
renal impairment confirmed | 0 
diffuse acute bilateral RCN confirmed | 0 
cortical necrosis confirmed | 0 
sepsis confirmed | -24 
septic shock confirmed | -24 
toxins confirmed | -24 
burns confirmed | -24 
trauma confirmed | -24 
hemorrhagic pancreatitis confirmed | -24 
abruptio placentae confirmed | -24 
vasoactive substances confirmed | -24 
cytotoxic substances confirmed | -24 
renal parenchymal damage confirmed | -24 
afferent arterioles confirmed | -24 
interlobular arteries confirmed | -24 
vasospasm confirmed | -24 
thrombosis confirmed | -24 
renal biopsy confirmed | 0 
percutaneous renal biopsy confirmed | 0 
CT scan confirmed | 0 
intensive care confirmed | 0 
dialysis confirmed | 0 
renal arteries patent confirmed | 0 
renal cortical enhancement confirmed | 0 
subcapsular areas confirmed | 0 
juxtamedullary areas confirmed | 0 
medulla confirmed | 0 
renal tubular necrosis confirmed | 0 
renal arterial occlusion confirmed | 0 
renal arterial thromboembolism confirmed | 0 
striated nephrogram confirmed | 0 
wedge-shaped defects confirmed | 0 
nephrographic defects confirmed | 0 
high-density striations confirmed | 0 
renal cortex not enhanced confirmed | 0 
renal medulla well enhanced confirmed | 0 
parenchymal phase confirmed | 0 
arterial phase confirmed | 0 
CT scan shows confirmed | 0 
characteristic finding confirmed | 0 
lack of renal cortical enhancement confirmed | 0 
thin rim of viable tissue confirmed | 0 
dialysis and intensive care confirmed | 0 
high mortality and morbidity confirmed | 0 
second and third decade confirmed | 0 
predominantly female confirmed | 0 
pregnancy-related cases confirmed | 0 
hypotension confirmed | 0 
advanced age confirmed | 0 
high mortality confirmed | 0 
high morbidity confirmed | 0 
rare confirmed | 0 
renal cortical necrosis confirmed | 0 
bilateral renal cortical necrosis confirmed | 0 
acute renal failure confirmed | 0 
renal impairment confirmed | 0 
diffuse acute bilateral RCN confirmed | 0 
cortical necrosis confirmed | 0 
sepsis confirmed | -24 
septic shock confirmed | -24 
toxins confirmed | -24 
burns confirmed | -24 
trauma confirmed | -24 
hemorrhagic pancreatitis confirmed | -24 
abruptio placentae confirmed | -24 
vasoactive substances confirmed | -24 
cytotoxic substances confirmed | -24 
renal parenchymal damage confirmed | -24 
afferent arterioles confirmed | -24 
interlobular arteries confirmed | -24 
vasospasm confirmed | -24 
thrombosis confirmed | -24 
renal biopsy confirmed | 0 
percutaneous renal biopsy confirmed | 0 
CT scan confirmed | 0 
intensive care confirmed | 0 
dialysis confirmed | 0 
renal arteries patent confirmed | 0 
renal cortical enhancement confirmed | 0 
subcapsular areas confirmed | 0 
juxtamedullary areas confirmed | 0 
medulla confirmed | 0 
renal tubular necrosis confirmed | 0 
renal arterial occlusion confirmed | 0 
renal arterial thromboembolism confirmed | 0 
striated nephrogram confirmed | 0 
wedge-shaped defects confirmed | 0 
nephrographic defects confirmed | 0 
high-density striations confirmed | 0 
renal cortex not enhanced confirmed | 0 
renal medulla well enhanced confirmed | 0 
parenchymal phase confirmed | 0 
arterial phase confirmed | 0 
CT scan shows confirmed | 0 
characteristic finding confirmed | 0 
lack of renal cortical enhancement confirmed | 0 
thin rim of viable tissue confirmed | 0 
dialysis and intensive care confirmed | 0 
high mortality and morb