72 years old | 0
man | 0
previously diagnosed colonic adenocarcinoma | 0
underwent aortic aneurysm surgery | -576
fever (37.8°C) | -576
blood collected for culture | -576
urine collected for culture | -576
meropenem plus colistin administered empirically | -576
transferred to intensive care unit | -528
septic shock | -528
gram-negative rods isolated from anaerobic blood culture bottles | 0
obligate anaerobes | 0
catalase-producing | 0
inhibited on Bacteroides bile aesculin agar | 0
resistant to vancomycin (5 μg) | 0
resistant to kanamycin (1 mg) | 0
resistant to colistin sulphate (10 μg) | 0
positive for β-galactosidase | 0
positive for N-acetyl-β-glucosaminidase | 0
positive for glutamic acid decarboxylase | 0
positive for indole | 0
positive for alkaline phosphatase | 0
positive for leucyl glycine | 0
positive for alanine | 0
positive for glutamyl glutamic acid | 0
positive for arylamidases | 0
positive for pyroglutamic acid arylamidase | 0
insufficient identification with Rapid ID 32A | 0
insufficient identification with VITEK MS | 0
16S rRNA gene sequence showing 99% identity to Butyricimonas virosa | 0
investigation of next closely related species | 0
ampicillin sensitivity | 0
sulbactam@ampicillin sensitivity | 0
amoxicillin@clavulanic acid sensitivity | 0
piperacillin@tazobactam sensitivity | 0
imipenem sensitivity | 0
meropenem sensitivity | 0
clindamycin sensitivity | 0
metronidazole sensitivity | 0
did not produce β-lactamase | 0
fever disappeared | 72
clinical condition improved | 72
followed up in intensive care unit | 72
died | 672
Acinetobacter septicaemia | 672
multi-organ failure | 672
positive for alkaline phosphatase |*→
fever (37.8°C) | 0
blood collected for culture | 0
urine collected for culture | 0
meropenem plus colistin administered empirically | 0
transferred to intensive care unit | 24
septic shock | 24
gram-negative rods isolated from anaerobic blood culture bottles | 72
obligate anaerobes | 72
catalase-producing | 72
inhibited on Bacteroides bile aesculin agar | 72
resistant to vancomycin (5 μg) | 72
resistant to kanamycin (1 mg) | 72
resistant to colistin sulphate (10 μg) | 72
positive for β-galactosidase | 72
positive for N-acetyl-β-glucosaminidase | 72
positive for glutamic acid decarboxylase | 72
positive for indole | 72
positive for alkaline phosphatase | 72
positive for leucyl glycine | 72
positive for alanine | 72
positive for glutamyl glutamic acid | 72
positive for arylamidases | 72
positive for pyroglutamic acid arylamidase | 72
insufficient identification with Rapid ID 32A | 72
insufficient identification with VITEK MS | 72
16S rRNA gene sequence showing 99% identity to Butyricimonas virosa | 72
investigation of next closely related species | 72
ampicillin sensitivity | 72
sulbactam@ampicillin sensitivity | 72
amoxicillin@clavulanic acid sensitivity | 72
piperacillin@tazobactam sensitivity | 72
imipenem sensitivity | 72
meropenem sensitivity | 72
clindamycin sensitivity | 72
metronidazole sensitivity | 72
did not produce β-lactamase | 72
