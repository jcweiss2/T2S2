70 years old | 0
male | 0
obstructive sleep apnea | 0
type 2 diabetes | 0
hypertension | 0
BCG instillation | -4
bladder surface tumor | 0
traumatic catheter placement | -4
hemorrhagic catheter placement | -4
deteriorated | 0
admitted to emergency department | 0
flu-like syndrome | 0
fever | 0
chills | 0
oliguric acute kidney injury | 0
liver failure | 0
thrombocytopenia | 0
sepsis biologic signs | 0
transferred to ICU | 0
amoxicillin-clavulanic acid initiated | 0
inflammatory syndrome | 0
hepatic cytolysis | 0
cholestasis | 0
negative sediment cultures | 0
negative urinary cultures | 0
blood cultures for mycobacteria | 0
empirical anti-tuberculous treatment started | 0
chest X-ray showed interstitial syndrome |
