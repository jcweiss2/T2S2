55 years old | 0
    woman | 0
    presented with fever | -168
    presented with dysuria | -168
    presented with malaise | -168
    urinary incontinence | -168
    difficulty ambulating due to worsening back pain | -168
    denied recent illness | 0
    denied hospitalization | 0
    denied back trauma | 0
    denied paraspinal injections | 0
    denied skin infection | 0
    denied weight loss | 0
    denied night sweats | 0
    past medical history of poorly-controlled diabetes mellitus type 2 | 0
    past medical history of hypertension | 0
    past medical history of hyperlipidemia | 0
    past medical history of chronic low back pain | 0
    denied tobacco use | 0
    denied alcohol use | 0
    denied illicit drug abuse | 0
    acutely ill appearance | 0
    diaphoretic | 0
    temperature 38.3°C | 0
    blood pressure 186/82 mmHg | 0
    pulse 114 beats per minute | 0
    respiratory rate 20 breaths per minute | 0
    oxygen saturation 98% on room air | 0
    normal chest examination | 0
    normal abdomen examination | 0
    mild confusion | 0
    lethargic | 0
    normal neurological exam | 0
    electrocardiography showing poor R-wave progression | 0
    electrocardiography showing left ventricular hypertrophy | 0
    chest X-ray no acute process | 0
    white blood cell count 15,600 per cubic millimeter | 0
    neutrophils 87% | 0
    normal comprehensive metabolic panel | 0
    normal coagulation studies | 0
    urine analysis 3+ bacteria | 0
    blood cultures obtained | 0
    urine cultures obtained | 0
    admitted for sepsis secondary to urinary tract infection | 0
    initial antibiotic ceftriaxone | 0
    antibiotic switched to piperacillin-tazobactam | 24
    persistent fever | 24
    worsening mentation | 24
    transferred to medical intensive care unit | 24
    encephalopathy | 24
    generalized weakness | 24
    diminished strength | 24
    diminished tone | 24
    diminished sensation in all extremities | 24
    absent patella tendon reflexes bilaterally | 24
    normal rectal tone | 24
    nuchal rigidity | 24
    moderate tenderness along entire spine | 24
    blood culture gram negative bacilli | 24
    urine culture gram negative bacilli | 24
    antimicrobials widened to vancomycin | 24
    antimicrobials widened to meropenem | 24
    emergent MRI spine with contrast | 24
    extensive posterior epidural fluid collection | 24
    internal air locules extending from C1 to L4 | 24
    mass effect on the cord | 24
    severe thecal sac stenosis in low cervical and mid thoracic levels | 24
    taken to operating room | 24
    underwent cervical decompression | 24
    underwent thoracic decompression | 24
    underwent lumbar decompression | 24
    evacuation of epidural abscess | 24
    aggressive irrigation of epidural abscess | 24
    blood cultures isolated ESBL-producing Klebsiella pneumoniae | 24
    urine cultures isolated ESBL-producing Klebsiella pneumoniae | 24
    abscess cultures isolated ESBL-producing Klebsiella pneumoniae | 24
    sensitive to fluoroquinolones | 24
    sensitive to gentamicin | 24
    sensitive to meropenem | 24
    fungal cultures negative | 24
    acid fast cultures negative | 24
    recovery painstakingly slow | 24
    intensive physical therapy | 24
    intensive occupational therapy | 24
    discharged to skilled nursing facility | 24
    continuation of physical therapy rehabilitation | 24
    remained on meropenem for 12 weeks | 24
    repeat MRI entire spine | 840
    complete resolution of epidural abscess | 840
    <|eot_id|>