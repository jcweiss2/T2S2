23 years old | 0
female | 0
admitted to the hospital | 0
2nd para | 0
P2L1 | 0
cuffed endotracheal tube | -336
ventilated with ambu bag and oxygen supplementation | -336
LUSCS | -408
intrauterine death | -408
oligohydramnios | -408
no fetal cardiac activity | -408
no fetal movement | -408
anterior placenta | -408
emergency LUSCS | -408
oliguric | -288
drowsy | -288
jaundice | -288
high-grade fever | -288
intubated and ventilated | -288
transfused four packed blood cells | -288
transfused 21 fresh frozen plasmas | -288
2½-year-old female baby | -1008
previous LUSCS | -1008
febrile | 0
temperature of 38.9°C | 0
pulse rate of 140/min | 0
blood pressure of 130/80 mmHg | 0
SpO2 of 99% | 0
icterus | 0
pallor | 0
generalized anasarca | 0
abdominal distention | 0
scattered rhonchi | 0
crepitations | 0
abdominal wound clean | 0
urinary catheter in place | 0
nasogastric tube in situ | 0
bleeding per vaginum | 0
intermittent positive pressure ventilation | 0
volume control | 0
pressure support | 0
total leukocyte count of 22,000 cu/mm | 0
polymorphonuclear leukocytosis | 0
hemoglobin of 9.3 g/dl | 0
Prothrombin Time of 17.4 seconds | 0
PTI Index of 74.7 | 0
renal function tests normal | 0
urea of 50 mg/dl | 0
liver function severely deranged | 0
serum glutamic-oxaloacetic transaminase 220 IU/L | 0
serum glutamic pyruvic transaminase 132 IU/L | 0
total bilirubin 3.4 mg/dl | 0
conjugated 2.1 mg/dl | 0
alkaline phosphatase 120 IU/L | 0
total proteins 4.5 g/L | 0
albumin 2.0 g/L | 0
viral markers nonreactive | 0
24 h urine for albumin 2+ positive | 24
samples sent for culture and sensitivity | 24
vasopressor noradrenaline | 48
inotropic dopamine | 48
exploratory laparotomy | 72
intraoperative findings insignificant | 72
collection of serosanguineous fluid | 72
Pantoea dispersa isolated | 96
sensitive to tigecycline | 96
sensitive to colistin | 96
injection colistimethate | 96
loading dose of 9 MU | 96
4.5 MU/day | 96
fibrin degradation products positive | 120
D-Dimer negative | 120
closed tracheal suctioning revealing blood-stained secretions | 120
frank blood | 120
urine showing growth of Candida spp. | 168
ARDS | 168
ventilator support | 168
vasopressors and inotropes | 168
renal failure | 168
multiple dialyses | 168
multiple packs of red blood cells | 168
fresh frozen plasma | 168
total parentral nutrition | 168
enteral nutrition | 168
albumin | 168
cardiac arrest | 432
resuscitated | 432
cardiopulmonary cerebral resuscitation | 432
inotropes and vasopressors | 432
cardiac arrest | 480
declared dead | 480