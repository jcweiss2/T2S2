48 years old | 0
male | 0
Asian | 0
admitted to the hospital | 0
fever | -216
tachycardia | -216
hypotension | -216
swollen right neck | -216
redness | -216
tenderness | -216
warmth | -216
headache | -96
coma | -96
emergency decompressive craniotomy | -96
CVC insertion | -216
CVC inserted through the right subclavian vein | -216
poorly controlled hypertension | -0
no diabetes | -0
no smoking | -0
no alcohol | -0
no drug abuse | -0
farmer | -0
acute fever | 0
hypotension | 0
tachycardia | 0
elevated respiratory rate | 0
septic shock | 0
leukocytosis | 0
elevated inflammatory markers | 0
elevated alanine aminotransferase | 0
elevated aspartate aminotransferase | 0
normal renal function parameters | 0
arterial blood gas measures | 0
POCUS | 0
thrombosis in the right internal jugular vein | 0
gas bubbles in the IJV | 0
misplaced CVC | 0
septic emphysematous thrombophlebitis | 0
CVC removal | 0
fluid resuscitation | 0
intravenous noradrenaline | 0
antibiotic treatment | 0
low-molecular-weight heparin | 0
contrast-enhanced CT scan | 24
swollen right IJV filled by a thrombus | 24
no gas bubbles | 24
CVC and peripheral venous blood cultures | 96
methicillin-resistant Staphylococcus cohnii | 96
sensitivity to vancomycin | 96
CVC-BSI caused by S. cohnii | 96
weaned off vasopressors | 168
symptoms of redness and swelling subsided | 168
left limb weakness | 168
stroke | 168
emphysematous thrombophlebitis | 168
transferred to a general ward | 168
neurological rehabilitation | 168
discharged | 216
full recovery | 216
right IJV thrombus organized | 744
blood flow stable | 744