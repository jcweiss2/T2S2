38 years old | 0
female | 0
referred from peripheral hospital | 0
gestation 32 weeks | 0
previous three pregnancies | -6720
fetal loss at 6-8th months of gestation | -6720
hypocellular bone marrow | 0
severe thrombocytopenia | 0
pregnancy induced hypertension (PIH) | 0
admitted to hospital | 0
hemodynamically stable | 0
blood pressure 140/90 mmHg | 0
methyldopa 250 mg | 0
total leukocyte count 7200/μL | 0
hemoglobin 8.5 g/dl | 0
hematocrit 22.6% | 0
platelet count 6000/mm3 | 0
blood group O negative | 0
pancytopenia | 0
hypoplastic marrow | 0
intrauterine growth retardation (IUGR) | 0
fetal well-being concerns | 0
received 20 units platelets | 0
received 2 units whole blood | 0
clinically very pale | 0
oral prednisolone 10 mg tid | 0
oral hematinic | 0
counts did not improve | 0
repeated platelet concentrate transfusion | 0
antiplatelet antibody negative | 0
ANA negative | 0
antigen test paroxysmal nocturnal hemoglobinopathies negative | 0
factor V mutation negative | 0
direct comb's test negative | 0
Fanconi anemia negative | 0
no abnormality on Hb electrophoresis | 0
advised transfuse single donor platelets peri-operatively | 0
leaking per vaginal | 0
USG Doppler IUGR | 0
intermittent absent end diastolic flow | 0
posted for emergency LSCS | 0
arranged adequate units blood | 0
arranged single donor platelets | 0
fasting status confirmed | 0
high-risk written informed consent | 0
emergency LSCS under general anesthesia | 0
blood pressure 210/100 mmHg | 0
heart rate 160 beats/min | 0
Hb 9.7 g/dl | 0
platelet count 7000/mm3 | 0
taken to Operation theatre | 0
Electrocardiogram attached | 0
Oxygen saturation monitored | 0
Non-invasive Blood Pressure monitors attached | 0
administered IV Nitroglycerine 60 μg | 0
administered IV metoprolol 1.5 mg | 0
transfused 6 units platelets prior induction | 0
pre-medication IV Ranitidine 50 mg | 0
pre-medication IV ondonsetron 4 mg | 0
pre-medication IV glycopyrrolate 0.2 mg | 0
pre-medication IV hydrocortisone 100 mg | 0
pre-oxygenated 100% oxygen | 0
anesthesia induced thiopentone sodium 300 mg | 0
tracheal intubation with succinylcholine 100 mg | 0
administered IV xylocard 50 mg | 0
anesthesia maintained nitrous oxide-oxygen-vecuronium | 0
delivered female infant 960 g | 0
poor Apgar scores ≤4 | 0
infant shifted to NICU | 0
administered Midazolam 1 mg | 0
administered fentanyl 100 μg | 0
stable hemodynamics intra-operatively | 0
total blood loss 1200 ml | 0
transfused 2 units blood | 0
transfused 10 units platelets | 0
reversed neuromuscular blockade neostigmine 0.25 mg | 0
reversed neuromuscular blockade glycopyrollate 0.8 mg | 0
trachea extubated | 0
shifted to PACU | 0
received 2 units blood | 0
received 3 units cryoprecipitates | 0
received 12 units platelets | 0
avoided intramuscular injections | 0
continued prophylactic antibiotics | 0
IV cefuroxime 1.2 gm 12 hourly | 0
IV metronidazole 500 mg 8 hourly |. 0
post-operative analgesia IV paracetamol 15 mg/kg 8 hourly | 0
post-operative persistent hypertension | 0
controlled Nitroglycerine infusion 0.5-1 μg/kg/h | 0
shifted oral antihypertensive Labetalol 100 mg 12 hourly | 0
continued oral prednisolone 10 mg 8 hourly | 0
Hb 9.8 gm | 48
platelet count 28000/mm3 | 48
shifted to ward | 72
discharged | 240
planned bone marrow transplant | 240
