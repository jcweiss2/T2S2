47 years old | 0
female | 0
hypertensive | 0
chronic kidney disease-5 | 0
on thrice weekly hemodialysis | 0
cough | -672
expectoration | -672
breathlessness | -672
fever | -240
amlodipine | -168
erythropoietin | -168
imipenem | -168
admitted to the hospital | 0
conscious | 0
well-oriented | 0
heart rate of 116 beats/min | 0
non-invasive blood pressure of 108/66 mmHg | 0
temperature of 100.2°F | 0
respiratory rate of 34/min | 0
accessory muscles being used | 0
bilateral normal vesicular breath sounds | 0
decreased air entry | 0
occasional coarse crepts in the right lower zone | 0
right lower lobe consolidation/collapse with pleural effusion | 0
blood cultures sent | 0
urine cultures sent | 0
managed in the medical intensive care unit | 0
injection imipenem 500 mg twice daily | 0
total leukocyte count (TLC) up to 28,600/mm3 | 72
repeat blood cultures sent | 72
injection teicoplanin | 72
injection caspofungin | 72
gram-negative coccobacilli in blood | 96
Acinetobacter baumannii | 96
injection colistin | 96
fever decreased | 144
TLC decreased | 144
caspofungin de-escalated | 240
imipenem stopped | 240
abnormal facial twitchings | 384
seizures | 384
injection midazolam | 384
injection phenytoin | 384
generalized tonic clonic seizures | 384
levirecetam | 384
laboratory workup reflected no acute metabolic derangements | 384
liver profile was normal | 384
neuroimaging of the brain | 384
electroencephalography | 384
nerve conduction velocity | 384
lumbar puncture | 384
cerebral spinal fluid (CSF) was clear | 384
CSF biochemistry was within normal limits | 384
colistin stopped | 384
fresh blood cultures sent | 432
blood cultures were sterile | 432
seizures did not recur | 432
antiepileptics tapered | 432
discharged | 792