68 years old | 0
male | 0
admitted to the hospital | 0
type 2 diabetes | 0
high blood pressure | 0
cholecystectomy | - hours unknown
dental extraction | - hours unknown
superior digestive tract hemorrhage | 0
bleeding at home | -1
rushed to the Emergency Room | -1
diagnostic endoscopy | 0
endoscopic hemostasis treatment | 0
lost consciousness | 0
orotracheal intubation | 0
admitted to Intensive Care Unit | 0
altered mental status | 0
ventilator support | 0
stable hemodynamic state | 0
blood pressure 100/60 mmHg | 0
hemoglobin 6.3 g/dL | 0
hematocrit 22% | 0
blood urea 94 mg/dL | 0
blood creatinine 0.7 mg/dL | 0
lactic acid 4.5 mmol/l | 0
glycemia 350 mg/dL | 0
activated partial thromboplastin time 38 seconds | 0
international normalized ratio 0.8 | 0
transaminases 9.9 U/L | 0
direct bilirubin 0.13 mg/dL | 0
total bilirubin 0.3 mg/dL | 0
serum total protein 5 g/dL | 0
serum albumin 28 g/L | 0
transfused with whole blood | 0
transfused with fresh frozen plasma | 0
continuous saline and colloid infusion | 0
hemostatic and prokinetic agents | 0
proton pump inhibitor continuous infusion | 0
osmotic diuretic therapy | 0
pulmonary congestion | 0
cerebral edema | 0
weaned from ventilator | 48
four more episodes of bleeding | 24-72
endoscopic hemostasis attempted | 24-72
chest CT angiography | 72
prolonged prothrombin time | 72
coagulometer test | 96
low plasma value of FVIII | 96
infusion of FVIII concentrate | 96
plasma value of FVIII increased | 108
endoscopic hemostasis | 108
cicatricial ulcer with clips | 120
peripheral blood smear analysis | 120
microcytic, hypochromic red blood cells | 120
hospital acquired infection | 72-120
broad-spectrum antibiotic therapy | 72-120
transferred to Department of Gastroenterology | 168
discharged | 168
mild hemophilia A | 96
esophageal ulcer | 0
digestive bleeding | 0
coagulopathy | 0
severe anemia | 0
cardiac failure | 0
sepsis | 72-120
soft tissue infection | 72-120
stress response | 0
immunosuppressant effect | 72-120
severe bleeding | 0
hypovolemic shock | 0
coagulation tests | 96
FVIII inhibitors | unknown
nephews with mild hemophilia A | unknown