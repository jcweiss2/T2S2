72 years old | 0
male | 0
colonic adenocarcinoma | -672
aortic aneurysm surgery | -576
fever | -576
blood culture | -576
urine culture | -576
meropenem | -576
colistin | -576
septic shock | -552
transferred to intensive care unit | -552
Gram-negative rods isolated | -504
anaerobic blood culture | -504
catalase-producing | -504
inhibited on Bacteroides bile aesculin agar | -504
resistant to vancomycin | -504
resistant to kanamycin | -504
resistant to colistin sulphate | -504
Rapid ID 32A | -504
matrix-assisted laser desorption/ionization time-of-flight | -504
16S rRNA gene sequence | -504
Butyricimonas virosa | -504
investigation of next most closely related species | -504
Butyricimonas paravirosa | -504
Butyricimonas faecihominis | -504
Butyricimonas synergistica | -504
no β-lactamase production | -504
antibiotic susceptibilities | -504
sensitive to ampicillin | -504
sensitive to sulbactam-ampicillin | -504
sensitive to amoxicillin-clavulanic acid | -504
sensitive to piperacillin-tazobactam | -504
sensitive to imipenem | -504
sensitive to meropenem | -504
sensitive to clindamycin | -504
sensitive to metronidazole | -504
fever disappeared | 72
improved clinical condition | 72
followed up in intensive care unit | 72
died | 672
Acinetobacter septicaemia | 672
multi-organ failure | 672