31 years old | 0
    man | 0
    admitted to a hospital | 0
    high fever | 0
    sore throat | 0
    previously healthy | -720
    no medications | -720
    lived with wife and 11-month-old baby boy | -720
    started keeping a dog | -720
    son suffered from high fever | -504
    strawberry tongue | -504
    desquamation of the fingertips | -504
    body temperature 39℃ | 0
    swollen and reddened pharynx | 0
    erythema of the trunk | 0
    erythema of the right thigh | 0
    negative streptococcal antibody tests | 0
    ampicillin/sulbactam | 0
    septic shock | 0
    noradrenalin support | 0
    referred to our hospital | 0
    no gastrointestinal symptoms | 0
    no abdominal pain | 0
    no diarrhea | 0
    well oriented | 0
    blood pressure 112/54 mmHg | 0
    heart rate 110 beats/min | 0
    respiratory rate 24 breaths/min | 0
    oxygen saturation 96% | 0
    body temperature 37.3℃ | 0
    conjunctival congestion | 0
    multiple areas of erythema | 0
    increased white blood cell count | 0
    elevated erythrocyte sedimentation rate | 0
    elevated C-reactive protein | 0
    elevated total bilirubin | 0
    elevated direct bilirubin | 0
    elevated serum ferritin | 0
    elevated soluble interleukin-2 receptor | 0
    elevated brain natriuretic peptide | 0
    elevated procalcitonin | 0
    decreased total protein | 0
    decreased albumin | 0
    normal platelet count | 0
    unremarkable blood cultures | 0
    unremarkable urine cultures | 0
    unremarkable cerebrospinal fluid cultures | 0
    bilaterally enlarged posterior cervical lymph nodes | 0
    pulmonary congestion | 0
    mild splenomegaly | 0
    no abdominal lymphadenopathy | 0
    no ileocecal lymphadenopathy | 0
    IV meropenem | 0
    gamma-globulin | 0
    levofloxacin | 48
    clindamycin | 48
    minocycline | 120
    fever resolution | 0
    general condition improved | 216
    moved to general ward | 216
    bilateral desquamation of fingertips | 216
    Kawasaki disease diagnosis | 216
    increased platelet count | 0
    maximum platelet count 869,000 /μL | 0
    coronary CT angiography | 384
    no coronary lesions | 384
    cardiac ultrasonography | 1440
    negative anti-leptospiral antibodies | 72
    negative anti-leptospiral antibodies | 408
    discharged | 480
    no recurrence | 480
    considered streptococcal toxic shock | 0
    considered staphylococcal toxic shock | 0
    positive Y. pseudotuberculosis antibody | 96
    diagnosed with FESLF | 480
    paired serum samples negative for anti-YPM antibodies | 480
    positive agglutination test for YP2a | 96
    elevated Y. pseudotuberculosis specific antibodies | 480
    