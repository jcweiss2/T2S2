29 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
complex regional pain syndrome | -8760 | 0 | Factual
sports-related injury | -8760 | -8760 | Factual
shoulder surgery | -8760 | -8760 | Factual
recurrent shoulder infections | -8760 | -120 | Factual
Pseudomonas aeruginosa | -120 | -120 | Factual
Sphingomonas paucimobilis | -120 | -120 | Factual
Candida colliculosa | -120 | -120 | Factual
Staphylococcus aureus | -120 | -120 | Factual
left shoulder tendon release | -720 | -720 | Factual
revision | -720 | -720 | Factual
CRPS symptoms | -720 | 0 | Factual
severe pain | -720 | 0 | Factual
allodynia | -720 | 0 | Factual
edema | -720 | 0 | Factual
muscle spasms | -720 | 0 | Factual
temperature changes | -720 | 0 | Factual
electromyography | -168 | -168 | Factual
brachial plexus injury | -168 | -168 | Factual
asthma | -720 | 0 | Factual
selective IgG3 deficiency | -720 | 0 | Factual
oral medical management | -168 | 0 | Factual
opioids | -168 | 0 | Factual
antidepressants | -168 | 0 | Factual
antispasmodics | -168 | 0 | Factual
left stellate ganglion blockade | -168 | -168 | Factual
continuous cervical epidural infusions | -168 | -168 | Factual
epidural catheter placement | 0 | 0 | Factual
fluoroscopic guidance | 0 | 0 | Factual
antibiotic prophylaxis | -1 | 0 | Factual
vancomycin | -1 | 120 | Factual
epidural infusion | 0 | 120 | Factual
bupivacaine | 0 | 120 | Factual
hydromorphone | 0 | 120 | Factual
clonidine | 0 | 120 | Factual
methadone | 0 | 120 | Factual
diazepam | 0 | 120 | Factual
baclofen | 0 | 120 | Factual
amitriptyline | 0 | 120 | Factual
decrease in pain | 24 | 24 | Factual
improved sleep | 48 | 48 | Factual
decrease in LUE spasms | 48 | 48 | Factual
decrease in edema | 48 | 48 | Factual
febrile | 120 | 120 | Factual
temperature 38.1°C | 120 | 120 | Factual
wean the infusion | 120 | 120 | Factual
remove the epidural catheter | 120 | 120 | Factual
headache | 126 | 126 | Factual
neck pain | 126 | 126 | Factual
temperature 40.0°C | 126 | 126 | Factual
neurological examination | 126 | 126 | Factual
blood cultures | 126 | 126 | Factual
urine cultures | 126 | 126 | Factual
chest x-ray | 126 | 126 | Factual
laboratory workup | 126 | 126 | Factual
increase in white count | 126 | 126 | Factual
cefepime | 126 | 216 | Factual
abatement of fever | 144 | 144 | Factual
decrease in white count | 144 | 144 | Factual
MRI | 150 | 150 | Factual
epidural collection | 150 | 150 | Factual
nerve roots compression | 150 | 150 | Factual
interstitial edema | 150 | 150 | Factual
transfer to NSICU | 150 | 150 | Factual
hourly neurological examination | 150 | 216 | Factual
intractable nausea | 216 | 216 | Factual
vomiting | 216 | 216 | Factual
left arm weakness | 216 | 216 | Factual
emergent decompression | 216 | 216 | Factual
evacuation | 216 | 216 | Factual
intraoperative cultures | 216 | 216 | Factual
P aeruginosa | 216 | 216 | Factual
cefepime | 216 | 432 | Factual
vancomycin | 216 | 216 | Factual
resolution of arm weakness | 240 | 240 | Factual
postoperative course | 240 | 432 | Factual
discharged home | 432 | 432 | Factual
intravenous cefepime | 432 | 1008 | Factual