63 years old | 0
woman | 0
relapsed AML | 0
diabetes mellitus | 0
admitted for induction chemotherapy | 0
cytarabine | 0
clofarabine |1
allogeneic stem cell transplantation | 0
developed loose stools | 144
developed diffuse abdominal pain | 144
Clostridium difficile infection | 144
oral metronidazole treatment | 144
abdominal pain persisted | 144
abdominal pain localized to right lower quadrant | 144
neutropenic | 144
afebrile | 144
abdominal CT scan | 144
pelvic CT scan | 144
segmental hypoenhancing area in mid appendix | 144
minimal surrounding fat stranding | 144
appendicitis | 144
no drainable fluid collections | 144
high risk of perioperative morbidity | 144
high risk of mortality | 144
treated with meropenem | 144
hemodynamically normal | 144
right lower quadrant abdominal pain continued | 144
developed localized peritoneal signs | 144
repeat CT scan | 216
stable inflammation of appendix | 216
adjacent loop of small bowel with thickened wall | 216
no extraluminal air | 216
no drainable fluid collections | 216
appendectomy | 216
laparoscopic approach | 216
necrotic appendix | 216
segmentally necrotic terminal ileum | 216
ileocecectomy | 216
primary stapled anastomosis | 216
fascia closed | 216
skin left open | 216
admitted to intensive care unit | 216
extubated on POD1 | 240
empiric meropenem | 240
empiric linezolid | 240
empiric fluconazole | 240
fever to 38.5°C on POD2 | 264
clinically deteriorated on POD4 | 312
re-intubated for tachypnea | 312
re-intubated for hypoxia | 312
chest CT scan | 312
peripheral cavitary lesions | 312
bronchoalveolar lavage | 312
pathological diagnosis of zygomycosis on POD5 | 336
H&E-stained sections | 336
ischemic changes | 336
hemorrhage | 336
thrombosed vessels | 336
broad irregular aseptate hyphae | 336
inflammatory cells rare | 336
GMS-stained sections | 336
wide ribbon-like aseptate hyphae | 336
hyphae branching at wide angles | 336
involving vessels | 336
involving submucosa | 336
invading muscularis propria of appendix | 336
antifungal therapy switched to amphotericin B | 336
fungal overgrowth in surgical wound on POD6 | 360
culture of bronchoalveolar lavage recovered Absidia spp. | 360
severe hypotension | 360
required increasing doses of vasopressors | 360
transitioned to comfort care | 360
expired on POD8 | 408
