61 years old | 0
male | 0
admitted to the hospital | 0
acute dyspnea | 0
productive cough | 0
health care–associated pneumonia | 0
chest x-ray opacities | 0
elevated procalcitonin level | 0
decrease in blood pressure | 24
end-stage renal disease (ESRD) | -10080
hemodialysis | -10080
peripheral artery disease (PAD) | -10080
prior right above-the-knee amputation | -10080
prior left below-the-knee amputation | -10080
type 2 diabetes mellitus | -10080
creation of an AV fistula | -10080
failure of AV fistula | -10080
placement of a tunneled right internal jugular vein hemodialysis catheter | -10080
severe sepsis due to pneumonia | 0
acute coronary syndrome complicated by cardiogenic shock | 0
acute pulmonary embolism | 0
new lateral T-wave inversions | 0
elevated cardiac biomarkers | 0
non-ST-segment elevation myocardial infarction (NSTEMI) | 0
admitted to the cardiac intensive care unit (CICU) | 0
norepinephrine | 0
mean arterial pressure >65 mm Hg | 0
right radial arterial line | 0
transthoracic echocardiography | 0
ejection fraction of 40% | 0
anterior, septal, and apical wall motion abnormalities | 0
absent bilateral femoral arterial pulses | 0
normal left radial pulse | 0
bounding left brachial pulse | 0
high-grade stenoses of the bilateral common iliac arteries | 0
left radial artery access | 0
counterpuncture approach | 0
6-F Glidesheath slender | 0
5-F JR 4 diagnostic catheter | 0
Baby-J guidewire | 0
radial arteriogram | 0
occlusion of the distal brachial artery | 0
patulous vein segment | 0
0.035-inch Wholey wire | 0
angled 0.035-inch Glidewire | 0
0.014-inch Runthrough coronary wire | 0
coronary angiography | 0
heavily calcified 99% lesion in the left anterior descending (LAD) | 0
first diagonal coronary arteries | 0
PCI | 0
6-F EBU 4 guide catheter | 0
exchange-length 0.035-inch J wire | 0
0.038-inch Amplatz Super Stiff guidewire | 0
5-F EBU 4 guide catheter | 0
balloon-assisted tracking (BAT) technique | 0
2.0 × 20-mm Euphora balloon | 0
PCI for the LAD lesion | 0
predilatation with sequential 1.0 × 15-mm, 2.0 × 15-mm, and 2.5 × 15-mm Sapphire balloons | 0
3.0 × 12-mm Resolute Onyx drug-eluting stent | 0
postdilated using a 3.0 × 12-mm Sapphire balloon | 0
PCI of the diagonal lesion | 0
1.0 × 15-mm Sapphire and 2.0 × 20-mm Euphora balloons | 0
2.25 × 22-mm Resolute Onyx stent | 0
transferred back to the CICU | 24
weaned off vasopressors | 24
discharged home | 336
doing well from a cardiac standpoint at 1 year of follow-up | 8760