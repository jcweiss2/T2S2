46 years old | 0
male | 0
admitted to the hospital | 0
fever | 0
hypotension | 0
asthenia | 0
history of arterial hypertension | -672
history of obesity | -672
cardiological examination | -672
electrocardiogram | -672
transthoracic echocardiography | -672
normal findings | -672
COVID-19 infection | -672
rhinitis | -672
mild cough | -672
admitted to ICU | 0
alert | 0
oriented | 0
cooperative | 0
asthenic | 0
blood pressure 85/55 mmHg | 0
heart rate 120 bpm | 0
arterial oxygen saturation 85% | 0
fever with body temperature 38.3 C° | 0
femoral central venous catheter positioned | 0
ECG showed sinus tachycardia | 0
diffuse low voltages | 0
absence of significant repolarization abnormalities | 0
neutrophilic leukocytosis | 0
white blood cell count 26800 x 1000/mm3 | 0
C-reactive protein elevation | 0
C-reactive protein 17.4 mg/dl | 0
Procalcitonin elevation | 0
Procalcitonin 11.7 ng/ml | 0
elevated high sensitivity Troponin | 0
high sensitivity Troponin 23000 ng/L | 0
elevated brain natriuretic peptide | 0
brain natriuretic peptide 6890 pg/ml | 0
elevated creatinine | 0
creatinine 1.8 mg/dl | 0
transaminases and total bilirubin | 0
reverse transcription-polymerase chain reaction (RT-PCR) nasopharyngeal swab for COVID-19 negative | 0
COVID-19 IgM antibody test high IgM levels | 0
transthoracic echocardiography | 0
normal left ventricular cavitary dimensions | 0
diffuse LV parietal thickening | 0
several areas of increased myocardial echogenicity | 0
severely reduced LV global systolic function | 0
ejection fraction 26% | 0
indexed stroke volume 11 ml/m2 | 0
cardiac index 1.3 l/min/m2 | 0
grade II LV diastolic dysfunction | 0
normal cavitary dimensions | 0
reversed global right ventricular systolic function | 0
basal end-diastolic diameter 37 mm | 0
mean diameter of 28 mm | 0
TAPSE 14 mm | 0
tricuspid S-wave velocity at tissue doppler imaging 7.3 cm/sec | 0
inferior vena cava dilated | 0
maximum diameter of 26 mm | 0
inspiratory collapse <50% | 0
right ventricular systolic pressure 41 mmHg | 0
absence of hemodynamically significant valvulopathy | 0
slight amount of pericardial effusion | 0
thoracic computed tomography scan | 0
perivascular aortic and pulmonary adipose tissue imbibition | 0
abdominal ultrasonography | 0
no significant findings | 0
blood cultures started | 0
broad-spectrum antibiotic therapy | 0
INN-daptomycin and piperacillin/tazobactam | 0
crystalloid hydration | 0
nasal cannula ventilatory therapy | 0
norepinephrine in continuous intravenous infusion | 0
therapy with levosimendan initiated | 0
bolus administration avoided | 0
continuous maintenance intravenous infusion | 0
levosimendan dosage 0.1 mcg/kg/min | 0
BP increased to 100/60 mmHg | 12
HR decreased to 110 bpm | 12
further hemodynamic improvement | 24
BP 125/70 mmHg | 24
HR 95 bpm | 24
diuresis 1800 ml | 24
control with TTE | 12
clear and progressive improvement of systolic performance indices | 12
LV EF 66% | 24
dP/dT ratio 1275 mmHg/sec | 24
TAPSE 23 mm | 24
tricuspid S-wave velocity at TDI 11.2 cm/sec | 24
SVi 27 ml/m2 | 24
CI 2.5 l/min/m2 | 24
LV diastolic function improved | 24
IVC maximum diameter 18 mm | 24
RVSP 28 mmHg | 24
diffuse parietal thickening persisted | 24
increased myocardial reflectivity | 24
no significant changes in LV and RV volumes | 24
inflammation indices showed no substantial differences | 24
blood culture results available, all negative | 24
CVC removed | 24
culture of its tip performed, also with negative results | 24
cardiac magnetic resonance imaging (CMR) | 24
normal LV and RV volumes and systolic function | 24
mild hypokinesia of the mid and basal segments | 24
increased signal intensity defined as the ratio of skeletal muscle intensity > 1.9 | 24
edema spread to almost all LV myocardial segments | 24
subendocardial localization at the basal and mid segments | 24
edema and EGE/LGE involving basal segments of the RV and the pericardium | 24
CMR findings defined a picture compatible with immune-mediated myocarditis | 24
endomyocardial biopsy performed | 48
lymphocytic myocarditis confirmed | 48
coronary arteriography | 48
normal coronary circulation | 48
discharged | 168
normal laboratory, electrocardiographic, and echocardiographic findings | 168
TTE performed at 1 and 3 months after discharge | 168