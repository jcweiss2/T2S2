45 years old | 0
woman | 0
semiurban area | 0
intermittent pain abdomen | -2160
loss of appetite | -168
mild breathlessness | -72
no jaundice | 0
no hematemesis | 0
no malena | 0
no nausea | 0
no vomiting | 0
no chest pain | 0
no systemic medical disease |1 0
previous exposure to general anesthesia |0 0
delayed emergence from anesthesia |0 0
heart rate 86/min |0 0
occasional missed beats |0 0
blood pressure 118/72 mmHg |0 0
decreased air entry over left lower zones |0 0
normal cardiovascular examinations |0 0
normal echocardiography |0 0
abnormal ECG with ventricular complexes |0 0
tenderness over left hypochondrium |0 0
tenderness over epigastric region |0 0
no organomegalies |0 0
Mallampati Score grade II |0 0
chest X-ray cystic lesion |0 0
air and fluid level at left lower zones |0 0
CT cystic lesion in hepatic segments |0 0
immunohemagglutination test positive |0 0
hydatid cyst of liver |0 0
hydatid cyst of lower lobe of left lung |0 0
cyst close proximity to heart |0 0
thoracoscopic drainage/excision of lung cyst |0 0
laparoscopic drainage/excision of liver cyst |0 0
albendazole started | -336
normal hemogram |0 0
normal renal function tests |0 0
normal hepatic function tests |0 0
normal blood glucose |0 0
normal viral markers |0 0
normal urine routine examination |0 0
increased SGOT |0 0
increased SGPT |0 0
incentive spirometry taught |0 0
written informed consent |0 0
ranitidine administered | -12
metoclopramide administered | -12
alprazolam administered | -12
general anesthesia planned |0 0
double lumen tube intubation planned |0 0
thoracic epidural analgesia planned |0 0
monitors attached |0 0
intravenous access secured |0 0
hydrocortisone injected |0 0
chlorpheniramine injected |0 0
adrenaline ready |0 0
theophylline ready |0 0
epidural catheter inserted |0 0
test dose lignocaine with adrenaline |0 0
ropivacaine injected |0 0
midazolam administered |0 0
glycopyrrolate administered |0 0
fentanyl administered |0 0
thiopentone sodium induction |0 0
suxamethonium muscle relaxation |0 0
double lumen tube intubation |0 0
bilateral equal air entry confirmed |0 0
ventilation checked |0 0
fiberoptic bronchoscopy confirmed |0 0
anesthesia maintained |0 0
vecuronium bromide maintained |0 0
atracurium avoided |0 0
right lateral decubitus position |0 0
bronchial lumen clamped |0 0
ventilation of right lung |0 0
surgical procedure stopped every 30 min |0 0
both lungs ventilated for 5 min |0 0
bradyarrhythmias observed |0 0
surgeon stopped surgery |0 0
lignocaine administered |0 0
amidarone administered |0 0
surgical procedure accomplished |0 0
supine position |0 0
both lungs ventilated |0 0
monitoring continued |0 0
ABG intermittently done |0 0
parameters within limits |0 0
neostigmine reversal |0 0
glycopyrrolate reversal |0 0
trachea extubated |0 0
shifted to ICU |0 0
epidural top-up ropivacaine |0 0
postoperative ECG normal |0 0
postoperative echocardiography normal |0 0
recovery uneventful |0 0
shifted to surgical ICU |24
