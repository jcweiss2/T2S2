Here is the table of events and timestamps:

39 years old | 0
female | 0
diagnosed with a palpable mass on her right breast | 0
Hodgkin lymphoma | -20016
treated with chemotherapy (6 courses of ABVD) | -20016
mantle field radiation | -20016
inflammatory colitis | -2016
treated with mesalazine | -2016
no specific therapy was ongoing | 0
family history of myxoid liposarcoma | 0
radiological examination of the breast | 0
nodular area of about 30 mm | 0
invasive ductal carcinoma, G3, with triple-negative phenotype and MIB1 85% | 0
staging CT scan of the thorax and abdomen | 0
negative for distant metastasis | 0
neoadjuvant chemotherapy with paclitaxel 80 mg/m2 plus carboplatin AUC2 d1-8-15 q28 for 4 cycles | 0
first cycle completed on April 19, 2017 | 0
port-à-cath insertion | 72
temperature of 38.8°C and normal vital signs | 96
subcutaneous cellulitis and colliquative necrosis | 96
elevated white blood cell count (21,000/mm3), with neutrophilia (16,470/mm3) and elevated C-reactive protein (250 mg/L) | 96
broad-spectrum i.v. antibiotic therapy with piperacillin/tazobactam and daptomycin | 96
PORT rimotion and necrosectomy | 96
defervescence and improvement in subcutaneous cellulitis and blood works | 96
febrile seizure with WBC rise (20,510/mm3) and worsening of skin lesion | 120
second necrosectomy | 120
negative for infection | 120
i.v. catheter tip showed positivity for Klebsiella pneumoniae sensitive to both meropenem and levofloxacin | 120
antibiotic therapy modified accordingly | 120
mediastinitis and bilateral pleural effusion with left pulmonary atelectasis | 120
left thoracoscopy with pleural and mediastinal drainage | 120
admitted to the Intensive Care Unit for observation and support | 120
sepsis | 120
broad-spectrum antibiotic and antifungal therapy, hemodynamic support and non-invasive ventilation | 120
specimens of skin and subcutaneous and muscular tissue from necrosectomy | 120
intensive inflammatory infiltrate including mainly neutrophils | 120
differential diagnosis included PG | 120
systemic methylprednisolone 20 mg/day and topical cyclosporine | 120
progressive resolution of mediastinitis and pleural effusion | 168
wound improvement with scar | 168
blood works indicated progressive normalization of blood count and flogosis index | 168
breast ultrasound | 168
no change in the dimension of the lump | 168
mastectomy and axillary dissection | 168
fibroelastosis and chronic inflammation, with isolated neoplastic cells for maximum 2 mm extension | 168
8 axillary nodes were negative | 168
restaging brain/chest/abdomen CT was negative for distant metastasis | 168
BRCA and p53 mutation tests were negative | 168
released from the hospital | 672
autologous skin graft | 672
PICC implant | 672
resumed chemotherapy with carboplatin and paclitaxel with dose reduction | 672
completed her fourth and last cycle | 672
follow-up | 672