61 years old | 0
male | 0
hypertension | -672
obesity | -672
hyperlipidemia | -672
body mass index: 33 kg/m2 | -672
emergency department presentation | -336
coronavirus disease 2019 pandemic | -336
2-week history of progressive shortness of breath | -336
cough | -336
generalized fatigue | -336
muscle aches | -336
denied chest pain | 0
denied arm pain | 0
denied jaw pain | 0
denied pressure | 0
past medical history negative for diabetes mellitus | 0
past medical history negative for cardiovascular disease | 0
past medical history negative for chronic lung disease | 0
past medical history negative for liver disease | 0
past medical history negative for kidney disease | 0
denied current tobacco use | 0
denied previous tobacco use | 0
visibly distressed | 0
tachypneic | 0
respiratory rate above 50 breaths per minute | 0
hypoxic | 0
blood oxygen saturation of 85% on 15 L oxygen via simple mask | 0
hypotensive | 0
blood pressure 68/42 mm-Hg | 0
tachycardic | 0
heart rate above 140 beats per minute | 0
alert | 0
diaphoretic | 0
significant respiratory distress | 0
weak peripheral pulses | 0
cool extremities | 0
suspected SARS-CoV-2 infection | 0
moved to negative pressure isolation room | 0
decision for early sedation | 0
intubation | 0
circulatory support with norepinephrine | 0
circulatory support with vasopressin | 0
circulatory support with dobutamine | 0
workup for sepsis | 0
workup for septic shock | 0
positive SARS-CoV-2 laboratory result | 0
negative other viral respiratory pathogens | 0
negative bacterial respiratory pathogens | 0
elevated D-dimer level (32 563 ng/mL) | 0
elevated cardiac troponin I level (7.457 ng/mL) | 0
WBC 15.7 (×103/µL) | 0
platelet 151 (×103/µL) | 0
hemoglobin 13.6 g/dL | 0
creatinine 1.16 mg/dL | 0
INR 1.5 | 0
CRP 306.8 mg/L | 0
LDH 707 U/L | 0
IL-6 23 pg/mL | 0
ferritin 2831.22 ng/mL | 0
CK 86 U/L | 0
new diffuse bilateral airspace opacities on chest X-ray | 0
pulmonary infection detected | 0
previous chest X-ray 2 weeks prior | -336
mild cough | -336
myalgia | -336
suspected pulmonary embolism | 0
started on heparin infusion | 0
transthoracic echocardiography performed | 0
hemodynamic instability | 0
risk for patient deterioration during transportation | 0
risk for disease transmission | 0
echocardiography revealed normal right ventricle size | 0
normal right ventricle systolic pressure | 0
mildly elevated pulmonary arterial pressure (31 mm Hg) | 0
moderate global hypokinesis of left ventricle | 0
reduced overall systolic function | 0
ejection fraction 30-35% | 0
previous echocardiography 4 months prior | -2688
LV systolic function normal | -2688
ejection fraction 62% | -2688
electrocardiogram demonstrated diffuse ST elevation (leads I, II, V2-V6) | 0
markedly abnormal ECG | 0
new ischemic changes | 0
previous ECG 2 weeks prior | -336
ECG findings consistent with STEMI | 0
suspicion of acute coronary syndrome | 0
acute coronary occlusion | 0
acute myocarditis | 0
extensive coronary microvascular thrombosis | 0
started on dual antiplatelet therapy (aspirin and ticagrelor) | 0
ongoing heparin infusion | 0
inotropic support with norepinephrine | 0
inotropic support with vasopressin | 0
inotropic support with dobutamine | 0
discussion with interventional cardiology team | 24
deferred coronary angiography | 24
deferred left heart catheterization | 24
suspicion for myocarditis | 24
severe inflammatory state | 24
septic shock | 24
risk of infection transmission | 24
thrombolytics not advised | 24
potential risk for pulmonary hemorrhage | 24
ECG revealed new ST elevation in lead aVF | 48
worsening ST elevation in lead II | 48
worsening ST elevation in anterolateral leads (I, V3-V6) | 48
diffuse ST elevation not confined to single coronary territory | 48
multiple episodes of ventricular tachycardia observed | 48
decision to proceed to emergent LHC | 48
coronary angiography performed | 48
patent left coronary arteries | 48
patent right coronary arteries | 48
no epicardial stenosis | 48
no thrombosis | 48
no delayed coronary filling | 48
left ventriculography negative for Takotsubo cardiomyopathy | 48
diffuse hypokinesis | 48
ejection fraction 40A45% | 48
left ventricular end-diastolic pressure 22 mm Hg | 48
excluded epicardial coronary thrombosis | 48
excluded STEMI | 48
excluded Takotsubo cardiomyopathy | 48
SARS-CoV-2-induced fulminant myocarditis as primary diagnosis | 48
prior thrombosis with distal emboli showering not ruled out | 48
COVID-related micro-thrombotic occlusions not ruled out | 48
started on steroid therapy | 48
cardiac arrest | 72
failed cardiopulmonary resuscitation | 72
expired | 72
autopsy revealed patent coronaries | 72
no significant atherosclerotic changes | 72
no acute myocardial infarct | 72
scattered focal ischemic changes on histopathological examination | 72
hyper-eosinophilic myocytes | 72
nuclear degeneration | 72
no inflammatory neutrophil infiltrates | 72
no myocarditis | 72
no pericarditis | 72
interstitial edema | 72
increased number of macrophages (CD68 staining) | 72
left atrial thrombus (1.5 cm) | 72
marked thromboembolism of left pulmonary artery | 72
diffuse pulmonary vascular microthrombi | 72
pulmonary consolidation | 72
hemorrhage with early hyaline membrane formation | 72
myocardial injury common in SARS-CoV-2 patients | 72
coagulopathy with arterial and pulmonary microthrombi | 72
elevated D-dimer predicts thrombotic complications | 72
cytokine storm contributing to coagulopathy | 72
elevated IL-6 levels | 72
autopsy findings of micro-thrombosis and macro-thrombosis | 72
scattered microscopic cardiomyocyte necrosis | 72
emboli showering from left atrial thrombus | 72
baseline ECG recommended for COVID-19 patients | 72
ST-segment elevation and cTnI as indicators | 72
conservative medical management implemented | 72
LHC demonstrated normal coronaries | 72
Takotsubo cardiomyopathy unlikely | 72
diffuse LV hypokinesis without apical ballooning | 72
definitive diagnosis of PE not made | 72
treated with heparin infusion | 72
plasmapheresis suggested | 72
intra-arterial thrombolysis considered | 72
thrombectomy considered | 72
myocardial injury multifactorial | 72
need for further research on SARS-CoV-2-induced coagulopathy | 72
verbal informed consent obtained | 72
