intrauterine pregnancy | 0
vaginal bleeding | 0
placental remnants in the uterus | 0
surgical evacuation of the uterus | 0
discharged | 0
readmitted | 24
temperature of 39.5°C | 24
abdominal pain | 24
severe endometritis | 24
metronidazole administration | 24
benzylpenicillin administration | 24
gentamicin administration | 24
deterioration | 48
saturation fell to 90% | 48
respiratory rate rose to around 40 breaths per minute | 48
oxygen given by mask | 48
temperature peaked at 40.7°C | 48
C-reactive protein rose to around 300 mg/L | 48
leukocytes to around 15 × 10^9/L | 48
intubated | 48
CT scan | 48
thrombophlebitis of the internal jugular vein | 48
hepatomegaly | 48
Lemierre's syndrome diagnosis | 48
benzylpenicillin discontinued | 48
gentamicin discontinued | 48
tazocin administration | 48
clindamycin administration | 48
metronidazole administration | 48
heparin injections | 48
recovered | 336
discharged | 336
F. necrophorum infection | -6
sore throat | -6
fever | -6
pulmonary infarcts | -6
respiratory dysfunction | -6
arthritic manifestations | -6
multiorgan failure | -6
death | -6 
no shortness of breath | 0
no symptoms from the oropharyngeal tract | 0
no chest pain | 0 
blood cultures showed infection with F. necrophorum | 48
F. necrophorum cultivated from the patient's cervix | 48 
infection originated from the cervix | 48