59 years old | 0
    white woman | 0
    no significant past medical history | 0
    presented as a transfer from an outside facility | 0
    complaining of shortness of breath | 0
    progressively worsening exertional dyspnea | -720
    cough | -720
    weakness in her legs | -720
    atrial fibrillation | 0
    rapid ventricular rate | 0
    started on amiodarone | 0
    started on anticoagulant | 0
    transferred for a higher level of care | 0
    four hospitalizations for worsening dyspnea | 0
    respiratory rate of 27 | 0
    SpO2 of 83% on room air | 0
    microscopic hematuria | 0
    diffuse alveolar hemorrhage | 0
    positive cytoplasmic anti-neutrophil cytoplasmic antibodies | 0
    high proteinase 3 IgG | 0
    Granulomatosis with Polyangiitis (GPA) | 0
    extensive infectious disease workup was negative | 0
    positive qualitative CMV PCR | 0
    lack of other features | 0
    low viral load in bronchoscopy | 0
    concern for active CMV infection was low | 0
    consulted Rheumatology | 0
    consulted Nephrology | 0
    treated with rituximab | 0
    high-dose steroids | 0
    started on 1 mg/kg of prednisone | 0
    plans to taper over six months | 0
    prophylaxis for Pneumocystis jirovecii pneumonia | 0
    received a dose of 1 gm of rituximab | 0
    started on ganciclovir | 0
    possible CMV reactivation prophylactically | 0
    experienced nausea | 0
    experienced chills | 0
    experienced rigors | 0
    resolved on slowing the infusion | 0
    as-needed IV hydrocortisone | 0
    second dose of rituximab (1 gm) | 744
    tolerated well | 744
    IgG level below normal | 768
    IgM level below normal | 768
    IgG 308 mg/dL | 768
    IgM 27 mg/dL | 768
    no fevers | 768
    no concern for infection | 768
    plan to monitor closely | 768
    presented again to Medical Intensive Care Unit | 1344
    intubated | 1344
    sedated | 1344
    acute respiratory failure | 1344
    septic shock with E. coli bacteremia | 1344
    aggressive management including ACLS protocol | 1344
    died | 1344
    no history of recurrent infections | 0
    no sinusitis | 0
    no bronchitis | 0
    no pneumonia | 0
    no organomegaly | 0
    no cytopenias | 0
    suspicion for primary hypogammaglobulinemia was low | 0
    baseline immunoglobulin levels not obtained | 0
    primary hypogammaglobulinemia not ruled out | 0
    