76 years old | 0
female | 0
diagnosed with mesenteric ischemia | 0
scheduled for emergency laparotomy | 0
oral airway assessed as Mallampati Class 2 | 0
no restriction of mouth opening noted | 0
no anticipated difficulty in intubation | 0
flexion and extension of the neck were normal | 0
blood pressure was 100/70 mmHg | 0
tachycardia | 0
tachypnea | 0
hypertensive | 0
diabetic | 0
past history of coronary artery disease | 0
ongoing mesenteric ischemia | 0
severe sepsis syndrome | 0
acute respiratory distress syndrome (ARDS) | 0
low hemoglobin value of 7.6 g/dL | 0
mild hyponatremia of 128 mmol/l | 0
general anesthesia with rapid sequence induction and intubation | 0
preoxygenated for 5 min | -5
Sellick's maneuver applied | 0
given 150 mg of pentothal sodium IV | 0
given 100 mg of rocuronium IV | 0
attempt to open the patient's mouth made | 1
teeth were firmly approximated | 1
mouth could not be opened | 1
no peripheral nerve stimulator | 1
second attempt to open the mouth failed | 2
mask ventilation attempted | 2
jaw was locked | 2
airway obstruction could not be relieved | 2
nasopharyngeal airway used | 2
blind nasal intubation attempted | 2
blind nasal intubation unsuccessful | 2
decision for tracheostomy made | 2
surgeon summoned | 2
tracheostomy performed | 2
patient progressively desaturating | 2
hemodynamics deteriorating | 2
cardiac arrest | 2
attempt to pull anteriorly on the jaw | 2
TMJ displacement suspected | 2
mouth opened to a small degree | 2
patient died | 2
no history of TMJ disorders | -672 
TMJ disease overlooked | -672 
fiberoptic bronchoscope not available | 0 
cricothyroidotomy not considered | 2 
ventilation feasible with nasopharyngeal airway | 2 
low preoperative oxygen reserve | 0 
hemodynamic instability | 0 
apnea period | 2 
tracheostomy attempted | 2 
patient could not be revived | 2