30 years old | 0
woman | 0
anorexia nervosa | 0
body mass index 11 kg/m² | 0
nausea | -72
vomiting | -72
diarrhea | -72
worsening abdominal pain | -72
emaciated | 0
dehydrated | 0
distended abdomen | 0
generalized peritonitis | 0
hypovolemic shock | 0
heart rate 92/min | 0
blood pressure 70/30 mmHg | 0
hypothermic 34.3°C | 0
tachypneic 30/min | 0
oxygen saturation 98% | 0
metabolic acidosis | 0
electrolyte derangement | 0
sodium 116 mmol/L | 0
potassium 3.9 mmol/L | 0
chloride 85 mmol/L | 0
bicarbonate 10 mmol/L | 0
blood urea nitrogen 94 mg/dL | 0
anion gap 21 mmol/L | 0
creatinine 3.01 mg/dL | 0
microcytic anemia | 0
white blood cell count 14,200/mm³ | 0
hemoglobin 10.7 g/dL | 0
hematocrit 31% | 0
mean corpuscular volume 73 fL | 0
platelets 546,000/mm³ | 0
abdominal X-ray portal venous gas | 0
CT scan bowel wall pneumatosis | 0
resuscitation with crystalloids | 0
sodium bicarbonate infusion | 0
nasogastric tube placement | 0
broad spectrum antibiotics | 0
admission to ICU | 0
unstable hemodynamic status | 3
vasoactive agents | 3
exploratory laparotomy | 6
necrosis of entire small bowel | 6
necrosis of right hemicolon | 6
patient expired | 6
previous hospitalizations for severe weakness | -672
previous hospitalizations for electrolyte disbalance | -672
previous hospitalizations for anemia | -672
