Here is the extracted table of clinical events and timestamps:

56 years old | 0
male | 0
janitor | 0
admitted to ICU | 0
diabetes mellitus | -672
hypertension | -672
hyperlipidemia | -672
obesity | -672
antihypertensive association | -672
metformin | -672
glimepiride | -672
atorvastatin | -672
inhaled fluticasone propionate/salmeterol | -672
intermittent fever | -336
muscle ache | -336
nonproductive cough | -168
dyspnea | -168
amoxicillin | -168
pristinamycin | -168
bacterial pneumonia | -168
heart rate 99 beats/min | 0
respiratory rate 34 breaths/min | 0
blood pressure 132/92 mmHg | 0
temperature 38 °C | 0
oxygen saturation 95% | 0
arterial blood gas | 0
pH 7.41 | 0
pCO2 27.9 mmHg | 0
pO2 87.9 mmHg | 0
PaO2/FiO2 87.9 | 0
white blood-cell count 10,720 cells per mm3 | 0
neutrophils 82.6% | 0
lymphocytes 12.7% | 0
lactate dehydrogenase 882 U per liter | 0
CRP 206 mg per deciliter | 0
ferritin 556 ng per milliliter | 0
D-Dimer 2390 ng per milliliter | 0
interleukin-6 93.6 pg per milliliter | 0
SOFA score 8 | 0
hypoxemic respiratory failure | 0
mechanical ventilation | 0
norepinephrine | 0
diabetic ketoacidosis | 0
continuous insulin infusion | 0
acute kidney failure | 0
creatinine level 2.76 mg per deciliter | 0
chest CT | 0
multiple bilateral ground-glass opacities | 0
crazy paving pattern | 0
pulmonary nodules | 0
nasopharyngeal swab | 0
SARS-CoV-2 positive | 0
dexamethasone | 0
eculizumab | 48
piperacillin-tazobactam | 0
cefotaxime | 0
spiramycin | 0
tracheal aspirate | 144
branching hyphae | 144
A. fumigatus culture | 144
A. fumigatus quantitative PCR | 144
serum galactomannan index | 0
serum β-D-Glucan | 0
transthoracic echocardiogram | 144
hypertrophy and dilation of the right ventricle | 144
D-dimer level >20000 ng per milliliter | 144
fibrinogen 3.85 g per liter | 144
cardiac arrest | 168
death | 168
antifungal susceptibility testing | 168
posaconazole resistant | 168
itraconazole resistant | 168
voriconazole resistant | 168
isavuconazole resistant | 168
TR34/L98H mutation | 168