59 years old | 0
woman | 0
hypertension | -120
diabetes | -120
admitted to the hospital | 0
fever | -120
cough | -120
nasal obstruction | -120
diarrhea | -120
denied dyspnea | 0
denied chest pain | 0
axillary temperature 38.5°C | 0
blood pressure 170/102 mmHg | 0
respiratory rate 20 breaths per minute | 0
oxygen saturation 93% | 0
breathing ambient air | 0
leukocytes 9260 per microliter | 0
D-dimer 2404 ng/mL | 0
fibrinogen 954 mg/dL | 0
positive SARS-CoV-2 test | 0
CT chest showed ground-glass opacities | 0
ceftriaxone | 0
azithromycin | 0
oseltamivir | 0
prophylactic low molecular weight heparin | 0
supplemental oxygen 2 L/m | 0
ROTEM performed | 0
hypercoagulability pattern | 0
developed tachypnea | 24
developed dyspnea at rest | 24
oxygen saturation decreased to 88% | 24
oxygen increased to 5 L/m | 24
intubation | 24
mechanical ventilation | 24
fibrinogen 729 mg/dL | 24
IL-6 149 | 24
antithrombin III 107% | 24
D-dimer 40130 ng/mL | 24
suspected pulmonary thromboembolism | 24
started high dose heparin | 24
CT angiography showed PE | 24
extubated after 7 days | 192
pain in right lower limb | 240
right second toe turned blue | 240
no palpable pulses | 240
suspected acute arterial occlusion | 240
femoral arterial line removed | 240
anticoagulation maintained | 240
venous Doppler negative for DVT | 240
echocardiogram showed mild tricuspid regurgitation | 240
arteriography showed stenosis | 240
angioplasty right lower limb | 240
anterior tibial pulse palpable | 240
posterior tibial pulse palpable | 240
persistent second toe pain | 240
amputation of right second toe | 288
discharged | 336
Apixaban 5 mg twice daily | 336
returned to vascular surgeon after 15 days | 552
amputation stump in good condition | 552
denying new complaints | 552
no respiratory symptoms | 552
