47 years old | 0
male | 0
driver | 0
motor vehicle collision | -192
subarachnoid hemorrhage | -192
bilateral lung contusions | -192
rib fractures | -192
blunt abdominal injury | -192
lumbar fractures | -192
open-book pelvic fracture | -192
abdominal CT scan | -192
injury severity score | -192
ascites | -144
diagnostic paracentesis | -144
emergency exploratory laparotomy | -144
mass intestinal fluid | -144
severe edema of the intestinal wall | -144
complete rupture of the jejunum | -144
primary anastomosis | -144
Gram-negative sepsis | -96
hypotension | -96
MODS | -96
acute kidney injury | -96
acute gastrointestinal injury | -96
hyperbilirubinemia | -96
hepatic dysfunction | -96
transfer to trauma referral center | -96
comatose | 0
Glasgow coma scale score 2T1 | 0
shock | 0
acidotic | 0
peritonitic | 0
skin and sclera turned yellow | 0
admitted to TICU | 0
hemodynamic monitoring | 0
abdominal examinations | 0
serial laboratories | 0
imaging | 0
organ support | 0
digestive juice-like fluid | 0
drainage tubes | 0
FAST | 0
mild amount of ascites | 0
CT | 0
extensive exudation | 0
dilated proximal jejunum | 0
multiple orthopedic injuries | 0
DCS | 48
open abdomen management | 48
temporary abdominal closure | 48
TDE | 48
bioelectrical impedance analysis-directed fluid restriction | 72
continuous renal replacement therapy | 72
ultrafiltration rate | 72
net negative fluid balance | 72
bedside dressing change | 72
open abdomen | 72
split-thickness skin grafting | 1872
EN | 120
nutrition support therapy | 120
chyme reinfusion | 192
CR | 192
jejunal feeding tube | 192
chyme reinfusion to distal portion of TDE | 192
distal portion EN | 216
short peptide formula | 216
supplemental enteral glutamine | 216
gut integrity | 216
home EN | 4320
staged reconstruction | 4320
abdominal wall reconstruction | 4320
TDE reversal | 4320
discharge | 4560