63 years old| 0
male | 0
married | 0
smoker | 0
non-drinker | 0
admitted to the hospital | 0
fever | 0
melena | 0
hematemesis | 0
generalized weakness | 0
constant fatigue | 0
shortness of breath | 0
no dysphagia | 0
no dyspepsia | 0
no abdominal pain | 0
no abnormal change of bowel habits | 0
no history of continuous use of NSAIDs | 0
anemia | -24
juxtarenal abdominal aortic aneurysm | -8760
synthetic grafting aortobifemoral bypass | -8760
hypertension | 0
type 2 diabetes mellitus | 0
glaucoma | 0
lens transplantation | 0
ischemic heart disease | 0
catheterization | -8760
stents | -8760
blood pressure medications | 0
diabetes medications | 0
lipid medications | 0
anticoagulant medications | 0
upper GI endoscopy | 0
CT angiogram | 0
opening in the second-third portion of the duodenum | 0
pus discharge | 0
blood coming out | 0
aortoenteric fistula | 0
caecal air bubbles | 0
transferred to Surgical ICU | 0
sepsis | 0
blood pressure 90/50 mmHg | 0
tachycardia 135 bpm | 0
temperature 38°C | 0
white blood cell 5.56 | 0
neutrophil 96.8 | 0
hemoglobin 11.41 | 0
ESR 35 mm/h | 0
CRP 185.4 mg/dl | 0
IV antibiotics | 0
referred to surgical ward | 0
exclusion aortic limb graft | 48
endarterectomy | 48
axillofemoral bypass | 48
femoro-femoral bypass | 48
PTFE graft | 48
transferred to ICU | 48
intestinal adhesion | 96
aorto-duodenal fistula | 96
aortocecal fistula | 96
severe inflammation | 96
unhealthy tissue | 96
infected aortobifemoral graft | 96
pus discharge | 96
large infrarenal AAA | 96
infrarenal aortic neck control | 96
removal of juxtarenal abdominal aortic aneurysm | 96
closure of infrarenal abdominal aorta | 96
fistula management | 96
primary repair of duodenum | 96
right hemicolectomy | 96
primary anastomosis | 96
transferred to SICU | 96
total parental nutrition | 96
stabilized | 96
transferred to surgical ward | 96
oral diet | 96
follow-up CT scan | 240
discharged | 240
afebrile | 240
stable vital signs | 240
