38 years old | 0
primigravida | 0
admitted to the hospital | 0
utero fibroids | 0
superimposed preeclampsia | 0
laparoscopic myomectomy | -5 years
no history of uterine instrumentation | 0
transvaginal ultrasonography | 0
uterine fibroid | 0
multiple other fibroids | 0
methyldopa | -16 weeks
chronic gestational hypertension | -16 weeks
blood pressure 220/120 mmHg | 0
pulse rate 100 bpm | 0
temperature 36.5 °C | 0
urine protein/creatinine ratio 7.39 g/gCr | 0
bilateral butterfly shadows | 0
calcium-channel antagonist | 0
magnesium sulfate | 0
unmanageable blood pressure | 0
emergency CS | 24
lower transverse uterine incision | 24
increased bleeding risk | 24
intensive care | 24
antihypertensive drugs | 24
diuretics | 24
body temperature rose to 38.2 °C | 216
shivering | 216
fever did not last for 2 h | 216
discharged | 336
fever and symptoms resolved | 336
urination | 336
uncomplicated cystitis | 336
high fever | 432
shivering | 432
tachycardia | 432
blood pressure 120/80 mmHg | 432
temperature 40.2 °C | 432
white blood cell count | 432
neutrophils 90% | 432
C-reactive protein 31 mg/dL | 432
internal examination | 432
no uterine tenderness | 432
no malodor of discharge | 432
computer tomography | 432
degenerated 8-cm-sized fibroid | 432
no apparent abscess formation | 432
piperacillin–tazobactam | 432
Gardnerella vaginosis | 432
vaginal discharge culture | 432
no organisms in blood and urine cultures | 432
fever remained | 492
blood urine and vaginal cultures | 492
lumbar spinal magnetic resonance imaging | 492
echocardiography | 492
pelvic MRI scan | 492
12-cm fibroid | 492
edematous changes | 492
increased diffusion-weighted image signal | 492
marginal zone of the degenerative fibroid | 492
myomectomy | 744
resolved fever | 744
WBC and CRP diminished | 744
surgery | 744
no abscess | 744
clear abdominal fluid | 744
uterine surface smooth | 744
incision at the bottom of the uterine fundus | 744
yellow-greenish odorless fluid | 744
1000-g dark red degenerated myoma | 744
histopathology | 744
degenerated leiomyoma | 744
neutrophilic invasion | 744
necrotic lesions | 744
Mycoplasma hominis | 744
mass spectrometry | 744
M. hominis not detected in intraoperative ascites fluid | 744
M. hominis not detected in normal myometrium tissue | 744
M. hominis not detected in degenerated myoma tissue | 744
excellent clinical course | 816
no fever | 816
discharged | 816
oral levofloxacin | 816
stable and symptom-free | 816
blood samples one month postpartum | 1008
no signs of infection | 1008
ultrasound examination | 1008
no abscess or hematoma formation | 1008