43 years old | 0
female | 0
abdominal pain | -720
lumbar pain | -720
nausea | -720
retching | -720
no fever | -720
cesarean sections | -720
cholecystectomy | -720
hiatoplasty for hiatal hernia | -5184
admitted to the hospital | 0
ill-looking appearance | 0
pained expression | 0
pale | 0
anicteric | 0
afebrile | 0
normal respiratory pattern | 0
blood pressure 124/82 mmHg | 0
pulse 84 regular beats per minute | 0
respiratory rate 20 respiratory movements per minute | 0
room air oximetry 98% | 0
normal cardiac examination | 0
normal pulmonary examination | 0
thoracic kyphosis | 0
painful abdominal palpation | 0
negative rebound tenderness test | 0
normal bowel sounds | 0
increased WBC count | 0
increased leucocytes | 0
increased bands | 0
increased eosinophil | 0
increased ALT | 0
increased AST | 0
increased total bilirubin | 0
increased glucose | 0
increased amylase | 0
increased lipase | 0
increased CRP | 0
increased PT | 0
increased urea | 0
abdominal computed tomography | 0
gastric volvulus | 0
organoaxial and mesenteroaxial rotation | 0
herniation of the stomach into the thoracic cavity | 0
splenic arteriovenous vascular pedicle pulled up | 0
pancreatic tail pulled up | 0
tachypnea | 2
decreased oxygen saturation | 2
hypotension | 2
urgent exploratory laparotomy | 4
herniation of the stomach into the chest | 4
gastric volvulus with necrosis and perforation | 4
gastroenteric contents in the left pleural cavity | 4
reduction of the stomach to the abdominal cavity | 4
vertical gastrectomy | 4
thoracic and mediastinal drainage | 4
intensive care unit | 4
sedated | 4
mechanical ventilatory support | 4
norepinephrine infusion | 4
multiple organ failure | 48
death | 48
autopsy | 48
foul-smelling enteric liquid in the pleural cavity | 48
thick brownish fibrinous material on the pericardial and left pleural surface | 48
congestion, edema, alveolar hemorrhage, pneumonia | 48
diffuse alveolar damage | 48
focal thrombosis with infarction of the subpleural parenchyma | 48
acute pleurisy with focal food debris | 48
petechiae on the anterior pericardial surface | 48
chronic myocarditis | 48
diaphragm laceration | 48
gastric serositis | 48
acute pancreatitis with steatonecrosis | 48
hepatic congestion with foci of lobular necrosis | 48
microvesicular steatosis | 48
acute tubular necrosis | 48
foci of recent mucosal and submucosal hemorrhage | 48