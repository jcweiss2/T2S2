37 years old | 0
female | 0
body mass index of 67 kg/m2 | 0
back pain | 0
gastroesophageal reflux disease | 0
obstructive sleep apnea | 0
hyperlipidemia | 0
hypertension | 0
admitted to the hospital | 0
Da Vinci-assisted laparoscopic one-stage single-anastomosis DS procedure | 0
terminal ileum identified | 0
duodeno-ileal anastomosis | 0
greater omentum taken | 0
window created for transection of the duodenum | 0
sleeve gastrectomy | 0
staple line oversewn | 0
duodenum transected | 0
duodenal stump oversewn | 0
two-layer hand sewn anastomosis | 0
anastomosis tested with methylene blue and air | 0
drain placed in left upper quadrant | 0
stomach removed | 0
upper gastrointestinal study on postoperative day 2 | 48
bariatric phase 1 diet started | 48
patient tolerated diet well | 48
discharged on postoperative day 3 | 72
persistent nausea | 264
fatigue | 264
severe abdominal pain | 264
tachycardic | 264
anemic | 264
leukocytosis | 264
abdominal distension | 264
guarding | 264
upper gastrointestinal study | 264
computed tomography of the abdomen | 264
free fluid suggestive of leak or bleeding | 264
diagnostic laparoscopy | 264
hemoperitoneum | 264
evacuation of hemoperitoneum | 264
no active bleeding source | 264
complete inspection of gastroileostomy anastomosis | 264
no leakage seen with methylene blue test | 264
attempt to explore duodenal stump | 264
unsuccessful exploration | 264
three large 19F Blake drains placed | 264
transfused with 2 units of packed red blood cells | 264
kept intubated | 264
sent to intensive care unit | 264
doing well | 288
transferred to step down | 288
hypotensive | 360
unresponsive to fluids | 360
increased sanguinous output | 360
frank bile | 360
elevated bilirubin | 360
elevated amylase | 360
tachycardic | 360
taken back to operating room | 360
exploratory laparotomy | 360
gastroduodenal artery bleeding | 360
over-sewn | 360
duodenal stump blowout | 360
Malecot tube placed | 360
purse-string suture | 360
abdomen closed | 360
drains placed | 360
blood loss | 360
received 5 units of PRBCs | 360
received 4 units of fresh frozen plasma | 360
transferred to ICU | 360
hemorrhagic fluid collections | 432
atelectasis | 432
acute thrombosis of left internal jugular and subclavian veins | 432
pulmonary embolism ruled out | 432
therapeutic Lovenox | 432
octreotide | 432
intravenous piperacillin/taxobactam | 432
changed to cefazolin | 432
discharged on postoperative day 17 | 408
home health care | 408
dressing changes | 408
total parenteral nutrition | 408