14 years old | 0
female | 0
admitted to the hospital | 0
fatigue | -168
nose bleeding | -168
generalized ecchymosis | -168
arthralgia | -168
pallor | 0
tachycardia | 0
dermal/mucosal petechiae | 0
ecchymosis | 0
liver 6 cm palpable | 0
spleen 4 cm palpable | 0
WBC 333,000/mm3 | 0
hemoglobin 4 g/dl | 0
platelet count 29,000/mm3 | 0
L1-type blasts 97% | 0
myeloperoxidase negative | 0
Pre-B-cell ALL | 0
transaminases normal | 0
blood urine nitrogen normal | 0
creatinine normal | 0
uric acid normal | 0
phosphor normal | 0
lactate dehydrogenase high | 0
leukopheresis | -24
leukopheresis | -24
lumbar punction | 96
no cells in cerebrospinal fluid | 96
benign cytology | 96
modified BFM protocol | 0
Turk ALL 2000 | 0
poor steroid response | 192
blast count 1,395/mm3 | 192
no hematologic remission | 360
blast rate 27% | 360
no hematologic remission | 792
blast rate 12% | 792
BCR-ABL fusion gene positive | 0
t(9;22) | 0
High Risk block therapy | 0
imatinib 400 mg/m2/day | 0
severe mucositis | 0
total parenteral nutrition | 0
severe gastrointestinal hemorrhage | 0
erythrocyte transfusion | 0
platelet transfusion | 0
severe neutropenia | 0
fever 39°C | 0
CRP positive | 0
remission | 888
depressive mood | 888
no verbal cooperation | 888
decreased muscle strength | 888
increased muscle tonus | 888
deep tendon reflex | 888
Babinski test positive | 888
cranial magnetic resonance imaging normal | 888
severe mucositis | 1032
hemorrhagic diarrhea | 1032
typhlitis | 1032
hyperemesis | 1032
total parenteral nutrition | 1032
unconsciousness | 1032
Glasgow coma score 7 | 1032
cardiac pulse 34/min | 1032
arterial blood pressure 70/30 mm Hg | 1032
capillary perfusion time 3 s | 1032
hypothermic | 1032
WBC 2,030/mm3 | 1032
absolute neutrophil count 1,640/mm3 | 1032
hemoglobin 5.09 g/dl | 1032
platelets 44,000/mm3 | 1032
CRP 6.8 mg/dl | 1032
urea 113 mg/dl | 1032
creatinine 0.9 mg/dl | 1032
glucose 136 mg/dl | 1032
AST 77 IU/l | 1032
ALT 91 IU/l | 1032
bilirubin 0.3 mg/dl | 1032
GGT 88 IU/l | 1032
prothrombin time 17.6 s | 1032
INR 1.4 | 1032
activated partial thromboplastin time 43 s | 1032
D-dimer 1,211 ng/ml | 1032
fibrinogen 190 mg/dl | 1032
metabolic acidosis | 1032
lactic acid 12.6 mmol/l | 1032
intensive fluid replacement | 1032
positive inotropic support | 1032
erythrocyte suspension | 1032
thrombocyte suspension | 1032
left ventricular ejection fraction 64% | 1032
broad spectrum antibiotherapy | 1032
encephalopathy | 1032
generalized tonic-clonic convulsions | 1032
intubation | 1032
mechanical ventilation | 1032
cranial computed tomography | 1032
bleeding region 9 mm | 1032
peripheral edema | 1032
lactic acidosis | 1032
hemodiafiltration | 1032
thiamine treatment | 1032
thiamine deficiency | 1032
lactic acidosis regression | 1032
remission | 1512
BCR-ABL gene fusion negative | 1512
mechanic ventilation | 1512
extubation | 1512
percutaneous endoscopic gastrostomy | 1512
swallowing dysfunction | 1512
cognitive functions normal | 2592
mucositis regression | 2592
physiotherapy | 2592
spastic tetraparesis | 2592
discharge | 3024
imatinib 400 mg/m2/day | 3024
no transfusion | 3024
bone marrow examination | 3024
morphological remission | 3024
molecular remission | 3024
no matched donor | 3024
morphological remission | 6480
molecular remission | 6480