34 years old | 0
African | 0
female | 0
emergency room | 0
fever | -168
blisters | -24
rash | -24
HIV infection | -87600
Combivir | -87600
lamivudine | -87600
zidovudine | -87600
Kaletra | -87600
lopinavir | -87600
ritonavir | -87600
supportive care | -120
vitamins | -120
micronutrients | -120
pain relieving medications | -120
acetylsalicylic acid | -120
acetaminophen | -120
general practitioner consultation | -120
bacterial infection concern | -120
cefuroxime | -120
azithromycin | -120
fluconazole | -120
rash onset | -96
blisters worsening | -48
fever increase | -48
malaise | -48
conscious | 0
oriented | 0
normotensive | 0
blood pressure 120/65 | 0
sinus tachycardia | 0
heart rate 124/min | 0
dry lips | 0
dry tongue | 0
dehydration | 0
conjunctival injection | 0
no chest abnormalities | 0
no abdominal abnormalities | 0
blisters size 0.5-4 cm | 0
blisters coverage 45% | 0
TEN suspicion | 0
dermatologist consultation | 0
burn surgeon consultation | 0
ICU transfer | 0
central venous access | 0
fluid resuscitation | 0
lactated Ringer's solution | 0
standard monitoring | 0
central venous pressure measurement | 0
arterial pressure measurement | 0
antimicrobial therapy discontinuation | 0
CRP increase | 0
leucocytes normal | 0
serum protein elevated | 0
LDH elevated | 0
no pathological findings | 0
chest X-ray normal | 0
blood culture negative | 0
urine culture negative | 0
wound culture negative | 0
blisters disinfection | 0
Octenisept | 0
Acticoat application | 0
dry sterile gauzes | 0
vital stability | 0
intermittent high fever | 0
bacterial screenings negative | 0
fungal screenings negative | 0
unclear infection focus | 0
infectious disease consultation | 0
Avalox | 0
moxifloxacin | 0
Ecalta | 0
anidulafungin | 0
continued HIV therapy | 0
dengue virus DNA detected | 72
denied recent travel | 0
recent visit to Kenya | 72
antimicrobials stopped | 72
fever decrease | 120
wound recovery | 0
discharge | 432
no secondary deficits | 432
TEN diagnosis | 0
DF diagnosis | 72
SCORTEN score 2 | 0
Nikolsky's sign | 0
mucosal involvement | 0
ocular involvement | 0
thermoregulatory disturbance | 0
no lung failure | 0
no renal failure | 0
no liver failure | 0
no heart failure | 0
mortality risk 40% | 0
drug reaction | 0
cefuroxime reaction | 0
azithromycin reaction | 0
HIV positive | 0
dengue fever | 72
Aedes aegypti exposure | -72
DENV infection | 72
febrile returning traveler | 0
interdisciplinary approach | 0
no conflict of interest | 0
