10 years old | 0
male | 0
admitted to the hospital | 0
persistent fever | -504
cough | -504
weight loss | -504
sepsis | 0
cardiac tamponade | 0
respiratory distress | 0
dyspnoea | 0
polypnea | 0
heart rate 108 beats/min | 0
temperature 38.7°C | 0
hepatomegaly | 0
distended neck veins | 0
muffled heart sounds | 0
thiamphenicol and clavulanic acid and amoxicillin | -504
chest X-ray normal | -504
thoracoabdominal sonogram | 0
left liver lobe abscess | 0
chest and abdominal computer tomography scan | 0
bilateral pleuropneumopathy | 0
diaphragmatic collection | 0
hepatosplenomegaly | 0
minor ascites | 0
amoebic serology normal | 0
IV antibiotic | 0
amoxicillin and clavulanic acid | 0
gentamicin | 0
pericardial effusion | 0
amediastinal abscess | 0
right mediastinal drainage | 24
500ml of frank greenish pus | 24
ceftriaxone | 72
metronidazole | 72
gentamicin | 72
blood transfusion | 72
severe anaemia | 72
thoracotomy | 96
pericardiectomy | 96
2 litres of frank pus | 96
Staphylococcus aureus | 120
HIV serology positive | 120
ciprofloxacin | 120
gentamicin stopped | 120
temperature subsided | 216
hemodynamic parameters improved | 216
persistent purulent drainage | 216
corticotherapy | 312
drains removed | 312
persistent bilateral lower lobe infiltrate | 312
mild cardiomegaly | 312
thickened pericardium | 312
no pericardial effusion | 312
no valvular anomaly | 312
discharged home | 576
per os ciprofloxacin | 576
iron treatment | 576
steroids stopped | 576
antiretroviral drugs | 672
cotrimoxazole | 672
CD4 count 14 cells/ml | 672
mother on antiretroviral treatment | 672