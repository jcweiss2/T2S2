60 years old | 0
female | 0
hypertension | 0
chronic obstructive pulmonary disease (COPD) | 0
admitted to the hospital | 0
fever | -48
cough | -48
dyspnea | -48
tachypnea | 0
hypotension | 0
confusion | 0
oxygen through nasal cannula | 0
IV fluids | 0
IV azithromycin | 0
IV ceftriaxone | 0
chest x-ray (CXR) | 0
no consolidations or infiltrates | 0
hypotensive | -12
transferred to the intensive care unit | -12
IV piperacillin-tazobactam | -12
levofloxacin | -12
vasopressors | -12
hydrocortisone | -12
febrile | 72
no improvement | 72
hypertriglyceridemia | 72
thrombocytopenia | 72
leukopenia | 72
hyperferritinemia | 72
hypofibrinogenemia | 72
normal coagulation profile | 72
normal procalcitonin | 72
negative work-up for connective tissue diseases | 72
negative work-up for viral infections | 72
peripheral blood smear unremarkable | 72
family history of malignancies | 0
computerized tomography scan | 72
moderate splenomegaly | 72
elevated soluble cluster differentiation 25 (CD-25) | 72
bone marrow aspirate | 72
hemophagocytosis | 72
IV methylprednisolone | 72
improved markedly | 120
no longer in septic shock | 120
flow cytometry testing | 168
cytogenetics results | 168
no lymphomas or leukemias | 168
switched to HLH-94 protocol | 168
high dose of dexamethasone | 168
etoposide | 168
mean arterial pressure maintained | 216
no episodes of fever | 216
transferred to medical floor | 216
discharged | 216
dexamethasone | 216
etoposide | 216
follow up with Hematology–Oncology Outpatient Clinics | 216