55 years old | 0
male | 0
alcohol abuse | -672
shortness of breath | -48
cough | -48
fever | -48
chills | -48
confusion | -48
altered mental status | -48
unconscious | -12
intubated | 0
assist-control mechanical ventilation | 0
sinus tachycardia | 0
hypotension | 0
vasopressors | 0
right-sided decreased air entry | 0
diffuse crackles | 0
leukopenia | 0
white blood cells 0.8 × 10^9/L | 0
absolute neutrophil count 360 mm^3 | 0
hemoglobin 8.1 g/L | 0
platelets 109,000 | 0
creatinine 3.5 mg/dl | 0
potassium 4.5 meq/L | 0
right lower lobe consolidation | 0
right pleural effusion | 0
Streptococcus pneumoniae | 0
vancomycin | 0
piperacillin/tazobactam | 0
remarkable recovery | 72
discharged | 72
alcoholic leukopenic pneumococcal sepsis (ALPS) syndrome | 0