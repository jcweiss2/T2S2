22 years old | 0
    male | 0
    5-year history of smoking | -43800
    20 cigarettes per day | -43800
    exposed to live poultry | -48
    high fever | 0
    chills | 0
    prescription of ibuprofen | 0
    prescription of azithromycin | 0
    progressed complaints | -72
    emergency department visit | -72
    lymphopenia | 0
    thrombocytopenia | 0
    normal white blood cell count | 0
    normal PaO2/FiO2 | 0
    patchy shadows in right lung | 0
    consolidation in right lung | 0
    treated with meropenem | 0
    treated with moxifloxacin | 0
    throat swab obtained | 0
    oseltamivir administered | 0
    PaO2/FiO2 declined to 84 | 144
    elevated aspartate aminotransferase | 144
    elevated alanine aminotransferase | 144
    elevated lactate dehydrogenase | 144
    elevated creatine kinase | 144
    elevated myoglobin | 144
    septic shock | 144
    SOFA score increased from 2 to 10 | 144
    H5N6 virus identified | 144
    transferred to ICU | 144
    invasive mechanical ventilation | 144
    BALF galactomannan >5 g/mL | 144
    increased oseltamivir dosage | 144
    peramivir administered | 144
    amphotericin B administered | 144
    low-dose corticosteroid administered | 144
    mediastinal emphysema | 168
    subcutaneous emphysema | 168
    rapid progression of lung consolidation | 240
    VV ECMO initiated | 240
    condition deteriorated | 240
    high tracheal aspirate viral titer | 288
    sirolimus administered | 288
    decreased viral titers | 312
    H5N6 undetectable in throat swab | 384
    improved clinical condition | 384
    PaO2/FiO2 increased to 278 | 384
    SOFA score decreased to 3 | 384
    increased white blood cell count | 384
    decreased aspartate aminotransferase | 384
    decreased alanine aminotransferase | 384
    decreased lactate dehydrogenase | 384
    decreased creatine kinase | 384
    decreased myoglobin | 384
    ECMO stopped | 528
    endotracheal tube removed | 600
    sirolimus discontinued | 600
    NAIs discontinued | 600
    antibiotics discontinued | 600
    resolution of bilateral lung infiltrations | 672
    discharged | 1560
    good condition at 2-year follow-up | 17352
    bilateral interstitial changes in lungs | 17352
    normal ventilation | 17352
    slightly decreased diffusion efficiency | 17352

    