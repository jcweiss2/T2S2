35 years old | 0
    male | 0
    autosomal dominant polycystic kidney disease | 0
    underwent kidney transplantation | 0
    end-stage renal failure | 0
    original bilateral polycystic kidneys not removed | 0
    donor brain death caused by hypertensive intracerebral hemorrhage | 0
    donor no confirmed infection | 0
    immune induction therapy | 0
    methylprednisolone | 0
    basiliximab | 0
    rabbit anti-human thymocyte immunoglobulin (ATG) | 0
    delayed graft function | 0
    maintenance immunosuppressive regimen | 0
    tacrolimus | 0
    mycophenolate mofetil | 0
    prednisone | 0
    tacrolimus concentration maintained at 6–8 ng/mL | 0
    hemodialysis before renal transplantation | -672
    urine output more than 3000 mL per day | 0
    no dialysis after surgery | 0
    Corynebacterium detected in donor kidney preservation solution | 0
    no drug sensitivity test | 0
    no Corynebacterium-related infection observed | 0
    absence of infection symptoms | 0
    no pathogens cultured from blood, urine, surgical site samples | 0
    ceftazidime prophylactically administered | 0
    oral trimethoprim/sulfamethoxazole for PJP prophylaxis | 0
    discharged | 336
    serum creatinine level 160–170 µmol/L | 0
    low fever 37.9°C | -672
    light hematuria | -672
    mild frequent urination | -672
    urgent urination | -672
    painful urination | -672
    white blood cell count 17.46×10⁹/L | 0
    hemoglobin level 95 g/L | 0
    C-reactive protein level 231.06 mg/L | 0
    serum creatinine level 196.1 µmol/L | 0
    prothrombin time 15.40 s | 0
    blood pressure 87/64 mmHg | 0
    partial intracapsular hemorrhage in bilateral polycystic kidneys | 0
    septic shock | 0
    disseminated intravascular coagulation | 0
    severe infection | 0
    intracapsular hemorrhage with infection of cysts | 0
    supportive treatment | 0
    vital signs remained stable | 0
    immunosuppressive regimen tapered | 0
    mycophenolate withdrawn | 0
    tacrolimus replaced by cyclosporin | 0
    meropenem administered | 0
    Corynebacterium found in blood | 0
    Enterococcus faecium found in urine | 0
    Pseudomonas putida found in urine | 0
    linezolid additionally administered | 0
    ultrasound examination performed | 168
    no special findings | 168
    tacrolimus used again | 168
    cyclosporin used for 3 days | 168
    patient intolerance | 168
    troponin T increased | 0
    atrial natriuretic peptide levels increased | 0
    chest pain | 192
    dyspnea | 192
    unable to lie in supine position | 192
    sinus tachycardia | 192
    premature ventricular beats | 192
    acute anuria | 192
    serum creatinine increased to 346 µmol/L | 192
    multiple thromboses in right external iliac artery | 192
    largest thrombosis around anastomotic orifice of transplanted renal artery | 192
    transferred to intensive care unit | 192
    continuous renal replacement therapy | 192
    meropenem adjusted | 192
    vancomycin used | 192
    sudden persistent angina pectoris | 216
    chest tightness | 216
    no sweating | 216
    increase in myocardial enzymes | 216
    cardiac murmur in each valve | 216
    grade 3/6 diastolic murmur in apical region | 216
    echocardiography revealed medium echoic mass at posterior mitral valve tip | 216
    moderate-to-severe mitral regurgitation | 216
    mild-to-moderate tricuspid regurgitation | 216
    chest tightness | 240
    significant increase in myocardial enzymes | 240
    non-ST segment elevation myocardial infarction | 240
    fraxiparin administered | 240
    cough with bloody sputum | 264
    fraxiparin stopped | 264
    scheduled operation | 336
    allograft nephrectomy planned | 336
    mitral valve replacement | 336
    vegetative resection | 336
    cardiac arrest | 336
    ventricular fibrillation | 336
    emergency external chest compression | 336
    electric defibrillation | 336
    endotracheal intubation | 336
    vital signs stabilized | 336
    large polypoid vegetation found on posterior leaflet of mitral valve | 336
    allograft nephrectomy not performed | 336
    patient died | 360
    no pathogens cultured from mitral valve or vegetation tissue | 336
    large polypoid excrescences in pathological sections | 0
    Gram staining revealed valvular and leukocyte necrosis | 0
    colonies of bacteria | 0
    mNGS performed | 0
    C. striatum confirmed | 0
    C. striatum endocarditis | 0
    <|eot_id|>