50 years old | 0
male | 0
admitted to the emergency department | 0
high spiking fever | 0
disorientation | 0
antiphospholipid syndrome | -672
deep vein thrombosis | -672
ischemic stroke | -672
warfarin | -672
prosthetic tissue aortic valve replacement | -672
aortic stenosis | -672
brainstem hemorrhage | -216
nosocomial pneumonia | -216
severe renal failure | -216
hemodialysis | -216
permacath | -216
enoxaparin | -216
permacath removal | -24
temperature of 39°C | 0
blood pressure of 80/50 mmHg | 0
pulse of 128 beats per minute | 0
36 breaths per minute | 0
oxygen saturation of 88% | 0
leukocytosis of 20,000 per cubic millimeter | 0
hemoglobin concentration of 12 g/dL | 0
platelets count of 550,000 per cubic millimeter | 0
blood urea nitrogen and creatinine levels were slightly elevated | 0
microscopic hematuria | 0
vancomycin | 0
piperacillin-tazobactam | 0
amikacin | 0
vasopressors | 0
ICU | 0
MRSA bacteremia | 0
MRSA susceptible to vancomycin | 0
MRSA susceptible to daptomycin | 0
MRSA susceptible to rifampin | 0
MRSA susceptible to TMP/SMX | 0
permacath extracted | 0
transthoracic echocardiogram | 24
normal function of the prosthetic valve | 24
fever persisted | 48
blood cultures grew MRSA | 48
vancomycin and rifampin | 48
MRSA resistant to rifampin | 48
vancomycin plus piperacillin-tazobactam | 72
transesophageal echocardiogram | 96
thrombus in the SVC | 96
daptomycin and oxacillin | 120
MRSA non-susceptible to daptomycin | 120
MRSA resistant to vancomycin | 120
daptomycin dose increased | 144
intravenous TMP/SMX | 144
clearance of MRSA bacteremia | 168
cardiac arrest | 192
death | 192
septic thrombus formation | -672
SVC thrombosis | 96
anticoagulation | 0
thrombectomy | -672
thrombolysis | -672
balloon angioplasty | -672
stent insertion | -672
SVC syndrome | -672
pulmonary embolism | 192
linezolid | -672
ceftaroline | -672
quinupristin/dalfopristin | -672
telavancin | -672
trimethoprim/sulfamethoxazole | -672