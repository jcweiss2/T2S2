62 years old | 0
female | 0
congestive heart failure | 0
type 1 diabetes | 0
hypertension | 0
admitted to the hospital | 0
dyspnea | 0
encephalopathy | 0
intubated | 0
influenza A | 0
bacterial pneumonia | 0
acute respiratory failure | 0
acute respiratory distress syndrome | -48
septic shock | -48
broad-spectrum antibiotics | -48
vasopressors | -48
ejection fraction of 20% | -48
cardiogenic shock | -48
Impella device | -48
extracorporeal membranous oxygenation | -48
systemic heparin | -48
transferred to the cardiac intensive care unit | -48
continuous renal replacement therapy | -192
anasarca | -192
oliguria | -192
hematochezia | -240
hemoglobin level 6.4 g/dL | -240
pantoprazole drip | -240
intravenous fluid resuscitation | -240
transfused packed red blood cells | -240
esophagogastroduodenoscopy | -240
superficial punctate esophageal ulcers | -240
oozing blood | -240
clotted blood | -240
metoclopramide | -228
repeat esophagogastroduodenoscopy | -228
Hemospray | -228
hematochezia stopped | -228
Hb stabilized | -228
crusted vesicular lesions | -228
upper lip | -228
lateral aspect of her tongue | -228
herpes simplex virus | -228
IV acyclovir | -228
buccal ulceration | -228
HSV polymerase chain reaction | -228
HSV-1 antibody IgG | -228
HSV IgM immunoglobulin | -228
Helicobacter pylori stool antigen | -228
serologies | -228
hematochezia slowly stopped | -192
blood counts stabilized | -192
finished acyclovir | -168
repeat EGD | -168
normal esophageal mucosa | -168
Impella support weaned off | -240
vasopressors weaned off | -240