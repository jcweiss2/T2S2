72 years old | 0
male | 0
hypertension | 0
atrial fibrillation | 0
alcoholic liver cirrhosis | 0
metastatic urothelial carcinoma | 0
admitted to the hospital | 0
rash | -48
erythematous rash | -48
skin sloughing | -48
enfortumab vedotin | -168
acetaminophen | 0
acyclovir | 0
metoprolol | 0
gabapentin | 0
discontinued enfortumab vedotin | 0
started on topical steroid | 0
biopsy | 24
interface dermatitis | 24
full-thickness epidermal necrosis | 24
oliguria | 24
acute kidney injury | 24
acute tubular necrosis | 24
started on continuous renal replacement therapy | 24
rash progressed | 48
diagnosed with TEN | 48
discussed intravenous immunoglobulin | 48
discussed cyclosporine | 48
discussed etanercept | 48
started on empiric vancomycin/meropenem | 48
hypotension | 72
started on norepinephrine | 72
started on vasopressin | 72
hyperbilirubinemia | 96
increased international normalized ratio | 96
multiorgan failure | 120
septic shock | 120
end-of-life measures discussed | 120
died | 480