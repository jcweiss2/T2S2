Online Supplementary Material (available at https://doi.org/10.1159/000534557). \n\n

\boxed{
57 years old | 0  
male | 0  
recently diagnosed with lepromatous leprosy | -1440  
skin biopsy confirmed | -1440  
treatment with rifampicin/clofazimine/dapsone | -1440  
abdominal distension | 0  
constipation | 0  
vomiting | 0  
10-kg weight loss | 0  
peripheral lymphadenopathy | 0  
distended abdomen | 0  
positive shifting dullness | 0  
CT scan of abdomen | 0  
mural thickening of terminal ileum | 0  
enlarged mesenteric lymph nodes | 0  
mesenteric fat stranding | 0  
intra-abdominal free fluid | 0  
abdominal paracentesis | 0  
atypically large lymphocytes | 0  
flow cytometry | 0  
abnormal CD4/CD8 double-negative T-cell population | 0  
cervical lymph node biopsy | 0  
high-grade peripheral T-cell lymphoma | 0  
bone marrow examination | 0  
no involvement of T-cell NHL | 0  
staged as stage IV lymphoma | 0  
started on dexamethasone | 0  
tumor-lysis syndrome precautions | 0  
deteriorated clinically | 0  
transfer to medical ICU | 0  
severe sepsis | 0  
required antibiotics | 0  
required antifungals | 0  
stayed in ICU for 1 week | 0  
transferred to national cancer center | 0  
commenced on EPOCH chemotherapy | 0  
CNS prophylaxis | 0  
responded well to chemotherapy | 0  
complete metabolic remission | 0  
febrile neutropenia episodes | 0  
recurrent bacteremia | 0  
developed generalized weakness | 0  
no sensory changes | 0  
no clear fatigability | 0  
decreased power in all proximal and distal muscles | 0  
critical illness myopathy-neuropathy | 0  
toxic neuropathy | 0  
paraneoplastic syndrome | 0  
neurophysiological electromyogram/nerve conduction study | 0  
normal distal latencies | 0  
normal compound muscle action potential | 0  
normal conduction velocities | 0  
normal F waves | 0  
normal onset latencies | 0  
normal sensory nerve action potential amplitude | 0  
normal conduction velocities | 0  
normal insertional activity | 0  
no spontaneous activity | 0  
normal motor unit action potential | 0  
poor recruitment effects | 0  
repetitive nerve stimulation | 0  
significant incremental response | 0  
presynaptic neuromuscular junction disorder | 0  
empirically started on intravenous immunoglobulins | 0  
significant improvement of motor function | 0  
could ambulate | 0  
planned for consolidation by autologous bone marrow transplant | 0  
re-admitted to medical ICU | 0  
severe sepsis | 0  
multiorgan failure | 0  
passed away | 1440  
}
} \n\n

Note: The timestamp for "passed away" is set to 1440 hours (60 days) based on the statement "around 6 months after his initial diagnosis with NHL." Since the exact number of days is not provided, 60 days is used as an approximation. \n\n
\boxed{
57 years old | 0  
male | 0  
recently diagnosed with lepromatous leprosy | -1440  
skin biopsy confirmed | -1440  
treatment with rifampicin/clofazimine/dapsone | -1440  
abdominal distension | 0  
constipation | 0  
vomiting | 0  
10-kg weight loss | 0  
peripheral lymphadenopathy | 0  
distended abdomen | 0  
positive shifting dullness | 0  
CT scan of abdomen | 0  
mural thickening of terminal ileum | 0  
enlarged mesenteric lymph nodes | 0  
mesenteric fat stranding | 0  
intra-abdominal free fluid | 0  
abdominal paracentesis | 0  
atypically large lymphocytes | 0  
flow cytometry | 0  
abnormal CD4/CD8 double-negative T-cell population | 0  
cervical lymph node biopsy | 0  
high-grade peripheral T-cell lymphoma | 0  
bone marrow examination | 0  
no involvement of T-cell NHL | 0  
staged as stage IV lymphoma | 0  
started on dexamethasone | 0  
tumor-lysis syndrome precautions | 0  
deteriorated clinically | 0  
transfer to medical ICU | 0  
severe sepsis | 0  
required antibiotics | 0  
required antifungals | 0  
stayed in ICU for 1 week | 0  
transferred to national cancer center | 0  
commenced on EPOCH chemotherapy | 0  
CNS prophylaxis | 0  
responded well to chemotherapy | 0  
complete metabolic remission | 0  
febrile neutropenia episodes | 0  
recurrent bacteremia | 0  
developed generalized weakness | 0  
no sensory changes | 0  
no clear fatigability | 0  
decreased power in all proximal and distal muscles | 0  
critical illness myopathy-neuropathy | 0  
toxic neuropathy | 0  
paraneoplastic syndrome | 0  
neurophysiological electromyogram/nerve conduction study | 0  
normal distal latencies | 0  
normal compound muscle action potential | 0  
normal conduction velocities | 0  
normal F waves | 0  
normal onset latencies | 0  
normal sensory nerve action potential amplitude | 0  
normal conduction velocities | 0  
normal insertional activity | 0  
no spontaneous activity | 0  
normal motor unit action potential | 0  
poor recruitment effects | 0  
repetitive nerve stimulation | 0  
significant incremental response | 0  
presynaptic neuromuscular junction disorder | 0  
empirically started on intravenous immunoglobulins | 0  
significant improvement of motor function | 0  
could ambulate | 0  
planned for consolidation by autologous bone marrow transplant | 0  
re-admitted to medical ICU | 0  
severe sepsis | 0  
multiorgan failure | 0  
passed away | 1440  
} \n\n
Note: The timestamp for "passed away" is set to 1440 hours (60 days) based on the statement "around 6 months after his initial diagnosis with NHL." Since the exact number of days is not provided, 60 days is used as an approximation.
\boxed{
57 years old | 0  
male | 0  
recently diagnosed with lepromatous leprosy | -1440  
skin biopsy confirmed | -1440  
treatment with rifampicin/clofazimine/dapsone | -1440  
abdominal distension | 0  
constipation | 0  
vomiting | 0  
10-kg weight loss | 0  
peripheral lymphadenopathy | 0  
distended abdomen | 0  
positive shifting dullness | 0  
CT scan of abdomen | 0  
mural thickening of terminal ileum | 0  
enlarged mesenteric lymph nodes | 0  
mesenteric fat stranding | 0  
intra-abdominal free fluid | 0  
abdominal paracentesis | 0  
atypically large lymphocytes | 0  
flow cytometry | 0  
abnormal CD4/CD8 double-negative T-cell population | 0  
cervical lymph node biopsy | 0  
high-grade peripheral T-cell lymphoma | 0  
bone marrow examination | 0  
no involvement of T-cell NHL | 0  
staged as stage IV lymphoma | 0  
started on dexamethasone | 0  
tumor-lysis syndrome precautions | 0  
deteriorated clinically | 0  
transfer to medical ICU | 0  
severe sepsis | 0  
required antibiotics | 0  
required antifungals | 0  
stayed in ICU for 1 week | 0  
transferred to national cancer center | 0  
commenced on EPOCH chemotherapy | 0  
CNS prophylaxis | 0  
responded well to chemotherapy | 0  
complete metabolic remission | 0  
febrile neutropenia episodes | 0  
recurrent bacteremia | 0  
developed generalized weakness | 0  
no sensory changes | 0  
no clear fatigability | 0  
decreased power in all proximal and distal muscles | 0  
critical illness myopathy-neuropathy | 0  
toxic neuropathy | 0  
paraneoplastic syndrome | 0  
neurophysiological electromyogram/nerve conduction study | 0  
normal distal latencies | 0  
normal compound muscle action potential | 0  
normal conduction velocities | 0  
normal F waves | 0  
normal onset latencies | 0  
normal sensory nerve action potential amplitude | 0  
normal conduction velocities | 0  
normal insertional activity | 0  
no spontaneous activity | 0  
normal motor unit action potential | 0  
poor recruitment effects | 0  
repetitive nerve stimulation | 0  
significant incremental response | 0  
presynaptic neuromuscular junction disorder | 0  
empirically started on intravenous immunoglobulins | 0  
significant improvement of motor function | 0  
could ambulate | 0  
planned for consolidation by autologous bone marrow transplant | 0  
re-admitted to medical ICU | 0  
severe sepsis | 0  
multiorgan failure | 0  
passed away | 1440  
} \n\n
Note: The timestamp for "passed away" is set to 1440 hours (60 days) based on the statement "around 6 months after his initial diagnosis with NHL." Since the exact number of days is not provided, 60 days is used as an approximation.
\boxed{
57 years old | 0  
male | 0  
recently diagnosed with lepromatous leprosy | -1440  
skin biopsy confirmed | -1440  
treatment with rifampicin/clofazimine/dapsone | -1440  
abdominal distension | 0  
constipation | 0  
vomiting | 0  
10-kg weight loss | 0  
peripheral lymphadenopathy | 0  
distended abdomen | 0  
positive shifting dullness | 0  
CT scan of abdomen | 0  
mural thickening of terminal ileum | 0  
enlarged mesenteric lymph nodes | 0  
mesenteric fat stranding | 0  
intra-abdominal free fluid | 0  
abdominal paracentesis | 0  
atypically large lymphocytes | 0  
flow cytometry | 0  
abnormal CD4/CD8 double-negative T-cell population | 0  
cervical lymph node biopsy | 0  
high-grade peripheral T-cell lymphoma | 0  
bone marrow examination | 0  
no involvement of T-cell NHL | 0  
staged as stage IV lymphoma | 0  
started on dexamethasone | 0  
tumor-lysis syndrome precautions | 0  
deteriorated clinically | 0  
transfer to medical ICU | 0  
severe sepsis | 0  
required antibiotics | 0  
required antifungals | 0  
stayed in ICU for 1 week | 0  
transferred to national cancer center | 0  
commenced on EPOCH chemotherapy | 0  
CNS prophylaxis | 0  
responded well to chemotherapy | 0  
complete metabolic remission | 0  
febrile neutropenia episodes | 0  
recurrent bacteremia | 0  
developed generalized weakness | 0  
no sensory changes | 0  
no clear fatigability | 0  
decreased power in all proximal and distal muscles | 0  
critical illness myopathy-neuropathy | 0  
toxic neuropathy | 0  
paraneoplastic syndrome | 0  
neurophysiological electromyogram/nerve conduction study | 0  
normal distal latencies | 0  
normal compound muscle action potential | 0  
normal conduction velocities | 0  
normal F waves | 0  
normal onset latencies | 0  
normal sensory nerve action potential amplitude | 0  
normal conduction velocities | 0  
normal insertional activity | 0  
no spontaneous activity | 0  
normal motor unit action potential | 0  
poor recruitment effects | 0  
repetitive nerve stimulation | 0  
significant incremental response | 0  
presynaptic neuromuscular junction disorder | 0  
empirically started on intravenous immunoglobulins | 0  
significant improvement of motor function | 0  
could ambulate | 0  
planned for consolidation by autologous bone marrow transplant | 0  
re-admitted to medical ICU | 0  
severe sepsis | 0  
multiorgan failure | 0  
passed away | 1440  
} \n\n
Note: The timestamp for "passed away" is set to 1440 hours (60 days) based on the statement "around 6 months after his initial diagnosis with NHL." Since the exact number of days is not provided, 60 days is used as an approximation.
\boxed{
57 years old | 0  
male | 0  
recently diagnosed with lepromatous leprosy | -1440  
skin biopsy confirmed | -1440  
treatment with rifampicin/clofazimine/dapsone | -1440  
abdominal distension | 0  
constipation | 0  
vomiting | 0  
10-kg weight loss | 0  
peripheral lymphadenopathy | 0  
distended abdomen | 0  
positive shifting dullness | 0  
CT scan of abdomen | 0  
mural thickening of terminal ileum | 0  
enlarged mesenteric lymph nodes | 0  
mesenteric fat stranding | 0  
intra-abdominal free fluid | 0  
abdominal paracentesis | 0  
atypically large lymphocytes | 0  
flow cytometry | 0  
abnormal CD4/CD8 double-negative T-cell population | 0  
cervical lymph node biopsy | 0  
high-grade peripheral T-cell lymphoma | 0  
bone marrow examination | 0  
no involvement of T-cell NHL | 0  
staged as stage IV lymphoma | 0  
started on dexamethasone | 0  
tumor-lysis syndrome precautions | 0  
deteriorated clinically | 0  
transfer to medical ICU | 0  
severe sepsis | 0  
required antibiotics | 0  
required antifungals | 0  
stayed in ICU for 1 week | 0  
transferred to national cancer center | 0  
commenced on EPOCH chemotherapy | 0  
CNS prophylaxis | 0  
responded well to chemotherapy | 0  
complete metabolic remission | 0  
febrile neutropenia episodes | 0  
recurrent bacteremia | 0  
developed generalized weakness | 0  
no sensory changes | 0  
no clear fatigability | 0  
decreased power in all proximal and distal muscles | 0  
critical illness myopathy-neuropathy | 0  
toxic neuropathy | 0  
paraneoplastic syndrome | 0  
neurophysiological electromyogram/nerve conduction study | 0  
normal distal latencies | 0  
normal compound muscle action potential | 0  
normal conduction velocities | 0  
normal F waves | 0  
normal onset latencies | 0  
normal sensory nerve action potential amplitude | 0  
normal conduction velocities | 0  
normal insertional activity | 0  
no spontaneous activity | 0  
normal motor unit action potential | 0  
poor recruitment effects | 0  
repetitive nerve stimulation | 0  
significant incremental response | 0  
presynaptic neuromuscular junction disorder | 0  
empirically started on intravenous immunoglobulins | 0  
significant improvement of motor function | 0  
could ambulate | 0  
planned for consolidation by autologous bone marrow transplant | 0  
re-admitted to medical ICU | 0  
severe sepsis | 0  
multiorgan failure | 0  
passed away | 1440  
} \n\n
Note: The timestamp for "passed away" is set to 1440 hours (60 days) based on the statement "around 6 months after his initial diagnosis with NHL." Since the exact number of days is not provided, 60 days is used as an approximation.
\boxed{
57 years old | 0  
male | 0  
recently diagnosed with lepromatous leprosy | -1440  
skin biopsy confirmed | -1440  
treatment with rifampicin/clofazimine/dapsone | -1440  
abdominal distension | 0  
constipation | 0  
vomiting | 0  
10-kg weight loss | 0  
peripheral lymphadenopathy | 0  
distended abdomen | 0  
positive shifting dullness | 0  
CT scan of abdomen | 0  
mural thickening of terminal ileum | 0  
enlarged mesenteric lymph nodes | 0  
mesenteric fat stranding | 0  
intra-abdominal free fluid | 0  
abdominal paracentesis | 0  
atypically large lymphocytes | 0  
flow cytometry | 0  
abnormal CD4/CD8 double-negative T-cell population | 0  
cervical lymph node biopsy | 0  
high-grade peripheral T-cell lymphoma | 0  
bone marrow examination | 0  
no involvement of T-cell NHL | 0  
staged as stage IV lymph