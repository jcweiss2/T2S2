46 years old| 0\
    male | 0\
    arterial hypertension | -672\
    obesity | -672\
    admitted | 0\
    fever | 0\
    hypotension | 0\
    marked asthenia | 0\
    cardiological examination | -672\
    electrocardiogram (ECG) | -672\
    transthoracic echocardiography (TTE) | -672\
    hypertension follow-up | -672\
    normal findings | -672\
    COVID-19 infection | -336\
    rhinitis | -336\
    mild cough | -336\
    alert | 0\
    oriented | 0\
    cooperative | 0\
    asthenic | 0\
    blood pressure (BP) 85/55 mmHg | 0\
    heart rate (HR) 120 bpm | 0\
    arterial oxygen saturation 85% | 0\
    fever 38.3°C | 0\
    femoral central venous catheter (CVC) placement | 0\
    ECG sinus tachycardia 122 bpm | 0\
    diffuse low voltages | 0\
    absence of significant repolarization abnormalities | 0\
    neutrophilic leukocytosis | 0\
    white blood cell count 26800 x 1000/mm³ | 0\
    C-reactive protein (CRP) 17.4 mg/dl | 0\
    Procalcitonin 11.7 ng/ml | 0\
    high sensitivity Troponin (hs-Tn) 23000 ng/L | 0\
    brain natriuretic peptide (BNP) 6890 pg/ml | 0\
    creatinine 1.8 mg/dl | 0\
    transaminases elevation | 0\
    total bilirubin elevation | 0\
    RT-PCR nasopharyngeal swab negative | 0\
    COVID-19 IgM high levels | 0\
    TTE normal LV cavitary dimensions | 0\
    indexed end-diastolic volume (EDVi) 41 ml/m² | 0\
    diffuse LV parietal thickening 15-16 mm | 0\
    increased myocardial echogenicity | 0\
    severely reduced LV global systolic function | 0\
    ejection fraction (EF) 26% | 0\
    dP/dT ratio 672 mmHg/sec | 0\
    indexed stroke volume (SVi) 11 ml/m² | 0\
    cardiac index (CI) 1.3 l/min/m² | 0\
    low output | 0\
    grade II LV diastolic dysfunction | 0\
    normal RV cavitary dimensions | 0\
    reduced RV global systolic function | 0\
    RV basal EDD 37 mm | 0\
    RV mid EDD 28 mm | 0\
    TAPSE 14 mm | 0\
    tricuspid S-wave velocity 7.3 cm/sec | 0\
    IVC dilated 26 mm | 0\
    inspiratory collapse <50% | 0\
    RVSP 41 mmHg | 0\
    absence of hemodynamically significant valvulopathy | 0\
    slight pericardial effusion | 0\
    thoracic CT perivascular aortic and pulmonary adipose tissue imbibition | 0\
    abdominal ultrasonography no significant findings | 0\
    blood cultures initiated | 0\
    broad-spectrum antibiotic therapy | 0\
    INN-daptomycin | 0\
    piperacillin/tazobactam | 0\
    crystalloid hydration | 0\
    nasal cannula oxygen 4 l/min | 0\
    norepinephrine 0.6 mcg/kg/min | 0\
    poor hemodynamic response | 0\
    norepinephrine increased to 0.9 mcg/kg/min | 0\
    BP 90-95/60 mmHg | 0\
    oliguria | 0\
    levosimendan initiated | 0\
    levosimendan 0.1 mcg/kg/min | 0\
    BP 100/60 mmHg at 12 hours | 12\
    HR 110 bpm at 12 hours | 12\
    BP 125/70 mmHg at 24 hours | 24\
    HR 95 bpm at 24 hours | 24\
    diuresis 1800 ml | 24\
    TTE control at 12 hours | 12\
    TTE control at 24 hours | 24\
    LV EF 66% at 24 hours | 24\
    dP/dT ratio 1275 mmHg/sec at 24 hours | 24\
    TAPSE 23 mm at 24 hours | 24\
    tricuspid S-wave velocity 11.2 cm/sec at 24 hours | 24\
    SVi 27 ml/m² at 24 hours | 24\
    CI 2.5 l/min/m² at 24 hours | 24\
    LV diastolic function normal at 24 hours | 24\
    IVC diameter 18 mm at 24 hours | 24\
    IVC complete collapse at 24 hours | 24\
    RVSP 28 mmHg at 24 hours | 24\
    blood culture results negative | 0\
    CVC removed | 24\
    CVC tip culture negative | 24\
    cardiac magnetic resonance imaging (CMR) | 24\
    SSFp-CINE sequences normal LV and RV volumes | 24\
    mild hypokinesia of LV lateral and inferolateral walls | 24\
    TIR/T2w increased signal intensity | 24\
    myocardial edema | 24\
    subendocardial localization | 24\
    EGE enhancement | 24\
    LGE enhancement | 24\
    RV free wall edema | 24\
    pericardium edema | 24\
    CMR compatible with immune-mediated myocarditis | 24\
    endomyocardial biopsy | 48\
    lymphocytic myocarditis | 48\
    coronary arteriography normal | 48\
    discharge after 21 days | 504\
    TTE at 1 month post-discharge | 720\
    TTE at 3 months post-discharge | 2160\
    normal hemodynamic compensation | 504\
    normal laboratory findings | 504\
    normal ECG findings | 504\
    normal echocardiographic findings | 504\
    negative blood cultures | 0\
    negative CVC tip culture | 24\
    no substantial inflammation index changes | 24\
    no LV/RV volume changes | 24\
    persistent myocardial inflammation signs | 24\
    absence of ischemic repolarization changes | 0\
    no new Q waves | 0\
    gradual ECG normalization | 24\