58 years old | 0
male | 0
pancreatogenic diabetes | 0
cholecystectomy | 0
bright red blood stool | -48
abdominal pain | -48
difficulty breathing | -48
dehydrated | 0
tachycardic | 0
hypotensive | 0
confused | 0
severe anemia | 0
lactate 5 mmol/L | 0
bicarbonate 12 meq/L | 0
creatinine level 3.5 mg/dl | 0
elevated liver chemistries | 0
normal coagulation profile | 0
admitted to ICU | 0
vigorous volume resuscitation | 0
transfused 4 units of blood | 0
vasopressors | 0
colonoscopy inconclusive | 0
enhanced abdominal CT | 0
left colic artery aneurysm | 0
angiography | 0
transcatheter arterial embolization | 0
bleeding controlled | 0
improved | 0
vasopressors phased out | 0
discharged | 0
high fever | 672
acute abdominal pain (upper left abdomen) | 672
diffuse abdominal tenderness | 672
leukocytosis | 672
neutrophilia | 672
elevated C-reactive protein | 672
increased serum procalcitonin | 672
contrast-enhanced abdominal CT | 672
enlarged spleen | 672
hypodense low-density lesion with gas | 672
free liquid in abdomen | 672
surgery | 672
laparotomy | 672
purulent fluid in abdomen | 672
splenic necrosis | 672
purulent discharge | 672
peritoneal lavage | 672
splenectomy | 672
drain placed | 672
readmitted to ICU | 672
Escherichia coli identified | 672
carbapenems treatment | 672
extensive necrosis of splenic tissue | 672
spleen abscess diagnosis | 672
postoperative recovery | 672
discharged after full diet | 672
drain removed | 672
