41 years old | 0
    female | 0
    admitted to the hospital | 0
    untreated hypertension | -336
    morbid obesity | -336
    chronic back pain | -336
    intravenous drug use | -336
    worsening low back pain | -336
    diffuse abdominal pain | -336
    lower extremity weakness | -336
    anorexia | -336
    fever | -336
    chills | -336
    shortness of breath | -336
    dizziness | -336
    constipation | -336
    recent use of acetaminophen | -336
    recent use of gabapentin | -336
    recent use of hydrocodone | -336
    recent use of methamphetamines | -336
    recent use of marijuana | -336
    blood pressure of 79/53 mmHg | 0
    heart rate of 149 bpm | 0
    lactic acid of 4.2 mg dl−1 | 0
    white blood cell count 37,500 u l−1 | 0
    erythrocyte sedimentation rate 75 mm h−1 | 0
    urine toxicology positive for cannabis | 0
    urine toxicology positive for amphetamines | 0
    midline tenderness of the lumbar spine | 0
    3/5 strength in bilateral lower extremities | 0
    bilateral shoulder warmth | 0
    bilateral shoulder erythema | 0
    bilateral shoulder tenderness | 0
    limited range of motion in shoulders | 0
    multiple needle puncture sites on antecubital fossas | 0
    unclear if needle sites from IVDU or medical procedures | 0
    smaller puncture wounds between toes of right foot | 0
    blood cultures collected | 0
    started on vancomycin | 0
    started on metronidazole | 0
    started on aztreonam | 0
    started on IV fluids | 0
    initial blood cultures grew MRSA | 0
    vancomycin MIC 1 mg l−1 | 0
    rifampin MIC ≤1 mg l−1 | 0
    levofloxacin MIC ≤1 mg l−1 | 0
    clindamycin MIC ≤0.5 mg l−1 | 0
    daptomycin MIC ≤0.5 mg l−1 | 0
    linezolid MIC 2 mg l−1 | 0
    bilateral shoulder plain radiographs showed no abnormalities | 0
    arthrocentesis of AC joints | 0
    WBC 93,137 u l–1 in one shoulder | 0
    WBC 32,043 u l–1 in other shoulder | 0
    aspirates cultured and grew MRSA | 0
    taken for emergent surgical debridement of shoulders | 0
    intubated | 0
    MRI lumbar spine showed L3–L5 osteomyelitis | 0
    facet septic arthritis | 0
    dorsal paraspinous myositis | 0
    L2–L5 epidural abscess | 0
    bilateral psoas myositis | 0
    bilateral psoas abscesses | 0
    MRI bilateral shoulders after debridement showed septic arthritis of AC joints | 0
    right distal trapezius abscess | 0
    left supraclavicular abscess | 0
    MRI brain showed no acute intracranial processes | 0
    transthoracic echocardiogram negative for valvular vegetations | 0
    cardiology deferred transoesophageal echocardiogram | 0
    repeat surgical debridement of shoulders | 24
    neurosurgery evaluation for epidural abscess debridement | 24
    recommendation for medical management | 24
    leukocytosis continued to rise | 24
    leukocytosis peaked at 52,100 u l–1 | 24
    trough levels of vancomycin monitored | 24
    repeat blood cultures positive for MRSA | 24
    antibiotics escalated to daptomycin | 240
    antibiotics escalated to ceftaroline | 240
    blood cultures became negative | 336
    rifampin added | 336
    critical care required until extubation | 336
    repeat MRI lumbar spine showed worsening epidural abscess | 432
    neurosurgery surgical drainage with drain placement | 432
    intravenous antimicrobials given for 14 days after negative cultures | 336
    intraoperative wound cultures positive for MRSA | 432
    intraoperative wound cultures positive for Proteus mirabilis | 432
    patient improved clinically | 672
    all drains removed | 672
    discharged | 672
    prescribed oral levofloxacin | 672
    prescribed oral rifampin | 672
    lost to follow-up after discharge | 672
    