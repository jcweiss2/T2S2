72 years old | 0
female | 0
admitted to the hospital | 0
primary biliary cholangitis | 0
general fatigue | 0
dyspnea on effort | 0
lumbar vertebral compression fracture | -8760
osteoporosis | -8760
heart failure | -8760
tachycardia-induced cardiomyopathy | -8760
persistent atrial fibrillation | -8760
paroxysmal atrial flutter | -8760
sinus bradycardia | -8760
radiofrequency catheter ablation | -8760
bisoprolol fumarate | -8760
enalapril maleate | -8760
rivaroxaban | -8760
ursodeoxycholic acid | -8760
Celestamine | -10980
sarcopenia | 0
blood pressure 90/42 mmHg | 0
regular pulse rate 60 beats/min | 0
normocytic anemia | 0
elevated serum brain natriuretic peptide | 0
elevated serum anti-mitochondrial antibody M2 | 0
mild generalized hypokinesis of the left ventricle | 0
bilateral atrial dilatation | 0
intact coronary arteries | 0
cardiogenic shock | 24
pericardiocentesis | 24
surgical closure | 24
percutaneous cardiopulmonary support | 24
dobutamine | 24
intubated | 24
discontinued medications | 24
biventricular Takotsubo cardiomyopathy | 48
progressive reduction in blood pressure | 72
progressive reduction in daily urine output | 72
systemic vascular resistance reduction | 72
low serum glucose | 72
suspected acute adrenal insufficiency | 72
hydrocortisone | 72
hemodynamic stabilization | 96
normalization of systemic vascular resistance | 96
elevated serum adrenocorticotropic hormone | 96
elevated serum cortisol | 96
tapered intravenous hydrocortisone | 168
oral hydrocortisone | 168
discharged | 168