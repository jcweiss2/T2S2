57 years old|0
    male|0
    kidney transplantation|-5040
    end-stage renal disease|-5040
    chronic hemodialysis treatment|-5040
    family history of proteinuria|-5040
    hypertension|-5040
    hypercholesterolemia|-5040
    asthma bronchiale|-5040
    protocol biopsy|-5040
    borderline acute rejection|-5040
    corticosteroids not withdrawn|-5040
    pneumocystis jirovecii prophylaxis|-5040
    trimethoprim-sulfamethoxazole stopped|-5040
    mycophenolate mofetil|-5040
    tacrolimus|-5040
    methylprednisolone|-5040
    cough|0
    hemoptysis|0
    right-sided pleuritic chest pain|0
    dyspnea on exertion|0
    general malaise|0
    denies direct exposure to livestock|0
    afebrile|0
    total leukocyte count 9.11 × 10⁹/L|0
    hemoglobin 10.6 g/dL|0
    elevated CRP 18.5 mg/L|0
    elevated LDH 378 U/L|0
    renal allograft function deteriorated|0
    glomerular filtration rate 21 mL/min|0
    transaminases normal|0
    bilirubin concentrations normal|0
    electrolyte panel normal|0
    chest radiographs|0
    CT scan|0
    roundish lung lesion 32 × 32 × 32 mm|0
    air bronchograms|0
    infracarinal lymphadenopathy|0
    bronchoscopy|0
    bronchoalveolar lavage|0
    empiric amoxicillin-clavulanate|0
    favorable clinical evolution|-5040
    no resolution of symptoms|0
    neutrophilic cellular pattern|0
    aerobic cultures negative|0
    anaerobic cultures negative|0
    mycobacterial cultures negative|0
    yeast cultures negative|0
    fungal cultures negative|0
    antigen tests negative|0
    immunofluorescent assay negative|0
    galactomannan test positive|0
    probable invasive aspergillosis|0
    peripheral biopsies|0
    voriconazole|0
    mycophenolate mofetil dose reduced|0
    tacrolimus dose reduced|0
    low blood pressure 95/40 mmHg|168
    sudden dizziness|168
    nausea|168
    atypical chest pain|168
    afebrile|168
    renal allograft function worsened|168
    CRP elevated 35.4 mg/L|168
    blood cultures|168
    chest radiographs unchanged|168
    abdominal ultrasound normal|168
    ST segment depression|168
    troponin I elevated 2.88 μg/L|168
    non-ST elevation myocardial infarction suspected|168
    low molecular weight heparin|168
    transferred to cardiac intensive care unit|168
    blood cultures positive for R. equi|168
    BAL cultures negative|168
    meropenem|168
    vancomycin|168
    mycophenolate mofetil stopped|168
    tacrolimus trough levels reduced|168
    voriconazole stopped|168
    clinical condition deteriorated|168
    high fever|168
    chills|168
    CRP rose to 252 mg/L|168
    crepitations over both lungs|168
    CT scan increased lung mass|168
    lymphadenopathy|168
    bilateral patchy pulmonary opacities|168
    blood cultures positive R. equi|168
    transferred to university hospital|168
    third bronchoscopy|168
    BAL|168
    levofloxacin added|168
    progressive hypoxic respiratory failure|168
    transferred to intensive care unit|168
    CRP 345 mg/L|168
    LDH 542 U/L|168
    HIV serology negative|168
    cytomegalovirus negative|168
    Epstein-Barr virus negative|168
    CT scan bilateral diffuse ground glass opacity|168
    trimethoprim-sulfamethoxazole added|168
    lung nodule smaller|168
    P. jirovecii PCR positive|168
    methylprednisolone added|168
    BAL fluid cytology negative|168
    levofloxacin withdrawn|168
    blood cultures cleared|168
    vital signs stable|168
    oxygen supply tapered|168
    hyperkalemia|168
    primaquine|168
    clindamycin|168
    meropenem continued|168
    vancomycin continued|168
    clinical improvement|168
    radiological improvement|168
    in vitro susceptibility testing|168
    oral moxifloxacin|672
    rifampicin|672
    chest CT persistence of lung lesion|672
    ground glass opacity diminished|672
    trimethoprim-sulfamethoxazole continued|672
    renal function restored|672
    CRP 9.9 mg/L|672
    discharged home|672
    mild exertional dyspnea persisted|672
    CT scans gradual diminution|672
    left lower lobe cavitation|672
    volume decreased|672
    moxifloxacin discontinued|2232
    rifampicin discontinued|2232
    outpatient follow-up|2232
    no recurrent infection|2232
    radiological resolution|2232
    <|eot_id|>
    