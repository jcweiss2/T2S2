42 years old | 0
female | 0
admitted to the hospital | 0
fever | -168
abdominal pain | -168
discomfort during intercourse | -168
abnormal area in the cervix | 0
abnormal cells | 0
cervical intraepithelial neoplasia (CIN) grade 3 | 0
squamous cell carcinoma | 0
chemotherapy | 0
radiotherapy | 0
discharged home | 168
diabetes mellitus | 8760
abdominal distension | 8760
appetite loss | 8760
hypoalbuminemia | 8760
intestinal sub occlusion | 8760
bowel resection | 8760
jejunostomy | 8760
parenteral nutrition | 8760
antibiotic therapy | 8760
adhesions between bowel loops | 9360
stenosis | 9360
mucous fistula | 9360
corrective enterectomy | 9360
intestinal evisceration | 9360
aponeurotic dehiscence | 9360
surgical wound infection | 9360
Pseudomonas aeruginosa | 9360
Citrobacter sp. | 9360
Acinetobacter sp. | 9360
sepsis | 9360
vancomycin | 9360
imipenem | 9360
metronidazole | 9360
fever episodes | 10920
severe abdominal pain | 10920
weakness | 10920
respiratory distress | 10920
elevated urea | 10920
elevated creatinine | 10920
leukopenia | 10920
low hemoglobin | 10920
low platelets | 10920
blood cultures | 10920
Cryptococcus laurentii | 10920
antifungal treatment | 10920
fluconazole | 10920
central venous catheter removal | 11280
discharged home | 11520