71 years old | 0
woman | 0
admitted | 0
left flank pain | 0
oliguria | 0
hypotension | 0
pyuria | 0
severe sepsis | 0
acute pyelonephritis | 0
abdominal computed tomography intravenous pyelogram | 0
normal-sized kidneys | 0
poorly determined differentiation between cortex and medulla | 0
amorphic low attenuation lesion | 0
incompletely malrotated kidneys | 0
anteriorly facing hila | 0
renal vessels and ureter located laterally | 0
renal ectopia | 0
mild dilation at proximal ureter of left kidney | 0
three-dimensional computed tomography reconstruction image | 0
anteriorly rotated kidneys | 0
piperacillin-tazobactam | 0
E. coli infection in bloodstream | 0
switched to cefotaxime | 0
improved hemodynamic state | 72
released from intensive care unit | 72
recurrent urinary tract infections | -720
ureteral deformation | -720
renal malrotation | -720
septic shock | 0
dilated left ureter | 0
mild obstruction | 0
ureteropyelic junction obstruction | -720
urolithiasis | -720 
discharged | 72