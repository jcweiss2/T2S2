64 years old | 0
female | 0
admitted to the hospital | 0
found unresponsive | 0
lethargic | 0
lack of interest in environment | 0
slow responses to stimulation | 0
tendency to fall asleep | 0
blood pressure 131/91 mm Hg | 0
pulse rate 78 beats/min | 0
respiratory rate 15 breaths/min | 0
oxygen saturation 99.8% | 0
afebrile | 0
no signs of meningeal irritation | 0
pupils 4 mm and equally reactive to light | 0
no evidence of ophthalmoplegia | 0
no facial asymmetry | 0
no cranial nerve deficits | 0
moved all extremities spontaneously | 0
biceps, triceps, brachioradialis, patellar, and ankle reflexes all 1+ | 0
no ankle clonus | 0
Babinski sign absent | 0
past history of atrial fibrillation | -8760
past history of right frontal ischemic stroke | -8760
survived cardiac arrest | -8760
received pacemaker/defibrillator | -8760
fully recovered | -8760
CT of the head showed encephalomalacia in the right frontal lobe | 0
electrocardiogram showed regular atrial-sensed ventricular-paced rhythm | 0
nonconvulsive seizures/status epilepticus ruled out by stat EEG | 0
blood counts, blood chemistry, and chest X-ray were normal | 0
tissue plasminogen activator not administered | 0
intubated for airway protection | 0
admitted to the intensive care unit | 0
repeat head CT 12 hours later revealed bilateral paramedian thalamic infarcts | 12
CT angiography showed filling defects at the top of the basilar artery and the P1 segments of the posterior cerebral arteries | 12
clopidogrel added to aspirin | 12
intravenous levetiracetam administered | 12
cEEG recording over a 48-hour period showed diffuse slowing and no signs of abnormal cortical hyperexcitability | 12
methylphenidate started on day 3 | 72
became progressively more alert | 72
started following simple commands | 72
extubation attempted on day 6 | 144
failed due to upper airway edema | 144
tracheostomy and percutaneous endoscopic gastrostomy on day 9 | 216
lapsed into stupor on day 12 | 288
blood pressure 144/95 mm Hg | 288
pulse rate 72 beats/min | 288
respiratory rate 18 breaths/min | 288
oxygen saturation 99.1% | 288
telemetry showed normal rate and rhythm | 288
blood test results were normal | 288
no clear evidence of a new stroke | 288
EEG recording showed sustained generalized epileptiform discharges | 288
convulsive seizure of the legs | 288
lorazepam 2 mg injected | 291
attenuation and dissipation of epileptiform discharges | 291
right third nerve palsy | 291
stat CT of the head showed extension of the infarct from the paramedian zones of the thalami to the paramedian zones of the midbrain | 291
cEEG showed waxing-waning generalized epileptiform discharges | 291
increasing the dose of levetiracetam and phenytoin and intermittent boluses of lorazepam temporarily suppressed NCSE | 291
adding sodium valproate to her antiepileptic regimen resulted in suppression of epileptiform activity | 291
became more alert and responsive | 291
remained nonverbal and only followed simple commands | 291
discharged to a long-term acute care facility on hospital day 33 | 792