15 years old | 0
male | 0
admitted to the hospital | 0
blurring of vision | -360
drowsy | 0
Glasgow coma scale 12/15 | 0
tubercular meningitis | -720
short stature | 0
height 140 cm | 0
weight 25 kg | 0
hypertelorism | 0
downslanting prominent eyes | 0
thick lips | 0
high palatal arch | 0
Mallampati score 3 | 0
limited neck extension | 0
mouth opening 4 cm | 0
scoliosis of dorsal spine | 0
reduced volume of thorax | 0
systolic murmur | 0
sinus tachycardia | 0
heart rate 140 beats/min | 0
systemic hypertension | 0
blood pressure 180/100 mm Hg | 0
high blood pressure during previous hospitalization | -720
untreated hypertension | -720
Cushing's reflex | -720
no family history of Noonan's syndrome | 0
no past medical or surgical history | 0
mild motor delay | 0
growth retardation | 0
physical deformities since birth | 0
no cardiac or respiratory decompensation symptoms | 0
hemoglobin 12.8 g/dl | 0
normal serum electrolytes | 0
normal glucose | 0
normal liver function tests | 0
normal renal function tests | 0
normal coagulation profile | 0
normal platelet count | 0
chest X-ray | 0
X-ray neck anterior-posterior and lateral view | 0
non-contrast computed tomography head | 0
magnetic resonance imaging of the brain | 0
basilar invagination | 0
atlantoaxial dislocation | 0
poor visualization of atlas and axis | 0
altered alignment of cervical spine | 0
sinus tachycardia on electrocardiogram | 0
left ventricular hypertrophy | 0
Q-waves in leads II, III, aVF, V5, V6 | 0
hypertrophic cardiomyopathy | 0
no left ventricular outflow tract obstruction | 0
no systolic anterior motion of mitral valve | 0
poor acoustic window due to scoliosis | 0
malalignment of ribs | 0
standard monitors attached | 0
heart rate 130 beats/min | 0
SpO2 100% | 0
antibiotic prophylaxis with cefuroxime | 0
resuscitation cart ready | 0
difficult airway cart ready | 0
premedication with midazolam 1.5 mg | 0
right radial artery cannulation | 0
high blood pressure | 0
systolic pressure 180-220 mm Hg | 0
diastolic pressure 100-120 mm Hg | 0
esmolol bolus 10 mg | 0
target 25% decrease in blood pressure | 0
esmolol infusion 500 μg/kg/min | 0
induction after blood pressure stabilization | 0
preoxygenation for 5 minutes | 0
induction with morphine 3 mg | 0
induction with thiopentone 100 mg | 0
successful bag-mask ventilation | 0
check laryngoscopy | 0
Cormack-Lehane Grade 2b | 0
vecuronium bromide 2.5 mg | 0
fentanyl 40 μg | 0
lignocaine 30 mg | 0
tracheal intubation with 6.5 mm tube | 0
left internal jugular vein cannulation | 0
anesthesia maintenance with O2/N2O | 0
sevoflurane 1.5 MAC | 0
small tidal volumes 4 ml/kg | 0
high respiratory rates | 0
end-tidal CO2 maintained at 30 mm Hg | 0
estimated blood loss 50 ml | 0
surgery duration 120 minutes | 0
normal intraoperative blood gas analysis | 0
pH 7.5 | 0
PaO2 97 mm Hg | 0
PaCO2 29 mm Hg | 0
HCO3 22 mmol/L | 0
urine output monitoring | 0
temperature monitoring | 0
reversal of paralysis with glycopyrrolate 0.2 mg | 0
neostigmine 1.5 mg | 0
successful extubation | 0
GCS 12 | 0
transfer to ICU | 0
shunt obstruction | 24
GCS deterioration to 7 | 24
reintubation | 24
septic shock | 360
multi-organ dysfunction syndrome | 360
death | 360
