27 years old | 0
female | 0
presented with hypotension | 0
presented with fever | 0
presented with pain | 0
presented with redness | 0
presented with swelling over both breasts | 0
bilateral liposuction of the thighs | -240
liposuction of the abdomen | -240
bilateral fat grafting to the breasts | -240
developed fever | -216
developed bilateral breast pain | -216
given paracetamol | -216
no antibiotic therapy initiated | -216
symptoms progressed to both upper arms | -168
affected skin became more erythematous | -168
affected skin became more swollen | -168
affected skin became more painful | -168
febrile | 0
in septic shock | 0
extensive erythema | 0
swelling present over chest wall | 0
swelling extending into both upper arms | 0
palpable subcutaneous crepitus | 0
clinical diagnosis of necrotizing fasciitis | 0
aggressive fluid resuscitation started | 0
inotropes started | 0
empirical intravenous penicillin G initiated | 0
clindamycin initiated | 0
ceftazidime initiated | 0
computed tomography scans revealed ill-defined masses | 0
computed tomography scans revealed large collections containing air-fluid level | 0
proceeded to surgery and debridement | 0
620 mL foul-smelling dishwater fluid evacuated | 0
435 mL fluid drained | 0
overlying skin was not necrotic | 0
breast tissue was still viable | 0
repeat debridement 24 hours after initial operation | 24
further unhealthy tissue removed | 24
planned third debridement extended into neck | 48
left sternocleidomastoid muscle involvement | 48
sepsis gradually improved | 0
bacterial cultures grew Proteus mirabilis | 0
bacterial cultures grew Enterobacter aerogenes | 0
bacterial cultures grew Enterococcus faecalis | 0
bacterial cultures grew Bacteroides fragilis | 0
antibiotic therapy adjusted to piperacillin-tazobactam | 0
required another four debridement operations | 24
wounds closed | 24
skin graft placed on right arm | 24
continues to receive regular follow-up | 0
hypertrophic scars | 0
