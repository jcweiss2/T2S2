35 years old | 0
    male | 0
    admitted to the cardiology unit | 0
    unremitting fever | -360
    chest pain | -360
    abdominal pain | -360
    palpitation | -360
    stable vitals | 0
    critical general conditions | 0
    unspecific ECG abnormalities | 0
    endocarditis | 0
    aortic valve involvement | 0
    mitral valve involvement | 0
    optimal medical therapy initiated | 0
    high risk for cardiac surgery | 0
    multiorgan failure | 0
    pulmonic failure | 0
    kidney failure | 0
    metabolic failure | 0
    septic condition | 0
    daily echocardiographic examination scheduled | 0
    CA on the 5th day | 120
    high-quality chest compressions | 120
    advanced cardiac life support procedures | 120
    ROSC in 16 min | 120
    echocardiographic check for cardiac function | 120
    right atrial thrombus formation | 120
    heparin administration 5000 IU | 120
    continued chest compressions | 120
    heparin administration 5000 IU (second bolus) | 120
    thrombus disappearance | 120
    moved to intensive care department | 120
    poor prognosis | 120
    spontaneous echo contrast | 120
    septic syndrome | 120
    hypercoagulability | 120
    acidosis | 120
    tissue hypoperfusion | 120
    