84 years old | 0
male | 0
admitted to the hospital | 0
edema on both legs | -720
diabetes mellitus | -131400
insulin | -131400
hypertension | -8760
angiotensin converting enzyme inhibitor | -8760
calcium channel blocker | -8760
right hand tremor | -61360
idiopathic Parkinsons disease | -61360
alcoholic liver cirrhosis | 0
small ascites around the liver | 0
serum albumin concentration 2.5 g/dL | 0
serum bilirubin concentration 2.4 mg/dL | 0
prothrombin time 88% | 0
Childs classification B | 0
thrombocytopenia | 0
platelets 79,000 /mm3 | 0
diabetic chronic renal failure | 0
creatinine 2.2 mg/dL | 0
mild cardiomegaly | 0
brain natriuretic peptide 193 pg/mL | 0
left ventricle ejection fraction 55% | 0
leg edema improved | 48
diuretics | 48
albumin | 48
dyspnea | 192
tachycardia 123 beats/min | 192
tachypnea 30 breaths/min | 192
hypoxemia SaO2 80% | 192
creatine kinase within normal range | 192
CK-MB within normal range | 192
troponin-I within normal range | 192
electrocardiography no significant ST depression or elevation | 192
lung perfusion scan eliminated pulmonary embolism | 192
oxygen supplementation | 192
SaO2 below 90% | 192
tachypnea 32 breaths/min | 192
septic shock | 192
endotracheal intubation | 192
transferred to intensive care unit | 192
hypotension blood pressure 75/40 mm Hg | 216
mean arterial pressure 48 mm Hg | 216
tachycardia 130 beats/min | 216
hypothermia 34℃ | 216
WBC 700/mm3 | 216
Hb 9.7 g/dL | 216
platelet count 59,000/mm3 | 216
BUN/Cr 57/2.2 mg/dL | 216
C-reactive protein 8.3 mg/dL | 216
lactic acid concentration 4.4 mmol/L | 216
urinalysis no nitrate or pyuria | 216
urine culture no growth | 216
chest radiograph no pneumonic consolidation | 216
diagnostic ascites tapping not performed | 216
hospital-acquired infection | 216
blood culture examination | 216
piperacillin/tazobactam | 216
ciprofloxacin | 216
intravenous fluid | 216
central venous pressure 12 mmHg | 216
systolic blood pressure 80 mmHg | 216
dobutamine 10 µg/kg/min | 216
dopamine 25 µg/kg/min | 216
norepinephrine 100 µg/min | 216
central venous catheter right subclavian vein | 216
anuria | 216
exacerbated azotemia | 216
continuous veno-venous hemodialysis | 216
norepinephrine infusion for 26 hours | 216
mean arterial pressure low | 216
skin necrosis not developed before vasopressin | 216
vasopressin infusion 0.02 unit/min | 216
systolic blood pressure increased to 120 mmHg | 216
mean arterial pressure increased to 80 mmHg | 216
multiple purpura on both wrists and lower legs | 220
skin necrosis expanded to both arms, thighs, abdomen | 220
superficial erosion | 220
bullous lesions | 220
low-dose vasopressin induced skin necrosis | 220
discontinued vasopressin infusion | 242
Escherichia Coli growth confirmed | 242
continuous dobutamine | 242
continuous norepinephrine | 242
hemodynamic instability | 242
died | 242
