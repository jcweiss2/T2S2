39 years old | 0
male | 0
intensive care unit admission | 0
ventilator-associated pneumonia | -1080
Acinetobacter baumannii infection | -1080
confusion | -1080
intra-abdominal trauma | -1080
traffic accident | -1080
pustular eruptions on erythematous areas (facial and neck region) | -96
pustular eruptions spread to upper and lower extremities | -96
fever (39.5℃) | -168
tigecycline 50 mg IV twice daily | -120
ventilator-associated nosocomial pneumonia | -120
sepsis | -120
mild erupted lesions | -48
tigecycline treatment stopped | -48
A. baumannii recovered from tracheal aspirate cultures | -24
tigecycline treatment restarted | -24
generalized erupted lesions (skin) | 0
erythema (face and neck) | 0
pustules (face, neck, legs) | 0
dermatologic examination | 0
oral examination (no pathologies) | 0
psoriasis (negative personal and family history) | 0
family history (no known allergies) | 0
fever | 0
leukocytosis | 0
pustule culture (negative) | 0
AGEP diagnosis | 0
pustular psoriasis differential diagnosis | 0
intravenous methylprednisolon 60 mg/d | 0
local moisturizers | 0
topical steroids | 0
new pustule appearance stopped | 24
healing with exfoliation | 24
dermatologic pathologies resolved (except facial area) | 360
death (sepsis and multiorgan failure) | 2160
