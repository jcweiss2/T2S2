69 years old | 0
    woman | 0
    labile blood pressure | 0
    recurrent headaches | 0
    paresthesias | 0
    lightheadedness | 0
    decreased hearing | 0
    garbled speech | 0
    word-finding difficulties | 0
    episodic thoracic back pain | 0
    dyspnea | 0
    hypertensive emergency | 0
    pulmonary edema | 0
    troponin 0.02 ng/mL | 0
    troponin peaked at 6.77 ng/mL | 0
    demand ischemia | 0
    recent angiogram with patent coronary arteries | -24
    ECG non-specific anterolateral and inferior ST changes | 0
    transient left bundle branch block | 0
    QT prolongation | 0
    echocardiogram moderate concentric left ventricular hypertrophy | 0
    wall motion abnormalities consistent with apical ballooning syndrome | 0
    akinesis of the mid1 to apical left ventricular myocardium | 0
    left ventricular ejection fraction 37% | 0
    hypertension | 0
    anxiety | 0
    former smoker | -302400
    quit smoking approximately 35 years ago | -302400
    denied alcohol use | 0
    denied illicit drug use | 0
    previously consumed 1–3 glasses of wine daily | -1440
    quit alcohol 2 months prior | -1440
    mother died from heart disease | 0
    father died from bladder cancer | 0
    brother had a stroke | 0
    family history negative for genetic syndromes | 0
    history of 3 prior episodes of reversible stress-induced cardiomyopathy | -26280
    labile hypertension | 0
    nonspecific neurological complaints | 0
    generalized anxiety disorder | 0
    intolerance to beta-blockers | 0
    first diagnosed with takotsubo cardiomyopathy 3 years prior | -26280
    presented with chest pain | -26280
    no trigger identified | -26280
    echocardiogram LVEF 20% | -26280
    apical dyskinesis | -26280
    coronary angiogram minimal non-obstructive CAD | -26280
    3-month follow-up echocardiogram | -25920
    complete resolution of wall motion abnormalities | -25920
    LVEF normalization to 55–65% | -25920
    second episode of cardiomyopathy 21 months later | -18240
    presented with hypertensive emergency | -18240
    pulmonary edema | -18240
    LVEF 20% | -18240
    new apical dyskinesis | -18240
    hyperkinetic base | -18240
    no cause found | -18240
    repeat echocardiogram 1 month later | -18000
    normal echocardiogram | -18000
    no wall motion abnormalities | -18000
    normal LVEF | -18000
    third hospital presentation 14 months later | -720
    nonspecific neurological complaints | -720
    decreased hearing | -720
    slurred speech | -720
    facial paresthesias | -720
    right upper extremity paresthesias | -720
    uncontrolled hypertension | -720
    pulmonary edema | -720
    blood pressure labile | -720
    echocardiogram LVEF 40% | -720
    severe basal hypokinesis | -720
    preserved function of the apical myocardium | -720
    reverse takotsubo | -720
    repeat angiogram unchanged | -720
    CT/CTA of the chest | -720
    no significant vascular abnormalities | -720
    irregular heterogenous lesion along the left adrenal gland | -720
    outpatient follow-up arranged | -720
    24-hour urine collection elevated epinephrine 230 µg | -720
    normal norepinephrine | -720
    normal cortisol | -720
    normal dopamine | -720
    home medications beta-blocker | 0
    home medications losartan/hydrochlorothiazide | 0
    not on alpha-blockade | 0
    self-discontinued carvedilol | 0
    intolerance to metoprolol | 0
    intolerance to nebivolol | 0
    believed beta-blockers caused neurological symptoms | 0
    blood pressure labile | 0
    multiple medication changes | 0
    admitted to intensive care unit | 0
    hypertensive emergency managed | 0
    severe anxiety managed | 0
    nicardipine drip | 0
    IV labetalol | 0
    lorazepam | 0
    elevated plasma metanephrines | 0
    confirmed adrenal mass | 0
    started on alpha-blocker prazosin | 0
    left laparoscopic adrenalectomy on hospital day 12 | 12
    pathology confirmed pheochromocytoma | 12
    postoperative hypotension | 12
    required norepinephrine | 12
    recovery with normalized blood pressure | 12
    resolution of neurological symptoms | 12
    ECG normalization | 12
    discharged on post-operative day 3 | 72
    metoprolol for cardiomyopathy | 72
    follow-up at 1 month | 720
    follow-up at 6 months | 4320
    follow-up at 12 months | 8640
    no recurrence of symptoms | 8640
    anxiety improved | 8640
    tolerating metoprolol | 8640
    repeat serum metanephrines normal | 8640
    repeat echocardiogram normalization | 8640
    no residual wall motion abnormalities | 8640
    ECG unremarkable | 8640
    pheochromocytoma-induced cardiomyopathy | 0
    recurrent reversible cardiomyopathy | 0
    plasma metanephrines elevated | 0
    CT abdomen/pelves left adrenal mass | 0
    laparoscopic adrenalectomy | 12
    pathology pheochromocytoma | 12
    postoperative recovery | 12
    normalization of blood pressure | 12
    resolution of neurological symptoms | 12
    ECG normalization | 12
    discharged post-operative day 3 | 72
    metoprolol at discharge | 72
    follow-up 1, 6, 12 months | 720
    6 months | 4320
    12 months | 8640
    no recurrence of symptoms | 8640
    anxiety improved | 8640
    tolerating metoprolol | 8640
    normal serum metanephrines | 8640
    repeat echocardiogram normalization | 8640
    no wall motion abnormalities | 8640
    unremarkable ECG | 8640