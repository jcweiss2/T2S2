48 years old | 0
female | 0
postmenopausal | 0
presented with lateral neck pain | -240
pain was gradual onset | -240
no associated fever | -240
no throat pain | -240
no trauma | -240
diabetic | -240
regular oral hypoglycemic medication | -240
skipped medication for last four days | -96
hypothyroidism | -240
hypertension | -240
works at private firm | 0
has three children | 0
drinks alcohol socially | 0
thyroxine 87.5 microgram daily | 0
liraglutide 5 mg daily | 0
repaglinide 1 mg thrice daily | 0
aspirin 75 mg daily | 0
atorvastatin 10 mg daily | 0
normal BMI | 0
conscious | 0
calm | 0
cooperative | 0
well-oriented | 0
stable vitals | 0
non-revealing general examinations | 0
non-revealing systemic examinations | 0
localized ill-defined area on left neck | 0
tender area | 0
local rise in temperature | 0
crepitations felt | 0
intact distal neurovascular status | 0
palpable draining lymph nodes | 0
total leukocyte count 30,330 | 0
87% neutrophils | 0
hemoglobin 12.5 g/dl | 0
platelets 166,000/ml | 0
random blood sugar 502 mg/dl | 0
serum urea 63 | 0
serum creatinine 3.5 | 0
normal serum sodium | 0
normal serum potassium | 0
urine sugar +++ | 0
urine protein + | 0
acetone positive | 0
serum protein 6.4 g/dl | 0
serum albumin 3.3 g/dl | 0
arterial pH 7.067 | 0
pCO2 8.7 | 0
pO2 77% | 0
serum bicarbonate 12.6 | 0
diagnosis of diabetic ketoacidosis | 0
diagnosis of neck abscess | 0
admitted to ICU | 0
insulin therapy | 0
IV fluids | 0
piperacillin and tazobactam started | 0
ultrasonography neck | 0
ill-defined mass on left neck | 0
posterior acoustic shadow | 0
separate from parotid and submandibular glands | 0
size 3x6 cm | 0
neck exploration | 24
debridement of wound | 24
general anesthesia | 24
wound swab culture | 24
pseudomonas aeruginosa | 24
sensitive to amikacin | 24
sensitive to ciprofloxacin | 24
changed to ciprofloxacin 200 mg twice daily | 24
changed to amikacin 500 mg thrice daily | 24
continued regular treatment | 24
histopathology report | 24
fibrofatty tissue | 24
inflammatory cells infiltrate | 24
neutrophils | 24
histiocytes | 24
focal necrosis | 24
crushed inflammatory cell profiles | 24
suggestive of necrotizing fasciitis | 24
daily dressing | 0
stayed for next week | 168
signs of recovery | 168
tolerated oral feeding | 168
normal hematological parameters | 168
normal renal function | 168
blood sugar 166 mg/dl | 168
wound healing | 168
anti-hyperglycemic medications prescribed | 168
advised regular dressing | 168
advised blood sugar monitoring | 168
discharged home | 168
subsequent visits | 168
doing well | 168
