41 years old | 0
male | 0
admitted to the hospital | 0
fever | -2160
fatigue | -2160
weight loss | -2160
disseminated skin lesions | -2160
low urine output | -2160
mental confusion | -2160
thoracic herpes zoster | -504
HIV infection | -504
antiretroviral therapy not initiated | -504
afebrile | 0
dehydrated | 0
blood pressure 109/72 mmHg | 0
pulse rate 130 beats/min | 0
oxygen saturation 97% | 0
mental confusion (GCS 14) | 0
clear lung sounds | 0
innocent abdomen | 0
no peripheral lymphadenopathy | 0
diffuse maculopapular skin lesions | 0
crusty skin lesions | 0
hemoglobin 13.9 g/dL | 0
white blood cell count 6,500/mm3 | 0
platelet count 82,000/mm3 | 0
C-reactive protein 26.1 mg/dL | 0
creatinine level 4.0 mg/dL | 0
sodium concentration 127 mg/dL | 0
lactate dehydrogenase 5,782 U/L | 0
aspartate aminotransferase 342 U/L | 0
alanine aminotransferase 340 U/L | 0
total bilirubin 3.9 mg/dL | 0
direct bilirubin 3.4 mg/dL |%3
