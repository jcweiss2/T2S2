25 years old | 0
primiparous | 0
healthy | 0
uneventful pregnancy | 0
presented to the labour ward | 0
spontaneous labour |.0
39 weeks pregnant | 0
normal vaginal delivery | 0
right medio-lateral episiotomy | 0
discharged home | 24
postpartum day 1 | 24
postpartum day 2 | 48
presented to the emergency room | 48
general weakness | 48
severe pain | 48
swelling at the episiotomy site | 48
tachycardia | 48
pulse rate of 110 BPM | 48
normal blood pressure | 48
125/80 mmHg | 48
perineal examination | 48
ecchymosis | 48
induration | 48
severe tenderness | 48
no crepitus | 48
elevated white blood count | 48
WBC 40 × 10^9/L | 48
elevated C-reactive protein | 48
CRP 170 mg/L | 48
intravenous fluids | 48
broad-spectrum antibiotics | 48
ceftriaxone | 48
metronidazole | 48
gentamicin | 48
urgent exploration of the episiotomy site | 48
general anaesthesia | 48
no obvious hematoma | 48
no pus collection | 48
viable tissues in the episiotomy bed | 48
culture swabs collected | 48
surgical drain sited | 48
episiotomy wound edges approximated with interrupted sutures | 48
clinical picture deteriorated rapidly | 72
tachycardia | 72
hypotension | 72
no response to IV fluids resuscitation | 72
transferred to the intensive care unit | 72
CRP rise to 200 mg/L | 72
WBC rise to 60 × 10^9/L | 72
pelvic CT scan | 72
bulky uterus | 72
pelvic ascites | 72
no evidence of tissue fluid or gas collection | 72
surgical consultation sought | 72
laparoscopy | 72
explore ascites | 72
exclude uterine rupture | 72
re-explore episiotomy site | 72
no evidence of uterine rupture | 72
no pelvic hematoma | 72
100 mL ascitic fluid drained | 72
culture swabs obtained | 72
incision lateral to episiotomy site | 72
unviable tissue | 72
tissue extending from right labia majora to upper medial thigh | 72
extensive tissue debridement | 72
healthy viable tissues reached | 72
wound left open | 72
iodine-soaked pack applied | 72
antibiotics adjusted | 72
clinical condition improved | 96
several debridements under anaesthesia | 96
viable tissues in wound | 96
V-Y advancement fascial flap | 168
complete closure of wound | 168
discharged | 168
followed up in outpatient department | 168
recovered completely | 168
pregnant again six months later | 168
regular antenatal care | 168
elective cesarean section | 168
39 weeks gestation | 168
Hailey-Hailey disease | 72
acantholysis | 72
dyskeratosis | 72
epidermal hyperplasia | 72
polymicrobial infection | 72
E. coli | 72
Enterococcus faecalis | 72
Bacteroides fragilis | 72
histopathological examination | 72
no Group A Streptococcus | 72
no Group B Streptococcus | 72
no Staphylococcus | 72
no Klebsiella | 72
no Pseudomonas | 72
no Peptostreptococcus | 72
no Peptococcus | 72
written consent obtained | 0
