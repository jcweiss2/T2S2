41 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
history of untreated hypertension | -672 | 0 | Factual
history of morbid obesity | -672 | 0 | Factual
history of chronic back pain | -672 | 0 | Factual
history of IVDU | -672 | 0 | Factual
low back pain | -336 | 0 | Factual
diffuse abdominal pain | -336 | 0 | Factual
lower extremity weakness | -336 | 0 | Factual
anorexia | -336 | 0 | Factual
fever | -336 | 0 | Factual
chills | -336 | 0 | Factual
shortness of breath | -336 | 0 | Factual
dizziness | -336 | 0 | Factual
constipation | -336 | 0 | Factual
recent use of acetaminophen | -168 | 0 | Factual
recent use of gabapentin | -168 | 0 | Factual
recent use of hydrocodone | -168 | 0 | Factual
recent use of methamphetamines | -168 | 0 | Factual
recent use of marijuana | -168 | 0 | Factual
blood pressure of 79/53 mmHg | 0 | 0 | Factual
heart rate of 149 bpm | 0 | 0 | Factual
lactic acid of 4.2 mg dl-1 | 0 | 0 | Factual
WBC 37 500 u l-1 | 0 | 0 | Factual
erythrocyte sedimentation rate 75 mm h-1 | 0 | 0 | Factual
urine toxicology positive for cannabis | 0 | 0 | Factual
urine toxicology positive for amphetamines | 0 | 0 | Factual
midline tenderness of the lumbar spine | 0 | 0 | Factual
3/5 strength in bilateral lower extremities | 0 | 0 | Factual
bilateral shoulder warmth | 0 | 0 | Factual
bilateral shoulder erythema | 0 | 0 | Factual
bilateral shoulder tenderness | 0 | 0 | Factual
limited range of motion | 0 | 0 | Factual
multiple needle puncture sites on the antecubital fossas | 0 | 0 | Factual
puncture wounds on the right foot | 0 | 0 | Factual
blood cultures collected | 0 | 0 | Factual
empirically started on vancomycin | 0 | 0 | Factual
empirically started on metronidazole | 0 | 0 | Factual
empirically started on aztreonam | 0 | 0 | Factual
empirically started on IV fluids | 0 | 0 | Factual
MRSA with sensitivities to vancomycin | 24 | 24 | Factual
MRSA with sensitivities to rifampin | 24 | 24 | Factual
MRSA with sensitivities to levofloxacin | 24 | 24 | Factual
MRSA with sensitivities to clindamycin | 24 | 24 | Factual
MRSA with sensitivities to daptomycin | 24 | 24 | Factual
MRSA with sensitivities to linezolid | 24 | 24 | Factual
bilateral shoulder plain radiographs showed no abnormalities | 24 | 24 | Factual
arthrocentesis of the AC joints | 48 | 48 | Factual
WBC of 93 137 u l-1 in one shoulder | 48 | 48 | Factual
WBC of 32 043 u l-1 in the other shoulder | 48 | 48 | Factual
aspirates cultured and grew MRSA | 48 | 48 | Factual
emergent surgical debridement of the shoulders | 72 | 72 | Factual
intubated | 72 | 72 | Factual
MRI of the lumbar spine showed L3-L5 osteomyelitis | 96 | 96 | Factual
MRI of the lumbar spine showed facet septic arthritis | 96 | 96 | Factual
MRI of the lumbar spine showed dorsal paraspinous myositis | 96 | 96 | Factual
MRI of the lumbar spine showed L2-L5 epidural abscess | 96 | 96 | Factual
MRI of the lumbar spine showed bilateral psoas myositis and abscesses | 96 | 96 | Factual
MRI of the bilateral shoulders after debridement showed septic arthritis of the AC joints | 120 | 120 | Factual
MRI of the bilateral shoulders after debridement showed right distal trapezius abscess | 120 | 120 | Factual
MRI of the bilateral shoulders after debridement showed left supraclavicular abscess | 120 | 120 | Factual
MRI of the brain showed no acute intracranial processes | 120 | 120 | Factual
TTE was negative for any valvular vegetations | 120 | 120 | Factual
cardiology deferred acquiring a transoesophageal echocardiogram | 120 | 120 | Factual
repeat surgical debridement of the shoulders | 144 | 144 | Factual
neurosurgery evaluated the patient for possible debridement of the epidural abscess | 144 | 144 | Factual
leukocytosis continued to rise and peaked at 52 100 u l-1 | 168 | 168 | Factual
trough levels of vancomycin were being monitored | 168 | 168 | Factual
repeat blood cultures continued to be positive for MRSA | 168 | 168 | Factual
antibiotics escalated to daptomycin and ceftaroline | 240 | 240 | Factual
blood cultures ultimately became negative | 336 | 336 | Factual
rifampin was added to the current antibiotic regimen | 336 | 336 | Factual
patient required critical care until she was stable for extubation | 336 | 336 | Factual
repeat MRI of the lumbar spine showed worsening epidural abscess | 432 | 432 | Factual
neurosurgery took the patient for surgical drainage with drain placement | 432 | 432 | Factual
intraoperative wound cultures were positive for MRSA and Proteus mirabilis | 432 | 432 | Factual
patient improved clinically | 504 | 504 | Factual
all drains were removed | 504 | 504 | Factual
patient was discharged | 672 | 672 | Factual
prescribed oral levofloxacin and rifampin | 672 | 672 | Factual
lost to follow-up | 672 | 672 | Factual