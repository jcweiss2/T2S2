38 years old | 0
female | 0
fever | -48
fatigue | -48
arthralgia | -48
furuncle-like skin lesion located on the inside of left arm | 0
admitted to the institution | 0
generalized abdominal pain | 0
nausea | 0
vomiting | 0
general discomfort | 0
nasogastric tube placement | 0
dyspnea grade IV | 0
desaturation | 0
CT scan | 0
right perirenal abscess | 0
thickening of the left renal vein | 0
bilateral pulmonary septic impacts | 0
bilateral mild pleural effusion | 0
intensive care unit admission | 0
bilateral hypoventilation | 0
jaundice | 0
oligoanuria | 0
low platelet count | 0
urine culture | 0
blood culture | 0
empirical treatment with vancomycin plus tazobactam | 0
anticoagulation treatment with Low Molecular Weight Heparin | 0
warfarin | 0
severe sepsis | 0
multi-organ failure | 0
mechanical respiratory assistance | 0
dialysis | 0
clindamycin | 0
fever persisted | 0
multi-organ failure persisted | 0
blood culture positive for methicillin-resistant Staphylococcus aureus | 0
gram-negative bacillus verified in alveolar fluid wash | 0
antibiotic scheme of vancomycin, daptomycin, and meropenem | 0
bacteremia | 12
persistent fever | 12
mechanical respiratory assistance continued | 12
inotropic drugs | 12
dialysis continued | 12
new thorax abdomen and pelvis tomography | 12
phleboectasia | 12
thrombus extending to inferior vena cava | 12
surgical exploration | 12
bilateral nephrectomy | 12
thrombectomy | 12
torpid evolution after surgery | 12
feverish records | 12
colistin started | 12
antibiotic scheme vanco-dapto-mero-colistin | 12
bronchoalveolar lavage | 12
Serratia + Kleb KPC culture | 12
culture of intra-surgical samples showed yeast | 12
fluconazole started | 12
antibiotic scheme vanco-dapto-mero-colistin-fluco | 12
improved after 11 days | 23
antibiotic scheme vanco-colistin-fluco | 23
left thoracentesis | 23
antibiotic scheme vanco + fluco + colistin + mero + metronidazole | 23
regular evolution persisted | 26
episodes of intermittently altered hemodynamic status | 26
vancomycin continued | 26
blood cultures x2 | 26
adrenal profile requested | 26
suprarenal insufficiency diagnosed | 26
hydrocortisone started | 26
improved general condition | 26
transferred to intermediate care unit | 63
urology division follow-up | 73
three-weekly dialysis | 73
discharged from hospital | 73
mental health follow-up | 73
decolonization treatment suggested | 73
body cleaning with chlorhexidine | 73
daily application of mupirocin in nostrils | 73
avoid sharing personal items | 73
