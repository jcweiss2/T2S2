75 years old | 0
male | 0
admitted to the hospital | 0
collapse | 0
seizures | 0
end stage renal disease (ESRD) | -672
intermittent dialysis | -672
left lacunar infarct in temporal lobe | -672
coronary artery bypass graft (CABG) | -2880
hypertension | -672
chronic obstructive pulmonary disease (COPD) | -672
atrial fibrillation | -672
warfarin | -672
confused | 0
pupils equal and reactive to light | 0
Glasgow coma scale of 12/15 | 0
tachycardic | 0
hypotensive | 0
tachypnoec | 0
raised renal parameters | 0
altered coagulation profile | 0
intubated | 0
mechanically ventilated | 0
right radial artery cannulated | 0
blood pressure and ABG measurements | 0
cannula in situ for 7 days | 0
cannula removed | 168
skin site inflamed | 168
wound swab grew MRSA | 168
inflammation settled | 168
distinct bulging of the radial artery | 216
ultrasound performed | 216
radial artery pseudoaneurysm diagnosed | 216
angiogram confirmed diagnosis | 216
radial artery compressed | 216
pseudoaneurysm ruptured | 280
surgical intervention | 280
surgical exploration of the radial artery | 280
pseudoaneurysm confirmed | 280