69 years old | 0
male | 0
admitted to the hospital | 0
septic shock | 0
bloody diarrhea | -72
hypertension | -672
cardiomyopathy | -672
chronic obstructive pulmonary disease | -672
laryngeal carcinoma | -672
amoxicillin/clavulanic acid | -672
confused mental state | 0
hypotension | 0
temperature | 0
diffuse abdominal tenderness | 0
increased inflammation parameters | 0
renal insufficiency | 0
low albumin | 0
normal lactate | 0
broad-spectrum antibiotics | 0
abdominal CT-scan | 0
diffuse colonic wall thickening | 0
mucosal enhancement pattern | 0
infiltration | 0
C. difficile | 0
vancomycin | 0
metronidazole | 0
vasopressor support | 216
progressive abdominal distension | 216
delirium | 216
metabolic acidosis | 216
surgical consultation | 216
colectomy | 216
FMT | 288
fidaxomicin | 288
nasoduodenal tube | 288
improvement | 432
decrease in abdominal distension | 432
negative feces polymerase chain reactions | 432
discharged from the ICU | 672
no recurrent CDI | 672