52 years old | 0\
male | 0\
admitted to the hospital | 0\
right upper quadrant pain | -168\
abdominal fullness | -168\
abdominal distention | -168\
paroxysmal pain | -168\
worsened after meals | -168\
diagnosed with hepatic abscess | -24\
treated with hepatic puncture and drainage | -24\
afebrile | 0\
pulse rate of 80 beats/minute | 0\
blood pressure of 118/73 mmHg | 0\
respiratory rate of 26 breaths/minute | 0\
leukocyte count of 16.4×10^9/L | 0\
haemoglobin level of 85 g/L | 0\
platelet count of 240×10^9/L | 0\
procalcitonin level of 2.3 ng/mL | 0\
plasma fibrinogen level of 7.48 g/L | 0\
serum glutamic oxalacetic transaminase level of 67 U/L | 0\
glutamic-pyruvic transaminase level of 83 U/L | 0\
cholinesterase level of 1360 U/L | 0\
total protein level of 50.8 g/L | 0\
albumin level of 21.5 g/L | 0\
blood urea nitrogen level of 10.8 mmol/L | 0\
creatinine level of 51.3 umol/L | 0\
negative for HIV | 0\
negative for syphilis | 0\
abdominal distension | 48\
mild bellyache | 48\
extreme thirst | 48\
right abdominal tenderness | 48\
temperature of 36.8 °C | 48\
drainage catheter yield of 150 mL of fulvous fluid | 48\
submitted to the microbiology laboratory for analysis | 48\
abdominal and pelvic computed tomography scan | 48\
irregular, slightly low-density lesion in the right posterior hepatic lobe | 48\
gas density shadow inside | 48\
liquid density shadow and high-density drainage tube shadow | 48\
round-like low-density lesion of about 0.8 cm in diameter | 48\
appendix thickened to about 20 mm in diameter | 48\
structure of the ascending colon near the ileocecal region became disorganised | 48\
multiple gas accumulation and dilation in the bowel | 48\
air-fluid levels inside the abdomen | 48\
hepatic abscesses | 48\
ileus | 48\
mild ascites | 48\
appendicitis | 48\
liver cyst | 48\
abdominal infection | 48\
peritonitis | 48\
pre-shock | 72\
insufficient blood pressure of 93/59 mmHg | 72\
taken to the operating room for urgent exploratory laparotomy | 72\
fulvous purulent exudate and necrotic tissue | 72\
partial postnecrotic defect in the peritoneum | 72\
massive epiploon adhesion in the right upper abdomen | 72\
two perforations | 72\
ileocecal resection | 72\
partial resection of the ascending colon | 72\
ileostomy | 72\
drainage of hepatic, abdominal and extraperitoneal abscesses | 72\
postoperative course was eventful | 72\
orotracheal intubation | 72\
hypotension | 72\
anemia | 72\
fever | 72\
transferred to the intensive care unit | 72\
noradrenaline | 72\
ventilator | 72\
intravenous hydration | 72\
nutritional support therapy | 72\
blood transfusion | 72\
empirically started on intravenous tigecycline and piperacillin/tazobactam | 72\
temperature went up to 39.3°C | 96\
pulse rate of 130 beats/minute | 96\
leukocyte count of 35.9×10^9 cells/L | 96\
PCT level of 8.15 ng/mL | 96\
CRP level of 174 mg/L | 96\
blood samples were taken for aerobic and anaerobic cultures | 96\
anaerobic blood culture vials were reported to be positive | 120\
Gram stain revealed short Gram-positive bacillus without spores | 120\
positive culture broth was inoculated onto blood agar base medium | 120\
anaerobically incubated for three more days | 120\
colony from the agar plate was identified as E. lenta | 120\
MALDI-TOF MS | 120\
antimicrobial susceptibility testing of E. lenta was not performed | 120\
plasma fibrinogen fell to 1.0 g/L | 120\
tigecycline was replaced by teicoplanin | 120\
piperacillin/tazobactam was discontinued | 120\
ertapenem was added to teicoplanin | 120\
cultures of the drainage fluid were obtained | 120\
isolation of organism as Escherichia coli | 120\
treated with ertapenem and teicoplanin | 120\
fever, leukocytosis, PCT level and CRP level promptly improved | 120\
transferred to the general ward | 120\
administered ertapenem and teicoplanin for another 14 days | 120\
debridement, dressing change and symptomatic supportive treatment | 120\
repeated blood cultures after the introduction of antibiotics were negative | 120\
repeat CT revealed that the size of the hepatic abscess and the amount of ascites decreased | 120\
symptoms achieved further alleviation | 216\
discharged from the hospital | 216\
prescription for oral antibiotics | 216\
follow-up with a six-week course of intravenous ertapenem | 216\
complete resolution of the abscess | 216