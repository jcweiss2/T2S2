75 years old | 0
female | 0
dementia | 0
left THA | -18000
osteaoarthritis | -18000
left hip pain | -72
inability to ambulate | -72
dislocation | -72
posterosuperior prosthetic hip dislocation | -72
internally rotated left leg | -72
shortened left leg | -72
left hip pain | -72
detailed neurovascular examination | -72
no neurovascular deficits | -72
closed reduction attempted | 0
general anesthesia | 0
paralytic agent | 0
axial traction | 0
90 degrees of flexion | 0
internal rotation | 0
adduction | 0
flexion | 0
external rotation | 0
radiographs | 0
difficult reduction | 0
dense sciatic nerve motor injury | 0
no motor function below the knee | 0
decreased sensation | 0
paresthesia | 0
peroneal nerve distribution | 0
tibial nerve distribution | 0
severe reaction to anesthesia | 0
florid acute pulmonary edema | 0
Takotsubo cardiomyopathy | 0
intensive care unit admission | 0
transfer to tertiary referral center | 72
closed reduction | 72
specialized traction table | 72
Hana table | 72
axial traction | 72
internal rotation | 72
external rotation | 72
leg adduction | 72
bone fragment | 72
ischium | 72
medial aspect of the acetabulum | 72
nerve exploration | 72
tenuous medical condition | 72
discharged home | 120
ankle foot orthosis | 120
recurrent dislocation | 504
bending over | 504
play with grandchildren | 504
persistent instability | 504
difficulty of prior closed reduction attempts | 504
ongoing sciatic nerve injury | 504
revision | 504
sciatic nerve exploration | 504
extensile posterior approach | 504
laceration of sciatic nerve | 504
60% of entire width | 504
neurolysis | 504
ceramic-on-polyethylene articulation | 504
dual-mobility liner | 504
primary cup | 504
7 mm of added head length | 504
22 + 7-mm inner-diameter ball | 504
41-mm polyethylene sphere | 504
peripheral nerve consult | 504
forgo sciatic nerve repair | 504
postoperative sensation | 504
diminished sensation | 504
abnormal sensation | 504
sciatic nerve distribution | 504
0/5 motor function | 504
sciatic nerve distribution | 504
dislocation event | 720
inability to maintain posterior hip precautions | 720
spinopelvic immobility | 720
stable | 1008
no further dislocation events | 1008
ambulating with walker | 1008
slap foot/steppage gait | 1008
no pain | 1008
discontinued ankle foot orthosis | 1008
heel ulcer | 1008
nerve injury | 1008
neuropathy | 1008