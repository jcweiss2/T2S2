65 years old | 0 | 0 
male | 0 | 0 
admitted to the hospital | 0 | 0 
no history of smoking | 0 | 0 
no underlying pulmonary diseases | 0 | 0 
not vaccinated against COVID-19 | 0 | 0 
shortness of breath | -96 | 0 
fever | -96 | 0 
dry cough | -96 | 0 
fatigue | -96 | 0 
reduced breath sounds | 0 | 0 
oxygen saturation 93% | 0 | 0 
bilateral peripheral ground-glass attenuation | 0 | 0 
patchy consolidation | 0 | 0 
lung involvement 60%-70% | 0 | 0 
nasopharyngeal SARS-CoV-2 RT-PCR test positive | 0 | 0 
negative SARS-CoV-2 RT-PCR test | 504 | 504 
increased temperature | 0 | 468 
decreased oxygen saturation | 0 | 468 
white cell count 7.93 х 109/ L | 0 | 0 
neutrophils 80% | 0 | 0 
lymphocytes 8% | 0 | 0 
monocytes 10% | 0 | 0 
plasma cell 2% | 0 | 0 
hemoglobin 159 g/l | 0 | 0 
platelet count 468 × 109/l | 0 | 0 
Westergren ESR 41 mm/h | 0 | 0 
interleukine 6 102 pg/ml | 0 | 0 
С-reactive protein 142 mg/l | 0 | 0 
ferritin 939.92 μg/ml | 0 | 0 
D-dimer 609 ng/ml | 0 | 0 
procalcitonin 0.11 ng/ml | 0 | 0 
treatment with dexamethason | 0 | 720 
treatment with heparin | 0 | 720 
treatment with tocilizumab | 0 | 720 
treatment with acetylcysteine | 0 | 720 
treatment with pantoprazole | 0 | 720 
treatment with nadroparin calcium | 0 | 720 
oxygen supplementation | 0 | 720 
air and pleural effusion in the right pleural cavity | 360 | 360 
collapse of the right lung | 360 | 360 
thoracentesis | 360 | 360 
thoracostomy | 360 | 360 
evacuation of 1400 ml of pleural fluid | 360 | 360 
linezolid therapy | 360 | 720 
imipenem/cilastatin therapy | 360 | 720 
increased oxygen supplementation | 360 | 720 
daily drainage volume 300-1000 ml | 360 | 720 
pleural effusion with gas bubbles | 432 | 432 
focal area of subpleural infiltration | 432 | 432 
central cavity of destruction | 432 | 432 
air layer along the anterior chest wall | 432 | 432 
hydropneumothorax | 432 | 432 
exudative lymphocytic-rich effusion | 432 | 432 
Acinetobacter baumannii in pleural fluid | 504 | 504 
Pseudomonas aeruginosa in pleural fluid | 504 | 504 
Klebsiella pneumonia in urine | 504 | 504 
needle thoracocentesis | 504 | 504 
new pleural drainage | 504 | 504 
air and creamy purulent mass | 504 | 504 
serofibrinous hemorrhagic fluid | 504 | 720 
pleural empyema | 576 | 576 
transfer to the Surgical Department | 576 | 576 
irrigation with antiseptic solutions | 576 | 720 
lung expansion by continuous vacuum aspiration | 576 | 720 
encapsulated pleural effusion | 624 | 624 
ultrasound-guided puncture | 624 | 624 
new drainage of the pleural cavity | 624 | 624 
colistimethatum natrium therapy | 576 | 720 
imipenem/cilastatin therapy | 576 | 720 
discharge from the hospital | 720 | 720 
oxygen saturation 97% | 720 | 720 
small amount of fluid in the right pleural cavity | 720 | 720 
normal lab test scores | 720 | 720 
С-reactive protein 11.7 mg/l | 720 | 720 
procalcitonin < 0.1 ng/ml | 720 | 720