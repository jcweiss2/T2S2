64 years old | 0
male | 0
hypertension | 0
tobacco consumption | 0
moderate obesity | 0
BMI 31 kg/m² | 0
weight 91 kg | 0
height 1.71 m | 0
moderate alcohol consumption | 0
30 g/day alcohol | 0
hepatocellular carcinoma | 0
right liver tumor | 0
appendicular syndrome | 0
abdominal pain | 0
right iliac fossa pain | 0
preoperative evaluation | 0
no liver cirrhosis | 0
no portal hypertension | 0
normal liver function | 0
prothrombin time 100% | 0
bilirubinemia 9 µmol/L | 0
albuminemia 43 g/L | 0
creatininemia 69 µmol/L | 0
platelet count 303 G/L | 0
CT | 0
MRI | 0
tumor extending into segment I | 0
tumor extending into segment IV | 0
close contact with inferior vena cava | 0
preoperative liver volumetry | 0
total liver volume 1924 cm³ | 0
tumor-free volume 204 cm³ | 0
left liver volume 484 cm³ | 0
future liver remnant-to-body weight ratio 0.5% | 0
right liver volume 1644 cm³ | 0
extended right hepatectomy | 0
segment I resection | 0
Dissectron device use | 0
remnant left liver fixation | 0
perioperative Doppler ultrasound control | 0
vascular patency | 0
intermittent portal clamping | 0
43 minutes portal clamping | 0
caval clamping | 0
20-minute caval clamping periods | 0
total operating time 10 hours | 0
no hemodynamic insufficiency | 0
amine drugs not required | 0
6 L crystalloids administered | 0
2 red blood cell transfusions | 0
R0 resection | 0
well-differentiated hepatocellular carcinoma | 0
Edmondson and Steiner grade II | 0
pT2 classification | 0
microvesicular steatosis | 0
macrovesicular steatosis | 0
50% non-tumoral parenchyma steatosis | 0
postoperative pulmonary embolism | 48
POD 2 pulmonary embolism | 48
non-severe pulmonary embolism | 48
remnant liver volume 711 cm³ | 48
33% initial total liver volume | 48
liver-to-body weight ratio 0.8% | 48
PHLF | 120
POD 5 PHLF | 120
PT 49% | 120
hyperbilirubinemia 125 µmol/L | 120
significant ascites | 120
2 L/24h ascites | 120
ascites infection | 120
Proteus mirabilis sepsis | 120
antibiotic treatment | 120
intensive care transfer | 120
ICU stay 14 days | 168
POD 9 remnant liver volume 916 cm³ | 216
43% initial total liver volume | 216
liver-to-body weight ratio 1% | 216
POD 18 contrasted-enhanced CT | 432
bilirubin 565 µmol/L | 432
PT 73% | 432
left hepatic vein stenosis | 432
DUS confirmation | 432
loss of triphasic flow | 432
stricture of left hepatic vein | 432
cavography confirmation | 432
LHV-IVC gradient 9 mmHg | 432
percutaneous transluminal angioplasty | 432
metallic stent placement | 432
diameter 10 mm | 432
length 6 cm | 432
LHV-IVC gradient decreased to 3 mmHg | 432
post-intervention recovery uneventful | 432
progressive bilirubinemia reduction | 432
discharge | 720
POD 30 discharge | 720
two months post-surgery bilirubin 230 µmol/L | 1440
normal PT | 1440
four months bilirubin normal | 2880
10-month follow-up | 7200
no late complications | 7200
normal liver function tests | 7200
no patient complaints | 7200
left remnant liver regeneration 1300 cm³ | 7200
post-hepatectomy remnant-to-body ratio 1.2% | 7200
satisfactory inflow | 7200
satisfactory outflow | 7200
no liver failure recurrence | 7200
metallic stent permeable | 7200
metallic stent in place | 7200
