56 years old | 0
female | 0
height 146 cm | 0
weight 74 kg | 0
arterial hypertension | -72
valsartan 80 mg/day | -72
hydrochlorothiazide 12.5 mg/day | -72
admitted to the hospital | 0
carpal tunnel release surgery | 0
general anesthesia | 0
induction of anesthesia with propofol 120 mg | 0
remifentanil 10 μ10i | 0
fentanyl | 0
rocuronium 50 mg | 0
oral intubation | 0
endotracheal tube 6.5 mm internal diameter | 0
cuff inflated with 4 ml of air | 0
anesthesia maintained with desflurane | 0
surgery lasted 25 minutes | 25
anesthesia discontinued | 25
endotracheal tube suctioned | 25
patient coughed vigorously | 25
violent neck movement | 25
extubated endotracheal tube not tinged with blood | 25
transferred to post-anesthesia care unit | 25
chest discomfort | 30
dyspnea | 30
swelling of the neck and upper anterior chest | 30
arterial blood gasses | 30
pH = 7.32 | 30
PCO2 = 51 mmHg | 30
PO2 = 78 mmHg | 30
HCO3 = 26.8 mmol/L | 30
SpO2 = 93% | 30
chest X-ray | 30
pneumomediastinum | 30
subcutaneous emphysema | 30
computed tomography scan | 30
tracheal laceration | 30
bronchoscopy | 30
tracheal defect 5 cm linear | 30
thoracic surgeon’s opinion | 30
thoracic surgical repair impossible | 30
intensive care unit | 30
7.5 mm ID cuffed endotracheal tube | 30
low-tidal-volume lung ventilation | 30
pressure-controlled mode | 30
tidal volume 250 - 350 ml/kg | 30
frequency 20 - 25/min | 30
pressure-limited ventilation | 30
permissive hypercapnia | 30
broad-spectrum intravenous antibiotics | 30
patient improved | 72
chest CT | 72
mediastinal and subcutaneous emphysema reduced | 72
bronchoscopy | 192
lesion healing | 192
endotracheal tube extubation | 312
patient discharged | 317