78 years old | 0
male | 0
Caucasian | 0
former smoker | 0
40 pack-year history of tobacco use | 0
chronic obstructive pulmonary disease (COPD) | 0
prostate cancer | 0
postradical prostatectomy | 0
radiation therapy | 0
radiation colitis | 0
admitted to the hospital | 0
shortness of breath | -48
altered mental status | -24
productive cough | -48
subjective fevers | -48
confusion | -24
inability to get into bed | -24
hypotensive | 0
blood pressure of 92/61 | 0
tachycardic | 0
heart rate of 130 | 0
tachypneic | 0
respiratory rate of 25 | 0
hypoxic | 0
oxygen saturation of 71% | 0
afebrile | 0
temperature of 99.9°F | 0
alert and oriented | 0
diminished breath sounds | 0
scattered crackles | 0
noninvasive positive pressure ventilation with BiPAP | 0
leukocytosis | 0
white blood cell 30.6 | 0
12% bands | 0
lactic acidosis | 0
lactic acid of 3.6 mmol/l | 0
acute kidney injury | 0
creatinine of 1.5 mg/dl | 0
baseline creatinine of 0.8 mg/dl | 0
left upper and lower lobe opacity | 0
pneumonia | 0
pneumonia severity index of 131 | 0
Class V management strategy | 0
intubation with mechanical ventilation | 12
broad-spectrum antibiotics | 12
vancomycin | 12
piperacillin-tazobactam | 12
azithromycin | 12
healthcare-associated pneumonia (HCAP) | 12
blood cultures positive for P. multocida | 48
ownership of five cats | -720
involvement in cat care and grooming | -720
switch to ampicillin-sulbactam | 48
clinical improvement | 96
extubation | 168
discharge | 432
amoxicillin-clavulanic acid | 432
completion of 14 days of antibiotic therapy | 720
recent hospitalization for COPD exacerbation | -1440
suspected bowel obstruction | -1440