48 years old | 0
female | 0
admitted to the hospital | 0
intractable migraine headaches | -14400
history of migraine headaches | -14400
DHE 0.5 mg × 1 | 0
DHE 1 mg every 8 h | 0
DHE for 8 doses | 0
DHE on days 1-3 | 0
DHE on days 7-9 | 168
obtunded | 192
minimally responsive | 192
hypotensive | 192
blood pressure 80/45 mm Hg | 192
abdomen moderately distended | 192
few bowel sounds | 192
lactate acid level 4.5 mmol/l | 192
white blood cell count 18.0 | 192
stool Clostridium difficile negative | 192
transferred to the intensive care unit | 192
intravenous fluid boluses | 192
vasopressors | 192
broad spectrum antibiotics | 192
intubation | 192
chest radiograph unremarkable | 192
abdominal x-rays mild prominence of the colon | 192
progressively acidotic | 216
worsening bandemia | 216
bedside colonoscopy | 216
diffuse ischemic colitis | 216
fecal impaction | 216
no pseudomembranes | 216
laparotomy | 240
peritoneal cavity filled with murky fluid | 240
gangrene of the descending colon | 240
necrosis in the area distal to the splenic flexure | 240
necrosis to the sigmoid colon | 240
impacted stool in the left colon | 240
vasculature intact | 240
audible Doppler signals | 240
removal of the gangrenous bowel | 240
condition improved | 240
final pathology | 264
surgical specimen | 264
86 cm of patchy dark green/black large bowel | 264
ischemic necrosis | 264
bowel wall intact | 264
gangrenous large bowel | 264
ischemic colitis | 264
thrombi or emboli | 264
hypercoaguable panel | 264
negative for clotting disorders | 264
discharged | 720