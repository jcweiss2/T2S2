18 years old | 0
male | 0
admitted to the hospital | 0
cough | -72
fevers | -72
shortness of breath | -72
pleuritic chest pain | -72
light-headedness | -72
near syncope | -72
acutely worsened dyspnoea | -72
obesity | -72
body mass index (BMI) 37 | -72
febrile | -72
tachycardic | -72
normotensive | -72
hypoxic saturating 82% on room air | -72
COVID-19 | -72
positive nasopharyngeal qualitative polymerase chain reaction (PCR) | -72
acute sub-massive pulmonary embolism (PE) | -72
unfractionated heparin (UFH) | -72
hypotensive | -48
massive PE | -48
catheter-directed thrombolysis (CDT) | -48
bilateral pulmonary arteries | -48
improved clinically | -24
discharged | -24
acute respiratory failure | 0
hypotension | 0
intubated | 0
cardiac arrest | 0
return of spontanous circulation (ROSC) | 0
vasopressors | 0
veno-arterial extracorporeal membrane oxygenation (ECMO) | 0
pulmonary artery angiogram | 0
interval worsening of bilateral pulmonary emboli | 0
recurrence of massive PE | 0
repeat CDT | 0
ventilation parameters improved | 24
vasopressors were discontinued | 24
ECMO weaned | 24
venous duplex ultrasound | 24
deep venous thrombus of the right femoral vein and right popliteal vein | 24
inferior vena cava (IVC) filter | 24
UFH transitioned to low-molecular weight heparin | 24
repeat pulmonary artery angiogram | 24
improvement in emboli burden | 24
successfully weaned from ECMO | 24
decannulated | 24
septic shock | 40
right thigh haematoma with compartment syndrome | 40
surgical debridement | 40
transitioned to rivaroxaban | 40
discharged | 52
returned home | 99
perform activities of daily living independently | 99
anticoagulated on rivaroxaban 20 mg daily | 99
no major adverse events | 99
COVID-19 | -72
SARS-CoV-2 infection | -72
coagulopathy | -72
pulmonary embolism (PE) | -72
sub-massive PE | -72
massive-PE | -48
catheter directed thrombolysis (CDT) | -48
extracorporeal membrane oxygenation (ECMO) | -48
repeat CDT | -48
recurrent massive PE | -48
septic shock | 40
treated with broad spectrum antibiotics | 40
right thigh haematoma and compartment syndrome | 40
surgical debridement | 40
transitioned to rivaroxaban | 40
discharged | 52
returned home | 99
perform activities of daily living independently | 99
anticoagulated on rivaroxaban 20 mg daily | 99
no major adverse events | 99