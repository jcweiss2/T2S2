9 years old | 0
female | 0
eastern Indian origin | 0
admitted to the emergency room | 0
abdominal pain | -72
fever | -72
nausea | -72
vomiting | -72
completed 2-dose Pfizer-BioNTech COVID-19 immunization series | -744
SARS-CoV-2 PCR test positive | -384
asymptomatic | -384
traveled to the US Virgin Islands | -384
returned to the United States | -168
persistent fever | -168
emesis | -168
nausea | -168
abdominal pain | -168
respiratory viral PCR panel negative | -72
oseltamivir | -72
painful area at the tip of her tongue | -72
presented to the emergency department | 0
persistently febrile | 0
maximum temperature of 40°C | 0
heart rate between 124 and 133 beats per minute | 0
respiratory rate between 20 and 30 breaths/min | 0
oxygen saturation 96% to 100% | 0
blood pressure 94 to 102/44 to 54 mm Hg | 0
mild conjunctival injection | 0
epigastric abdominal tenderness | 0
mild hyponatremia | 0
leukopenia | 0
thrombocytopenia | 0
lymphopenia | 0
elevated inflammatory markers | 0
IVIG treatment started | 0
empiric ceftriaxone and doxycycline started | 0
antibiotics discontinued | 72
macular, nonpruritic, nonpetechial rash | 5
bilateral conjunctival injection | 24
afebrile | 24
prednisone started | 24
intermittent episodes of confusion and agitation | 24
DVT prophylaxis with low-molecular weight heparin started | 24
anticoagulation discontinued | 48
aspirin not started | 48
inflammatory markers trended downward | 48
pancytopenia persisted | 48
hemoglobin 9.7 g/dL | 72
red blood cell count 3.61 M/uL | 72
platelet count 30,000/uL | 72
white blood cell count 2580 cells/uL | 72
absolute lymphocyte count 240 | 72
BNP increased to 4114 pg/mL | 72
echocardiography remained normal | 72
complement levels normal | 96
anti-nuclear antibody positive | 96
proinflammatory markers IL-6 and CXCL-9 elevated | 96
direct antibody test negative | 96
bone marrow aspiration not performed | 96
thrombocytopenia began to improve | 168
platelet count 104 000/uL | 168
discharged | 168
follow-up laboratories showed platelet count recovering | 1008
ALC, WBC, and Hgb recovering | 1008
mild persistent fatigue | 1008
closely followed by cardiology, rheumatology, hematology and oncology, and infectious disease specialists | 1008
no evolution of an alternative diagnosis | 1008