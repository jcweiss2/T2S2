13 years old | 0
female | 0
admitted to the hospital | 0
marked hepatomegaly | 0
laparoscopy | 0
liver biopsy | 0
large and typically orange-yellow liver | 0
greatly elevated hepatic content of cholesteryl esters | 0
lysosomal enzyme defect in the fibroblast culture | 0
headaches | 0
feeling of pressure in the right epigastrium | 0
increasing jaundice | 0
bilirubin 6.0 mg/dL | 0
total cholesterol 316 mg/dL | 0
HDL cholesterol 26 mg/dL | 0
triglycerides 178 mg/dL | 0
alpha1-antitrypsin 363 mg/dL | 0
hospitalized in 2013 | -262080
laparoscopic cholecystectomy | -262080
symptomatic gallstones | -262080
chronic and florid fibroplastic cholecystitis | -262080
Child-Pugh A/B cirrhosis | -262080
Lab-MELD 14 cirrhosis | -262080
esophageal varices grade III | -262080
solitary fundal varix | -262080
hepatosplenomegaly | -262080
thrombocytopenia | -262080
vitamin D deficiency | -262080
calcium deficiency | -262080
discharged without medication | -262080
readmitted in July 2016 | -1728
subjective increase in abdominal circumference | -1728
tiredness | -1728
scleral jaundice | -1728
nausea | -1728
pruritus | -1728
lack of appetite | -1728
Child-Pugh C cirrhosis | -1728
Lab-MELD score 18 | -1728
increased NSAIDs use | -1728
axillary herpes zoster | -1728
hepatic encephalopathy occurred twice | -1728
rifaximin given for 4 months | -1728
esophageal varices | -1728
fundal varices | -1728
Histoacryl treatment | -1728
elevated transaminases | -1728
pancytopenia | -1728
abnormal clotting tests | -1728
early discharge | -1728
readmitted for acute onset of epigastric pain | -720
rapid improvement in symptoms | -720
prompt discharge requested | -720
re-hospitalized with febrile urinary tract infection | -480
E. coli sepsis | -480
parenteral antibiotics treatment | -480
admitted in September 2016 | 0
compensated cirrhosis | 0
splenomegaly | 0
planned repeat ligature of esophageal varices | 0
exclusion of relevant fundal varices | 0
vomited blood | 24
emergency endoscopy | 24
Histoacryl treatment of esophageal varix | 24
bleeding stopped temporarily | 24
transfer to intensive care ward | 24
intubated and ventilated | 24
emergency transfusion of erythrocytes | 24
ROTEM-based clotting factor replacement | 24
bleeding arrested by esophageal stent | 24
clipping of acute Forrest Ia bleed in the cardia | 24
severe coagulopathy | 24
hemorrhagic shock developed | 24
laboratory abnormalities indicated infection | 24
antibiotics given | 24
replacement treatment for severe hypoalbuminemia | 24
diffuse nosebleed | 24
tamponade treatment | 24
inability to stabilize patient | 24
Hb-relevant diffuse bleeding tendency persisted | 24
dried blood test on September 9, 2016 | 168
reduced acid lipase 0.03 nmol/spot*3 hours | 168
reduced beta-galactosidase 0.08 nmol/spot*21 hours | 168
apoptosis marker M30 rose | 144
overall cell death marker M65 rose | 144
progressive hepatic decompensation | 144
clotting situation not stabilized | 144
multiorgan failure | 144
liver transplant not possible | 144
no further escalation of intensive medical therapy | 144
patient died | 360
multiorgan failure as sequelae of advanced liver disease | 360
increased troponin I | 360
increased myoglobin | 360
pathological cardiovascular changes | 360
