18 years old | -672
female | -672
gravida one | -672
fever | -168
prolonged premature rupture of membranes (PPROM) | -168
betamethasone | 0
ampicillin | 0
gentamicin | 0
mechanical ventilation | 0
emergency cesarean section delivery | 0
birth | 0
mechanical ventilation | 0
intravenous ampicillin | 0
intravenous gentamicin | 0
extubated | 24
noninvasive ventilation | 24
less active | 72
temperature instability | 72
bradycardia | 72
vancomycin | 72
cefotaxime | 72
multiple episodes of apnea | 72
deteriorating bradycardic spells | 72
desaturation | 72
hypercarbia | 72
re-intubated | 72
synchronized intermittent mandatory ventilation | 72
cefepime | 72
fluconazole | 72
acyclovir | 72
increasing metabolic acidosis | 96
worsening respiratory failure | 96
high frequency oscillating ventilation | 96
hypotensive | 96
poor perfusion | 96
vasopressors | 96
blood products | 96
patent ductus arteriosus | 96
left-to-right shunt | 96
pulmonary hypertension | 96
small pericardial effusion | 96
moderately decreased left ventricular function | 96
low cardiac output | 96
sepsis | 96
severe metabolic acidosis | 96
disseminated intravascular coagulation | 96
cardiopulmonary arrest | 120
death | 120
mucocutaneous culture sampled | 72
HSV positive | 120
placental pathology report | 0
third-trimester placenta | 0
moderate intervillous fibrosis | 0
no chorioamnionitis | 0
no funisitis | 0
autopsy | 120
normally developed premature female infant | 120
no dysmorphic features | 120
no congenital anomalies | 120
serous fluid in the right pleural cavity | 120
serous fluid in the left pleural cavity | 120
serosanguineous ascites | 120
normal-sized heart | 120
unremarkable immature myocardium | 120
ductus arteriosus open | 120
foramen ovale open | 120
hemorrhagic right upper and middle lobes | 120
thickened septa | 120
saccular stage of development | 120
disorganized large cells | 120
viral nuclear inclusions | 120
HSV-infected cell | 120
multinucleated cell | 120
margination of chromatin | 120
molding | 120
viral nuclear inclusion | 120
diffuse fibrin plugs | 120
diffuse alveolar hemorrhage | 120
bloody mucus | 120
normal mucosa | 120
centrilobular congestion | 120
hemorrhage around portal areas | 120
hemorrhage under the capsule | 120
hepatocyte nuclei | 120
viral inclusions | 120
margination of chromatin | 120
wine red appearance | 120
immunohistochemistry for HSV-1 and HSV-2 | 120
positive | 120
peripelvic hemorrhage | 120
no herpetic infection | 120
karyorrhexis | 120
perivascular cell fragments | 120
microglial nodules | 120
thalamus | 120
midbrain | 120
HSV isolated from postmortem lung cultures | 120
disseminated HSV infection | 120
resolving hyaline membrane disease | 120
ascites | 120
pleural effusion | 120
persistent ductus arteriosus | 120
involution of thymus | 120
medullary congestion | 120
pelvic hemorrhage of the kidneys | 120