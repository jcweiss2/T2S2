42 years old | 0
female | 0
admitted to the hospital | 0
elective parathyroidectomy | 0
stag horn calculus | -672
hyperparathyroidism | -672
morbid obesity | -672
BMI 75 | -672
limited exercise tolerance | -672
obstructive sleep apnea (OSA) | -672
hypertension | -672
diabetes | -672
acid reflux disease | -672
hepatitis C | -672
smoker | -672
postoperative nausea and vomiting (PONV) | -672
insulin | -672
lisinopril | -672
hydrochlorthiazide | -672
atorvastatin | -672
aspirin | -672
venlafaxine | -672
trazadone | -672
rosuvastatin | -672
premedicated with sodium citrate | -3
premedicated with ranitidine | -3
intravenous canula placed | -2
arterial line placed | -2
preoxygenated | -1
anesthesia induced with propofol | -1
anesthesia induced with suxamethonium | -1
trachea intubated | -1
anesthesia maintained with oxygen/air | 0
anesthesia maintained with sevoflurane | 0
rocuronium given | 0
neck explored | 0
parathyroid adenoma resected | 4.5
parathyroid hormone levels normalized | 4.75
transferred to ICU | 4.5
propofol infusion started | 4.5
propofol dose escalated | 5
failed spontaneous breathing test (SBT) | 24
respiratory failure | 24
basal atelectasis | 24
ventilator-associated pneumonia | 24
rhabdomyolysis | 72
myoglobin levels elevated | 72
urine output declined | 72
creatinine levels elevated | 72
BUN levels elevated | 72
acute renal failure | 72
septic shock | 72
metabolic acidosis | 72
norepinephrine given | 72
propofol infusion stopped | 72
lorazepam given | 72
fentanyl given | 72
dialyzed | 72
rhabdomyolysis resolved | 240
renal failure resolved | 240
tracheostomy | 384
decubitus ulcer | 384
died | 1560