56 years old| 0
    male | 0
    admitted to the hospital | 0
    prosthetic aortic graft infection | 0
    aortobifemoral graft | 0
    lifestyle-limiting claudication | 0
    hypertension | 0
    transient ischemic attack | 0
    acute occlusion of left limb of graft | -8760
    thrombectomy attempt | -8760
    femoral crossover graft | -8760
    acute right groin pain | -4344
    swelling | -4344
    erythema | -4344
    abscess around right limb of graft | -4344
    Proteus mirabilis infection | -4344
    Staphylococcus epidermidis infection | -4344
    Enterococcus faecalis infection | -4344
    intravenous daptomycin | -4344
    intravenous teicoplanin | -4344
    oral ciprofloxacin | -4344
    explant of aortobifemoral graft | -4344
    explant of femoral crossover graft | -4344
    rifampicin-bonded graft | -4344
    omental wrap | -4344
    severe systemic inflammatory response | 0
    pyrexia | 0
    tachycardia | 0
    large right groin abscess | 0
    anterior abdominal wall cellulitis | 0
    groin cellulitis | 0
    inflammatory changes around aortic anastomosis | 0
    inflammatory changes around left limb of graft | 0
    right common iliac artery patent | 0
    right internal iliac artery patent | 0
    common femoral arteries patent | 0
    profunda femoris arteries patent | 0
    right superficial femoral artery occlusion | 0
    left superficial femoral artery severe stenosis | 0
    small bowel fistulae onto graft | 0
    infrarenal aortic clamp placement | 0
    Dacron graft excision | 0
    arteriosclerosis of aortic wall | 0
    use of previous aortotomy | 0
    sartorius flaps | 0
    vasopressor support | 72
    renal replacement therapy | 72
    sepsis | 72
    major surgery | 72
    lower limb ischemia/reperfusion injury | 72
    left leg compartment syndrome | 48
    four-compartment fasciotomy | 48
    venous hypertension | 48
    severe abdominal pain | 264
    back pain | 264
    hypovolemic shock | 264
    aortic anastomotic pseudoaneurysm | 264
    endovascular salvage | 264
    left axillary artery exposure | 264
    GORE Dry Seal sheath placement | 264
    Amplatzer vascular plugs placement | 264
    Medtronic flared limb stent graft | 264
    completion angiography | 264
    exclusion of pseudoaneurysm | 264
    discharge | 240
    intravenous ertapenem | 240
    intravenous daptomycin | 240
    multidrug-resistant E coli infection | 240
    vancomycin-resistant Enterococcus infection | 240
    oral doxycycline | 240
    oral trimethoprim | 240
    white cell count normal | 2160
    C-reactive protein normal | 2160
    albumin normal | 2160
    surveillance CT angiogram | 2160
    no inflammatory change around aortic reconstruction | 2160
