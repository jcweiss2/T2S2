51 years old | 0
male | 0
admitted to the hospital | 0
gas gangrene suspicion | 0
emphysema | 0
warm skin | 0
local tenderness | 0
septic shock | 0
blood pressure 100/50mmHg | 0
mean arterial pressure 68mmHg | 0
heart rate 110bpm | 0
body temperature 39.0°C | 0
fluid resuscitation | -3
tobacco abuse | -6720
nickel allergy | -6720
sciatica | -6720
cortisone injections | -6720
non-steroidal anti-inflammatory drugs | -6720
emergency surgery | 0
muscles incised | 0
grey muscles | 0
malodor | 0
right hemipelvectomy | 0
double-transverse transversostoma | 0
debridement | 0
histology | 0
soft tissue necrosis | 0
muscle necrosis | 0
phlegmonous inflammation | 0
empirical antibiotic therapy | 0
Meropenem | 0
Linezolid | 0
Penicillin G | 0
Clindamycin | 0
postoperative CT scan | 2
acicular foreign body | 2
rectoscopy | 4
toothpick perforation | 4
sigmoid colon perforation | 4
rectoscopy | 4
toothpick removal | 4
second control CT examination | 12
peritonitis | 12
free intraabdominal air | 12
laparotomy | 12
sigmoid colon resection | 12
transversostoma rearranged | 12
proctosigmoidectomy | 12
clinical improvement | 24
wound revisions | 48
plastic coverage | 72
ESBL-Escherichia coli | 72
antibiotic therapy deescalation | 120
Meropenem monotherapy | 120
Levofloxacin | 150
discontinued | 180
mobilization | 432
transfer to rehabilitation | 504