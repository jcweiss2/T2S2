70 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
emergency esophageal diversion | -1300 | -1300 | Factual
injury to the cervical esophagus | -1300 | -1300 | Factual
spinal surgery | -1300 | -1300 | Factual
gastric pull-up procedure | -504 | -504 | Factual
postoperative anastomotic leakage | -504 | -504 | Factual
endoscopy | -504 | -504 | Factual
esophageal stent | -504 | -504 | Factual
local cervical infection | -378 | -378 | Factual
sepsis | -378 | -378 | Factual
arterial hypertonus | 0 | 0 | Factual
non-active smoking status | 0 | 0 | Factual
ischemic stroke | 0 | 0 | Factual
incomplete senso-motoric hemiparesis | 0 | 0 | Factual
thyroidectomy | 0 | 0 | Factual
open prostatectomy | 0 | 0 | Factual
prostate cancer | 0 | 0 | Factual
malnutrition | 0 | 0 | Factual
systemic inflammation | 0 | 0 | Factual
jugular and cervical phlegmon | 0 | 0 | Factual
hemoglobin level of 6.7 g/dL | 0 | 0 | Factual
white blood cell count of 6400 cells/μL | 0 | 0 | Factual
platelet count of 210 × 10^3/μL | 0 | 0 | Factual
creatinine level of 0.76 mg/dL | 0 | 0 | Factual
unremarkable liver and cholestasis parameters | 0 | 0 | Factual
albumin level of 2.8 g/dL | 0 | 0 | Factual
dislodged esophageal stent | 0 | 0 | Factual
esophageal perforation | 0 | 0 | Factual
infected cavity | 0 | 0 | Factual
esophageal stenosis | 0 | 0 | Factual
endoscopic vacuum therapy | 0 | 336 | Factual
EsoSponge system | 0 | 336 | Factual
jugular and cervical phlegmon resolved | 168 | 336 | Factual
repeated endoscopic balloon dilatation | 168 | 336 | Factual
subtotal esophageal resection | 336 | 336 | Factual
reconstruction using a free-jejunal graft interposition | 336 | 336 | Factual
CT angiography | 336 | 336 | Factual
partial sternotomy | 336 | 336 | Factual
laparotomy | 336 | 336 | Factual
harvesting of a jejunal segment | 336 | 336 | Factual
implantation of the graft | 336 | 336 | Factual
cervical anastomosis | 336 | 336 | Factual
upper mediastinal gastro-jejunostomy | 336 | 336 | Factual
resection of the upper sternum | 336 | 336 | Factual
coverage with a sternocleidomastoid muscle flap | 336 | 336 | Factual
abdominal reconstruction | 336 | 336 | Factual
end-to-end jejunojejunostomy | 336 | 336 | Factual
postoperative course uneventful | 336 | 672 | Factual
oral alimentation reestablished | 336 | 672 | Factual
daily speech therapy | 336 | 672 | Factual
anastomotic healing confirmed | 672 | 672 | Factual
transfer to a rehabilitation clinic | 672 | 672 | Factual
cervical esophagocutaneous fistula | 0 | 336 | Factual
anastomotic stenosis | 0 | 336 | Factual
chronic malnutrition | 0 | 672 | Factual
systemic inflammation | 0 | 672 | Factual