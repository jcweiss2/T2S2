50 years old | 0
male | 0
admitted to the hospital | 0
progressive dyspnea | -72
cough | -72
cold sweats | -72
night sweating | -8760
15 kilograms weight loss | -8760
human immunodeficiency virus (HIV) infection | -156384
double-sided pneumonia | 0
Pneumocystis jirovecii | 0
acquired immunodeficiency syndrome (AIDS) | 0
antiretroviral therapy | -156384
undetectable viral load | -157680
stopped taking medication | -8760
lived in a homeless shelter | -8760
no (intravenous) drug use | 0
no alcohol use | 0
quit smoking | -131040
physical examination | 0
non-acutely ill | 0
tachypneic | 0
oxygen saturation of 88% | 0
blood pressure 130/80 mm Hg | 0
heart rate 132 per minute | 0
temperature 38.2°C | 0
percussion of the lungs | 0
no dullness | 0
auscultation normal breath sounds | 0
left lower side abnormality | 0
hemoglobin 7.2 mmol/L | 0
white blood cell count 6.6 × 10^9/L | 0
platelets 214 × 10^9/L | 0
C-reactive protein (CRP) 64 mg/L | 0
no renal insufficiency | 0
no hepatic insufficiency | 0
CD4: 0.039 × 10^9/L | 0
CD8: 1.2 × 10^9/L | 0
CD4/CD8 ratio: 0.033 | 0
chest X-ray bilateral cloudy infiltrates | 0
treated with local sepsis protocol | 0
gentamicin 280 mg | 0
amoxicillin/clavulanic acid 1200 mg | 0
cotrimoxazole 3 × 1920 mg | 24
prednisolone 2 × 40 mg | 24
suspected PJP | 24
bronchoscopy with bronchoalveolar lavage (BAL) | 48
dyspneic | 48
low oxygen saturations (82%) | 48
subcutaneous emphysema | 48
progressive respiratory insufficiency | 48
endotracheal intubation | 48
mechanical ventilation | 48
bronchoscopy-guided intubation | 48
computed tomography (CT) scan | 48
subcutaneous and mediastinal emphysema | 48
no pneumothorax | 48
severe air bronchograms | 48
bilateral infiltrations | 48
admitted to the intensive care unit (ICU) | 48
subcutaneous emphysema increased | 72
mediastinal emphysema increased | 72
swelling of the entire face | 72
swelling of the arms | 72
swelling of the torso down to the scrotum | 72
several bronchoscopies | 72
no tracheal injury | 72
lung protective ventilation | 72
low tidal volumes | 72
low airway pressures | 72
emphysema continued to increase | 72
new CT scan | 168
severe subcutaneous emphysema | 168
severe mediastinal emphysema | 168
treatment with skin incisions (blow holes) considered | 168
discarded due to high HIV viral load | 168
fear of viral spreading | 168
severity of symptoms | 168
no obvious tracheal injury | 168
search for treatment options | 168
two infraclavicular skin incisions | 168
VAC therapy initiated | 168
subcutaneous emphysema started to improve | 216
gradual clinical improvement | 216
VAC therapy ended | 240
subcutaneous emphysema continued to decrease | 240
inflammatory markers decreased | 408
pulmonary infiltrations decreased | 408
extubated | 408
significant ICU-acquired weakness | 408
dysphonia | 408
discharged to general ward | 600
antiretroviral medicine restarted | 600
discharged to rehabilitation center | 600
