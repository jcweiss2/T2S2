56 years old | 0
    male | 0
    admitted to the hospital | 0
    intermittent headache | -72
    fever | -72
    transsphenoidal pituitary adenoma resection | -26280
    gamma knife stereotactic radiosurgery (first) | -26280
    gamma knife stereotactic radiosurgery (second) | -8760
    body temperature 38.2°C | 0
    heart rate 85 bpm | 0
    blood pressure 125/78 mm Hg | 0
    respiratory rate 18 breaths/min | 0
    doubtful neck resistance | 0
    right pupil slightly larger | 0
    asthenocoria | 0
    white blood cell count 10.12×10^9/L | 0
    neutrophil ratio 59.9% | 0
    CRP 12.9 mg/L | 0
    blood glucose 6.63 mmol/L | 0
    D-dimer 860 μg/L | 0
    serum pituitary hormone tests normal | 0
    ECG normal | 0
    chest CT normal | 0
    abdominal ultrasonography normal | 0
    residual pituitary adenoma 25mm×24mm | 0
    acute residual tumor hemorrhage diagnosis | 0
    dehydration therapy | 0
    hemostasis therapy | 0
    progressive headache | 3
    sudden loss of left eye vision | 3
    loss of consciousness | 3
    arrest of spontaneous heartbeat | 3
    arrest of spontaneous breath | 3
    cardiopulmonary resuscitation | 3
    spontaneous heartbeat recovery | 3
    head CT scan | 3
    magnetic resonance imaging | 3
    MR venography | 3
    mechanical ventilation | 3
    intensive care unit transfer | 3
    endotracheal intubation | 3
    pupils equally dilated 4mm | 24
    no light reflex | 24
    GCS score 1+1+1 | 24
    highest body temperature 37.6°C | 24
    blood pressure unstable | 24
    hemodynamic unstable | 24
    lumbar puncture | 24
    intracranial pressure 400 mm H2O | 24
    CSF yellow and thick | 24
    CSF white blood cells 2520/μL | 24
    CSF neutrophils 90% | 24
    CSF red blood cells 34000/μL | 24
    CSF protein 2570 mg/L | 24
    CSF glucose 0.03 mmol/L | 24
    CSF chloride 112.7 mmol/L | 24
    lateral ventricular drainage | 24
    purulent meningitis diagnosis | 24
    septic shock diagnosis | 24
    daptomycin | 24
    linezolid | 24
    voriconazole | 24
    aerobic blood culture | 24
    anaerobic blood culture | 24
    CSF culture | 24
    Gram-negative Klebsiella pneumoniae identification | 24
    repeat CT scan | 72
    meropenem | 24
    vancomycin | 24
    bilateral ventricular irrigation suggestion | 24
    family refusal of invasive treatment | 24
    vital signs deterioration | 24
    cardiac arrest | 24
    death | 24
    