58 years old | 0
woman | 0
presented | 0
productive cough | -120
fatigue | -120
fever | -120
diarrhea | -120
diffuse rhonchi | 0
blood pressure 156/95 mm Hg | 0
heart rate 130 beats/min | 0
oxygen saturation 82% | 0
respiratory rate 24 breaths/min | 0
temperature 38.7°C | 0
chest radiograph showed bilateral infiltrates | 0
intubated | 0
hypoxic respiratory failure | 0
acute respiratory distress syndrome | 0
ECG showed sinus tachycardia | 0
ST-segment elevations in leads I and aVL | 0
PR interval depressions | 0
ST-T wave changes | 0
troponin I level negative | 0
troponin I level peaked at 11.02 ng/ml | 24
leukopenia | 0
absolute lymphocyte count 1.04 K/mm³ | 0
SARS-CoV-2 RNA detected | 0
COVID-19 positive | 0
diabetes mellitus type 2 | 0
hypertension | 0
dyslipidemia | 0
father ill with similar symptoms | 0
STEMI | 0
stress cardiomyopathy | 0
myopericarditis | 0
transthoracic echocardiogram | 0
akinetic segments | 0
hypokinetic segments | 0
hyperdynamic segments | 0
apical ballooning | 0
LV ejection fraction 20% | 0
RV akinetic | 0
RV hyperdynamic | 0
RV function mildly reduced | 0
admitted to ICU | 0
takotsubo syndrome | 0
wall motion abnormalities | 0
deferred coronary angiography | 0
dual antiplatelet therapy | 0
anticoagulation | 0
heparin | 0
hydroxychloroquine therapy | 0
discontinued hydroxychloroquine | 48
azithromycin | 0
shock | 0
cardiogenic shock | 0
septic shock |, 0
central venous oxygen saturation 42% | 0
dobutamine | 0
central venous oxygen saturation 65% | 72
dobutamine de-escalating | 72
repeat echocardiogram | 144
LV ejection fraction 55% | 144
ECG no Q-wave myocardial infarction | 144
acute respiratory distress syndrome | 144
venovenous ECMO | 144
LV function improved | 144
ECG no active ischemia | 144
ECG no infarction | 144
