42 years old | 0
male | 0
chronic alcoholism | 0
severe shock | 0
febrile (tympanic temperature 38°C) | 0
sedated with propofol | 0
invasive mechanical ventilation |4 0
blood pressure 60/40 mm Hg | 0
heart rate 120 beats/min | 0
vasopressor support (noradrenaline 0.5 μg/kg/min) | 0
ionotropic support (dobutamine 5 μg/kg/min) | 0
systolic heart murmur | 0
soft abdomen | 0
no tenderness to deep palpation | 0
leukocytosis (leukocytes 13,100/µL) | 0
anemia (hemoglobin 11.2 g/dL) | 0
mean corpuscular volume 88.2 fL | 0
prolonged international normalized ratio 5.86 | 0
high prothrombin time 71.9 s | 0
acute kidney injury (creatinine 2.3 mg/dL, urea 124 mg/dL) | 0
elevated aminotransferases (GPT 2822 U/L, GOT 5068 U/L) | 0
hyperbilirubinemia (4.8 mg/dL) | 0
elevated lactate dehydrogenase 4,245 U/L | 0
pro-calcitonin (4.47 ng/ml) | 0
N-terminal pro b-type natriuretic peptide (8,018 pg/mL) | 0
troponin (1.10 ng/mL) | 0
metabolic acidemia | 0
high lactate levels (14 mmol/L) | 0
left ventricle hypertrophy | 0
moderate-to-severe depression of global systolic function | 0
severe auricular dilatation | 0
thrombus in left auricular appendix | 0
native aortic valve vegetation | 0
severe septic shock | 0
multiple-organ dysfunction secondary to endocarditis | 0
empirical broad-spectrum antibiotics | 0
transferred to intensive care unit | 0
unknown drug abuse history | 0
negative secondary causes of immunosuppression | 0
negative syphilis | 0
blood cultures positive for Corynebacterium jeikeium | 0
initial clinical improvement | 216
severe hypotension | 216
vasopressor support re-introduced (noradrenaline 1.9 μg/kg/min) | 216
blood seen on nasogastric tube | 240
urgent upper endoscopy | 240
circumferential hemorrhagic mucosa | 240
fibropurulent plaques | 240
violaceus areas of elevated mucosa in lower third of esophagus | 240
loss of vascular pattern | 240
areas of pale mucosa | 240
hemorrhagic mucosa | 240
violaceus mucosa | 240
multiple erosions | 240
fibropurulent plaques in gastric fundus, body, antrum, duodenum | 240
biopsies consistent with extensive hemorrhagic necrosis | 240
acute kidney failure | 240
probable ischemic pancreatitis | 240
probable ischemic hepatitis | 240
contrast-enhanced abdominal computed tomography | 192
no alterations suggestive of intestinal ischemia | 192
no alterations suggestive of chronic liver disease | 192
died due to refractory multiple-organ dysfunction | 240
