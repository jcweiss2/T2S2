54 years old | 0 | 0 
male | 0 | 0 
admitted to the hospital | 0 | 0 
pre-syncope | -0.1 | 0 
syncope | -0.1 | 0 
left-sided chest tightness | -0.1 | 0 
generalized fatigue | -336 | 0 
weight loss | -336 | 0 
diffuse erythematous rash | 0 | 0 
unremarkable cardiac examination | 0 | 0 
unremarkable respiratory examination | 0 | 0 
normal sinus rhythm | 0 | 0 
raised troponin concentration | 0 | 0 
eosinophil count | 0 | 0 
referred to cardiology | 0 | 0 
myocarditis | 0 | 0 
cardiac magnetic resonance imaging | 24 | 24 
eosinophilic myocarditis | 24 | 24 
coronary angiography | 24 | 24 
no coronary artery disease | 24 | 24 
skin biopsy | 24 | 24 
cardiac biopsy | 24 | 24 
edoxaban | 48 | 744 
prednisolone | 48 | 744 
follow-up in the rheumatology clinic | 336 | 336 
missed appointment | 744 | 744 
neck swelling | 744 | 744 
urgently admitted to hospital | 744 | 744 
rise in eosinophil count | 744 | 744 
increase the dose of prednisolone | 744 | 744 
computed tomography of neck | 744 | 744 
lymphadenopathy | 744 | 744 
T-cell lymphoma | 744 | 744 
cyclophosphamide | 744 | 1200 
sepsis | 1200 | 1200 
cholecystitis | 1200 | 1200 
new onset of seizures | 1200 | 1200 
reduction in consciousness | 1200 | 1200 
Glasgow Coma Scale | 1200 | 1200 
head CT | 1200 | 1200 
multiple bilateral acute infarctions | 1200 | 1200 
transferred to the intensive care unit | 1200 | 1200 
hepatitis B | -10000 | 0 
asthma | -10000 | 0 
intravenous drug use | -10000 | 0 
excessive use of alcohol | -10000 | 0 
ischemic stroke | 1200 | 1200 
reduced GCS score | 1200 | 1200 
intracranial bleeding | 1200 | 1200 
malignancy | 744 | 744 
intracerebral infection | 1200 | 1200 
diffuse subendocardial late gadolinium enhancement | 24 | 24 
mild LV systolic impairment | 24 | 24 
eczematous changes | 24 | 24 
no increase in eosinophils | 24 | 24 
T-cell lymphoma | 744 | 744 
infarcts involving the frontal, parietal, and left temporo-occipital regions | 1200 | 1200 
apical tear | 1200 | 1200 
intramural myocardial tear | 1200 | 1200 
small apical cavity | 1200 | 1200 
small mobile structures | 1200 | 1200 
diastolic flow in the apical cavity | 1200 | 1200 
systolic flow out of the apical cavity | 1200 | 1200 
cyclophosphamide therapy | 1200 | 1200 
partial response | 1200 | 1200 
reduction of the eosinophil count | 1200 | 1200 
palliation | 1200 | 1200 
deterioration | 1200 | 1200 
poor prognosis | 1200 | 1200 
multidisciplinary team meeting | 1200 | 1200 
LV wall tear | 1200 | 1200 
EM | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
delay in diagnosis | 0 | 1200 
noncardiology specialists | 1200 | 1200 
transthoracic echocardiography | 1200 | 1200 
apical view | 1200 | 1200 
color flow Doppler | 1200 | 1200 
pulse wave Doppler | 1200 | 1200 
Glasgow Coma Scale score | 1200 | 1200 
seizures | 1200 | 1200 
reduction in consciousness | 1200 | 1200 
bilateral cerebral infarcts | 1200 | 1200 
eosinophilic myocarditis | 0 | 1200 
hypereosinophilic syndrome | 744 | 1200 
T-cell lymphoma | 744 | 1200 
eosinophil count | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
cyclophosphamide | 744 | 1200 
palliation | 1200 | 1200 
deterioration | 1200 | 1200 
poor prognosis | 1200 | 1200 
multidisciplinary team meeting | 1200 | 1200 
LV wall tear | 1200 | 1200 
EM | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
delay in diagnosis | 0 | 1200 
noncardiology specialists | 1200 | 1200 
transthoracic echocardiography | 1200 | 1200 
apical view | 1200 | 1200 
color flow Doppler | 1200 | 1200 
pulse wave Doppler | 1200 | 1200 
Glasgow Coma Scale score | 1200 | 1200 
seizures | 1200 | 1200 
reduction in consciousness | 1200 | 1200 
bilateral cerebral infarcts | 1200 | 1200 
eosinophilic myocarditis | 0 | 1200 
hypereosinophilic syndrome | 744 | 1200 
T-cell lymphoma | 744 | 1200 
eosinophil count | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
cyclophosphamide | 744 | 1200 
palliation | 1200 | 1200 
deterioration | 1200 | 1200 
poor prognosis | 1200 | 1200 
multidisciplinary team meeting | 1200 | 1200 
LV wall tear | 1200 | 1200 
EM | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
delay in diagnosis | 0 | 1200 
noncardiology specialists | 1200 | 1200 
transthoracic echocardiography | 1200 | 1200 
apical view | 1200 | 1200 
color flow Doppler | 1200 | 1200 
pulse wave Doppler | 1200 | 1200 
Glasgow Coma Scale score | 1200 | 1200 
seizures | 1200 | 1200 
reduction in consciousness | 1200 | 1200 
bilateral cerebral infarcts | 1200 | 1200 
eosinophilic myocarditis | 0 | 1200 
hypereosinophilic syndrome | 744 | 1200 
T-cell lymphoma | 744 | 1200 
eosinophil count | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
cyclophosphamide | 744 | 1200 
palliation | 1200 | 1200 
deterioration | 1200 | 1200 
poor prognosis | 1200 | 1200 
multidisciplinary team meeting | 1200 | 1200 
LV wall tear | 1200 | 1200 
EM | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
delay in diagnosis | 0 | 1200 
noncardiology specialists | 1200 | 1200 
transthoracic echocardiography | 1200 | 1200 
apical view | 1200 | 1200 
color flow Doppler | 1200 | 1200 
pulse wave Doppler | 1200 | 1200 
Glasgow Coma Scale score | 1200 | 1200 
seizures | 1200 | 1200 
reduction in consciousness | 1200 | 1200 
bilateral cerebral infarcts | 1200 | 1200 
eosinophilic myocarditis | 0 | 1200 
hypereosinophilic syndrome | 744 | 1200 
T-cell lymphoma | 744 | 1200 
eosinophil count | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
cyclophosphamide | 744 | 1200 
palliation | 1200 | 1200 
deterioration | 1200 | 1200 
poor prognosis | 1200 | 1200 
multidisciplinary team meeting | 1200 | 1200 
LV wall tear | 1200 | 1200 
EM | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
delay in diagnosis | 0 | 1200 
noncardiology specialists | 1200 | 1200 
transthoracic echocardiography | 1200 | 1200 
apical view | 1200 | 1200 
color flow Doppler | 1200 | 1200 
pulse wave Doppler | 1200 | 1200 
Glasgow Coma Scale score | 1200 | 1200 
seizures | 1200 | 1200 
reduction in consciousness | 1200 | 1200 
bilateral cerebral infarcts | 1200 | 1200 
eosinophilic myocarditis | 0 | 1200 
hypereosinophilic syndrome | 744 | 1200 
T-cell lymphoma | 744 | 1200 
eosinophil count | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
cyclophosphamide | 744 | 1200 
palliation | 1200 | 1200 
deterioration | 1200 | 1200 
poor prognosis | 1200 | 1200 
multidisciplinary team meeting | 1200 | 1200 
LV wall tear | 1200 | 1200 
EM | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
delay in diagnosis | 0 | 1200 
noncardiology specialists | 1200 | 1200 
transthoracic echocardiography | 1200 | 1200 
apical view | 1200 | 1200 
color flow Doppler | 1200 | 1200 
pulse wave Doppler | 1200 | 1200 
Glasgow Coma Scale score | 1200 | 1200 
seizures | 1200 | 1200 
reduction in consciousness | 1200 | 1200 
bilateral cerebral infarcts | 1200 | 1200 
eosinophilic myocarditis | 0 | 1200 
hypereosinophilic syndrome | 744 | 1200 
T-cell lymphoma | 744 | 1200 
eosinophil count | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
cyclophosphamide | 744 | 1200 
palliation | 1200 | 1200 
deterioration | 1200 | 1200 
poor prognosis | 1200 | 1200 
multidisciplinary team meeting | 1200 | 1200 
LV wall tear | 1200 | 1200 
EM | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
delay in diagnosis | 0 | 1200 
noncardiology specialists | 1200 | 1200 
transthoracic echocardiography | 1200 | 1200 
apical view | 1200 | 1200 
color flow Doppler | 1200 | 1200 
pulse wave Doppler | 1200 | 1200 
Glasgow Coma Scale score | 1200 | 1200 
seizures | 1200 | 1200 
reduction in consciousness | 1200 | 1200 
bilateral cerebral infarcts | 1200 | 1200 
eosinophilic myocarditis | 0 | 1200 
hypereosinophilic syndrome | 744 | 1200 
T-cell lymphoma | 744 | 1200 
eosinophil count | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
cyclophosphamide | 744 | 1200 
palliation | 1200 | 1200 
deterioration | 1200 | 1200 
poor prognosis | 1200 | 1200 
multidisciplinary team meeting | 1200 | 1200 
LV wall tear | 1200 | 1200 
EM | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
delay in diagnosis | 0 | 1200 
noncardiology specialists | 1200 | 1200 
transthoracic echocardiography | 1200 | 1200 
apical view | 1200 | 1200 
color flow Doppler | 1200 | 1200 
pulse wave Doppler | 1200 | 1200 
Glasgow Coma Scale score | 1200 | 1200 
seizures | 1200 | 1200 
reduction in consciousness | 1200 | 1200 
bilateral cerebral infarcts | 1200 | 1200 
eosinophilic myocarditis | 0 | 1200 
hypereosinophilic syndrome | 744 | 1200 
T-cell lymphoma | 744 | 1200 
eosinophil count | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
cyclophosphamide | 744 | 1200 
palliation | 1200 | 1200 
deterioration | 1200 | 1200 
poor prognosis | 1200 | 1200 
multidisciplinary team meeting | 1200 | 1200 
LV wall tear | 1200 | 1200 
EM | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
delay in diagnosis | 0 | 1200 
noncardiology specialists | 1200 | 1200 
transthoracic echocardiography | 1200 | 1200 
apical view | 1200 | 1200 
color flow Doppler | 1200 | 1200 
pulse wave Doppler | 1200 | 1200 
Glasgow Coma Scale score | 1200 | 1200 
seizures | 1200 | 1200 
reduction in consciousness | 1200 | 1200 
bilateral cerebral infarcts | 1200 | 1200 
eosinophilic myocarditis | 0 | 1200 
hypereosinophilic syndrome | 744 | 1200 
T-cell lymphoma | 744 | 1200 
eosinophil count | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
cyclophosphamide | 744 | 1200 
palliation | 1200 | 1200 
deterioration | 1200 | 1200 
poor prognosis | 1200 | 1200 
multidisciplinary team meeting | 1200 | 1200 
LV wall tear | 1200 | 1200 
EM | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
delay in diagnosis | 0 | 1200 
noncardiology specialists | 1200 | 1200 
transthoracic echocardiography | 1200 | 1200 
apical view | 1200 | 1200 
color flow Doppler | 1200 | 1200 
pulse wave Doppler | 1200 | 1200 
Glasgow Coma Scale score | 1200 | 1200 
seizures | 1200 | 1200 
reduction in consciousness | 1200 | 1200 
bilateral cerebral infarcts | 1200 | 1200 
eosinophilic myocarditis | 0 | 1200 
hypereosinophilic syndrome | 744 | 1200 
T-cell lymphoma | 744 | 1200 
eosinophil count | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
cyclophosphamide | 744 | 1200 
palliation | 1200 | 1200 
deterioration | 1200 | 1200 
poor prognosis | 1200 | 1200 
multidisciplinary team meeting | 1200 | 1200 
LV wall tear | 1200 | 1200 
EM | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
delay in diagnosis | 0 | 1200 
noncardiology specialists | 1200 | 1200 
transthoracic echocardiography | 1200 | 1200 
apical view | 1200 | 1200 
color flow Doppler | 1200 | 1200 
pulse wave Doppler | 1200 | 1200 
Glasgow Coma Scale score | 1200 | 1200 
seizures | 1200 | 1200 
reduction in consciousness | 1200 | 1200 
bilateral cerebral infarcts | 1200 | 1200 
eosinophilic myocarditis | 0 | 1200 
hypereosinophilic syndrome | 744 | 1200 
T-cell lymphoma | 744 | 1200 
eosinophil count | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
cyclophosphamide | 744 | 1200 
palliation | 1200 | 1200 
deterioration | 1200 | 1200 
poor prognosis | 1200 | 1200 
multidisciplinary team meeting | 1200 | 1200 
LV wall tear | 1200 | 1200 
EM | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
delay in diagnosis | 0 | 1200 
noncardiology specialists | 1200 | 1200 
transthoracic echocardiography | 1200 | 1200 
apical view | 1200 | 1200 
color flow Doppler | 1200 | 1200 
pulse wave Doppler | 1200 | 1200 
Glasgow Coma Scale score | 1200 | 1200 
seizures | 1200 | 1200 
reduction in consciousness | 1200 | 1200 
bilateral cerebral infarcts | 1200 | 1200 
eosinophilic myocarditis | 0 | 1200 
hypereosinophilic syndrome | 744 | 1200 
T-cell lymphoma | 744 | 1200 
eosinophil count | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
cyclophosphamide | 744 | 1200 
palliation | 1200 | 1200 
deterioration | 1200 | 1200 
poor prognosis | 1200 | 1200 
multidisciplinary team meeting | 1200 | 1200 
LV wall tear | 1200 | 1200 
EM | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
delay in diagnosis | 0 | 1200 
noncardiology specialists | 1200 | 1200 
transthoracic echocardiography | 1200 | 1200 
apical view | 1200 | 1200 
color flow Doppler | 1200 | 1200 
pulse wave Doppler | 1200 | 1200 
Glasgow Coma Scale score | 1200 | 1200 
seizures | 1200 | 1200 
reduction in consciousness | 1200 | 1200 
bilateral cerebral infarcts | 1200 | 1200 
eosinophilic myocarditis | 0 | 1200 
hypereosinophilic syndrome | 744 | 1200 
T-cell lymphoma | 744 | 1200 
eosinophil count | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
cyclophosphamide | 744 | 1200 
palliation | 1200 | 1200 
deterioration | 1200 | 1200 
poor prognosis | 1200 | 1200 
multidisciplinary team meeting | 1200 | 1200 
LV wall tear | 1200 | 1200 
EM | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
delay in diagnosis | 0 | 1200 
noncardiology specialists | 1200 | 1200 
transthoracic echocardiography | 1200 | 1200 
apical view | 1200 | 1200 
color flow Doppler | 1200 | 1200 
pulse wave Doppler | 1200 | 1200 
Glasgow Coma Scale score | 1200 | 1200 
seizures | 1200 | 1200 
reduction in consciousness | 1200 | 1200 
bilateral cerebral infarcts | 1200 | 1200 
eosinophilic myocarditis | 0 | 1200 
hypereosinophilic syndrome | 744 | 1200 
T-cell lymphoma | 744 | 1200 
eosinophil count | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
cyclophosphamide | 744 | 1200 
palliation | 1200 | 1200 
deterioration | 1200 | 1200 
poor prognosis | 1200 | 1200 
multidisciplinary team meeting | 1200 | 1200 
LV wall tear | 1200 | 1200 
EM | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
delay in diagnosis | 0 | 1200 
noncardiology specialists | 1200 | 1200 
transthoracic echocardiography | 1200 | 1200 
apical view | 1200 | 1200 
color flow Doppler | 1200 | 1200 
pulse wave Doppler | 1200 | 1200 
Glasgow Coma Scale score | 1200 | 1200 
seizures | 1200 | 1200 
reduction in consciousness | 1200 | 1200 
bilateral cerebral infarcts | 1200 | 1200 
eosinophilic myocarditis | 0 | 1200 
hypereosinophilic syndrome | 744 | 1200 
T-cell lymphoma | 744 | 1200 
eosinophil count | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
cyclophosphamide | 744 | 1200 
palliation | 1200 | 1200 
deterioration | 1200 | 1200 
poor prognosis | 1200 | 1200 
multidisciplinary team meeting | 1200 | 1200 
LV wall tear | 1200 | 1200 
EM | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
delay in diagnosis | 0 | 1200 
noncardiology specialists | 1200 | 1200 
transthoracic echocardiography | 1200 | 1200 
apical view | 1200 | 1200 
color flow Doppler | 1200 | 1200 
pulse wave Doppler | 1200 | 1200 
Glasgow Coma Scale score | 1200 | 1200 
seizures | 1200 | 1200 
reduction in consciousness | 1200 | 1200 
bilateral cerebral infarcts | 1200 | 1200 
eosinophilic myocarditis | 0 | 1200 
hypereosinophilic syndrome | 744 | 1200 
T-cell lymphoma | 744 | 1200 
eosinophil count | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
cyclophosphamide | 744 | 1200 
palliation | 1200 | 1200 
deterioration | 1200 | 1200 
poor prognosis | 1200 | 1200 
multidisciplinary team meeting | 1200 | 1200 
LV wall tear | 1200 | 1200 
EM | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
delay in diagnosis | 0 | 1200 
noncardiology specialists | 1200 | 1200 
transthoracic echocardiography | 1200 | 1200 
apical view | 1200 | 1200 
color flow Doppler | 1200 | 1200 
pulse wave Doppler | 1200 | 1200 
Glasgow Coma Scale score | 1200 | 1200 
seizures | 1200 | 1200 
reduction in consciousness | 1200 | 1200 
bilateral cerebral infarcts | 1200 | 1200 
eosinophilic myocarditis | 0 | 1200 
hypereosinophilic syndrome | 744 | 1200 
T-cell lymphoma | 744 | 1200 
eosinophil count | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
cyclophosphamide | 744 | 1200 
palliation | 1200 | 1200 
deterioration | 1200 | 1200 
poor prognosis | 1200 | 1200 
multidisciplinary team meeting | 1200 | 1200 
LV wall tear | 1200 | 1200 
EM | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
delay in diagnosis | 0 | 1200 
noncardiology specialists | 1200 | 1200 
transthoracic echocardiography | 1200 | 1200 
apical view | 1200 | 1200 
color flow Doppler | 1200 | 1200 
pulse wave Doppler | 1200 | 1200 
Glasgow Coma Scale score | 1200 | 1200 
seizures | 1200 | 1200 
reduction in consciousness | 1200 | 1200 
bilateral cerebral infarcts | 1200 | 1200 
eosinophilic myocarditis | 0 | 1200 
hypereosinophilic syndrome | 744 | 1200 
T-cell lymphoma | 744 | 1200 
eosinophil count | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
cyclophosphamide | 744 | 1200 
palliation | 1200 | 1200 
deterioration | 1200 | 1200 
poor prognosis | 1200 | 1200 
multidisciplinary team meeting | 1200 | 1200 
LV wall tear | 1200 | 1200 
EM | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
delay in diagnosis | 0 | 1200 
noncardiology specialists | 1200 | 1200 
transthoracic echocardiography | 1200 | 1200 
apical view | 1200 | 1200 
color flow Doppler | 1200 | 1200 
pulse wave Doppler | 1200 | 1200 
Glasgow Coma Scale score | 1200 | 1200 
seizures | 1200 | 1200 
reduction in consciousness | 1200 | 1200 
bilateral cerebral infarcts | 1200 | 1200 
eosinophilic myocarditis | 0 | 1200 
hypereosinophilic syndrome | 744 | 1200 
T-cell lymphoma | 744 | 1200 
eosinophil count | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
cyclophosphamide | 744 | 1200 
palliation | 1200 | 1200 
deterioration | 1200 | 1200 
poor prognosis | 1200 | 1200 
multidisciplinary team meeting | 1200 | 1200 
LV wall tear | 1200 | 1200 
EM | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
delay in diagnosis | 0 | 1200 
noncardiology specialists | 1200 | 1200 
transthoracic echocardiography | 1200 | 1200 
apical view | 1200 | 1200 
color flow Doppler | 1200 | 1200 
pulse wave Doppler | 1200 | 1200 
Glasgow Coma Scale score | 1200 | 1200 
seizures | 1200 | 1200 
reduction in consciousness | 1200 | 1200 
bilateral cerebral infarcts | 1200 | 1200 
eosinophilic myocarditis | 0 | 1200 
hypereosinophilic syndrome | 744 | 1200 
T-cell lymphoma | 744 | 1200 
eosinophil count | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
cyclophosphamide | 744 | 1200 
palliation | 1200 | 1200 
deterioration | 1200 | 1200 
poor prognosis | 1200 | 1200 
multidisciplinary team meeting | 1200 | 1200 
LV wall tear | 1200 | 1200 
EM | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
delay in diagnosis | 0 | 1200 
noncardiology specialists | 1200 | 1200 
transthoracic echocardiography | 1200 | 1200 
apical view | 1200 | 1200 
color flow Doppler | 1200 | 1200 
pulse wave Doppler | 1200 | 1200 
Glasgow Coma Scale score | 1200 | 1200 
seizures | 1200 | 1200 
reduction in consciousness | 1200 | 1200 
bilateral cerebral infarcts | 1200 | 1200 
eosinophilic myocarditis | 0 | 1200 
hypereosinophilic syndrome | 744 | 1200 
T-cell lymphoma | 744 | 1200 
eosinophil count | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
cyclophosphamide | 744 | 1200 
palliation | 1200 | 1200 
deterioration | 1200 | 1200 
poor prognosis | 1200 | 1200 
multidisciplinary team meeting | 1200 | 1200 
LV wall tear | 1200 | 1200 
EM | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
delay in diagnosis | 0 | 1200 
noncardiology specialists | 1200 | 1200 
transthoracic echocardiography | 1200 | 1200 
apical view | 1200 | 1200 
color flow Doppler | 1200 | 1200 
pulse wave Doppler | 1200 | 1200 
Glasgow Coma Scale score | 1200 | 1200 
seizures | 1200 | 1200 
reduction in consciousness | 1200 | 1200 
bilateral cerebral infarcts | 1200 | 1200 
eosinophilic myocarditis | 0 | 1200 
hypereosinophilic syndrome | 744 | 1200 
T-cell lymphoma | 744 | 1200 
eosinophil count | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
cyclophosphamide | 744 | 1200 
palliation | 1200 | 1200 
deterioration | 1200 | 1200 
poor prognosis | 1200 | 1200 
multidisciplinary team meeting | 1200 | 1200 
LV wall tear | 1200 | 1200 
EM | 0 | 1200 
corticosteroids | 48 | 744 
anticoagulation | 48 | 744 
delay in diagnosis | 0 | 1200 
noncardiology specialists | 1200 | 1200 
transthoracic echocardiography | 1200 | 1200 
apical view | 1200 | 1200 
color flow Doppler | 1200 | 1200 
pulse wave Doppler | 1200 | 1200 
Glasgow Coma Scale score | 1200 | 1200 
seizures | 1200 | 1200 
reduction in consciousness | 1200 | 1200 
bilateral cerebral infarcts | 1200 | 1200 
eosinophilic myocard