18 years old | 0
female | 0
35 weeks of gestation | 0
pregnancy | 0
in vitro fertilization | 0
facial nerve paresis | 0
healthy twins | 0
cesarean section | 0
severe headache | -24
generalized tonic-clonic seizures | -24
loss of consciousness | -24
hypertension | -24
heart rate 120 beats/min | -24
eclampsia | -24
magnesium sulphate | -24
ebrantil | -24
manitol | -24
diazepam | -24
bilateral vision loss | -24
proteinuria 2+ | -24
normal complete blood count | -24
normal liver function tests | -24
normal clotting parameters | -24
normal electrocardiogram | -24
normal other system examinations | -24
cortical blindness | -24
normal pupillary responses | -24
normal fundus findings | -24
mild right-sided facial nerve paresis | -24
hypodensity of the posterior white matter | -24
vasogenic edema | -24
MRI | -24
T2- and fluid-attenuated inversion recovery (FLAIR)-weighted images | -24
hyperintense signals in the white matter | -24
enalapril maleate | -24
methyldopa | -24
human albumin | -24
significant bilateral improvement of the visual function | -5
best-corrected visual acuity 1.0 | -5
peripheral relative scotoma | -5
depressed sensitivity of the paracentral left visual field | -5
discrete residual changes over the posterior horns of the side ventricles | -5
oral antihypertensive therapy | -5
physical therapy for the paresis of the facial nerve | -5
discharged from the clinic | -3
follow-up MRI | -3
significant regression of the edema | -3
persistent discrete residual changes over the posterior horns of the side ventricles | -3