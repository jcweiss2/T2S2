63 years old | 0
female | 0
past medical history of psychiatric disorders | -672
mild traumatic brain injury | -72
fall | -72
aspiration pneumonia | -72
no initial loss of consciousness | -72
computed tomography (CT) | -72
normal CT | -72
no sign of bleeding | -72
thin ventricles | -72
median structure in place | -72
pneumonia evolved toward ARDS | -48
prone positioning | -48
deep sedation by midazolam | -48
deep sedation by sufentanil | -48
electrical brain activity monitored by bispectral index (BIS) | -48
low BIS values | -48
discontinuation of sedative drugs | 0
recovered spontaneous ventilation | 72
no sign of waking up | 72
low BIS values | 72
sluggish reaction to painful stimuli on the left arm | 72
intermediate and reactive pupils | 72
ultrasonography | 72
transcranial Doppler (TCD) | 72
pulsatility Index = 1.09 | 72
end diastolic velocity = 52.11 cm/s | 72
ONSD measurements | 72
elevated ICP | 72
osmotherapy | 72
blood pressure elevation | 72
head elevation | 72
control of temperature | 72
control of carbon dioxide | 72
control of glycemia | 72
new brain CT | 96
multiple deep parenchymal hematomas | 96
bilateral cerebellar ischemia | 96
diffuse cerebral edema | 96
brain coning | 96
emergent treatment | 96
unfavorable evolution | 120
brain death | 192
TCD demonstrated a backflow in MCA | 192
brain death confirmed by electroencephalograms | 192