76 years old | 0
female | 0
abdominal pain | -24
fever | -24
systolic blood pressure 70 mmHg | -24
referred to hospital | 0
alert | 0
body temperature 37.9°C | 0
blood pressure 83/52 mmHg | 0
heart rate 103 beats/min | 0
respiratory rate 30/min | 0
oxygen saturation 80% | 0
abdomen soft and flat | 0
tenderness on the entire abdomen | 0
rebound tenderness on the entire abdomen | 0
autoimmune hepatitis | 0
oral steroid | 0
osteoporosis | 0
compression fracture of the spine | 0
spinal canal stenosis | 0
chronic kidney dysfunction | 0
fracture of the left hand | 0
fracture of the femur | 0
pneumonia | 0
temporomandibular joint myelitis | 0
cesarean birth with median incision at the lower abdomen | 0
elevation of WBC | 0
elevation of CRP | 0
elevation of BUN | 0
elevation of serum creatinine | 0
purulent urine | 0
rich bacteria in urine | 0
WBC in urine | 0
admitted to hospital | 0
diagnosis of ileus | 0
diagnosis of septic state | 0
Sequential Organ Failure Assessment Score 2 points | 0
ileus tube insertion | 0
transnasal endoscopy | 0
antibiotic meropenem | 0
abdominal pain worsened | 24
elevation of inflammation reaction values | 24
free air in abdominal cavity | 24
fluid collection in anterior space of bladder | 24
emergency laparotomy | 24
digestive tract perforation | 24
hole at the dome of the urinary bladder | 24
hole at the peritoneum | 24
thick pus extruded into abdominal cavity | 24
sutured the hole | 24
sutured the bladder | 24
permanent urinary catheter placement | 24
bladder drainage | 24
bladder decompression | 24
postoperative course uneventful | 24
inflammation reaction improved | 120
discharged | 504
no recurrence | 504