89 years old | 0
female | 0
admitted to the hospital | 0
loss of consciousness | 0
LOC | 0
dry cough | -48
body aches | -48
vaccinated with Sinopharm vaccine | -672
Glasgow Coma Scale score was three | 0
oral temperature was 36.5 | 0
oxygen saturation was 98% | 0
elevated lactate dehydrogenase | 0
elevated C-reactive protein level | 0
elevated ESR | 0
elevated CPK | 0
elevated Urea | 0
elevated blood sugar | 0
low hemoglobin | 0
partial dilatation of the ventricles | 0
senile parenchymal atrophy | 0
severe small vessel disease | 0
ground glass patches | 0
consolidation areas | 0
bilateral minimal pleural effusion | 0
SARS-CoV-2 nucleic acid detected | 0
treated based on routine COVID-19 therapy | 0
fever | 24
severe lymphopenia | 24
condition worsened | 24
admitted to the ICU | 72
intubated | 72
decline in respiration | 72
sudden drop in O2sat | 72
lymphopenia corrected | 480
inflammatory biomarkers corrected | 480
O2sat deficiency corrected | 480
respiratory distress corrected | 480
discharged | 624
partial recovery | 624
negative PCR testing | 624
living without any particular problem | 7776