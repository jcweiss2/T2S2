21 years old | 0
pregnant | 0
admitted to Shalkar Medical Center | 0
primigravida | 0
severe PE | 0
intrauterine fetal death (IUFD) | 0
abruptio-placentae | 0
delivered by cesarean section (CS) | 0
placenta totally separated | 0
Couvelaire uterus | 0
atonic postpartum hemorrhage (PPH) | 0
B-Lynch | 0
intravenous carbetocin | 0
tranexamic acid | 0
misoprostol | 0
blood loss during CS and PPH | 0
received fresh frozen plasma | 0
received packed red blood cells (RBCs) | 0
magnesium sulfate (MgSO4) for 24 hours | 0
transferred to West Kazakhstan University (WKU) maternal intensive care unit (ICU) | 0
severe PE complicated by IUFD due to abruptio-placentae and renal failure (anuria) | 0
monitored in WKU-ICU using central venous pressure (CVP) | 0
fluid chart | 0
laboratory investigation | 0
anemic (hemoglobin 7.8 gm/dl) | 0
generalized edema | 0
anuria | 0
160/110 mmHg blood pressure | 0
thrombocytopenia (21 × 1000/mm3 platelet count) | 0
normal coagulation profile | 0
normal bilirubin | 0
normal liver function tests | 0
HELLP syndrome excluded | 0
evidence of hemolysis excluded | 0
elevated total leucocyte count (15.000/mm3) | 0
maternal sepsis excluded | 0
managed by multidisciplinary team approach | 0
correction of anemia using packed RBCs | 0
correction of thrombocytopenia using platelet concentrate | 0
control of blood pressure | 0
renal dialysis | 0
human albumin to correct hypoalbuminemia | 0
laboratory investigations every 3 days | 0
tonic colonic convulsions on the 5th day postpartum | 120
comatosed (11-12 Glasgow coma scale) | 120
brain computerized tomography (CT) showed right partial lobe intracranial hemorrhage (ICH) | 120
carbamazepine for control of convulsions | 120
thrombocytopenia added to final diagnosis | 120
anemia added to final diagnosis | 120
ICH added to final diagnosis | 120
postpartum eclampsia added to final diagnosis | 120
renal failure managed by five sessions of dialysis | 240
urine output normal with normal renal function tests | 240
ICH size decreased and resolved on the 16th postpartum day | 384
discharged from hospital on the 20th postpartum day | 480