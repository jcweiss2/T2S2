44 years old | 0
male | 0
heart transplant | -6720
tacrolimus | -6720
End-Stage Renal Disease (ESRD) | -6720
hemodialysis | -6720
CMV viremia | -168
necrotizing pancreatitis | -168
chills | -96
decreased appetite | -96
worsening non-bloody emesis | -96
dull left upper quadrant abdominal pain | -96
admitted to the hospital | 0
scleral icterus | 0
decreased bibasilar breath sounds | 0
moderate abdominal tenderness | 0
1+ bilateral pedal edema | 0
sinus tachycardia | 0
mild pulmonary edema | 0
WBC 8.3 k/uL | 0
hemoglobin 10.2 g/dL | 0
platelet count 90 k/uL | 0
BUN/creatinine 45/5.8 | 0
elevated high sensitivity troponin level | 0
elevated brain natriuretic peptide (BNP) | 0
elevated AST | 0
elevated ALT | 0
elevated ALP | 0
elevated lipase | 0
elevated total and conjugated bilirubin | 0
reduced left ventricular size | 0
hyperdynamic systolic function | 0
numerous new pulmonary nodules | 0
ring-enhancing lesions within the liver | 0
hyper-enhancement of the pancreas | 0
walled-off necrosis | 0
splenomegaly | 0
positive CMV serologies | 0
absent viral load on PCR | 0
started on broad-spectrum antibiotics | 0
started on vasopressors | 0
elevated CA19-9 levels | 24
liver biopsy | 24
poorly differentiated adenocarcinoma of pancreatic origin | 24
elevated ferritin | 48
elevated triglycerides | 48
elevated fibrinogen | 48
elevated soluble IL-2 R levels | 48
suspected HLH | 48
died | 168