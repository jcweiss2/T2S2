24 years old | 0
female | 0
26 weeks pregnant | 0
admitted to the emergency department | 0
abdominal pain | -120
distension | -120
constipation | -120
preterm delivery | -120
dehydrated | 0
hypotension | 0
tachycardia | 0
tachypnea | 0
asymmetrically distended abdomen | 0
tenderness all over | 0
empty rectum | 0
foetal viability | 0
vaginal examination | 0
threatened preterm labour | 0
labouratory investigations | 0
elevated white cell count | 0
urine analysis | 0
clear | 0
ultrasound scan | 0
distended bowel loop | 0
free fluid in the peritoneal cavity | 0
single viable foetus | 0
clinical diagnosis of IO | 0
abdominal X-ray | 0
dilated large bowel | 0
abnormal gas pattern | 0
coffee bean appearance | 0
sigmoid volvulus | 0
sigmoidoscopy | 0
twisted sigmoid colon | 0
foetal distress | 0
caesarean section | 0
laparotomy | 0
enormously distended sigmoid loop | 0
ischemic and gangrenous changes | 0
necrotic colon | 0
lower segment caesarean section | 0
male preterm infant | 0
mechanical ventilation | 0
lung immaturity | 0
Hartmann’s procedure | 0
end colostomy | 0
closure of the rectal stump | 0
post-operative course | 0
discharged home | 9
reversal of Hartmann’s | 174
colo-rectal anastomosis | 174
sigmoid volvulus in pregnancy | 0
diagnostic challenges | 0
clinical examination | 0
radiological modality | 0
abdominal X-ray | 0
radiation exposure | 0
foetal viability | 0
ultrasound examination | 0
MRI | 0
non-ionizing radiation modality | 0
abdominal pain | 0
gynaecologic emergencies | 0
gynaecological examination | 0
threatened preterm delivery | 0
management of IO | 0
aggressive resuscitation | 0
nasogastric decompression | 0
fluids and electrolytes correction | 0
tocolytics | 0
steroids | 0
surgical intervention | 0
bowel viability | 0
bowel resection | 0
stoma formation | 0
Hartmann’s procedure | 0
primary anastomosis | 0
colonic washout | 0
elective sigmoidectomy | 0
endoscopy | 0
detorsion and decompression | 0
gastroscope | 0
vaginal delivery | 0
obstetric intervention | 0
uterine contamination | 0
puerperal sepsis | 0