58 years old | 0
male | 0
admitted to the hospital | 0
syncope | -2
sore throat | -72
fever | -72
flu-like symptoms | -72
haemoconcentration | -8760
oedema of lower extremities | -8760
myopericarditis | -105120
normotensive | 0
normal heart rate | 0
normal oxygen saturation | 0
sinus rhythm | 0
normal ventricular repolarization | 0
decreased left ventricular ejection fraction | 0
mild concentric remodelling | 0
diffuse mild pericardial effusion | 0
moderate leukocytosis | 0
polyglobulia | 0
decreased serum albumin concentration | 0
mildly increased C-reactive protein | 0
elevated high sensitivity troponin T | 0
elevated NT-pro-B natriuretic peptide | 0
hospitalized for suspected myopericarditis | 0
hypotension | 48
pulmonary oedema | 48
signs of hypoperfusion | 48
cold extremities | 48
oliguria | 48
raise of blood lactates | 48
repeated echocardiography | 48
LVEF of 20% | 48
increased LV wall thickness | 48
restrictive transmitral filling pattern | 48
admitted to ICU | 48
mechanical ventilation | 48
high dosage of vasoactive drugs | 48
coronary angiography | 48
endomyocardial biopsy | 48
active myocarditis | 48
polymerase chain reaction assay | 48
positive for parvovirus B19 | 48
blood cultures | 48
negative blood cultures | 48
mechanical support with intra-aortic balloon pump | 72
pulmonary artery catheter | 72
right heart catheterization | 72
mixed hypovolemic-cardiogenic shock | 72
high doses of i.v. methylprednisolone | 72
diagnosis of SCLS triggered by PVB19 infection | 72
circulatory support | 96
shock persisted | 96
rhabdomyolysis | 96
acute kidney injury | 96
continuous renal replacement therapy | 96
cytokine adsorber haemofilter | 96
improved | 120
LVEF raised to 35% | 120
weaned from IABP | 168
weaned from inotropes and vasopressors | 264
haemofiltration stopped | 168
ventilatory weaning postponed | 168
ventilatory-associated pneumonia | 168
ventilatory weaning accomplished | 288
CMRI performed | 480
improvement of biventricular performance | 480
complete resolution of myocardial oedema | 480
late gadolinium enhancement images | 480
intramyocardial mild, widespread enhancement | 480
pre-discharge echocardiography | 720
restored LVEF of 52% | 720
reduced LV wall thickness | 720
tests for autoimmune diseases | 720
negative tests for autoimmune diseases | 720
further investigations on polyglobulia | 720
excluded JAK 2 mutation | 720
infection and organ failure resolved | 720
discharged | 720
restoration of normal haematocrit values | 720
restoration of renal function | 720
new ISCLS flare | 2160
hypotension | 2160
syncope | 2160
haemoconcentration | 2160
rhinovirus infection | 2160
admitted to ICU | 2160
haemodynamically stable | 2160
myocardial dysfunction did not occur | 2160
prophylactic regimen of intravenous immunoglobulin | 2160
no new syncopal episode | 8760
good clinical condition | 8760
no new SCLS flare | 8760