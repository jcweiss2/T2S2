67 years old | 0
female | 0
rheumatoid arthritis | 0
hydroxychloroquine | -3456
denies diabetes mellitus | 0
denies high blood pressure | 0
denies smoking | 0
denies alcohol consumption | 0
traveled to Italy | -336
returned to Brazil | -336
unverified fever | -336
dry cough | -336
malaise | -336
RT-qPCR test | -336
fever | -336
chills | -336
nausea | -336
admitted to the hospital | 0
COVID-19 diagnosis | 24
chest CT | 24
extensive ground-glass opacities | 24
consolidations | 24
oseltamivir | 24
enoxaparin | 48
respiratory failure | 72
SARS diagnosis | 72
azithromycin | 72
piperacycline with tazobactam | 72
mechanical ventilation | 72
septic shock | 72
pulmonary focus | 72
meropenem | 216
chest CT scan | 696
radiological improvement | 696
hearing loss | 696
discharged from ICU | 720
discharged from hospital | 816
audiometry | 816
isolated hearing loss | 816
tinnitus | 816
corticosteroid therapy | 816
prednisolone | 816
intratympanic applications | 816
dexamethasone | 816
blood pressure increased | 816
normalized blood pressure | 816
brain magnetic resonance imaging | 888
microhemorrhagic lesions | 888
magnetic resonance angiography | 888
no changes | 888
audiometry | 1056
improvement in hearing thresholds | 1056
tinnitus | 1056