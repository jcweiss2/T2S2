60 years old | 0
woman | 0
presented for elective percutaneous nephrolithotomy | 0
right-sided staghorn calculus | 0
pre-diabetes | 0
chronic obstructive pulmonary disease | 0
morbid obesity | 0
body mass index (BMI)=42 | 0
obstructive sleep apnea | 0
heart failure with preserved ejection fraction | 0
febrile (39.2°C) | 24
tachycardic (120–140 beats per minute) | 24
leukocytosis (17.6 x 10^9/L) | 24
vancomycin | 24
piperacillin/tazobactam | 24
meropenem | 24
presumed urosepsis | 24
respiratory distress | 48
hypoxemia refractory to non-invasive positive pressure ventilation | 48
endotracheal intubation | 48
lung protective ventilation (LPV) | 48
postoperative day 2 (POD2) chest X-ray | 48
CT angiogram | 48
bilateral pulmonary ground glass opacities | 48
infectious process | 48
acute respiratory distress syndrome (ARDS) | 48
pulmonary edema | 48
no evidence of pulmonary embolism | 48
transthoracic echocardiogram | 48
normal ejection fraction | 48
normal ventricular size | 48
early paralysis for ventilator desynchrony | 72
refractory hypoxemia | 72
bronchoalveolar lavage samples from POD6 | 144
negative for infectious pathogens | 144
nasopharyngeal swob on POD6 | 144
rhinovirus pneumonia | 144
antibiotics discontinued | 144
no antivirals administered | 144
continued requirement for higher airway pressures | 144
PaO2 to FiO2 ratio of 110 | 144
moderate to severe ARDS | 144
transitioned from LPV to APRV | 144
mechanical ventilation settings adjusted | 144
weaned to extubation on POD9 | 216
discharged home on POD13 | 312
