68 years old | 0
male | 0
carcinoma of pyriform fossa | -672
admitted to ICU | 0
hypoxemic respiratory failure | 0
septic shock | 0
trachea intubated | 0
fluid resuscitation | 0
vasopressor support | 0
7 Fr sized triple lumen central venous catheter inserted | 0
right IJV catheterization | 0
acute renal failure | 24
anuria | 24
metabolic acidosis | 24
HCO3 of 12 mEq/L | 24
hyperkalemia | 24
K + of 6.8 mEq/L | 24
urgent hemodialysis planned | 24
consent for hemodialysis | 24
left IJV chosen for dialysis catheter insertion | 24
patient positioned | 24
head slightly lower than the rest of the body | 24
left side of the neck cleaned | 24
2% w/v chlorhexidine gluconate | 24
draped | 24
local anesthesia | 24
4 ml of 2% lignocaine | 24
IJV located using ultrasound | 24
linear probe | 24
5 MHz frequency | 24
Sonosite Edge II | 24
vein punctured | 24
45° angle | 24
introducer needle | 24
free aspiration of blood | 24
guidewire threaded | 24
resistance felt | 24
guidewire removed | 24
syringe connected to needle hub | 24
free blood aspiration | 24
guidewire reinsertion attempted | 24
resistance felt again | 24
bilateral normal breath sounds | 24
normal respiratory rate | 24
oxygen saturation of 98% | 24
no subcutaneous emphysema | 24
no hematoma | 24
no venous congestion | 24
no limb ischemia | 24
senior ICU registrar called for help | 24
guidewire and needle scanned | 24
loop of guidewire visualized | 24
dual-point echogenicity | 24
introducer needle retracted | 24
guidewire pulled out | 24
loop disappeared | 24
guidewire advanced caudally | 24
dilatation | 24
dialysis catheter railroaded | 24
guidewire removed | 24
correct intraluminal placement confirmed | 24
ultrasonography | 24
blood aspirated | 24
free flow confirmed | 24
bedside chest X-ray | 24
correct placement of hemodialysis catheter | 24
discharged | 48