50 years old | 0
female | 0
admitted to the hospital | 0
history of celiac disease | -672
iron deficiency anemia | -672
hypothyroidism | -672
chronic febrile illness | -24
drenching night sweats | -24
fungal esophagitis | -24
antifungal medication | -24
nausea | -24
normal bowel motion | -24
CT scan | 0
tumor | 0
liver lesions | 0
mild pericardial effusion | 0
echocardiogram | 0
normal ejection fraction | 0
tissue biopsy | 0
GIST | 0
medical oncologist | 0
systemic therapy | 0
imatinib | 24
generalized fatigability | 168
symptomatic anemia | 168
bleeding tumor | 168
transfusions | 168
follow-up CT scan | 168
tumor progression | 168
sunitinib | 168
echocardiography | 168
persistent tachycardia | 168
small pericardial effusion | 168
high ejection fraction | 168
abdominal pain | 192
vomiting | 192
no bowel motion | 192
tachycardia | 192
tachypnea | 192
oxygenation | 192
nasal cannula | 192
abdominal tenderness | 192
guarding | 192
rigid abdomen | 192
lactate level | 192
electrocardiography | 192
sinus tachycardia | 192
CT scan | 192
ischemic changes | 192
jejunal loops | 192
pneumoperitoneum | 192
emergency laparotomy | 216
turbid intraperitoneal fluid | 216
large mass | 216
mid-jejunum | 216
perforation | 216
edematous bowel | 216
mass resection | 216
small bowel resection | 216
side-to-side anastomosis | 216
hypotension | 216
resuscitation | 216
pericardial window | 216
serous fluid | 216
intraoperative | 216
intraperitoneal drains | 216
abdomen closure | 216
extubation | 216
intensive care unit | 216
postoperative monitoring | 216
Regorafenib | 240
Pazopanib | 240
adjuvant chemotherapy | 240
liver metastasis | 240
obstructive phenomena | 240
percutaneous transhepatic cholangiography | 240
deteriorated condition | 240
death | 312
histopathological examination | 312
GIST | 312
mitotic activity rate | 312
safety margins | 312
lymph nodes | 312
negative mesenteric lymph node | 312
CD117 | 312
DOG1 | 312
immunoreactive | 312
anaplastic features | 312
necrosis | 312