73 years old | 0
male | 0
admitted to the hospital | 0
splenomegaly | -672
polycythaemia vera | -672
myelofibrosis | -672
mild valvular heart disease | -672
scheduled for splenectomy | 0
negative real-time PCR test for CoV-2 | 0
splenectomy | 0
exposure to an infected patient | 24
CoV-2 positive | 24
non-severe CoV-2 disease | 24
transferred to the surgical CoV-2 unit | 48
dyspnoea | 72
elevation in D-dimer | 72
chest CT scan | 72
multiple bilobar ground-glass opacities | 72
massive left pleural effusion | 72
left chest tube insertion | 72
improvement of dyspnoea | 96
severe hypotension | 168
massive drop in haemoglobin levels | 168
mild prolongation of prothrombin time | 168
re-surgery | 168
diffuse peritoneal bleeding spots | 168
abdominal lavage | 168
haemostatic patches positioning | 168
admitted to the intensive care unit | 192
extubated | 216
re-posted to the surgical CoV-2 unit | 216
fever | 240
hypoxaemia | 240
high-flow oxygen support | 240
mechanical ventilation | 264
sequential organ failure assessment score | 264
blood cultures | 264
pleural liquid sample | 264
cytomegalovirus DNA | 264
Staphylococcus epidermidis | 264
Bacillus licheniformis | 264
S. hominis | 264
deterioration of general conditions | 312
death | 528
CoV-2 DIC-like syndrome | 168 
thrombosis in the remnant of the splenic vein | 168
large blood collection in the left hypochondrium | 168 
abdomen CT scan | 168 
support with packed red blood cells | 168
support with platelets | 168 
urgent surgical exploration | 168 
no signs of active bleeding | 168 
no signs of pulmonary embolism | 72 
no parameters of multiple organ failure | 168 
no shortness of breath | -672 
no chest pain | -672 
no active bleeding | 168 
no pulmonary embolism | 72 
no multiple organ failure | 168 
no cytomegalovirus DNA | 264 
no improvement of general conditions | 312 
no difference in haemorrhagic or infectious complications | 528 
no specific grant for this research | 528 
next of kin consent obtained | 528 
not commissioned | 528 
externally peer-reviewed | 528