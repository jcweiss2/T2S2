3 years old | 0
female | 0
admitted to the hospital | 0
fever | 0
diarrhea | 0
abdominal pain | 0
severe dehydration | 0
tachypnea | 0
rapid shallow breathing | 0
hypotension | 0
blood pressure 60/40 mmHg | 0
evidence of severe dehydration | 0
purpuric eruption | 0
no organomegaly | 0
no lymphadenopathy | 0
pancytopenia | 0
absolute neutropenia | 0
renal impairment | 0
electrolyte imbalance | 0
hyperuricemia | 0
coagulopathy | 0
disseminated intravascular coagulation | 0
high inflammatory markers | 0
gram-negative Bacilli Escherichia coli | 0
intravenous fluid therapy | 0
blood components transfusion | 0
correction of electrolyte disturbance | 0
antibiotic therapy | 0
provisional diagnosis of acute infectious gastroenteritis | 0
sepsis | 0
severe dehydration | 0
acute renal failure | 0
disseminated intravascular coagulation | 0
pelvi-abdominal ultrasound normal | 0
bone marrow aspirate | 0
hypocellular bone marrow | 0
no abnormal cells | 0
discharged | 336
unexplained irritability | 504
abnormal behavior | 504
hallucinations | 504
failure to recognize parents | 504
vital stability | 504
normal hematological indices | 504
normal coagulation parameters | 504
normal renal panel | 504
normal serum electrolytes | 504
brain imaging studies | 504
magnetic resonance imaging | 504
magnetic resonance arteriography | 504
magnetic resonance venography | 504
thrombosis in left sigmoid and transverse sinuses | 504
workup of thrombophilia | 504
no thrombocytosis | 504
normal coagulation profile | 504
normal protein C and S | 504
antithrombin III | 504
genetic testing for thrombophilia mutations panel | 504
low molecular weight heparin | 504
improved | 504
discharged | 528
follow-up appointment | 528
fever | 672
pallor | 672
abdominal enlargement | 672
leukocytosis | 672
anemia | 672
thrombocytopenia | 672
peripheral smear | 672
many blast cells | 672
abdominal ultrasonography | 672
hepatosplenomegaly | 672
bone marrow examination | 672
hypercellular bone marrow | 672
blast cells | 672
immunophenotyping | 672
positive CD10 | 672
positive CD20 | 672
positive CD79a | 672
diagnosis of Common ALL | 672
induction therapy | 672
consolidation | 672
thrombophilia mutations panel result | 696
positive factor XIII V34L | 696
MTHFR A1298C homozygous mutations | 696
heterozygous positive factor V Leiden mutation | 696
follow-up MRV | 720
complete recanalization of thrombosed sinuses | 720
no new thrombi | 720
complete remission | 720
regular follow-up | 720
no thrombotic events | 720
no leukemia relapses | 720