23 years old | 0
man | 0
presented to hospital | 0
right thigh swelling | -720
draining sinus | -720
skin changes | -720
no history of fever | -720
no systemic symptoms | -720
past medical history unremarkable | -720
no regular medications | -720
non-smoker | -720
denied alcohol use | -720
denied illicit substance use | -720
closed midshaft fracture of the right femur | -43800
motorbike accident | -43800
intramedullary fixation | -43800
surgical site infection | -34560
hardware removed | -34560
two-week course of antibiotics | -34560
migrated to Australia | -720
hemodynamically stable | 0
afebrile | 0
body mass index 19 kg/m² | 0
difficulty gaining weight | 0
weight bearing with minimal pain | 0
right thigh swollen | 0
scaly skin discoloration | 0
draining sinus on posterolateral aspect of distal thigh | 0
neurovascular status intact | 0
preserved tone | 0
preserved power | 0
preserved range of motion | 0
elevated white cell count 11.5 × 10⁹/L | 0
raised CRP 46 mg/L | 0
raised ESR 17 mm/h | 0
normal electrolytes | 0
normal liver function tests |5 0
CT scan demonstrating united right femur fracture | 0
intramuscular collection within vastus intermedius | 0
non-specific bony changes | 0
MRI revealing COM of right femur | 0
extensive intramedullary involvement | 0
extensive cortical involvement | 0
extensive surrounding soft tissue involvement | 0
bone scintigraphy confirming osteomyelitis | 0
confined to right thigh | 0
punch biopsy showing chronic spongiotic tissue reaction | 0
lichen simplex chronicus | 0
ultrasound-guided aspiration of sinus | 0
culture yielding multi-resistant A. xylosoxidans | 0
sinus tract excision | 168
drainage of intramuscular collection | 168
soft tissue samples confirming A. xylosoxidans | 168
bone samples revealing S. aureus co-infection | 168
debridement of medullary canal using RIA technique | 192
systemic sepsis | 192
transferred to ICU | 192
intravenous fluid resuscitation | 192
transfusion of 2 units packed red blood cells | 192
vasopressor support with noradrenaline | 192
hemodynamic stability restored | 192
commenced on intravenous flucloxacillin | 192
commenced on intravenous meropenem | 192
blood cultures positive for methicillin-sensitive S. aureus | 216
repeat blood cultures negative | 264
remained alert | 192
remained oriented | 192
respiring spontaneously on room air | 192
discharged to ward after four days ICU | 432
negative blood cultures | 432
transthoracic echocardiogram excluding infective endocarditis | 432
intravenous antibiotics for one month | 432
transitioned to oral flucloxacillin | 1080
transitioned to oral co-trimoxazole | 1080
asymptomatic after one month oral antibiotics | 1440
weight bearing with no pain | 1440
full ROM in right hip and knee | 1440
intact neurovascular status | 1440
surgical wound healed | 1440
no sign of infection | 1440
hyperpigmentation persisted | 1440
successful weight gain | 1440
intermittent mild gastrointestinal discomfort | 1440
no impact on appetite | 1440
no medical intervention required | 1440
CRP within normal limits at six months | 4320
leukocyte counts within normal limits at six months | 4320
skin changes resolved | 4320
returned to full function | 4320
no pain reported | 4320
CRP within normal limits at one year | 8760
leukocyte counts within normal limits at one year | 8760
no clinical evidence of infection at one year | 8760
follow-up radiograph showing no residual disease | 8760
discharged from services | 8760
