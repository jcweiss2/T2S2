25 years old | 0
female | 0
admitted to the hospital | 0
diabetes | 0
headache | -168
right-side neck pain | -168
shoulder pain | -168
intermittent fever | -48
dry cough | -48
odynophagia | -48
exudative tonsillitis | 0
right-side neck tenderness | 0
WBC count 7.7 | 0
haemoglobin 10.9 | 0
thrombocytopaenia | 0
elevated C reactive protein | 0
toxic granulation on blood film | 0
normal electrolytes | 0
normal BUN | 0
normal creatinine | 0
normal liver function tests | 0
mild direct hyperbilirubinaemia | 0
sinus tachycardia | 0
bilateral infiltrates on chest X-ray | 0
right pleural effusion on repeat chest X-ray | 48
thrombosis of the right internal jugular vein | 0
septic emboli to the lungs | 0
commenced ceftriaxone treatment | 0
transferred to intensive care unit | 24
ventilatory support | 24
meropenem and vancomycin antibiotics | 24
vasopressors | 24
anticoagulated with rivaroxaban | 24
acute kidney injury | 48
rise in creatinine | 48
recovery | 480
discharged | 480
oral anticoagulants | 480
oral antibiotics | 480
insulin therapy | 480