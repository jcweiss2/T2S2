44 years old | 0
    woman | 0
    presented to the hospital emergency room | 0
    severe chest pain | -1
    pain radiating to her back | -1
    pain lasted for an hour | -1
    resolved in the emergency department | -1
    5 months postpartum | -1440
    vaginal delivery | -1440
    recovery period complicated by endometritis | -1440
    endometritis treated with cephalexin | -1440
    endometritis treated with metronidazole | -1440
    hypertension | -1440
    asthma | -1440
    tachycardic | 0
    hemodynamically stable | 0
    blood pressure 142/57 mm Hg | 0
    heart rate 99 beats per minute | 0
    respiration rate 16 breaths per minute | 0
    oxygen saturation 100% | 0
    first heart sound | 0
    second heart sound | 0
    no aortic regurgitation murmur | 0
    normal complete blood count | 0
    normal kidney function | 0
    normal electrolytes | 0
    D-dimer negative | 0
    elevated high-sensitivity troponin levels | 0
    electrocardiogram showed sinus tachycardia | 0
    no ST-segment changes | 0
    chest radiograph unremarkable | 0
    computed tomography chest revealed splenic aneurysm | 0
    splenic infarct | 0
    pulmonary edema | 0
    dilated pulmonary arteries | 0
    no acute aortic dissection | 0
    computed tomography angiogram ruled out aortic dissection | 0
    D-dimer ruled out pulmonary embolism | 0
    rising troponin levels | 0
    non-ST segment elevation myocardial infarction considered | 0
    recent stress due to daughter's illness | -1440
    recent stress due to financial strains | -1440
    differential diagnosis acute coronary syndrome | 0
    differential diagnosis stress-induced cardiomyopathy | 0
    differential diagnosis peripartum cardiomyopathy | 0
    differential diagnosis spontaneous coronary artery dissection | 0
    treated for acute coronary syndrome | 0
    transthoracic echocardiogram demonstrated masses on aortic valve | 0
    vegetation on right coronary cusp | 0
    vegetation on noncoronary cusp | 0
    severe aortic regurgitation | 0
    pan-diastolic flow reversal | 0
    mildly dilated left ventricle | 0
    moderate eccentric hypertrophy | 0
    dilated atria | 0
    elevated atrial pressure | 0
    moderate mitral regurgitation | 0
    mild pulmonary hypertension suspected | 0
    coronary angiography showed left main lesion | 0
    no angiographic coronary artery disease | 0
    assessed by cardiac surgeon | 0
    accepted for emergent operative intervention | 0
    vegetation at left coronary artery ostium | 0
    vegetation removed | 0
    infected aortic valve removed | 0
    annulus debrided | 0
    aortic root enlarged | 0
    mechanical prosthesis replacement | 0
    transferred to intensive care unit | 0
    sent to ward on postoperative day 5 | 120
    repeat angiography confirmed lesion removal | 120
    culture results negative | 120
    antibiotics continued | 120
    discharged home | 240
    intravenous vancomycin | 240
    intravenous ceftriaxone | 240
    follow-up with cardiac surgery | 240
    follow-up with infectious diseases | 240
    echocardiogram ordered in 6 weeks | 1008
    no traditional risk factors for IE | 0
    no fever | 0
    postpartum endometritis history | -1440
    aspiration of septic emboli during surgery | 0
    no distal vascular embolization | 0
    mechanical valve deployed | 0
    risks of future pregnancies discussed | 0
    contraceptive plans discussed | 0