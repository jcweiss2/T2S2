13 years old | 0
    male | 0
    electric burn over the right arm | -120
    electric burn over the right axilla | -120
    electric burn over the right-sided thoracic and abdominal region | -120
    post-burn contracture release | 0
    restriction of routine activity | 0
    electric burns over the right arm in 2013 | -120
    electric burns over the right axillary region in 2013 | -120
    electric burns over the right and left foot in 2013 | -120
    debridement of burnt area | -120
    amputation of the right great toe | -120
    amputation of the 4th and 5th toes of the left foot | -120
    skin grafting in 2013 | -120
    operated in June 2014 | -1464
    operated in June 2015 | -2928
    difficulty in extension of arm | -2928
    contracture release of right axillary region | -1464
    skin grafting in June 2014 | -1464
    restriction of movements | -120
    hospitalized for 1 month in 2013 | -120
    admitted for 15 days during subsequent surgeries | -1464
    received multiple blood transfusions | -1464
    vegetarian diet | 0
    weight loss of 2 kg over the last three months | 0
    reduced appetite | 0
    felt tired all the time | 0
    felt weaker | 0
    wounds taking a long time to heal | 0
    poor concentration | 0
    feeling cold most of the time | 0
    BMI of 12.9 | 0
    underweight | 0
    chest X-ray normal | 0
    electrocardiogram normal | 0
    informed consent from guardian | 0
    preoperative vitals: heart rate 94/min | 0
    preoperative vitals: BP 104/62 mm Hg | 0
    preoperative vitals: SpO2 98% | 0
    premedicated with glycopyrrolate | 0
    premedicated with ondansetron | 0
    premedicated with midazolam | 0
    premedicated with fentanyl | 0
    preoxygenated with 100% oxygen | 0
    anesthesia induced with propofol | 0
    anesthesia induced with atracurium | 0
    intubated with cuffed ET tube | 0
    anesthesia maintained with sevoflurane | 0
    anesthesia maintained with O2:N2O | 0
    intraoperative monitoring | 0
    intraoperative tachycardia | 0
    intraoperative hypotension | 0
    SpO2 dropped to 84% | 0
    pink frothy secretions in ET tube | 0
    bilateral crepitations on auscultation | 0
    procedure stopped | 0
    FiO2 increased to 100% | 0
    furosemide administered | 0
    positive pressure ventilation | 0
    deeper plane of anesthesia | 0
    atracurium administered | 0
    noradrenaline infusion | 0
    arterial blood gas analysis | 0
    hypoxia | 0
    decreased PaO2/FiO2 ratio | 0
    lactate level 4.5 mmol/l | 0
    saturation became 100% | 0
    BP 90/50 mm Hg | 0
    heart rate decreased to 130 beats/min | 0
    surgery completed | 0
    spontaneous respiratory attempts | 24
    reversed with neostigmine | 24
    reversed with glycopyrrolate | 24
    extubated | 24
    O2 support 6 L/min | 24
    shifted to ICU | 24
    bedside transthoracic 2D echo | 24
    LVEF 20% | 24
    global LV hypokinesia | 24
    dilated LV | 24
    mild MR/TR | 24
    acute decompensated heart failure due to thiamine deficiency | 24
    thiamine infusion started | 24
    carvedilol administered | 24
    spironolactone + furosemide administered | 24
    enalapril administered | 24
    chest X-ray showed pulmonary edema | 24
    IV fluid restricted | 24
    urine output measured hourly | 24
    vasopressor requirement decreased | 72
    vasopressor stopped | 24
    oxygen requirement decreased | 72
    repeat ABGA improved PaO2/FiO2 ratio | 72
    air entry equal and clear | 72
    repeat 2D echo after four days | 168
    LVEF 50% | 168
    fair LV function | 168
    normal-sized cardiac chambers | 168
    no MR/TR | 168
    discharged after seven days | 168
    follow up after six weeks | 168
    thiamine rich diet advised | 168
    weight loss guided nutritional assessment | 0
    vitamin B1 deficiency suspected | 0
    Shoshin beriberi diagnosis | 0
    pulmonary edema confirmed | 24
    hypovolemia excluded | 0
    fluid overload excluded | 0
    blood transfusion-related complications excluded | 0
    pulmonary embolism excluded | 0
    anemia-induced heart failure excluded | 0
    lighter planes of anesthesia excluded | 0
    hypoxia-induced heart failure excluded | 0
    multivitamin deficiency considered | 0
    blood transfusion reaction excluded | 0
    severe sepsis considered | 0
    burns considered | 0
    unexplained heart failure considered | 0
    lactic acidosis considered | 0
    neurological disorder considered | 0
    alcoholism considered | 0
    starvation considered | 0
    chronic malnutrition considered | 0
    long-term parenteral feeding considered | 0
    hyperemesis gravidarum considered | 0
    bariatric surgery considered | 0
    thiamine deficiency confirmed | 24
    financial support nil | 0
    no conflicts of interest | 0
    