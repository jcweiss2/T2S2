67 years old | 0
    African American | 0
    woman | 0
    obesity | 0
    body mass index 38 kg/m2 | 0
    chronic active smoker | 0
    chronic obstructive pulmonary disease | 0
    obstructive sleep apnea | 0
    continuous positive airway pressure therapy | 0
    severe pulmonary hypertension | 0
    atrial fibrillation | 0
    anticoagulation | 0
    well-controlled type 2 diabetes | 0
    hypertension | 0
    dyslipidemia | 0
    discharged to rehabilitation facility | -672
    hypercapnic hypoxic respiratory failure | -672
    mechanical ventilation | -672
    sudden-onset generalized weakness | 0
    light-headedness | 0
    shortness of breath | 0
    dry cough | 0
    discharged from rehabilitation center | -24
    physical therapy/hydrotherapy sessions | -24
    distress | 0
    denied subjective fevers | 0
    denied chills | 0
    denied headache | 0
    denied photophobia | 0
    denied sputum production |0
    denied nausea |0
    denied vomiting |0
    denied diarrhea |0
    denied dysuria |0
    denied vaginal discharge |0
    denied recent travel |0
    denied exposure to pets |0
    simvastatin |0
    metformin |0
    glipizide |0
    valsartan |0
    labetalol |0
    diltiazem |0
    warfarin |0
    fluticasone/salmeterol |0
    albuterol |0
    hypotension |0
    epinephrine drip |0
    tachypnea |0
    O2 saturation 78% |0
    2 liters per nasal cannula |0
    91% on biphasic positive airway pressure |0
    pulse 110/min |0
    temperature 98.9°F |0
    alert |0
    oriented to person |0
    oriented to place |0
    oriented to time |0
    conjunctival pallor |0
    dry mucous membranes |0
    arrhythmic heart sounds |0
    2/6 pansystolic tricuspid murmur |0
    bilateral crackles at bases |0
    wheezing |0
    nontender abdomen |0
    ascetic wave |0
    2+ edema in lower extremities |0
    decreased peripheral pulses |0
    no evidence of skin ulcers |0
    no meningeal signs |0
    no focal deficits |0
    empiric therapy cefepime |0
    empiric therapy vancomycin |0
    leukocyte count 15.6 cells/mL |0
    neutrophils 85% |0
    no bandemia |0
    platelets 877000/mL |0
    acute kidney injury |0
    creatinine 1.3 mg/dL |0
    hyperglycemia 183 mg/dL |0
    lactate level 3 mmol/L |0
    international normalized ratio 3 |0
    HIV test negative |0
    urinalysis negative for blood |0
    urinalysis negative for nitrates |0
    urinalysis negative for leukocyte esterase |0
    5 to 10 white blood cells |0
    many bacteria |0
    right pleural effusion |0
    right-sided atelectasis |0
    cardiomegaly |0
    moderate ascites |0
    enlarged caliber hepatic veins |0
    ejection fraction 60% |0
    severe pulmonary hypertension |0
    severe tricuspid regurgitation |0
    mild mitral regurgitation |0
    no signs of endocarditis |0
    cytology negative for malignant cells |0
    blood culture samples |0
    urine culture samples |0
    pleural fluid culture samples |0
    peritoneal fluid culture samples |0
    no longer required vasopressors |24
    two sets of blood culture Gram-negative bacilli |24
    vancomycin discontinued |24
    final identification blood cultures Sphingobacterium multivorum |96
    resistant to ceftazidime |96
    resistant to trimethoprim/sulfamethoxazole |96
    intermediate susceptibility meropenem |96
    intermediate susceptibility piperacillin/tazobactam |96
    cefepime switched to ciprofloxacin |96
    gram stain urine not reported |96
    urine culture negative |96
    peritoneal fluid cultures negative |96
    pleural fluid cultures negative |96
    clinically stable for discharge |96
    total 10 days ciprofloxacin |96
    repeated blood cultures negative |120
    repeated urine cultures negative |120
    followed up 2 weeks after discharge |672
    followed up 4 weeks after discharge |1344
    clinically stable |672
    clinically stable |1344
<|eot_id|>
