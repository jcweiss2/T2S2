73 years old | 0
male | 0
admitted to the hospital | 0
altered mental status | -168
decreased appetite | -168
poor oral intake | -168
hepatocellular carcinoma | -6720
history of alcohol use | -8760
congestive heart failure | -8760
coronary artery disease | -8760
chronic kidney disease | -8760
history of alcohol abuse | -72000
cigarette smoking | -144000
stopped alcohol abuse | -720
stopped cigarette smoking | -1440
afebrile | 0
hypotensive | 0
hypoxic | 0
mild tenderness in right upper quadrant | 0
shock | 0
admitted to intensive care unit | 0
hemodynamic support | 0
mildly elevated liver transaminases | 0
blood cultures obtained | 0
empiric antibiotic therapy with vancomycin | 0
empiric antibiotic therapy with cefepime | 0
empiric antibiotic therapy with metronidazole | 0
chest X-ray unremarkable | 0
urinalysis unremarkable | 0
CT of abdomen | 0
interval increase in intrahepatic metastatic disease | 0
multiple new and enlarging metastases | 0
diagnosed with hepatocellular carcinoma | -672
imaging at diagnosis | -672
well-defined solid-appearing mass in left liver lobe | -672
biopsy | -672
moderately differentiated hepatocellular carcinoma | -672
transarterial chemoembolization (TACE) | -672
second TACE procedure | -112
post-procedure admission for chest pain | -112
post-procedure admission for sepsis | -112
CT abdomen | -112
embolized left hepatic mass | -112
ill-defined hypodensities in left liver | -112
hepatic infarcts | -112
abdominal CT | 0
multiple new and enlarging masses | 0
liver abscesses | 0
blood cultures grew Raoultella planticola | 24
intermediate sensitivity to ampicillin | 24
sensitive to cephalosporins | 24
sensitive to quinolones | 24
antibiotics narrowed to ceftriaxone | 24
antibiotics narrowed to metronidazole | 24
two drains placed by Interventional Radiology | 96
fluid revealing elevated white blood cells | 96
no growth on culture | 96
repeat imaging showed decrease in size of masses | 120
overall clinical status significantly improved | 120
discharged on IV ceftriaxone | 168
discharged on oral metronidazole | 168
re-admitted | 672
progressively worsening lesions | 672
overall decompensation | 672
pursued a more comfort-based approach | 696
expired | 720