57 years old | 0
male | 0
presented with 4-day history of increasing breathlessness | -96
presented with 4-day history of abdominal discomfort | -96
40-pack year smoking history | 0
no regular medications | 0
febrile (temperature 39°C) | 0
tachycardic (heart rate 120 beats/min) | 0
lactate of 4 mmol/l | 0
underwent surveillance colonoscopy with biopsy of splenic flexure polyp | -120
histology was benign | -120
diverticular disease noted | -120
admitted | 0
possible abdominal perforation | 0
sepsis | 0
suddenly deteriorated | 24
developed painful cold legs | 24
became hypotensive (blood pressure 70/50 mmHg) | 24
agitated | 24
sweaty | 24
peripheral mottling | 24
massive hepatomegaly | 24
arterial blood gas demonstrated lactate of 14 mmol/l | 24
marked hypoglycaemia (glucose 0.8 mmol/l) | 24
resuscitated with crystalloid | 24
resuscitated with dextrose | 24
transferred to ICU | 24
colonic perforation was unlikely | 24
no clinical finding of peritonism | 24
cardiac arrest in ICU | 24
pulseless electrical activity | 24
intubated | 24
required 2 min of CPR | 24
return of spontaneous circulation | 24
central venous catheter inserted | 24
right internal jugular vein large and non-compressible | 24
central venous pressure 31 mmHg | 24
INR 5.9 | 24
fibrinogen 0.2 g/l | 24
platelets 38×10^9/l | 24
transthoracic echo performed | 24
massive pericardial effusion | 24
right ventricular collapse | 24
electrocardiogram (ECG) showed electrical alternans | 0
chest X-ray showed enlarged heart shadow | 0
pericardial effusion drained | 24
700 ml of fluid aspirated | 24
stabilized haemodynamically | 24
pericardial fluid heavily blood stained | 24
possible type A dissection | 24
possible metastatic bowel cancer | 24
CT of chest, abdomen, and pelvis performed | 24
CT aortogram performed | 24
CT showed haematoma in distal arch of aorta | 24
CT showed haematoma in descending aorta | 24
CT angiography images poor quality | 24
CT angiogram repeated | 36
two transoesophageal echocardiograms performed | 48
type A dissection excluded | 48
case management discussion | 48
dissection manageable medically | 48
serial echocardiograms performed | 168
moderate recurrence of pericardial effusion | 168
no significant haemodynamic compromise | 168
developed paraplegia | 168
pleural effusion evolved | 168
pleural effusion drained | 168
pleural fluid consistent with metastatic adenocarcinoma | 168
suspicious spiculate lesion in left upper lobe | 168
died | 1440
no post mortem | 1440
symptomatic pericardial effusion related to lung cancer | 0
acute type B aortic dissection | 0
