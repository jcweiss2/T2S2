66 years old | 0
male | 0
admitted to the hospital | 0
SARS-CoV-2 infection | -1440
septic shock | -1440
hemodynamic instability | -1440
orotracheal intubation | -1344
pulmonary insufficiency | -1344
renal failure | -1344
arterial hypertension | -6720
moderate alcoholism | -6720
coronary disease | -6720
placement of 2 stents | -6720
Dieulafoy gastric lesion | 0
esophageal ulcers | 0
cytomegalovirus (CMV) infection | 0
hepatomegaly | 0
no bile duct dilatation | 0
blood transfusions | 0
antibiotics | 0
corticosteroids | 0
ganciclovir | 0
pulmonary function improvement | 24
acute kidney injury | 0
hemodialysis | 0
cholestatic enzymes increase | 504
metabolic and genetic markers negative | 504
antibodies against autoimmune hepatic diseases negative | 504
serologies negative | 504
PCRs for hepatotropic and non-hepatotropic viruses negative | 504
serum immunoglobulin IgG normal | 504
serum immunoglobulin IgA normal | 504
serum immunoglobulin IgM normal | 504
gamma globulin levels normal | 504
magnetic resonance cholangiopancreatography (MRCP) | 504
diffuse irregularity of the intra-and extrahepatic bile ducts | 504
multiple focal strictures | 504
mild focal dilations of the biliary tree | 504
sclerosing cholangiopathy | 504
transjugular liver biopsy | 504
biliary cast | 504
hematic thrombus | 504
retrograde chol-angiography | 504
serum ammonia >250 | 504
neurological symptoms | 504
continuous hemo-dialysis | 504
sodium benzoate | 504
ursodeoxycholic acid | 504
corticosteroids | 504
serum ammonia decrease | 528
neurological function partial recovery | 528
liver function deterioration | 528
liver transplantation not performed | 528
liver biopsy | 504
prominent bile ductular reaction | 504
cholangiocyte injury | 504
inflammatory infiltrate rich in neutrophils | 504
biliary infarctions | 504
marked cholestasis | 504
portal fibrosis | 504
degenerative cholangiocyte injury | 504
extreme cholangiocyte cytoplasmic vacuolization | 504
bile ductular proliferation | 504
neutrophils | 504
discharged | 2880