51 years old | 0
male | 0
history of severe alcoholism | 0
high daily consumption of alcohol over 30 years | -262800
consumed rum | -262800
consumed cognac | -262800
consumed wines | -262800
refused to treat his addiction | 0
decrease in short-term memory | -8760
complained of paresthesias of lower limbs | -8760
complained of paresthesias of upper limbs | -8760
ingestion of large amounts of alcohol | -24
excessive drowsiness | -24
torpor | -24
coma | -24
Glasgow coma score 7 | 0
no signs of meningeal irritation | 0
no focal deficits | 0
no cranial nerve abnormalities | 0
IV thiamine 500 mg/day | 0
high doses of parenteral B vitamins | 0
hypodensity in corpus callosum on CT | 0
MRI involvement of cortical regions | 0
MRI involvement of subcortical white matter of both frontal lobes | 0
MRI involvement of post-central gyri | 0
MRI involvement of superior temporal gyri | 0
no signs of disruption of blood-brain barrier | 0
mild improvement in level of consciousness | 168
Glasgow coma score 10 | 168
mechanical ventilatory support | 168
multiple pulmonary infectious complications | 168
respiratory insufficiency dependent on mechanical ventilation | 168
tracheostomy | 168
sepsis | 1680
fever | 1680
worsening of respiratory status | 1680
hemodynamic condition deteriorated over 24 hours | 1680
vasoactive drugs | 1680
broad-spectrum IV antibiotics | 1680
cultures of blood | 1680
cultures of tracheal secretions | 1680
Rhodotorula mucilaginosa infection | 1680
amphotericin B treatment | 1680
no significant response to amphotericin B | 1680
septic shock | 1680
death | 1680
