25 years old | 0
female | 0
autoimmune hepatitis | -672
acetaminophen | -672
ibuprofen | -672
azathioprine | -672
prednisone | -672
unprotected sexual intercourse | -336
fever | -72
chills | -72
nausea | -72
dizziness | -72
heavy menorrhagia | -72
bilateral lower extremity pain | -72
edema | -72
ascites | -72
influenza vaccination | -672
COVID-19 vaccination | -672
admitted to the hospital | 0
hemodynamically unstable | 0
blood pressure 67/39 mmHg | 0
heart rate 129 beats per minute | 0
respirations 33 per minute | 0
temperature 35.1 degrees Celsius | 0
jaundice | 0
scleral icterus | 0
abdominal ascites with fluid wave | 0
anasarca | 0
erythematous vaginal vault | 0
minimal discharge | 0
no vesicles | 0
no lesions | 0
no retained foreign objects | 0
fine reticular violaceous patches | 0
lactic acidosis | 0
lactic acid 13.1 mmol/L | 0
creatinine 1.49 mg/dL | 0
aspartate transaminase 56 units/L | 0
alanine transaminase 62 units/L | 0
total bilirubin 3.7 mg/dL | 0
direct bilirubin 3.19 mg/dL | 0
alkaline phosphatase 213 units/L | 0
total protein 5.3 g/dL | 0
albumin 1.4 g/dL | 0
hemoglobin 5.2 g/dL | 0
leukocytes 1.3 k/uL | 0
platelets 90 k/uL | 0
prothrombin time 37.9 s | 0
international normalized ratio 3.9 | 0
beta-human chorionic gonadotropin test negative | 0
occasional schistocytes | 0
paracentesis | 0
peritoneal fluid analysis | 0
leukocyte count 9821 | 0
neutrophilic predominance | 0
CT angiography | 0
cirrhosis | 0
portal hypertension | 0
large volume abdominal ascites | 0
splenomegaly | 0
generalized edematous wall thickening | 0
intubation | 0
labored breathing | 0
tachypnea | 0
intravenous fluids | 0
blood products | 0
vasopressors | 0
broad-spectrum antibiotic therapy | 0
vancomycin | 0
piperacillin-tazobactam | 0
doxycycline | 0
clindamycin | 0
intravenous immunoglobulin | 0
large violaceous non-blanching ecchymoses | 16
flaccid bullae | 16
dusky and violaceous skin | 36
bullae | 36
lactate dehydrogenase 298 units/L | 36
fibrinogen 187 mg/dL | 36
D-dimer > 20 mcg/mL | 36
urinalysis | 36
salicylate level negative | 36
acetaminophen level negative | 36
Chlamydia trachomatis negative | 36
Neisseria gonorrhea negative | 36
urine toxicology screen negative | 36
peritoneal fluid culture negative | 36
blood culture positive for Streptococcus pneumoniae | 36
progressive hypoxia | 48
shock | 48
death | 48
autopsy | 48
cirrhotic liver | 48
diffuse alveolar damage | 48
serous fluid in abdominal compartment | 48