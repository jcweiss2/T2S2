71 years old | 0
male | 0
admitted to the hospital | 0
productive cough | -168
fever | -168
endoscopic removal of a fish bone | -168
symptoms suggestive of mediastinitis | -168
no mucosal defect found | -168
conservatively managed with nothing by mouth | -168
antibiotics | -168
productive cough progressed | -24
fever progressed | -24
chest computed tomography (CT) scan | -24
wide esophageal perforation | -24
mediastinal abscess | -24
right pleural empyema | -24
blood pressure was steady | 0
tachypneic | 0
gastrografin esophagogram | 0
perforation in the middle thoracic esophagus | 0
aspiration pneumonia progressed | 24
history of traumatic hemothorax | -720
pleural drainage for empyema | -720
calcified pleural lesions | 0
posterior mediastinal drainage | 48
Barovac PS400L | 48
incision on the left side of the neck | 48
drainage seemed insufficient | 72
esophageal endoscopy | 72
multiple sites of wall injuries | 72
perforation site | 72
laceration | 72
Levin tubes inserted | 72
internal mediastinal drainage | 72
gastric drainage | 72
Stenotrophomonas maltophilia identified | 72
antibiotic regimen adjusted | 72
continuous suction | 72
internal mediastinal drainage improved | 120
gastric drainage improved | 120
jejunostomy | 216
gastrostomy | 216
sufficient nutritional support | 216
extubated | 264
moved to the general ward | 432
suction turned off | 456
natural drainage started | 456
microbiologic culture | 312
no pathologic microorganism | 312
Levin tube removed | 600
follow-up endoscopic examination | 624
injury sites nearly healed | 624
defect | 624
follow-up chest CT scan | 696
notable decrease in the extent of the mediastinal abscess | 696
follow-up esophagogram | 936
no evidence of leakage | 936
oral diet started | 936
discharged | 1104
follow-up esophagogram | 3024
no abnormal findings | 3024
endoscopic examination | 3024
esophageal injury completely healed | 3024