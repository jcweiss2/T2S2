32 years old | 0
female | 0
Raynaud's phenomenon | -672
recurrent urinary tract infection (UTI) | -672
UTI symptoms | -120
shortness of breath | -48
hypotensive | 0
altered | 0
pressors | 0
broad spectrum antibiotics | 0
vancomycin | 0
cefepime | 0
metronidazole | 0
E. coli bacteremia | 0
enterobacter | 0
anemia | 0
thrombocytopenia | 0
coagulopathy | 0
transfusion of 3 units of platelets | 0
transfusion of 2 units of red blood cells | 0
transfusion of fresh frozen plasma | 0
hyponatremic | 0
sodium of 117 mmol/L | 0
brain MRI | 0
lumbar puncture | 0
unremarkable brain MRI | 0
unremarkable lumbar puncture | 0
acute respiratory distress | 24
intubation | 24
elevated creatinine | 24
creatinine of 6.4 mg/dL | 24
urinalysis | 24
3+ blood | 24
3+ leukocytes | 24
3+ protein | 24
4+ bacteria | 24
continuous renal replacement therapy | 24
improvement in renal function | 48
CT of the abdomen and pelvis | 48
enlarged kidneys | 48
hepatosplenomegaly | 48
persistent agitation | 72
transfer to the medical intensive care unit | 72
anemic | 72
thrombocytopenic | 72
hemoglobin of 7.6 g/dL | 72
platelet count of 15,000 k/cu mm | 72
leukocytosis | 72
white blood cell count of 30.78k/cu mm | 72
anion gap metabolic acidosis | 72
bicarbonate of 20 mmol/L | 72
anion gap of 18 | 72
elevated lactate | 72
lactate of 5.6 mmol/L | 72
hyponatremic | 72
sodium of 128 mmol/L | 72
elevated creatinine | 72
creatinine of 1.8 mg/dL | 72
differential considerations | 72
infiltrative diseases | 72
idiopathic Castleman disease | 72
malignancy | 72
IgG4-related disease | 72
granulomatous disease | 72
repeat CT of the abdomen and pelvis | 96
bilateral nephromegaly | 96
heterogeneous renal parenchymal enhancement | 96
loss of corticomedullary differentiation | 96
focal wedge-shaped hypodensities | 96
superimposed necrosis | 96
cinematic rendering | 96
3D renderings | 96
multifocal renal abscesses | 96
infiltrative bilateral renal disease | 96
glomerulonephritis | 96
lymphoma | 96
renal cell carcinoma | 96
renal biopsy | 120
diffuse infiltration by histiocytic cells | 120
focal abscesses | 120
Gram stain | 120
Gram Weigert stains | 120
Von Kossa stain | 120
Michaelis-Gutman bodies | 120
immunostain for CD163 | 120
infiltration of macrophages or histiocytes | 120
diagnosis of pyelonephritis | 120
focal micro-abscesses | 120
malakoplakia | 120
ultrasound imaging | 120
left greater than right nephromegaly | 120
multiple renal abscesses | 120
MRI | 144
bilateral nephromegaly | 144
intrarenal and perinephric fluid collections | 144
mild left hydronephrosis | 144
thickening of the left renal pelvis | 144
thickening of the left perinephric fascia | 144
extension to the retroperitoneal soft tissues | 144
tigecycline | 144
ceftriaxone | 144
bethanechol | 144
vitamin C | 144
minocycline | 168
liver biopsy | 168
no evidence of hepatic malakoplakia | 168
nephrectomy | 168
normal creatinine | 192
leukocytosis | 192
low-grade fevers | 192
progression of the disease | 192
extension to the left perinephric space | 192
extension to the retroperitoneum | 192
radical left nephrectomy | 216