35 years old | 0 | 0 
female | 0 | 0 
gave birth to healthy twins | -24 | -24 
in vitro fertilization | -280 | -280 
facial nerve paresis | -672 | 0 
severe headache | 24 | 24 
generalized tonic–clonic seizures | 24 | 26 
loss of consciousness | 24 | 26 
arterial blood pressure 195/110 mmHg | 24 | 24 
heart rate 120 beats/min | 24 | 24 
eclampsia | 24 | 24 
antihypertensive therapy | 24 | 120 
intravenous infusion of magnesium sulphate | 24 | 24 
ebrantil | 24 | 24 
20% manitol | 24 | 24 
diazepam | 24 | 24 
bilateral vision loss | 48 | 48 
proteinuria 2+ | 48 | 48 
cortical blindness | 48 | 48 
mild right-sided facial nerve paresis | 48 | 120 
hypodensity of the posterior white matter | 72 | 72 
vasogenic edema | 72 | 72 
T2- and fluid-attenuated inversion recovery-weighted images | 72 | 72 
hyperintense signals in the white matter | 72 | 72 
parietal and occipital regions | 72 | 72 
junctions of vascular watershed zones of the brain | 72 | 72 
stabilization of the general condition | 120 | 120 
oral antihypertensive medication | 120 | 216 
enalapril maleate | 120 | 216 
methyldopa | 120 | 216 
human albumin | 120 | 120 
normalization of the concentration of proteins in the plasma | 120 | 120 
bilateral improvement of the visual function | 168 | 168 
best-corrected visual acuity 1.0 | 168 | 168 
peripheral relative scotoma | 168 | 168 
depressed sensitivity of the paracentral left visual field | 168 | 168 
regression of the edema | 216 | 216 
discrete residual changes over the posterior horns of the side ventricles | 216 | 216 
discharge from the clinic | 216 | 216 
physical therapy for the paresis of the facial nerve | 216 | 504 
oral antihypertensive therapy | 216 | 504 
enalapril | 216 | 504