65 years old | 0
female | 0
admitted to the hospital | 0
nausea | -24
vomiting | -24
loss of appetite | -8760
weight loss | -8760
open cholecystectomy | -258384
cure for eventration | -262080
midline vertical scar | 0
extrinsic compression of the lesser curvature | 0
erythematous mucosa | 0
mixed dense lymphoid infiltrate | 0
heterogeneous formation | 0
disappearance of the separation border | 0
multiple parietal and central calcifications | 0
CA 19-9 slightly raised | 0
ACE normal | 0
irregular contour mass | 0
segment 3 of liver | 0
release of the mass from the duodenum | 0
biopsies of the duodenal edges | 0
atypical segmental hepatectomy | 0
kellyclasia | 0
surgical sponge | 0
necrotic textiloma | 0
extubated | 6
respiratory distress | 72
thoraco-abdominal CT | 72
lesion related to infection lung | 72
transferred to intensive care unit | 72
intubated | 72
ventilated | 72
hypotension | 72
tachycardia | 72
died | 240
unrecovered cardio-respiratory arrest | 240
resuscitation measures | 240
