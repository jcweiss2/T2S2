83 years old|0
    female|0
    presented to the emergency department|0
    accident involving her wheelchair|0
    subcutaneous abscess located on her abdomen|0
    flung from her wheelchair|0
    fully immobilized|0
    on a backboard|0
    taken off the backboard|0
    passing Nexus criteria for cervical spine immobilization|0
    no complaints of pain other than in her left lower quadrant|0
    full physical examination|0
    blood pressure of 124/59|0
    heart rate of 107|0
    respiratory rate of 18|0
    temperature of 97.5°F|0
    pulse oximetry of 95% on room air|0
    lungs clear bilaterally in all fields|0
    cardiac auscultation found normal S1 and S2|0
    no murmurs|0
    no gallops|0
    no rubs|0
    bowel sounds in all 4 quadrants|0
    pain elicited upon palpation of her left lower quadrant|0
    18 × 8-cm subcutaneous abscess|0
    fluctuant abscess|0
    central area of black necrotic skin measuring 8 × 3 cm|0
    oozing centrally|0
    Parkinson disease|0
    dementia|0
    primary historian|0
    noticed the mass in the previous 2 days|-48
    central black necrosis present since the previous day|-24
    complaining of increasing pain over the past few days|-72
    pain worsened with bowel movements|-72
    history of gastroesophageal reflux|0
    hypertension|0
    hypothyroidism|0
    renal failure|0
    pulmonary hypertension|0
    diastolic heart failure|0
    recently hospitalized for acute diverticulitis with perforation|0
    treated medically|0
    ordered complete blood count|0
    ordered basic metabolic panel|0
    ordered urinalysis|0
    ordered abdominal computed tomography with IV contrast|0
    surgical consult|0
    white blood cell count of 27.9 × 1,000/uL|0
    hemoglobin of 9.4 g/dL|0
    hematocrit of 27.6%|0
    platelet count of 446|0
    serum sodium of 134 mmol/L|0
    potassium of 3.4 mmol/L|0
    blood urea nitrogen of 23 mg/dL|0
    creatinine of 1.1 mg/dL|0
    urinalysis positive for nitrites|0
    microscopy showing 1+ leukocytes|0
    microscopy showing 4+ bacteria|0
    CT revealed inflamed colon|0
    fistulous tract winding into the left lower quadrant|0
    large subcutaneous abscess|0
    inflammatory changes|0
    pockets of gas|0
    subcutaneous air|0
    history indicative of necrotizing fasciitis|0
    physical examination indicative of necrotizing fasciitis|0
    laboratory findings indicative of necrotizing fasciitis|0
    CT findings indicative of necrotizing fasciitis|0
    surgical consultant evaluation|0
    agreement with findings of possible necrotizing infectious process|0
    given broad-spectrum antibiotics|0
    given IV fluids|0
    presurgical laboratory tests performed|0
    admitted to the ICU|0
    underwent surgical intervention|0
    debridement of pus and fluid|0
    mixed anaerobic infection|0
    complete survey of the abscess|0
    numerous areas of necrosis within the subcutaneous fat|0
    small opening at the base of the abscess|0
    emanated pus from the abdominal cavity|0
    enlarged for further examination|0
    distal right sigmoid colon inflamed|0
    tiny microperforation found|0
    examination of the rest of the large bowel|0
    no other signs of infection|0
    sigmoid microperforation ruled the source|0
    underwent sigmoid resection|0
    placement of a diverting colostomy|0
    wound vacuum placement|0
    wound site cultured during surgery|0
    grew Proteus mirabilis|0
    grew Escherichia coli|0
    grew E faecalis|0
    grew Bacillus fragilis|0
    grew coagulase-negative staphylococcus|0
    transferred to the ICU on ventilatory support|0
    received medical therapy for sepsis|0
    hospitalization complicated by failure to wean from ventilatory support|0
    multiple bouts of fever secondary to sepsis|0
    underwent 3 other surgeries for further abscess debridement|0
    transferred to a long-term acute care hospital|0
    long-term care|0
    rehabilitation|0
    