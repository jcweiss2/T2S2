66 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
dual-chamber pacemaker | -10512 | -10512 | Factual
sick sinus syndrome | -10512 | 0 | Factual
paroxysmal atrial fibrillation | -10512 | 0 | Factual
severe lumbar back pain | -24 | 0 | Factual
mental status changes | -24 | 0 | Factual
hypotension | -24 | 0 | Factual
acute renal failure | -24 | 0 | Factual
hypoxemic respiratory failure | -24 | 0 | Factual
emergent intubation | -24 | 0 | Factual
severe sepsis | -24 | 0 | Factual
hemodynamic support | -24 | 0 | Factual
vasopressin | -24 | 0 | Factual
norepinephrine | -24 | 0 | Factual
blood cultures | -24 | -24 | Factual
methicillin-sensitive Staphylococcus aureus | -24 | 0 | Factual
vancomycin | -24 | -12 | Factual
nafcillin | -12 | 0 | Factual
transthoracic echocardiogram | -12 | -12 | Factual
left ventricular ejection fraction | -12 | -12 | Factual
patent foramen ovale | -12 | 0 | Factual
computed tomography scan | -12 | -12 | Factual
osteomyelitis | -12 | 0 | Factual
magnetic resonance imaging | -12 | -12 | Factual
septic emboli | -12 | 0 | Factual
transesophageal echocardiogram | -6 | -6 | Factual
vegetation | -6 | 0 | Factual
pacemaker lead | -6 | 0 | Factual
tricuspid valve | -6 | 0 | Factual
cardiothoracic surgery | -6 | -6 | Factual
surgical intervention | -6 | -6 | Factual
laser lead extraction | -2 | 0 | Factual
Indigo Thrombectomy System | -1 | 1 | Factual
intracardiac echocardiography | -1 | 1 | Factual
vacuum-assisted vegetation removal | -1 | 1 | Factual
femoral veins | 0 | 0 | Factual
GORE DrySeal Flex introducer sheath | 0 | 0 | Factual
CARTO SoundStar | 0 | 0 | Factual
Indigo CAT8 XTORQ | 0 | 0 | Factual
aspiration | 0 | 1 | Factual
vegetation extraction | 0 | 1 | Factual
lead extraction | 1 | 2 | Factual
pocket inspection | 2 | 2 | Factual
hemostasis | 2 | 2 | Factual
procedure time | 0 | 2 | Factual
blood loss | 0 | 2 | Factual
pathology | 2 | 2 | Factual
gram-positive cocci | 2 | 2 | Factual
culture-positive | 2 | 2 | Factual
methicillin-sensitive Staphylococcus aureus | 2 | 2 | Factual
condition improved | 2 | 50 | Factual
tissue necrosis | 50 | 50 | Factual
lactic acidosis | 50 | 50 | Factual
renal failure | 50 | 50 | Factual
withdraw care | 50 | 50 | Factual
extubated | 50 | 50 | Factual
died | 50 | 50 | Factual