70 years old | 0
    woman | 0
    presented to the emergency department | 0
    acute epigastric pain | -1
    diabetes mellitus | 0
    cholecystectomy | 0
    heterozygote alpha-1 antitrypsin deficiency | 0
    epigastric tenderness | 0
    no fever | 0
    pulse rate 82 beats/min | 0
    blood pressure 128/68 mmHg | 0
    normal respiratory rate | 0
    normal oxygen saturation | 0
    total bilirubin 0.28 mg/dL | 0
    glutamic oxaloacetic transaminase 45 U/L | 0
    glutamic pyruvic transaminase 30 U/L | 0
    γ-glutamyltransferase 91 U/L | 0
    alkaline phosphatase 99 U/L | 0
    lipase 3518 U/L | 0
    complete blood count normal | 0
    C-reactive protein normal | 0
    coagulation normal | 0
    renal function normal | 0
    electrocardiogram normal | 0
    cardiac enzymes normal | 0
    acute pancreatitis suspected | 0
    intravenous fluid resuscitation | 0
    pain relief | 0
    deteriorated rapidly | 0
    severe septic shock | 0
    transferred to intensive care unit | 0
    mechanical ventilation | 0
    aggressive hemodynamic support | 0
    computed tomography scan showing large air-filled cavity | 0
    bile duct mildly dilated | 0
    nonradiopaque choledocholithiasis could not be ruled out | 0
    no apparent inflammation surrounding pancreas | 0
    diagnosis of emphysematous hepatitis | 0
    broad-spectrum intravenous antibiotics (meropenem, vancomycin, amikacin) | 0
    CT-guided percutaneous pigtail catheter drainage | 0
    no significant fluid or pus | 0
    pigtail drain flushed with continuous saline irrigation | 0
    elevated serum lipase | 0
    mildly dilated bile duct | 0
    endoscopic retrograde cholangiopancreatography performed | 0
    cholangiogram normal biliary anatomy | 0
    clear bile after endoscopic sphincterotomy | 0
    antibiotics rationalized to ceftriaxone and metronidazole | 0
    blood cultures revealed Escherichia coli | 0
    Streptococcus anginosus | 0
    Klebsiella oxytoca | 0
    continuous pigtail irrigation stopped after 3 days | 72
    drain removed after 5 days | 120
    weaned from ventilator | 168
    transferred to ward after 2 weeks | 336
    continued recovery favorably | 0
    discharged 1 month after admission | 720
    colonoscopy performed | 0
    transthoracic echocardiogram performed | 0
    CT scan showed liquefied collection in segment VII | 720
    magnetic resonance imaging performed 6 weeks later | 1008
    MRI showed 10 cm cystic formation | 1008
    positron emission tomography performed 9 weeks later | 1512
    PET scan showed no metabolic activity in large collection | 1512
    2 cm PET-positive nodule detected | 1512
    surgical drainage performed | 1512
    laparoscopic deroofing and debridement | 2160
    partial hepatectomy of 2 cm lesion | 2160
    no malignancy found | 2160
    microbiological cultures sterile | 2160
    antibiotics discontinued after 14 weeks | 2352
    uneventful recovery | 2160
    hospitalized again for COVID-19 infection | 2160
    asymptomatic | 2160
    no recurrence on follow-up imaging | 2160

  