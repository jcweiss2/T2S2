87 years old | 0
female | 0
admitted to the emergency unit | 0
abdominal pain | -24
diarrhea | -24
dizziness | -24
lower abdominal pain | -24
watery stool | -24
right-sided pelvic pain | -24
hypertension | 0
third-degree atrioventricular block | 0
pacemaker | 0
fallen at home | -24
tenderness over the pubic bone | 0
tenderness over the lower abdomen | 0
no peritoneal reaction | 0
right hip region swollen | 0
right hip region tender | 0
rectal examination normal | 0
hemoglobin 6.5 mmol/l | 0
white blood cell count 10.6 × 10^9/l | 0
platelets 102 × 10^9/l | 0
creatinine 196 µmol/l | 0
C-reactive protein 29 mg/l | 0
arterial blood gas analysis showed pH 7.16 | 0
lactate 13.6 mmol/l | 0
right-sided nondisplaced pubic ramus fracture | 0
arterial blood gas repeated | 9
pH 7.42 | 9
lactate 2.7 | 9
severe dehydration | 0
severe abdominal pain | 21
C-reactive protein increased to 123 mmol/l | 21
suspicion of intestinal ischemia | 21
exploratory laparotomy | 21
necrosis of the sigmoid colon | 21
necrosis of the proximal part of rectum | 21
flexible sigmoidoscopy | 21
non-vital mucosa 10–25 cm from anus | 21
non-vital ileum 20 cm from the ileocecal region | 21
retroperitoneal hematomas | 21
resection of non-vital intestinal segments | 21
ileostomy | 21
sigmoideostomy | 21
severe sepsis | 21
discharged | 240
histopathology of the resected tissue | 240
necrosis due to ischemia | 240
no sign of vasculitis | 240
no sign of thrombosis | 240