20 years old | 0
female | 0
pharyngitis | -336
exposure to group A beta-hemolytic streptococcus | -336
exposure to Epstein-Barr virus (EBV) | -336
azithromycin | -336
travel to Florida | -336
attended social events | -336
shared utensils and beverages | -336
dental cleaning | -720
persistent fever | -120
cough | -120
swollen glands | -120
worsening sore throat | -120
shortness of breath | -120
increased work of breathing | -120
rash on left wrist | -120
scleral icterus | -120
bright blurry vision | -120
admitted to outside hospital | -120
diagnosis of respiratory distress | -120
possible sepsis | -120
diagnosis of pharyngitis | -120
blood culture | -120
COVID-19 PCR tests | -120
complete blood count | -120
C-reactive protein | -120
ferritin | -120
procalcitonin | -120
chest x-ray | -120
CT scan of the chest | -120
bilateral cavitary pneumonia | -120
left pleural effusion | -120
doxycycline | -120
ceftriaxone | -120
transferred to BMSCH PICU | -96
admission to BMSCH PICU | 0
mild acute respiratory distress | 0
tachypnea | 0
suprasternal retractions | 0
rashes along ulnar side of the left hand | 0
swelling | 0
tenderness | 0
diminished breath sounds | 0
high-flow nasal cannula | 0
IV vancomycin | 0
cefepime | 0
metronidazole | 0
blood culture growing gram-negative rods | 24
Fusobacterium nucleatum | 24
cefepime changed to ceftriaxone | 24
vancomycin and metronidazole continued | 24
left wrist pain | 24
limited mobility of the left shoulder | 24
platelets decreased | 24
plasma and platelet transfusions | 24
echocardiogram | 24
fractional shortening | 24
ejection fraction | 24
synchronized intermittent mandatory ventilation (SIMV) | 48
inotropes | 48
left pleurocentesis | 48
video-assisted bilateral thoracoscopic surgery (VATS) | 48
bilateral chest tubes | 48
pleural fluid | 48
surgical pathology report | 48
repeat pleural fluid cultures | 48
high flow nasal cannula (HFLNC) | 72
procalcitonin and C-reactive protein trended down | 72
hemodynamic status improved | 72
additional chest tubes | 96
repeat echocardiogram | 96
tissue near the tricuspid valve | 96
small pericardial effusion | 96
MR of left upper extremity | 120
musculoskeletal edema | 120
proximal humeral osteomyelitis | 120
T12 vertebral body emphysematous osteomyelitis | 120
bilateral duplex venous ultrasounds | 120
duplex ultrasound of the bilateral carotids | 120
discharged from PICU | 168
follow-up care | 240