40 years old | 0
    man | 0
    admitted to the hospital | 0
    shock | 0
    flu-like illness | -72
    nausea | -72
    general malaise | -72
    lower abdominal pain | -72
    severe diarrhea | -72
    5% albumin administered | -72
    saline administered | -72
    consciousness deteriorated | -48
    right hemiparesis | -48
    temperature of 36.0°C | 0
    blood pressure of 95/72 mm Hg | 0
    pulse of 160 beats/min | 0
    respiratory rate of 25 breaths/min | 0
    SpO2 100% | 0
    jugular vein collapsed | 0
    bilateral radial artery pulses insufficiently palpable | 0
    extremities cold | 0
    whole-blood sample coagulated easily | 0
    hyperviscosity | 0
    polycythemia | 0
    hypoalbuminemia | 0
    severe leukocytosis | 0
    elevated creatinine | 0
    serum electrolytes normal | 0
    severe metabolic acidosis | 0
    influenza virus types A and B positive | 0
    pericardial effusion | 0
    collapsed inferior vena cava | 0
    occlusion of left M2 segment of MCA | 0
    high signal intensity in MCA territory | 0
    acute cerebral infarction | 0
    midline shift of the head | 20
    external decompression surgery performed | 20
    internal decompression surgery performed | 20
    postoperative intracranial pressure 9 mm Hg | 20
    cerebral edema progression | 20
    excessive cerebral edema developed | 20
    internal decompression added | 32
    hypoproteinemia | 0
    hemoconcentration | 0
    intravascular volume depletion | 0
    increased vascular permeability | 0
    extravasation of albumin | 0
    mechanical ventilation | 0
    massive fluid resuscitation (10 liters/day) | 0
    swelling in lateral surfaces of legs | 0
    redness in lateral surfaces of legs | 0
    heat sensation in lateral surfaces of legs | 0
    pretibial compartment syndrome | 0
    bilateral calf fasciotomy performed | 0
    pan cultures negative | 0
    toxic shock syndrome considered | 0
    sepsis considered | 0
    anaphylaxis considered | 0
    acute adrenal insufficiency considered | 0
    drug reactions considered | 0
    polycythemia vera considered | 0
    severe right hemiparesis persisted | 1464
    Broca's aphasia persisted | 1464
    unable to walk without assistance | 1464
    theophylline administered | 1464
    prophylaxis against ISCLS | 1464
    7 attacks of ISCLS documented | 8760
    2 severe episodes requiring fasciotomy | 8760
    appropriate fluid resuscitation | 8760
    no observed stroke recurrence | 8760
    monoclonal immunoglobulin (IgG kappa) found | 8760
    intravenous infusion of immunoglobulins | 8760
    corticosteroids administered | 8760
    immunosuppressive therapy administered | 8760