74 years old | 0
    white | 0
    woman | 0
    presented to the Emergency Department | 0
    low-grade fever | -48
    dry cough | -48
    shortness of breath | -48
    admitted to another hospital for an elective right total knee replacement | -168
    uneventful post-operative course | -168
    went to the hospital in a healthy state | -168
    stayed in a private room | -168
    denied any recent sick contacts | 0
    denied any travel history | 0
    pain in the right knee | -168
    redness in the right knee | -168
    swelling in the right knee | -168
    essential hypertension | 0
    obesity | 0
    myasthenia gravis in remission | 0
    osteoarthritis | 0
    body temperature of 37.3°C | 0
    blood pressure of 121/82 | 0
    pulse of 87 beats per minute | 0
    respiratory rate of 16 breaths per minute | 0
    oxygen saturation of 87% while breathing ambient air | 0
    lung auscultation revealed bilateral rhonchi | 0
    lung auscultation revealed rales | 0
    chest radiography performed | 0
    patchy air space opacity in the right upper lobe suspicious for pneumonia | 0
    remainder of the examination unremarkable | 0
    rapid NAAT for influenza A and B negative | 0
    nasopharyngeal swab specimen obtained | 0
    SARS-CoV-2 detection sent to state laboratory | 0
    admitted to the airborne-isolation unit | 0
    started on broad-spectrum antibiotics with cefepime | 0
    started on levofloxacin | 0
    blood cultures drawn | 0
    sputum cultures drawn | 0
    supportive care with 2 L of supplemental oxygen | 0
    developed mild diarrhea | 72
    developed generalized weakness | 72
    developed fatigue | 72
    evaluated by Neurology | 72
    started on 1 g/kg intravenous immunoglobulin for 4 days | 72
    mild MG exacerbation | 72
    pending MG crises | 72
    ABGs monitored | 0
    complete blood count monitored | 0
    basic metabolic profile monitored | 0
    mild absolute lymphopenia | 0
    anemia | 0
    ABGs revealed pH of 7.46 | 0
    ABGs revealed pCO2 of 44.6 mmHg | 0
    ABGs revealed pO2 of 94.7 mmHg | 0
    ABGs revealed bicarbonate of 31.4 mmol/L | 0
    creatinine kinase normal | 144
    lactic acid normal | 144
    lactate dehydrogenase elevated | 144
    ferritin elevated | 144
    interleukin-6 elevated | 144
    progressively increasing SOB | 24
    progressively increasing SOB | 72
    progressively increasing SOB | 96
    oxygen requirements increased up to 10 L high-flow nasal cannula | 96
    nasopharyngeal swab results positive for SARS-CoV-2 | 96
    started on oral hydroxychloroquine 400 mg once | 96
    started on hydroxychloroquine 200 mg twice a day | 96
    started on azithromycin 500 mg once a day intravenously | 96
    started on zinc sulfate 220 mg 3 times a day | 96
    started on oral vitamin C 1 g twice a day | 96
    blood cultures negative | 96
    sputum cultures negative | 96
    broad-spectrum antibiotics discontinued | 96
    SOB worsened rapidly | 144
    oxygen requirements went up to 15 L | 144
    drowsy | 144
    moderate distress | 144
    unable to protect the airways | 144
    blood pressure of 78/56 mmHg | 144
    heart rate of 112 beats per minute | 144
    temperature 38°C | 144
    respiratory rate of 28 breaths per minute | 144
    CXR revealed bilateral alveolar infiltrates due to pneumonia | 144
    CXR revealed interstitial edema consistent with ARDS | 144
    intubated | 144
    started on pressure-regulated volume-controlled mechanical ventilation | 144
    started on norepinephrine 0.02 mcg/kg/min | 144
    titrated to maintain mean arterial pressure more than 65 mmHg | 144
    started on colchicine 0.6 mg twice a day | 144
    elevated interleukin-6 levels | 144
    started on high-dose vitamin C 11 g per 24 h as a continuous intravenous infusion | 168
    clinical condition started to improve slowly | 168
    norepinephrine support stopped | 192
    CXR showed significant improvement of the pneumonia | 240
    CXR showed significant improvement of the interstitial edema | 240
    spontaneous breathing trial with CPAP/PS successfully tolerated | 240
    ABGs revealed pH of 7.49 mmHg | 240
    ABGs revealed pCO2 of 40.2 mmHg | 240
    ABGs revealed pO2 of 77.1 mmHg | 240
    ABGs revealed bicarbonate of 30.2 mmol/L | 240
    extubated to 4 L of oxygen with a nasal cannula | 240
    breathing status continued to improve | 240
    oxygen saturation of 92% on day 16 of illness while breathing ambient air | 384
    CXR revealed almost complete resolution of the infiltrates | 384
    received 5 days of treatment with hydroxychloroquine | 384
    received azithromycin | 384
    received 4 days of colchicine | 384
    high-dose vitamin C infusion continued for 10 days | 384
    oral zinc sulfate continued for 10 days | 384
    inpatient physical rehabilitation | 384
    inpatient occupational rehabilitation | 384
    transferred from the Critical Care Unit to an isolation room | 384
    still positive by RT-PCR for SARS-CoV-2 | 384
    discharged from the hospital | 384
    additional 14 days of quarantine | 384
    septic shock | 144
    ARDS | 144
    MV initiation | 144
    cytokine storm | 144
    ICU stay | 144
    mechanical ventilation duration | 144
    recovered from the disease | 240
    almost complete resolution of the infiltrates | 384
    discharged in stable condition | 384
    <|eot_id|>
    