46 years old | 0
male | 0
arterial hypertension | -672
obesity | -672
admitted to the hospital | 0
fever | -336
hypotension | 0
asthenia | 0
cardiological examination | -672
electrocardiogram (ECG) | -672
transthoracic echocardiography (TTE) | -672
COVID-19 infection | -336
rhinitis | -336
mild cough | -336
alert | 0
oriented | 0
cooperative | 0
asthenic | 0
blood pressure (BP) 85/55 mmHg | 0
heart rate (HR) 120 bpm | 0
arterial oxygen saturation 85% | 0
fever 38.3 C° | 0
femoral central venous catheter (CVC) | 0
sinus tachycardia | 0
diffuse low voltages | 0
absence of significant repolarization abnormalities | 0
neutrophilic leukocytosis | 0
C-reactive protein (CRP) elevation | 0
Procalcitonin elevation | 0
elevated high sensitivity Troponin (hs-Tn) | 0
elevated brain natriuretic peptide (BNP) | 0
elevated creatinine | 0
transaminases and total bilirubin | 0
reverse transcription-polymerase chain reaction (RT-PCR) nasopharyngeal swab for COVID-19 negative | 0
COVID-19 IgM antibody test positive | 0
normal left ventricular (LV) cavitary dimensions | 0
diffuse LV parietal thickening | 0
severely reduced LV global systolic function | 0
grade II LV diastolic dysfunction | 0
normal cavitary dimensions and reduced global right ventricular (RV) systolic function | 0
inferior vena cava (IVC) dilated | 0
right ventricular systolic pressure (RVSP) 41 mmHg | 0
absence of hemodynamically significant valvulopathy | 0
slight amount of pericardial effusion | 0
blood cultures started | 0
broad-spectrum antibiotic therapy | 0
INN-daptomycin | 0
piperacillin/tazobactam | 0
crystalloid hydration | 0
nasal cannula ventilatory therapy | 0
norepinephrine therapy | 0
poor hemodynamic response | 0
levosimendan therapy | 0
bolus administration avoided | 0
continuous maintenance intravenous infusion | 0
BP increased to 100/60 mmHg | 12
HR decreased to 110 bpm | 12
further hemodynamic improvement | 24
BP 125/70 mmHg | 24
HR 95 bpm | 24
diuresis 1800 ml | 24
control TTE performed | 12
control TTE performed | 24
LV EF 66% | 24
dP/dT ratio 1275 mmHg/sec | 24
TAPSE 23 mm | 24
tricuspid S-wave velocity at TDI 11.2 cm/sec | 24
SVi 27 ml/m2 | 24
CI 2.5 l/min/m2 | 24
LV diastolic function improved | 24
IVC diameter 18 mm | 24
IVC collapse 100% | 24
RVSP 28 mmHg | 24
diffuse parietal thickening persisted | 24
increased myocardial reflectivity | 24
blood culture results negative | 24
CVC removed | 24
culture of CVC tip negative | 24
cardiac magnetic resonance imaging (CMR) | 48
steady-state free precession-CINE (SSFp-CINE) | 48
double inversion recovery/T1 weighted (DIR/T1w) | 48
triple inversion recovery/T2 weighted (TIR/T2w) | 48
early gadolinium enhancement (EGE) | 48
late gadolinium enhancement (LGE) | 48
normal LV and RV volumes and systolic function | 48
mild hypokinesia of the mid and basal segments | 48
increased signal intensity defined as the ratio of skeletal muscle intensity > 1.9 | 48
edema spread to almost all LV myocardial segments | 48
subendocardial localization | 48
endomyocardial biopsy | 72
lymphocytic myocarditis | 72
coronary arteriography | 72
normal coronary circulation | 72
discharged | 504
excellent hemodynamic compensation | 504
normal laboratory findings | 504
normal electrocardiographic findings | 504
normal echocardiographic findings | 504
TTE performed at 1 month after discharge | 744
normal findings | 744
TTE performed at 3 months after discharge | 2232
normal findings | 2232