66 years old | 0
    woman | 0
    presented to the emergency department | 0
    positive blood cultures | -72
    Staphylococcus epidermidis | -72
    chills | -2160
    leukocytosis | -72
    20,000/mm3 | -72
    complete blood count | -72
    intermittent chills | -2160
    burning chest pain | -2160
    past 3 months | -2160
    rigors | -72
    denied objective fever | 0
    denied shortness of breath | 0
    denied cough | 0
    denied dysuria | 0
    denied indwelling catheters | 0
    denied intravenous drug use | 0
    febrile | 0
    temperature 102.2℉ | 0
    well-healed median sternotomy incision | 0
    grade 3 early systolic murmur | 0
    early diastolic sound | 0
    essential hypertension | -26280
    dyslipidemia | -26280
    severe aortic stenosis | -26280
    atherosclerotic coronary artery disease | -26280
    coronary artery bypass grafting | -26280
    surgical aortic valve replacement | -26280
    21 mm bioprosthetic valve | -26280
    3 years earlier | -26280
    infective endocarditis | 0
    sepsis of unknown etiology | 0
    intravenous antibiotics | 0
    chest x-ray | 0
    electrocardiogram | 0
    urinalysis | 0
    sputum cultures | 0
    transthoracic echocardiogram | 0
    large mobile hyperechoic mass | 0
    tricuspid valve | 0
    right ventricle | 0
    transesophageal echocardiography | 0
    large (3.0 × 1.6 cm) multilobed mobile hyperechoic mass | 0
    mild to moderate tricuspid regurgitation | 0
    moderately elevated right ventricular systolic pressure | 0
    sessile hyperechoic mass (3.0 × 1.7 cm) | 0
    right atrial appendage | 0
    vegetations | 0
    admitted to the cardiac unit | 0
    collaborative decision | 0
    AngioVac System | 0
    fluoroscopic guidance | 0
    TEE guidance | 0
    mechanical thrombectomy | 0
    tricuspid valve | 0
    right atrium | 0
    reduced vegetation burden | 0
    tricuspid leaflet integrity | 0
    remnant leads | 0
    nidus of infection | 0
    transferred to the intensive care unit | 0
    cardiac computed tomography | 0
    3D reconstruction | 0
    atrial epicardial wires | 0
    ventricular epicardial wires | 0
    postoperative period | 0
    migrated and perforated the right atrium | 0
    percutaneous lead removal | 24
    right femoral vein access | 24
    6 French 55 cm sheath | 24
    EN Snare three-loop system | 24
    CloverSnare | 24
    multipurpose guide catheter | 24
    Amplatz Goose Neck Snare | 24
    successful snaring | 24
    remnant lead removal | 24
    echocardiogram | 24
    no pericardial effusion | 24
    peripherally inserted central catheter | 24
    intravenous antibiotics | 24
    infectious disease specialist follow-up | 24
    no recurrent bacteremia | 168
    afebrile | 168
    repeat transthoracic echocardiogram | 1008
    no vegetations | 1008
    mild regurgitation | 1008
    