64 years old | 0
female | 0
diabetes mellitus | - (no timestamp provided)
admitted to the intensive care unit | 0
septic shock | 0
acute left pyelonephritis | 0
CT scan | 0
lower mass syndrome of the left kidney | 0
necrosis | 0
calcifications | 0
wide nephrectomy with adrenalectomy | 0
gross examination | 0
fleshy well-defined tumor | 0
patchy hemorrhagic areas | 0
necrotic areas | 0
histological examination | 0
dual carcinomatous proliferation | 0
clear cells | 0
eosinophilic cells | 0
lobular growth pattern | 0
tubulo-cystic growth pattern | 0
no vascular invasion | 0
renal capsule spared | 0
adrenal gland spared | 0
sarcomatoid differentiation | 0
spindle-shaped cells | 0
immunohistochemical study | 0
tumor cells negative for CD117 | 0
tumor cells negative for CD10 | 0
tumor cells negative for racemase | 0
tumor cells negative for vimentin | 0
septic shock uncontrolled | 0
patient state deteriorated | 0
died | 24 (assuming "a few days after admission" translates to ~24 hours)
diabetes mellitus | 0
eosinophilic cells |3 0
died | 24
