36 years old | 0
male | 0
IgA nephropathy | 0
hemo-dialysis | 0
left forearm AVF | 0
hepatitis B | 0
hypertension | 0
Charcot-Marie-Tooth disease | 0
left flank pain | 0
fever denied | 0
chest pain denied | 0
shortness of breath denied | 0
cough denied | 0
vomiting denied | 0
diarrhea denied | 0
dysuria denied | 0
prior problems with AVF denied | 0
temperature 98.5°F | 0
temperature 102.3°F | 24
pulse 108 beats per min | 0
respiratory rate 17 cycles per min | 0
blood pressure 106/64 mmHg | 0
99% oxygen saturation | 0
mild distress | 0
abdomen soft and non-tender | 0
costovertebral angle tenderness not elicited | 0
AVF site not tender | 0
electrocardiogram normal sinus rhythm | 0
WBC 10.2 k/ul | 0
WBC 41.9 k/ul | 192
WBC 36.5 k/ul | 192
WBC 10.2 k/ul | 456
hemoglobin 10.9 g/dl | 0
platelets 197 k/ul | 0
erythrocyte sedimentation rate 48 | 0
procalcitonin greater than 200 ng/dl | 0
C-reactive protein 4.81 mg/dl | 0
sodium 134 mmol/l | 0
potassium 4.2 mmol/l | 0
chloride 91 mmol/l | 0
bicarbonate 27 mmol/l | 0
blood urea nitrogen 66 mg/dl | 0
creatinine 12.4 mg/dl | 0
urinalysis WBC count 1/HPF | 0
urinalysis absence of bacteria | 0
urinalysis absence of leukocyte esterase | 0
urinalysis absence of nitrate | 0
CXR clear lungs | 0
CT abdomen and pelvis no evidence of acute appendicitis | 0
CT abdomen and pelvis no evidence of diverticulitis | 0
CT abdomen and pelvis no evidence of mechanical bowel obstruction | 0
CT abdomen and pelvis no ascites | 0
CT abdomen and pelvis no evidence of portal hypertension | 0
CT abdomen and pelvis both kidneys atrophic | 0
open wound at AVF fistula | 24
wound swabbed and sent for cultures | 24
wound examined and dressed regularly | 24
wound grew Streptococcus group A | 48
hypotensive | 24
vancomycin administration | 24
meropenem administration | 24
right internal jugular hemodialysis catheter inserted | 24
transferred to Medical Intensive Care Unit | 24
CXR moderate left pleural effusion | 24
chest CT large left pleural effusion | 48
CXR near-complete opacification of left lung | 48
pigtail chest tube inserted | 48
CXR left-sided pigtail catheter in situ | 48
pleural fluid analysis | 48
pleural fluid cloudy | 48
pleural fluid WBC 15 762/cumm | 48
pleural fluid red blood cell 3556/cumm | 48
pleural fluid polynuclear white blood cell 84% | 48
pleural fluid glucose 2 mg/dL | 48
pleural fluid total protein 4.2 | 48
pleural fluid lactate dehydrogenase 9208 u/L | 48
serum protein 5.1 g/dl | 48
serum lactate dehydrogenase 150 u/l | 48
clindamycin administration | 48
CXR small residual left effusion | 168
left pigtail catheter removed | 168
CXR re-accumulation of pleural fluid | 192
VATS with pleural drainage and decortication | 192
chest tubes inserted | 192
CXR improved left hemithorax | 240
left anterior and lateral chest tubes removed | 288
left posterior chest tube removed | 360
sepsis | 24
sepsis resolved | 72
vital signs improved | 72
blood cultures negative | 0
pleural fluid cultures negative | 0
transthoracic echocardiogram no valvular vegetations | 0
regular dialysis | 24
AVF revised and repaired | 240
meropenem discontinued | 288
ceftriaxone administration | 288
vancomycin administration | 0
discharged | 648
explosive pleuritis | 48