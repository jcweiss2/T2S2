61 years old | 0
    male | 0
    presented to a community hospital | 0
    transient loss of consciousness | 0
    acute chest discomfort | 0
    upper respiratory tract infection | -336
    subjective fever | -24
    rigors | -24
    apyrexic | 0
    normal physical examination | 0
    normal serum leukocyte count | 0
    normal chest radiograph | 0
    inferior ST-segment elevation myocardial infarction | 0
    no stigmata of endocarditis | 0
    no signs of aortic dissection | 0
    intravenous thrombolysis | 0
    transferred to a tertiary care hospital | 0
    coronary angiography | 0
    occlusion of the distal left-dominant posterior descending artery | 0
    no other significant lesions | 0
    angioplasty not possible | 0
    transthoracic echocardiography | 0
    left ventricular apical-inferior hypokinesis | 0
    no valve lesions |) 0
    cranial computed tomography | 0
    small cerebellar hemorrhage | 0
    clinically stable | 0
    transferred to cardiac intensive care unit | 0
    onset of polymorphic ventricular tachycardia storm | 24
    profound shock | 24
    admission blood cultures grew methicillin-sensitive Staphylococcus aureus | 0
    intravenous antibiotics | 0
    maximum supportive therapy | 0
    died | 48
    autopsy | 48
    acute bacterial myocarditis | 48
    multifocal suppuration of the lower interventricular septum | 48
    inferior ventricles | 48
    unremarkable cardiac valves | 48
    intramyocardial abscesses | 48
    gram-positive cocci | 48
    posterior descending artery exhibited acute bacterial vasculitis | 48
    adjacent abscess | 48
    microabscesses in the brain | 48
    microabscesses in the spinal cord | 48
    
    61 years old | 0
    male | 0
    presented to a community hospital | 0
    transient loss of consciousness | 0
    acute chest discomfort | 0
    upper respiratory tract infection | -336
    subjective fever | -24
    rigors | -24
    apyrexic | 0
    normal physical examination | 0
    normal serum leukocyte count | 0
    normal chest radiograph | 0
    inferior ST-segment elevation myocardial infarction | 0
    no stigmata of endocarditis | 0
    no signs of aortic dissection | 0
    intravenous thrombolysis | 0
    transferred to a tertiary care hospital | 0
    coronary angiography | 0
    occlusion of the distal left-dominant posterior descending artery | 0
    no other significant lesions | 0
    angioplasty not possible | 0
    transthoracic echocardiography | 0
    left ventricular apical-inferior hypokinesis | 0
    no valve lesions | 0
    cranial computed tomography | 0
    small cerebellar hemorrhage | 0
    clinically stable | 0
    transferred to cardiac intensive care unit | 0
    onset of polymorphic ventricular tachycardia storm | 24
    profound shock | 24
    admission blood cultures grew methicillin-sensitive Staphylococcus aureus | 0
    intravenous antibiotics | 0
    maximum supportive therapy | 0
    died | 48
    autopsy | 48
    acute bacterial myocarditis | 48
    multifocal suppuration of the lower interventricular septum | 48
    inferior ventricles | 48
    unremarkable cardiac valves | 48
    intramyocardial abscesses | 48
    gram-positive cocci | 48
    posterior descending artery exhibited acute bacterial vasculitis | 48
    adjacent abscess | 48
    microabscesses in the brain | 48
    microabscesses in the spinal cord | 48