48 years old | 0  
    female | 0  
    weight loss | -720  
    fever | -720  
    general weakness | -720  
    admitted to another hospital | -720  
    diagnosed with hyperparathyroidism | -720  
    febrile shock | -720  
    transferred to our hospital | 0  
    blood pressure of 86/54 mmHg | 0  
    pulse rate of 136/min | 0  
    body temperature of 38.5℃ | 0  
    respiratory rate of 28/min | 0  
    coarse breathing sounds | 0  
    crackles in both lower lung zones | 0  
    severe dyspnea | 0  
    serum urea 37 mg/dL | 0  
    creatinine 2.3 mg/dL | 0  
    calcium 14.1 mg/dL | 0  
    ionized calcium 7.8 mg/dL | 0  
    phosphorus 2.3 mg/dL | 0  
    intact PTH 635.30 pg/mL | 0  
    WBC 24,460/mm3 |8  
    arterial blood gas analysis pH 7.235 | 0  
    PaCO2 61.8 mmHg | 0  
    PaO2 75.9 mmHg | 0  
    HCO3 25.6 mmol/L | 0  
    O2 saturation 94% | 0  
    admission chest radiograph bilateral airspace consolidation | 0  
    precontrast chest CT airspace consolidation | 0  
    multifocal patchy ground-glass opacities | 0  
    neck CT parathyroid adenoma | 0  
    diagnosed hyperparathyroidism-associated hypercalcemia | 0  
    diagnosed pneumonia-complicated septic shock | 0  
    moved to intensive care unit | 0  
    mechanical ventilator care | 0  
    continuous renal replacement therapy | 0  
    bronchoscopy | 0  
    bronchoalveolar lavage | 0  
    MRSA | 0  
    parathyroidectomy | 168  
    improved from sepsis | 168  
    weaned from mechanical ventilation | 168  
    bilateral pulmonary airspace consolidations remained | 168  
    HRCT performed | 168  
    follow-up CT geographic high7.3attenuation consolidation | 168  
    ground-glass opacities | 168  
    bone scintigraphy dense accumulation bilateral lower lung zones | 168  
    diffusely increased uptake along stomach wall | 168  
    exertional dyspnea | 168  
    severely restrictive physiology | 168  
    low diffusion capacity | 168  
    percutaneous lung biopsy | 168  
    histologic specimen metastatic pulmonary calcification | 168  
    surgical resection of parathyroid | 648  
    serum calcium level normal | 648  
    pulmonary function test nearly complete recovery | 648  
    recovered health without symptoms | 648  
    metastatic pulmonary calcification | 168  
    dense airspace consolidation bilateral lower lobes | 168  
    pneumonia | -720  
    sepsis | -720  
    hypercalcemia | -720  
    chronic renal failure | -720  
    increased tissue alkalinity | -720  
    patchy bilateral airspace consolidation lower lung zones | 0  
    airspace consolidation bilateral lower lobes | 0  
    multifocal patchy ground-glass opacities | 0  
    right infrathyroid area parathyroid adenoma | 0  
    hyperparathyroidism | -720  
    mechanical ventilator care ACMV | 0  
    continuous renal replacement therapy CRRT | 0  
    bronchoscopy bronchoalveolar lavage BAL | 0  
    methicillin-resistant Staphylococcus aureus MRSA | 0  
    parathyroidectomy | 168  
    improved from sepsis | 168  
    weaned from mechanical ventilation | 168  
    bilateral pulmonary airspace consolidations remained | 168  
    HRCT performed | 168  
    follow-up CT high-attenuation consolidation | 168  
    ground-glass opacities | 168  
    bone scintigraphy Tc-99m MDP bilateral lower lung zones | 168  
    diffusely increased uptake along stomach wall | 168  
    exertional dyspnea | 168  
    severely restrictive physiology | 168  
    low diffusion capacity | 168  
    percutaneous lung biopsy | 168  
    histologic specimen metastatic pulmonary calcification | 168  
    surgical resection parathyroid | 648  
    serum calcium normal | 648  
    pulmonary function test recovery | 648  
    recovered health | 648  
    metastatic pulmonary calcification | 168  
    dense airspace consolidation bilateral lower lobes | 168  
    pneumonia | -720  
    sepsis | -720  
    hypercalcemia | -720  
    chronic renal failure | -720  
    increased tissue alkalinity | -720  
    patchy bilateral airspace consolidation lower lung zones | 0  
    airspace consolidation bilateral lower lobes | 0  
    multifocal patchy ground-glass opacities | 0  
    right infrathyroid area parathyroid adenoma | 0  
    hyperparathyroidism | -720  
    mechanical ventilator care ACMV | 0  
    continuous renal replacement therapy CRRT | 0  
    bronchoscopy bronchoalveolar lavage BAL | 0  
    methicillin-resistant Staphylococcus aureus MRSA | 0  
    parathyroidectomy | 168  
    improved from sepsis | 168  
    weaned from mechanical ventilation | 168  
    bilateral pulmonary airspace consolidations remained | 168  
    HRCT performed | 168  
    follow-up CT high-attenuation consolidation | 168  
    ground-glass opacities | 168  
    bone scintigraphy Tc-99m MDP bilateral lower lung zones | 168  
    diffusely increased uptake along stomach wall | 168  
    exertional dyspnea | 168  
    severely restrictive physiology | 168  
    low diffusion capacity | 168  
    percutaneous lung biopsy | 168  
    histologic specimen metastatic pulmonary calcification | 168  
    surgical resection parathyroid | 648  
    serum calcium normal | 648  
    pulmonary function test recovery | 648  
    recovered health | 648  
    