65 years old | 0
woman | 0
presented to the emergency room | 0
right flank pain | 0
fever | 0
diabetes | -175200
oral hypoglycemic agents | -175200
blood pressure 80/50 mmHg | 0
temperature 39°C | 0
pulse 130 beats/minute | 0
respiration rate 20 breaths/minute | 0
knocking tenderness on the right flank area | 0
WBC count 23400/μL | 0
hemoglobin 9.7 g/dL | 0
platelet count 97000/μL | 0
C-reactive protein 21.97 mg/dL | 0
blood urea nitrogen 35.3 mg/dL | 0
creatinine 2.21 mg/dL |:0
sodium 142 mEq/L | 0
potassium 3.7 mEq/L | 0
total protein 4.8 g/dL | 0
albumin 2.4 g/dL | 0
LDH 472 U/L | 0
HbA1c 9.8% | 0
PT 17.5 seconds | 0
INR 1.63 | 0
aPTT 52.8 seconds | 0
antithrombin III 70.5% | 0
FDPs 49.2 μg/mL | 0
fibrinogen 429.3 mg/dL | 0
urinalysis specific gravity 1.028 | 0
urinalysis pH 5.0 | 0
traces of protein | 0
10–19 WBCs per high power field | 0
0–1 RBCs per high power field | 0
sinus tachycardia | 0
KUB finding nonspecific | 0
contrast-enhanced abdominal CT | 0
focal wedge-shaped perfusion defect in the upper pole of right kidney | 0
no evidence of intravascular filling defect in renal vessels | 0
Escherichia coli isolated from blood and urine cultures | 0
right acute pyelonephritis | 0
sepsis | 0
intravenous ceftriaxone 2 g per day | 0
mental status became drowsy | 120
blood pressure fell to 80/60 mmHg | 120
fever developed | 120
chest X-ray increased haziness on both lower lung fields | 120
WBC count 27800/μL | 120
platelet count 26000/μL | 120
Cr 0.8 mg/dL | 120
chest CT scan | 120
passive atelectasis in both lungs | 120
no evidence of pneumonia | 120
echocardiography | 120
decreased cardiac wall motion | 120
left ventricular dysfunction | 120
ejection fraction 47% | 120
no evidence of thrombus in cardiac chambers | 120
septic shock | 120
acute heart failure | 120
diuretics | 120
inotropes | 120
antibiotics changed to piperacillin and tazobactam | 120
clinical course gradually improved | 120
sudden onset of severe right flank pain | 312
tenderness | 312
urinalysis 1–4 WBCs per high power field | 312
urinalysis 5–9 RBCs per high power field | 312
LDH 1768 U/L | 312
abdominal CT | 312
large perfusion defect in the upper to mid portion of the right kidney | 312
intravascular filling defect in the right renal artery | 312
PT 12.3 seconds | 312
INR 1.14 | 312
aPTT 23.8 seconds | 312
antithrombin III 84.7% | 312
FDP 19.5 μg/mL | 312
fibrinogen >500 mg/dL | 312
factor assay V 81% | 312
proteins C normal | 312
proteins S normal | 312
lupus anticoagulant Ab not found | 312
flank pain resolved | 384
hematuria disappeared | 384
follow-up abdominal CT | 384
perfusion defect partially regressed | 384
right renal artery thrombus partially regressed | 384
discharged | 528
