66 years old | 0
male | 0
admitted to the hospital | 0
dyspnoea on exertion | -720
orthopnoea | -720
paroxysmal nocturnal dyspnoea | -720
unintentional weight loss | -720
blood pressure 103/81 mmHg | 0
heart rate 90 b.p.m. | 0
respiratory rate 20 b.p.m. | 0
oxygen saturation 98% | 0
elevated jugular venous pressure | 0
bilateral peripheral oedema | 0
pansystolic murmur | 0
third heart sound | 0
bilateral crackles | 0
elevated N-terminal pro-brain natriuretic peptide | 0
normal troponin I | 0
sinus rhythm | 0
left axis deviation | 0
inferior Q-waves | 0
no ST changes | 0
dilated left and right ventricles | 0
moderate mitral and tricuspid regurgitation | 0
pulmonary artery systolic pressure 34 mmHg | 0
estimated mean right atrial pressure 10-15 mmHg | 0
masses in both apices | 0
masses in the right atrium | 0
type B thrombi | 0
cardiac magnetic resonance imaging | 48
ischaemic scars | 48
intracardiac masses | 48
high signal intensity on T1- and T2-weighted sequences | 48
low-signal on first pass imaging following gadolinium administration | 48
LV and RV end-diastolic volumes | 48
LVEF 19% | 48
RVEF 20% | 48
fluid overload | 48
small bilateral pleural effusions | 48
IVC diameter 29 mm | 48
near full thickness scars | 48
severe triple vessel disease | 192
occlusion of the left circumflex and right coronary arteries | 192
severe stenosis of the mid-left anterior descending artery | 192
elevated liver enzymes | 0
hyperbilirubinemia | 0
prolonged prothrombin time | 0
prothrombin ratio | 0
activated partial thromboplastin time | 0
warfarin therapy | 0
lisinopril 10 mg daily | 240
frusemide 40 mg daily | 240
carvedilol 12.5 mg twice daily | 240
discharged home | 240
out of hospital cardiac arrest | 672
percutaneous coronary intervention | 720
implantable cardioverter defibrillator inserted | 720
patient discharged home | 864
complete resolution of intracardiac masses | 720
LVEF 22% | 720
RVEF 46% | 720