18 years old | 0
male | 0
admitted to the hospital | 0
fever | 0
rash | 0
acne | -672
minocycline | -672
increased WBC count | 0
eosinophilia | 0
systemic involvement | 0
diffuse erythematous or maculopapular eruption | 0
pruritis | 0
DRESS syndrome | 0
fever persisted | 0
rash persisted | 0
discharged | 24
left lower quadrant abdominal pain | -672
pelvic heaviness | -672
urinary frequency | -672
tubal ligation | -672
active smoker | -672
large and painful mass | -672
pelvic MRI | -672
mass measuring 18 × 17 × 12 cm | -672
well-delimited, polylobed, poorly vascularized, with central fluid component | -672
located on the left ovary, extending up to the umbilicus | -672
no lymphadenopathy, ascites or peritoneal implants | -672
uterus and adnexa were normal | -672
serum tumor markers were negative | -672
surgical pelvic exploration | -672
30-centimeter mass of the left broad ligament | -672
no ascites or peritoneal carcinomatosis | -672
uterus and right adnexa were normal | -672
total hysterectomy with adnexectomy and removal of the mass | -672
leiomyosarcoma | -672
isolated fever of 39 °C | 2
major inflammatory syndrome | 2
leukocytes 15,000/μL | 2
C-reactive protein 317 mg/dL | 2
contrast-enhanced computed tomography scan of the abdomen and pelvis | 2
bilobed air and fluid collection | 2
abscess, located in the retroperitoneum and extending along the left psoas muscle | 2
sudden drop in blood pressure | 2
vasopressor therapy | 2
noradrenaline | 2
blood pressure stabilization | 2
emergency revision surgery | 2
peritoneal cavity exploration | 2
moderately abundant non-purulent serosanginous peritoneal fluid | 2
adhesions to the Douglas pouch | 2
peritonitis | 2
antibacterial treatment with piperacillin/tazobactam and gentamicin | 2
microbiological samples were taken | 2
extubated in the postoperative recovery room | 2
hemodynamic support with noradrenaline | 2
transferred to the intensive care unit | 2
clinical improvement | 2
decrease in inflammatory markers | 2
noradrenaline requirement decreased | 3
noradrenaline discontinued | 3
microbiological analysis of the peritoneal fluid | 2
Gardnerella vaginalis | 2
gentamicin discontinued | 2
metronidazole added | 2
Atopobium vaginae | 4
preoperative blood cultures remained sterile | 2
antibacterial susceptibility testing of Garderella vaginalis | 2
resistance to metronidazole and ciprofloxacin | 2
susceptibility to penicillin G, amoxicillin/clavulanate, cefotaxim, clindamicin and vancomycin | 2
antibacterial susceptibility testing of Atopobium vaginae | 4
susceptibility to all tested antibacterials, including metronidazole | 4
piperacillin/tazobactam was active against both bacteria | 2
final diagnosis | 2
early postoperative peritonitis-induced septic shock caused by Gardnerella vaginalis and Atopobium vaginae | 2
discharged from the intensive care unit | 5
antibacterial therapy was stopped | 7