31 years old | 0\
female | 0\
SLE | -8760\
lupus nephritis | -8760\
stroke | -8760\
intravenous drug use | -8760\
cardiogenic shock | 0\
mental status changes | 0\
elevated jugular venous pressure | 0\
prominent v wave | 0\
body temperature 36.3°C | 0\
blood pressure 95/66 mm Hg | 0\
heart rate 94 beats/min | 0\
hemoglobin 10.3 g/dL | 0\
white blood cell count 18.9 × 10^9/L | 0\
platelet count 64 × 10^9/L | 0\
international normalized ratio 3.6 | 0\
creatinine level 1.7 mg/dL | 0\
drug studies positive for narcotics | 0\
drug studies positive for cannabis | 0\
negative antiphospholipid serology | 0\
negative blood cultures | 0\
dehisced mitral valve prosthesis | 0\
severe mitral regurgitation | 0\
intervalvular fibrosa dehiscence | 0\
cavity at the intervalvular fibrosa | 0\
loculated cavity | 0\
perivalvular regurgitation | 0\
mitral valve prosthesis displaced to the mid atrium | 0\
two dominant jets of periprosthetic regurgitation | 0\
posterior annulus dehiscence | 0\
pseudoaneurysm | 0\
fourth sternotomy | 24\
mitral valve annulus reconstruction | 24\
integration of 33-mm bioprosthesis | 24\
reconstruction of the left atrial dome | 24\
reconstruction of the interatrial septal incision | 24\
well-seated mitral valve bioprosthesis | 24\
mean gradient 3 mm Hg | 24\
no regurgitation | 24\
extracorporeal membrane oxygenation | 24\
multiple blood product transfusions | 24-48\
layered thrombus in the left atrium | 120\
surgical clot removal | 120\
thrombus reaccumulation | 120\
withdrawal of extracorporeal membrane oxygenation support | 120\
death | 120