38 weeks gestational age | 0
female | 0
birth weight 3.2 kg | 0
born to a 26-year-old primigravida mother | 0
cesarean section | 0
breech presentation | 0
fine until the age of 15 days | -360
developed signs of respiratory distress | -336
tachypnea | -336
fever | -336
feeding refusal | -336
admitted to the neonatal intensive care unit | -336
provisional diagnosis pneumonia | -336
provisional diagnosis septicemia | -336
left lung consolidation | -336
right lung cysts | -336
oxygen therapy | -336
intra-venous antibiotics | -336
chest X-ray performed | -288
aggravating cystic lesions in the right lung | -288
referred to our hospital | -288
admitted to our neonatal intensive care unit | -288
mild respiratory distress | -288
family members COVID-19-positive | -672
nasopharyngeal swab for SARS‐CoV‐2 RNA | -288
positive SARS‐CoV‐2 RNA | -264
tachypnea | -264
respiratory rate 72 breaths/min | -264
subcostal/intercostal retractions | -264
absent breath sounds on the right side of the chest | -264
heart sounds better audible on the right side | -264
normal white blood cells count | -264
Hb level 13 gm/dL | -264
blood gas analysis | -264
pH 7.25 | -264
pO2 55 | -264
bicarbonate 18 | -264
base deficit 4 | -264
pCo2 55 | -264
O2 Saturation 90-95% | -264
nasal flow cannula | -264
chest X-ray | -264
chest tomography | -264
left lung opacities | -264
left lung consolidation | -264
right cystic lesions | -264
diagnosis of congenital pulmonary airway malformation | -264
echocardiogram | -264
normal echocardiogram | -264
blood culture | -264
sterile blood culture | -264
multidisciplinary team discussion | -264
decision to monitor closely | -264
indication of surgical resection | -264
low-flow nasal oxygen | -264
50% fraction of inspired oxygen | -264
intravenous antibiotics | -264
clinical improvement | -216
taken off oxygen | -216
signs respiratory distress disappeared | -216
normal feeding resumed | -216
discharge | -216
out-patient follow-up | 576
reassessment | 576
control chest-CT | 576
complete resolution of cystic lesions | 576
post-pneumonia healing changes | 576