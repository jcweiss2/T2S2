28 years old | 0
female | 0
gravida 1 | 0
para 0 | 0
singleton pregnancy | 0
conceived through in vitro fertilization and embryo transfer | 0
referred to hospital | 0
10 weeks of gestation | -560
no prior chorionic villous sampling | -560
no amniocentesis | -560
sudden uterine contraction | -72
genital bleeding | -72
watery discharge | -72
speculum examination | -72
watery discharge with a small amount of blood | -72
test for monoclonal antibodies against insulin-like growth factor-binding protein 1 positive | -72
premature rupture of the membrane suspected | -72
clinical chorioamnionitis diagnosed | -72
temperature over 38 °C | -72
tachycardia | -72
uterine tenderness | -72
intravenous ampicillin and gentamicin started | -72
amniocentesis performed | -72
blood and vaginal discharge cultures examined | -72
elevated white blood cell count | -72
elevated C-reactive protein level | -72
amniotic fluid showed numerous inflammatory cells | -72
Candida glabrata in amniotic fluid | -72
Candida glabrata in vaginal discharge | -72
persistent temperature over 38 °C | -48
blood test for 1,3-β-D-glucan negative | -48
termination of pregnancy decided | -24
fever resolved after delivery | 72
delivery at 18 weeks and 5 days of gestation | 72
Candida glabrata detected in blood culture | 144
re-admitted | 144
intravenous fluconazole administered | 144
no fever | 144
no uterine tenderness | 144
no elevated inflammatory markers in blood | 144
no systemic candidiasis | 144
chorioamnionitis confirmed by histological examination | 144
maternal inflammatory response stage II, grade I | 144
fetal inflammatory response stage I, grade I | 144
Candida spp. identified by Grocott-Gomori methenamine silver stain | 144