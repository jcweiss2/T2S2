65 years old | 0 | 0 
female | 0 | 0 
admitted to the hospital | 0 | 0 
stage IIIA lung cancer | -648 | -648 
smoking history | -648 | 0 
hypertension | -648 | 0 
hypothyroidism | -648 | 0 
dyslipidemia | -648 | 0 
spiculated suprahilar RUL nodule | -648 | -648 
lung-RADS 4X | -648 | -648 
PET/CT scan | -648 | -648 
bronchoscopy | -648 | -648 
NSCLC | -648 | -648 
adenocarcinoma | -648 | -648 
lymph node sampling | -648 | -648 
surgical resection | -648 | -648 
carboplatin | -216 | -168 
paclitaxel | -216 | -168 
radiation therapy | -216 | -168 
CT scan | -120 | -120 
adjuvant immunotherapy | -84 | -56 
durvalumab | -84 | -56 
pneumonitis | -56 | -56 
steroid taper | -56 | -28 
staging chest CT | -28 | -28 
RUL mass increase | -28 | -28 
follow-up chest CT | 0 | 0 
abdominal pain | 0 | 0 
pancreatic head lesion | 0 | 0 
abdominal and pelvic CT scan | 0 | 0 
constipation | 0 | 0 
loss of appetite | 0 | 0 
weight loss | 0 | 0 
epigastric pain | 0 | 0 
endoscopic ultra-sound-guided biopsy | 0 | 0 
pancreatic mass | 0 | 0 
tumor cells | 0 | 0 
CK7 | 0 | 0 
TTF-1 | 0 | 0 
Napsin-A | 0 | 0 
CDX-2 | 0 | 0 
KOC | 0 | 0 
synaptophysin | 0 | 0 
Smad-4 | 0 | 0 
lung adenocarcinoma | 0 | 0 
metastasized to the pancreas | 0 | 0 
liver enzymes | 0 | 0 
AST | 0 | 0 
ALT | 0 | 0 
ALP | 0 | 0 
total bilirubin | 0 | 0 
direct bilirubin | 0 | 0 
CA 19.9 | 0 | 0 
PET/CT scan | 24 | 24 
brain MRI scan | 24 | 24 
palliative radiation therapy | 168 | 168 
carboplatin | 168 | 168 
pemetrexed | 168 | 168 
chemotherapy | 168 | 168 
generalized weakness | 168 | 168 
dyspnea | 168 | 168 
electrolyte derangements | 168 | 168 
acute anemia | 168 | 168 
hemoglobin nadir | 168 | 168 
transfusion | 168 | 168 
CT scan of the chest | 168 | 168 
new left lower lobe nodule | 168 | 168 
staging PET/CT scan | 240 | 240 
metabolic activity | 240 | 240 
treatment continuation | 240 | 240 
pulmonology clinic | 288 | 288 
rapid response | 288 | 288 
oxygen supplementation | 288 | 288 
bilevel-positive airway pressure | 288 | 288 
broad-spectrum antibiotics | 288 | 288 
vancomycin | 288 | 288 
azithromycin | 288 | 288 
cefepime | 288 | 288 
acute hypoxic respiratory failure | 288 | 288 
sepsis | 288 | 288 
pneumonia | 288 | 288 
altered mentation | 288 | 288 
worsening hypoxemia | 288 | 288 
vasopressor support | 288 | 288 
palliative medicine team | 288 | 288 
inpatient hospice care | 288 | 288 
death | 288 | 288