46 years old | 0
African American | 0
male | 0
admitted to the hospital | 0
uncontrolled diabetes mellitus | -672
hypertension | -672
chronic kidney disease | -672
polysubstance abuse | -672
alcohol abuse | -672
tobacco abuse | -672
marijuana abuse | -672
cocaine abuse | -672
confusion | 0
difficulty speaking | 0
temperature 37.6 | 0
blood pressure 154/93 | 0
oriented to self | 0
expressive aphasia | 0
non-fluent speech | 0
impaired naming | 0
impaired repetition | 0
good comprehension | 0
dysarthria | 0
right-sided hemiparesis | 0
leukocytosis | 0
computer tomography | 0
left thalamic mass | 0
midline shift | 0
magnetic resonance imaging | 0
empiric intravenous antimicrobial therapy | 0
vancomycin | 0
meropenem | 0
stereotactic aspiration | 0
purulent material | 0
Gram stain | 0
Gram positive cocci | 0
Streptococcus anginosus | 0
negative blood cultures | 0
transthoracic echocardiogram | 0
no valvular vegetations | 0
computer tomography imaging | 0
sigmoid colitis | 0
ceftriaxone | 24
switched antibiotic regimen | 24
left against medical advice | 360
outpatient follow-up | 720
persistent hemiparesis | 720
no documentation of aphasia | 720