33 years old | 0
unmarried | 0
nullipara | 0
family history of brother with testicular cancer | 0
explorative laparoscopy | -43800
nonspecific abdominal pain | -43800
gelatinous tumor spread detected | -43800
biopsy specimens confirming disseminated peritoneal adenomucinosis (DPAM) | -43800
peritoneal lesions originated from perforated mucinous cystadenoma of the appendix | -43800
advised peritonectomy | -43800
advised bilateral oophorectomy | -43800
referred for fertility preservation consultation | -43800
decided to undergo IVF and embryo cryopreservation | -43800
20 oocytes retrieved | -43800
18 embryos fertilized with donor sperm | -43800
embryo cryopreservation at 2 pronuclear stage | -43800
PMP surgery performed by multidisciplinary team | -43800
extended spread of disease in Douglas pouch | -43800
disease over omentum | -43800
disease underneath diaphragm | -43800
disease over spleen | -43800
two large masses on both ovaries | -43800
mass on appendix | -43800
lesions over surface of uterus | -43800
parietal peritoneum resected | -43800
omentectomy | -43800
appendectomy | -43800
splenectomy | -43800
bilateral adnexectomy | -43800
lesions peeled off over uterus | -43800
uterus left intact | -43800
postoperative heated intraperitoneal infusions of mitomycin C | -43800
disease relapse 18 months later | 12960
moderate elevation of carcinoembryonic antigen (CEA) | 12960
intra-abdominal fluid accumulation | 12960
multiple peritoneal lesions by CT | 12960
explorative laparotomy | 12960
numerous small lesions over peritoneum | 12960
lesion over left diaphragm | 12960
lesion over posterior wall of uterus | 12960
cytoreduction | 12960
peritonectomy | 12960
