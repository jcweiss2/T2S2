71 years old | 0
woman | 0
admitted | 0
left flank pain | 0
oliguria | 0
hypotension | 0
pyuria | 0
severe sepsis | 0
acute pyelonephritis | 0
abdominal computed tomography intravenous pyelogram | 0
normal-sized kidneys | 0
poorly determined differentiation between cortex and medulla | 0
left kidney amorphic low attenuation lesion | 0
acute pyelonephritis (Fig. 1A) | 0
incompletely malrotated kidneys | 0
anteriorly facing hila | 0
laterally located renal vessels and ureter | 0
right kidney 5 cm lower than left kidney |-24
renal ectopia | 0
mild dilation at proximal ureter of left kidney | 0
three-dimensional computed tomography reconstruction image | 0
anteriorly rotated kidneys (Fig. 1B) | 0
piperacillin-tazobactam | 0
cefotaxime | 0
E. coli infection in bloodstream | 0
improved hemodynamic state | 72
released from intensive care unit | 72
malrotation of kidney | 0
partial obstruction of ureteropyelic junction | 0
increased incidences of urolithiasis and infection | 0
dilated left ureter | 0
mild obstruction due to ureteral deformation and renal malrotation | 0
recurrent urinary tract infections | -168
septic shock | 0
Wait, there's an error in the line: "right kidney 5 cm lower than left kidney |-24". That should be at 0, as it's part of the CT findings during admission. Correcting that:
right kidney 5 cm lower than left kidney | 0
partial obstruction of ureteropyelic junction |
