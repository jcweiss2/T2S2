48 years old | 0
female | 0
admitted to the hospital | 0
ERCP | 0
sphincter of Oddi dysfunction | 0
recent acute pancreatitis | -72
episodic abdominal pain | -72
Lehman perfusion aspiration manometry catheter | 0
common bile duct cannulated | 0
pancreatic duct cannulated | 0
basal sphincter pressures measured | 0
cholangiography | 0
pancreatography | 0
cystic duct cannulated | 0
cholecystokinin infusion | 0
bile aspirated | 0
microlithiasis analysis | 0
mild post-procedure discomfort | 0
chest pain | 2
white blood cell count 14.5 × 1,000/μL | 2
hematocrit 32.9% | 2
aspartate aminotransferase (AST) 176 U/L | 2
alanine aminotransferase (ALT) 32 U/L | 2
total bilirubin 0.46 mg/dL | 2
serum lipase 93 U/dL | 2
serum troponin 2.3 ng/mL | 2
non-ST elevation myocardial infarction | 2
medically treated | 2
abdominal pain | 24
peritoneal signs | 24
AST 250 U/L | 24
ALT 55 U/L | 24
total bilirubin 3.34 mg/dL | 24
direct bilirubin 2.85 mg/dL | 24
lipase 192 U/dL | 24
CT scan | 24
air in gallbladder | 24
air in lesser sac | 24
air in retroperitoneum | 24
air in intraperitoneal cavity | 24
air in bile duct | 24
loculated area of air in right hepatic lobe | 24
emphysematous cholecystitis | 24
bowel perforation suspected | 24
broad spectrum antibiotics | 24
ampicillin/sulbactam | 24
laparotomy | 48
gangrenous gallbladder | 48
cholecystectomy | 48
no gallstones | 48
common hepatic duct inflamed | 48
possible gangrene | 48
histopathologic examination | 48
gangrenous cholecystitis | 48
gram-positive rods | 48
gallbladder wall | 48
cultures from gallbladder | 48
Clostridium perfringens | 48
cultures from blood | 48
discharged home | 168
abdominal pain | 192
fever | 192
CT scan | 192
liver abscesses | 192
percutaneous drainage catheter | 192
bilious fluid | 192
cholangiography | 192
communication between abscess and left intrahepatic biliary system | 192
extravasation of contrast | 192
disruption of intrahepatic ducts | 192
necrosis of intrahepatic ducts | 192
trans-hepatic 8F locking loop draining catheter | 192
antibiotics | 192
supportive measures | 192
CHD drain exchanged | 216
internal external percutaneous drain | 216
discharged home | 216
abdominal pain | 504
fever | 504
septic shock | 504
broad spectrum antibiotics | 504
supportive measures | 504
revision of biliary drain catheters | 504
recurrent hospital admissions | 1008
cholangitis | 1008
hepatic abscesses | 1008
sepsis | 1008
Enterococcus | 1008
Pseudomonas | 1008
Klebsiella | 1008
Candida | 1008
hypotension | 1008
renal failure | 1008
respiratory failure | 1008
percutaneous drains | 1008
antibiotics | 1008
supportive care | 1008
ERCP | 1296
multiple strictures | 1296
beading in intra- and extra-hepatic biliary tree | 1296
biliary stents | 1296
placement and exchange of biliary stents | 1296
sclerosing cholangitis | 1296
end-stage liver disease | 1296
living donor liver transplantation | 1814
explant histopathology | 1814
secondary biliary cirrhosis | 1814
bile duct necrosis | 1814
fungal hyphae | 1814
bacterial organisms | 1814
normal hepatobiliary function | 2592
feeling well | 2592