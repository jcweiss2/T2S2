23 weeks gestational age | -672
female | -672
HELLP syndrome | -672
cesarean section | 0
birthweight 485 grams | 0
Apgar scores 3 at 1 minute | 0
Apgar scores 8 at 5 minutes | 0
intubated | 0
received surfactant | 0
mechanical ventilation | 0
white blood cells 2.1×10^9/L | 0
hematocrit 39.6% | 0
hemoglobin 12.6 g/100 mL | 0
platelet 186×10^3 mL | 0
differential 9% segmental WBC | 0
differential 1% bands | 0
differential 60% lymphocytes | 0
differential 26% monocytes | 0
603 nucleated red blood cells per 100 WBC | 0
C-reactive protein less than 0.3 mg/dL | 0
neutropenia | 0
thrombocytopenia | 0
bandemia | 0
hemodynamically significant hypotension | 0
vasopressors | 0
ampicillin | 0
gentamicin | 0
blood sample sent for culture | 0
anaerobic gram-positive branching rods | 96
Actinomyces species | 96
ampicillin switched to penicillin | 96
penicillin | 96
antimicrobial course of therapy | 0
subsequent blood culture had no growth | 120
Actinomyces viscosus | 624
16S ribosomal RNA gene sequencing | 624
Matrix-assisted laser desorption ionization-time of flight spectrometry | 624
persistent neutropenia | 0
persistent thrombocytopenia | 0
disseminated intravascular coagulation | 0
transient hypoglycemia | 0
electrolyte imbalance | 0
adrenal insufficiency | 0
acute renal failure | 0
endotracheal aspirate grew Staphylococcus aureus | 744
urine culture grew Enterococcus faecalis | 744
central line grew Staphylococcus epidermidis | 744
vancomycin | 744
ampicillin/sulbactam | 744
discharged | 2160