26 years old | 0
    male | 0
    no medical history | 0
    no family history of cancer | 0
    presented to local hospital | 0
    abdominal pain | 0
    night sweats | 0
    fever | 0
    intra-abdominal mass | 0
    referred to our centre | 0
    low-grade sarcoma | 0
    mixed epithelioid and spindle cell morphology | 0
    mucin 4-positive tumour | 0
    EWSR1 gene rearrangement | 0
    Sclerosing epithelioid fibrosarcoma (SEF) | 0
    extensive peritoneal carcinomatosis | 0
    doxorubicin-ifosfamide chemotherapy | 0
    maximum response of stable disease | 0
    radiological evidence of disease progression | -144
    clinical evidence of disease progression | -144
    cytoreductive surgery (CRS) | -96
    hyperthermic intraperitoneal chemotherapy (HIPEC) | -96
    cisplatin | -96
    doxorubicin | -96
    intravenous ifosfamide | -96
    remission | -72
    recurrence | -36
    CRS | -36
    HIPEC | -36
    remission | 0
    recurrence | 48
    gemcitabine | 48
    docetaxel | 48
    radiological progression | 72
    symptomatic treatment recommended | 72
    admitted with symptomatic COVID-19 | 216
    multiple enterocutaneous fistulas | 216
    nil-by-mouth status | 216
    parenteral nutrition | 216
    PET revealed further disease progression | 216
    multiple admissions to ICU | 288
    sepsis | 288
    intra-abdominal collections | 288
    trial of nivolumab | 336
    no clinical response | 336
    presented to molecular tumour board | 360
    next-generation sequencing (NGS) | 360
    ALK mutation | 360
    ALK inhibitor crizotinib | 360
    CT abdomen and pelvis showed disease progression | 360
    crizotinib 250 mg started | 432
    CT abdomen and pelvis showed significant size regression | 456
    hepatic metastases | 456
    no new metastatic lesions | 456
    further clinical improvement in tumour response | 480
    delayed third cycle due to grade 3 haematological toxicity | 528
    fatigue | 528
    third cycle administered at 200 mg | 528
    reduced dose of crizotinib | 528
    medically stable | 528
    moderate health | 528
    significant reduction in tumour size | 528
    enterocutaneous fistulas improvement | 528
    