61 years old | 0  
    male | 0  
    continuous high-grade intermittent fever | -192  
    chills | -192  
    rigor | -192  
    hiccup | -192  
    nausea | -24 to -48  
    breathlessness | -24  
    hypertension | -113568  
    cerebrovascular accident | -113568  
    right-sided hemiparesis | -113568  
    atenolol | -113568  
    amlodipine | -113568  
    amiloride | -113568  
    aspirin | -113568  
    confused | 0  
    temperature 104°F | 0  
    pulse 110/min | 0  
    blood pressure 130/80 mmHg | 0  
    respiration rate 40/min | 0  
    SPO2 96% | 0  
    pallor | 0  
    normal blood sugar | 0  
    ultrasonography of whole abdomen | 0  
    increased serum urea (76 mg/dl) | 0  
    increased serum creatinine (3.2 mg/dl) | 0  
    increased serum glutamic oxaloacetic transaminase (40 IU/L) | 0  
    increased serum glutamic pyruvic transaminase (49 IU/L) | 0  
    increased total leukocytic count (10600) | 0  
    negative tests for Plasmodium vivax | 0  
    negative tests for Plasmodium falciparum | 0  
    negative tests for Hepatitis C Virus | 0  
    negative tests for Australian antigen | 0  
    sepsis | 0  
    acute renal failure | 0  
    ceftriaxone | 0  
    tazobactam | 0  
    arteether 150 mg i.v. | 0  
    no relief in symptoms | 96  
    increased serum urea | 96  
    increased serum creatinine | 96  
    normal urine output | 96  
    teicoplanin | 120  
    meropenem | 120  
    hemodialysis | 144  
    symptoms start abated | 168  
    serum urea 116 mg/dl | 168  
    serum creatinine 4.3 mg/dl | 168  
    TLC 11900/cumm | 168  
    serum urea 168 mg/dl | 240  
    serum creatinine 4.34 mg/dl | 240  
    TLC 21600/cumm | 240  
    stopped ceftriaxone | 240  
    stopped tazobactam | 240  
    stopped arteether | 240  
    furosemide 40 mg twice daily | 240  
    torsemide 20 mg twice daily | 240  
    metolazone 5 mg once daily | 240  
    cefotaxime 1 g twice daily | 240  
    hemodialysis once every 3–4 days | 240  
    TLC 31000 | 288  
    serum urea 219 mg/dl | 288  
    serum creatinine 4.64 mg/dl | 288  
    hemodialysis | 288  
    decreased urea and creatinine | 288  
    increased urea and creatinine | 288  
    tigecycline 50 mg twice daily | 408  
    caspofungin 50 mg once daily | 576  
    TLC decreased | 696  
    doripenem 250 mg twice daily | 696  
    TLC 11000/cumm | 840  
    stopped all antibiotics | 840  
    serum urea 400 mg/dl | 840  
    serum creatinine 3.6 mg/dl | 840  
    chronic renal failure | 840  
    dialysis at regular intervals | 840  
    stopped torsemide | 984  
    stopped metolazone | 984  
    serum urea 208 mg/dl | 1008  
    serum creatinine 2.2 mg/dl | 1008  
    stopped furosemide | 1032  
    decreased serum urea | 1032  
    decreased serum creatinine | 1032  
    normal TLC 7700/cumm | 1440  
    normal urea 27 mg/dl | 1440  
    normal creatinine 1.1 mg/dl | 1440  
    dialysis not required | 1440  
