13 years old | 0
male | 0
atopic dermatitis | -672
not fully vaccinated | 0
admitted to the hospital | 0
progressive fatigue | -96
hypoactivity | -96
slurred speech | -48
lower extremity weakness | -96
multiple episodes of choking | -48
urinary incontinence | -48
fecal incontinence | -48
difficulty breathing | 0
drooling of saliva | 0
ascending weakness | 0
inability to bear weight | 0
conscious | 0
alert | 0
pale | 0
hypoactive | 0
T: 36.4 | 0
P: 110 | 0
SBP: 70 | 0
cold extremities | 0
poor perfusion | 0
respiratory distress | 0
Silverman score 5/10 | 0
Saturation: 89 | 0
bilateral decreased air entry | 0
diffuse crackles | 0
GCS was 15/15 | 0
decreased in motor power bilaterally in lower limbs | 0
absent deep tendon reflexes | 0
negative Babinski reflex | 0
septic shock | 0
IV fluid boluses | 0
systolic blood pressure became 100 | 0
arterial blood gases showed hypoxemia | 0
metabolic acidosis | 0
chest x-ray revealed right upper lobe collapse | 0
pneumonia with diffuse infiltrates in both lung fields | 0
early ARDS | 0
non-invasive ventilation | 0
decreasing level of consciousness | 12
urgent CT scan of brain | 12
no bleeding or any mass | 12
intubated | 12
mechanical ventilation | 12
urgent MRI Brain | 12
normal | 12
broad spectrum antibacterial stat doses | 12
transferred to the pediatric intensive care unit | 12
WBC 6000 | 12
Bands 29 | 12
Neutrophils 47 | 12
Lymphocytes 13 | 12
elevated inflammatory markers | 12
CRP: 22 | 12
ESR: 110 | 12
disseminated intravascular coagulopathy | 12
Platelets: 57,000 | 12
INR: 1.4 | 12
Fibrinogen: 456 | 12
D-dimer: 0.36 | 12
Guillain-Barre syndrome | 12
IVIG | 12
blood cultures were positive for Streptococcus pneumonia | 48
Mycoplasma pneumonia serology negative | 48
nasal wash for influenza negative | 48
severe ARDS | 96
hypoxia | 96
respiratory acidosis | 96
deteriorating condition | 96
died | 96