57 years old | 0
female | 0
admitted to the hospital | 0
generalized anxiety disorder | -672
choreiform movements | -180
oral and vaginal bleeding | 0
anxiety worsening | -168
diagnosed with chorea | -46
levetiracetam | -46
VPA | -21
traumatic subacute right frontoparietal subdural hematoma | -504
methicillin-susceptible Staphylococcus aureus bacteremia | -504
Glasgow Coma Scale (GCS) 15 | -504
choreiform type movements | -504
involuntary movements started | -180
family history of abnormal movements | -180
clonazepam | -504
levetiracetam 250 mg twice daily | -504
valproic acid 250 mg 3 times daily | -21
platelet count 139 000 μL | -504
platelet count 90 000 μL | -21
discharged | -483
GCS 15 | -483
platelet count 122 000 μL | -483
blood pressure 131/91 mm Hg | 0
heart rate 120 beats/min | 0
respiratory rate 16 breaths/min | 0
temperature 36.5°C | 0
GCS 15 | 0
atraumatic contusions and ecchymosis | 0
CT head without contrast | 0
left temporal frontal subdural hematoma | 0
acute subdural hematoma | 0
mass effect on the right lateral ventricle | 0
midline shift | 0
white blood cells 14.6×10^6/µL | 0
red blood cells 2.75×10^6/µL | 0
platelets 4000/μL | 0
hemoglobin 7.3 g/dL | 0
hematocrit 23.1% | 0
prothrombin time (PT) 15.7 secs | 0
partial thromboplastin time (PTT) 30.4 s | 0
fibrinogen 467 mg/dL | 0
VPA level 26.3 μg/mL | 0
valproic acid held | 0
thrombocytopenia | 0
heparin-induced thrombocytopenia | 0
heparin-platelet factor 4 (heparin-PF4)-related antibody | 0
serotonin release assay | 0
VPA level <10 μg/mL | 24
fibrinogen level 367 mg/dL | 24
hemoglobin 5.3 g/dL | 24
repeat CT of the head | 24
methylprednisolone 60 mg intravenous 3 times daily | 24
intravenous immune globulin 1 g/kg | 96
VPA discontinued | 0
clonazepam not re-initiated | 0
levetiracetam continued | 0
platelet counts improved | 504
hospitalized for 21 days | 504
altered mental status | 504
urinary tract infection | 504
Escherichia coli bacteremia | 504
sepsis | 504
discharged | 504
platelet count 108 000 | 504
GCS 14 | 504