64 years old | 0
male | 0
hypertension | -25920
arthritis | -25920
seizure disorder | -25920
Parkinson's disease | -25920
hiatal hernia | -25920
chronic anemia | -25920
non-bloody vomiting | -2160
non-bilious vomiting | -2160
decreased oral intake | -2160
progressive generalized weakness | -720
new-onset dyspnea | -720
dyspnea worsened | -24
not getting out of bed | -24
taking excessive NSAIDs | -720
chronic anemia | 0
gastritis | -26208
severe diverticulosis | -26208
1 cm tubular adenoma of the splenic flexure | -26208
hemorrhoids | -26208
blood pressure 65/30 mmHg | 0
heart rate 84 bpm | 0
oxygen saturation 96% on 4L oxygen | 0
afebrile | 0
ill-appearing | 0
labored breathing | 0
tachypnea (20-22 breaths per minute) | 0
decreased breath sounds on right lung | 0
mild ALT/AST elevations | 0
normal bilirubin | 0
white cell count 25.5 k/uL | 0
neutrophils 22.6 k/uL | 0
RBC 1.58 k/uL | 0
hemoglobin 2.3 g/dL | 0
hematocrit 10.9% | 0
platelets 652 u/L | 0
PT/INR 2.3 | 0
APTT 26 seconds | 0
lactate 13 ng/mL | 0
troponin 0.04 ng/mL | 0
sodium 141 mEq/L | 0
potassium 5.2 mEq/L | 0
chloride 107 mmol/L | 0
HCO3 13 mmol/L | 0
anion gap 21 | 0
glucose 114 mg/dL | 0
calcium 7.4 mg/dL | 0
creatinine 2.0 mg/dL | 0
eGFR 34 mL/min | 0
BUN 24 mg/dL | 0
protein 4.6 g/dL | 0
albumin 2.3 g/dL | 0
lactate dehydrogenase 774 units/L | 0
chest x-ray right-sided pneumothorax | 0
moderate right-sided pleural effusion | 0
compressive atelectasis of right lower lobe | 0
metabolic acidosis | 0
respiratory compensation | 0
high anion gap | 0
CT abdomen/pelvis sigmoid diverticulosis | 0
descending colon diverticulosis | 0
CT chest air and fluid in right pleural cavity | 0
volume resuscitation | 0
packed red blood cells | 0
transferred to intensive care | 0
blood cultures obtained | 0
sputum cultures obtained | 0
urine cultures obtained | 0
cefepime started | 0
chest tube placed | 0
drainage of 1L air | 0
drainage of purulent fluid | 0
respiratory status decline | 0
intubation | 0
pleural fluid straw color | 0
nucleated cell count 11,133/mm3 | 0
RBC 93,000/mm3 | 0
cloudy appearance | 0
pH 5.6 | 0
lymphocytes 2% | 0
monocytes/macrophages 7% | 0
segmented neutrophils 91% | 0
adenosine deaminase 7.3 | 0
lactate dehydrogenase 14,898 | 0
protein 3.1 g/dL | 0
glucose <2 mg/dL | 0
albumin 0.8 g/dL | 0
pleural fluid negative for malignant cells | 0
Candida tropicalis culture | 0
Candida glabrata culture | 0
Stenotrophomonas maltophilia culture | 0
broadened antibiotic coverage to meropenem | 0
caspofungin started | 0
polymicrobial flora | 0
elevated amylase >10,000 u/L | 0
esophageal tear suspected | 0
upper endoscopy 5-10 mm defect in posterior distal esophagus | 0
Boerhaave syndrome diagnosis | 0
gastric ulcers | 0
tissue fibrosis | 0
friability | 0
esophageal stenting | 0
biopsies obtained | 0
negative for malignant cells | 0
acute inflammation | 0
Candida species in biopsies | 0
ejection fraction 61% | 0
moderate to severe tricuspid regurgitation | 0
mitral regurgitation | 0
moderate pulmonary hypertension | 0
clinical improvement | 192
extubation | 192
CT-guided pigtail catheter placed | 192
pleural drainage | 192
decompensation | 216
Lactobacillus culture | 216
Staphylococcus lugdunensis culture | 216
antibiotic change to vancomycin | 216
ceftazidime | 216
metronidazole | 216
caspofungin | 216
worsening infiltrates bilaterally | 216
mediastinitis | 216
evolving ARDS | 216
re-intubation declined | 240
acute hypoxic respiratory failure | 240
death | 240
