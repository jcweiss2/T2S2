69 years old | 0  
    male | 0  
    paraumbilical hernia | -24  
    worsening abdominal distension | -24  
    diarrhoea | -24  
    weight loss | -24  
    lung fibrosis | 0  
    obstructive airway disease | 0  
    atrial fibrillation | 0  
    cardiomyopathy | 0  
    heart failure | 0  
    systemic sclerosis | 0  
    steroids | 0  
    methotrexate | 0  
    CT scan showing free air and fluid | -24  
    CT scan showing possible area of bowel necrosis | -24  
    admitted to the hospital | 0  
    cardiovascularly stable | 0  
    elevated CRP | 0  
    arterial lactate 1.2 mmol/L | 0  
    emergency laparotomy | 0  
    pockets of air on surface of small bowel | 0  
    short admission to intensive care | 0  
    prolonged stay on the ward | 0  
    ileus | 0  
    discharged | 0  
    oral antibiotics | 0  
    outpatient review with Rheumatology team | 0  
    systemic sclerosis as causative factor for PI | 0  
    represented one month later | 672  
    severe epigastric pain | 672  
    metabolic acidosis (pH 7.33) | 672  
    lactate of 4.6 mmol/L | 672  
    tachycardic (106 bpm) | 672  
    tachypneic (respiratory rate 34) | 672  
    normotensive | 672  
    white cell count 14 109/L | 672  
    haemoglobin 168 g/L | 672  
    creatinine 133 μmol/L | 672  
    INR 5.3 | 672  
    CT confirmed ongoing PI | 672  
    diffuse areas of hypoperfusion | 672  
    free air within the abdomen | 672  
    conservative approach | 672  
    p-possum score morbidity 99% | 672  
    p-possum score mortality 67.5% | 672  
    deteriorated | 672  
    pH 7.1 | 672  
    lactate 10.2 mmol/L | 672  
    decision to re-operate | 672  
    died | 672  
    post mortem findings confirmed small bowel perforation | 672  

