70 years old | 0
    female | 0
    lower abdominal pain | -24
    fever | -24
    nausea | -24
    vomiting | -24
    diaphoresis | -24
    right ovarian cyst | 0
    acute appendicitis | 0
    elective operation | 0
    hypertension | -43800
    congestive heart failure | -43800
    atrial fibrillation | -43800
    right coronary artery 90% stenosis | -43800
    digoxin | -43800
    dilatrend | -43800
    nitrate | -43800
    telmisartan | -43800
    thiazide | -43800
    AF with ventricular response 90-100 times/min | 0
    left ventricular hypertrophy | 0
    cardiomegaly | 0
    pleural effusion | 0
    ejection fraction 55% | 0
    left atrial enlargement | 0
    right atrial enlargement | 0
    eccentric hypertrophy | 0
    decreased mobility of the inferior wall of the left ventricle | 0
    moderate aortic valve insufficiency | 0
    aortic valve sclerosis | 0
    mild aortic stenosis | 0
    severe posterior mitral valve leaflet calcification | 0
    mitral valve width 1.92 cm2 | 0
    chronic cerebral infarction | 0
    dysarthria | 0
    dehydration | 0
    prerenal azotemia | 0
    FeNa 0.1% | 0
    serum creatinine 1.7 mg/dl | 0
    fluid therapy | 0
    serum creatinine 1.3 mg/dl | 0
    glycopyrrolate 0.2 mg IM | -0.5
    blood pressure 130/50 mmHg | 0
    ventricular response 90-100 times/min | 0
    arterial oxygen saturation 97% | 0
    right radial artery cannulation | 0
    induction of anesthesia | 0
    lidocaine 2 ml | 0
    propofol | 0
    remifentanil | 0
    unconscious | 0
    rocuronium 40 mg | 0
    endotracheal intubation | 0
    ventilation with 100% O2 | 0
    central venous catheterization | 0
    systolic BP 130-150 mmHg | 0
    diastolic BP 40-60 mmHg | 0
    ventricular response 100-110 times/min | 0
    CVP 8-9 mmHg | 0
    propofol effect site concentration 2.5-3.0 µg/ml | 0
    remifentanil effect site concentration 2.0 ng/ml | 0
    laparotomy | 0
    right ovary cystectomy | 0
    small bowel infarction | 0
    mesenteric arterial embolism | 0
    transesophageal echocardiography | 0
    spontaneous echo contrast (SEC) in left atrium | 0
    thrombus in left atrial appendage | 0
    segmental resection | 0
    intestinal anastomosis | 0
    hemodynamic stability | 0
    transferred to ICU | 0
    endotracheal tube | 0
    awareness confirmed | 0
    no neurologic disorder | 0
    extubation | 0
    low molecular weight heparin | 72
    warfarin | 120
    cardioversion | 672
    