10 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
Silver-Russell syndrome | -672 | 0 | Factual
Duchenne muscular dystrophy | -672 | 0 | Factual
birth weight 2100 g | -672 | -672 | Factual
birth length 48 cm | -672 | -672 | Factual
prominent forehead | -672 | 0 | Factual
relative macrocephaly | -672 | 0 | Factual
limb asymmetry | -672 | 0 | Factual
5th finger clinodactyly | -672 | 0 | Factual
2/3 toe syndactyly | -672 | 0 | Factual
hypomethylation of the 11p15 region | -504 | -504 | Factual
genetic examination | -504 | -504 | Factual
delayed motor development | -384 | 0 | Factual
hepatic dysfunction | -336 | -336 | Factual
increased alanine aminotransferase | -336 | -336 | Factual
increased aspartate aminotransferase | -336 | -336 | Factual
increased creatine kinase | -336 | -336 | Factual
genetic test | -252 | -252 | Factual
mutation of the maternal DMD gene | -252 | -252 | Factual
corticosteroids treatment | -192 | 0 | Factual
prednisone | -192 | -96 | Factual
deflazacort | -96 | 0 | Factual
G-CSF treatment | -72 | 0 | Factual
sepsis | -72 | -72 | Factual
hypoglycaemia | -72 | -72 | Factual
neurological symptoms | -72 | -72 | Factual
low glucose level | -72 | -72 | Factual
urological care | -72 | 0 | Factual
hypospadias | -72 | 0 | Factual
cardiological diagnostics | -12 | -12 | Factual
sinus tachycardia | -12 | -12 | Factual
heart murmur | -12 | -12 | Factual
propranolol | -12 | 0 | Factual
growth hormone deficiency | 0 | 0 | Negated
rhGH treatment | 0 | 18 | Factual
improved auxological parameters | 12 | 18 | Factual
increased height velocity | 12 | 18 | Factual
elevated IGF-1 | 12 | 18 | Factual
impaired glucose tolerance | 12 | 18 | Factual
insulin resistance | 12 | 18 | Factual
weight gain | 12 | 18 | Factual
reduced muscle mass | 12 | 18 | Factual
high content of fat tissue | 12 | 18 | Factual
discontinuation of rhGH therapy | 18 | 18 | Factual
progressive muscle weakness | 18 | 18 | Factual
low bone mineral density | 18 | 18 | Factual
scoliosis | 0 | 0 | Negated