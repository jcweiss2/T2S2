35 years old | 0
female | 0
pregnant | 0
admitted to the hospital | 0
fever | -240
cough | -240
dyspnoea | -120
aggravated dyspnoea | -120
cyanosis of the lip | 0
thick breathing sounds in both lungs | 0
dry and wet rales in the right lower lung | 0
tachycardia | 0
respiratory rate of 20 times/min | 0
COVID-19 infection | -240
S. aureus infection | -240
respiratory failure | 0
pregnancy with 34 + 4 wk | 0
G2P1 | 0
left occiput anterior | 0
elderly second parturient women | 0
maternal lower weight | 0
oligohydramnion | 0
premature live baby | 0
electrolyte disturbance | 0
hypoproteinaemia | 0
caesarean section | 24
oxyhemoglobin saturation decreased | 24
foetal distress | 24
dead foetus in utero | 24
oxygen therapy | 24
high-flow nasal cannula oxygen therapy | 24
fraction of inspired oxygen at 100% | 24
flow rate of 50 L/min | 24
improved oxyhemoglobin saturation | 48
assisted ventilation by endotracheal intubation | 48
empirical antibiotic therapy | 48
meropenem | 48
vancomycin | 48
symptomatic treatment | 48
metagenomic next-generation sequencing (mNGS) | 48
S. aureus detected | 48
2019-nCoV detected | 48
bacterial resistance gene test | 72
antibiotic resistance | 72
adjusted antibiotics | 216
sitafloxacin | 216
discharged from the hospital | 264
follow-up chest CT | 720
improved lung inflammation | 720
absorbed pleural effusion | 720