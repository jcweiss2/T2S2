56 years old | 0
    Hispanic | 0
    female | 0
    presented to the clinic | 0
    blurred vision | -336
    floaters | -336
    hospitalized in intensive care unit | -720
    septic shock | -720
    bilateral pneumonia | -720
    leptospirosis | -720
    elevated bilirubin | 0
    elevated liver enzymes | 0
    anemia | 0
    severe thrombocytopenia | 0
    platelet count of 37,000 | 0
    treated for Weil's disease | 0
    blood transfusions | 0
    intravenous ceftriaxone | 0
    retinal hemorrhages | -720
    visual loss | -720
    examination one month following initial diagnosis | 0
    visual acuity 20/200 OD | 0
    visual acuity 20/30 OS | 0
    intraocular pressure 14 OU | 0
    anterior segment quiet | 0
    2+ nuclear sclerosis noted bilaterally | 0
    sub-ILM hemorrhage concentrated in macula | 0
    dot hemorrhages in superior retina OD | 0
    retinal hemorrhage in macula OS | 0
    dot hemorrhages in superior and inferior retina OS | 0
    posterior vitreous detachment OU | 0
    OCT confirmed findings | 0
    fluorescein angiography confirmed findings | 0
    examined bi-weekly | 0
    no improvement in visual acuity | 0
    minimal hemorrhage resolution | 0
    sub-ILM hemorrhage surgically treated | 720
    pars-plana vitrectomy | 720
    internal limiting membrane removal | 720
    blood aspiration OD | 720
    improved BCVA 20/60 OD | 2400
    resolved dot hemorrhages OU | 2400
    last follow-up 8 months post vitrectomy | 8640
    BCVA remained 20/60 OD | 8640
    