3 years old | 0\
female | 0\
fever | -336\
diarrhea | -336\
abdominal pain | -336\
severe dehydration | -336\
tachypnea | -336\
rapid shallow breathing | -336\
hypotension | -336\
purpuric eruption | -336\
severe pancytopenia | -336\
absolute neutropenia | -336\
renal impairment | -336\
electrolyte imbalance | -336\
hyperuricemia | -336\
coagulopathy | -336\
disseminated intravascular coagulation | -336\
high inflammatory markers | -336\
positive stool culture for gram-negative Bacilli Escherichia coli | -336\
positive blood culture for gram-negative Bacilli Escherichia coli | -336\
intravenous fluid therapy | -336\
blood components transfusion | -336\
correction of electrolyte disturbance | -336\
antibiotic therapy | -336\
provisional diagnosis of acute infectious gastroenteritis with sepsis | -336\
severe dehydration | -336\
acute renal failure | -336\
disseminated intravascular coagulation | -336\
normal pelvi-abdominal ultrasound | -336\
hypocellular bone marrow | -336\
no abnormal cells in bone marrow | -336\
discharged | -336\
unexplained irritability | -168\
abnormal behavior | -168\
hallucinations | -168\
failure to recognize parents | -168\
thrombosis in both the left sigmoid and the transverse sinuses | -168\
normal coagulation profile | -168\
normal protein C and S | -168\
normal antithrombin III | -168\
initiation of low molecular weight heparin | -168\
improvement | -168\
discharged | -168\
fever | 0\
pallor | 0\
abdominal enlargement | 0\
leukocytosis | 0\
anemia | 0\
thrombocytopenia | 0\
blast cells in peripheral smear | 0\
hepatosplenomegaly | 0\
hypercellular bone marrow | 0\
blast cells in bone marrow | 0\
positive CD10 | 0\
positive CD20 | 0\
positive CD79a | 0\
diagnosis of Common ALL | 0\
induction therapy | 0\
consolidation therapy | 0\
positive factor XIII V34L mutation | 14\
positive MTHFR A1298C mutation | 14\
positive factor V Leiden mutation | 14\
complete recanalization of the thrombosed sinuses | 14\
no new thrombi | 14\
complete remission | 28