47 years old | 0
male | 0
admitted to the hospital | 0
decreased mentality | 0
diabetes mellitus | -672
diagnosed with diabetes mellitus | -672
blood pressure 60/30 mm Hg | 0
body temperature 38.5 | 0
white blood cell 13.150×10^9/L | 0
neutrophils 90.7% | 0
lymphocytes 8.5% | 0
hemoglobin 14.3 g/dL | 0
platelet count 507×10^9/L | 0
glucose levels 443 mg/dL | 0
blood urea nitrogen 52.5 mg/dL | 0
serum creatinine concentrations 1.9 mg/dL | 0
aspartate aminotransferase 69 IU/L | 0
alanine transaminase 38 IU/L | 0
sodium 125.7 mmol/L | 0
potassium 5.4 mmol/L | 0
C-reactive protein 19.42 mg/dL | 0
ketone bodies in the blood 3 positive | 0
HbA1c 18.20% | 0
arterial blood gas analysis | 0
pH 7.032 | 0
pCO2 21.8 mm Hg | 0
pO2 83.3 mm Hg | 0
HCO3 5.8 mmol/L | 0
chest X-ray | 0
computed tomography scans | 0
multiple consolidation | 0
ground glass opacities | 0
diabetic ketoacidosis | 0
severe pneumonia | 0
hydration | 0
insulin therapy | 0
piperacillin and tazobactam sodium | 0
mechanical ventilator therapy | 0
admitted to the intensive care unit | 0
ketoacidosis improved | 24
diuretic-resistant pulmonary edema | 48
continuous renal replacement therapy | 48
Klebsiella pneumonia | 48
sputum cultures | 48
lung lesions regressed | 192
moved to the general ward | 192
vague abdominal pain | 240
abdominal pain aggravated | 240
severe tenderness | 240
erect abdominal X-ray | 240
gaseous distention of small bowel loops | 240
stepladder sign | 240
mechanical obstruction | 240
abdominal CT | 240
multiple perforation of the transverse colon | 240
panperitonitis | 240
emergency laparotomy | 240
necrotic intestines | 240
resected specimen | 240
Periodic Acid Schiff | 240
Grocott's methenamine silver staining | 240
septated fungal hyphae | 240
acute angle branching | 240
aspergillus species | 240
colonic IA | 240
intravenous liposomal amphotericin-B | 240
discharged | 576
oral voriconazole | 576
abdominal discomfort | 576
mildly elevated CRP levels | 576
voriconazole discontinued | 624
abdominal discomfort relieved | 624
CRP levels normalized | 624