38 years old | 0
female | 0
gravida 2 | 0
para 1 | 0
admitted to the hospital | 0
heavy vaginal bleeding | 0
hypovolaemic shock | 0
caesarean section | -1092
viable intrauterine pregnancy | -672
cystic structure in the lower uterine cavity | -672
heterotopic pregnancy | -672
ultrasound | -672
vaginal bleeding | 0
unstable | 0
resuscitation | 0
emergency examination under anaesthesia | 0
dilation and curettage | 0
laparotomy | 0
hysterectomy | 0
viable fundal intrauterine pregnancy | 0
lower uterine segment distension | 0
large blood clot | 0
ongoing bleeding | 0
ultrasound-guided suction curettage | 0
thrombus removal | 0
products of conception removal | 0
Foley catheter insertion | 0
bilateral uterine artery ligation | 0
massive transfusion | 0
packed red blood cells | 0
fresh frozen plasma | 0
haemoglobin 96 g/L | 0
intensive care unit | 0
Foley catheter removal | 72
ultrasound at 9+4 weeks of gestation | 96
blood clot in the lower segment of the uterus | 96
single live fetus | 96
heterogenous area in the lower segment of the uterus | 96
antenatal care | 168
shortened cervix | 504
vaginal progesterone | 504
cervical shortening | 504
preterm rupture of membranes | 504
emergency lower-segment caesarean section | 504
antenatal steroids | 504
magnesium sulphate | 504
liveborn male infant | 504
neonatal intensive care unit | 504
neonate death | 528
extreme prematurity | 528
respiratory distress syndrome | 528
bilateral grade three intraventricular haemorrhages | 528
placenta percreta | 8760
elective laparotomy | 8760
classical caesarean section | 8760
total abdominal hysterectomy | 8760
intra-operative haemorrhage | 8760
neonate in good condition | 8760
intensive care unit | 8760
mother and baby discharged | 8784