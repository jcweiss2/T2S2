26 years old | 0
female | 0
vaginal deliveries | -672
complete prenatal care | -672
three doses of tetanus, diphtheria, and pertussis (DTaP) | -672
one dose of tetanus and diphtheria (Tdap) vaccine | -672
last dose of Tdap | -56
postpartum hemorrhage | 48
hypotension | 48
tachycardia | 48
altered sensorium | 48
flaccid uterus | 48
pelvic ultrasound | 48
retention of placental tissue | 48
uterine curettage | 48
discharged | 96
headache | 320
nausea | 320
general malaise | 320
fever | 320
scant lochia | 320
absence of vaginal bleeding | 320
hematocrit 24 % | 320
hemoglobin 7.3 g/dL | 320
white blood cells 14,000 m/mm3 | 320
creatinine 104 μmol/L | 320
urinalysis | 320
positive urine culture for E. coli | 320
hospitalized | 320
treatment with ceftriaxone | 320
treatment with iron saccharate | 320
treatment with hydration | 320
altered mental status | 344
no response to external stimuli | 344
Glasgow Coma Scale score of seven | 344
nuchal stiffness | 344
limb stiffness | 344
intubation | 344
transferred to a more equipped hospital | 344
laboratory exam | 344
non-contrast cerebral computed tomography | 344
lumbar puncture | 344
blood cultures | 344
admitted to the intensive care unit (ICU) | 344
empiric treatment for meningitis | 344
ceftriaxone | 344
vancomycin | 344
acyclovir | 344
severe trismus | 368
increased respiratory rate | 368
spasms of the upper and lower extremities and trunk | 368
passive motion of the limbs caused diffuse spasms | 368
clinical diagnosis of severe tetanus | 368
vaginal cultures | 368
treatment with penicillin G | 368
treatment with anti-tetanus immunoglobulin | 368
extubated | 432
clinical improvement | 432
discharged | 648
gait disorder | 648
mild long-term memory impairment | 648