46 years old | 0
female | 0
admitted to the Emergency Department | 0
headache | 0
vomiting | 0
neurological deterioration | 0
hyposthenia of the left hemysome | 0
cerebral CT scan showed intraparenchymal hemorrhage | 0
MRI of the brain showed rupture of internal carotid artery aneurysm | 0
emergency evacuation of the hematoma | 0
clipping of the aneurysm | 0
transferred to the ICU | 0
developed fever up to 38.5°C | 144
treated with intravenous gentamicin | 144
Escherichia coli urinary tract infection | 144
fever up to 39°C reappeared | 264
neutropenic leukocytosis | 264
thrombocytopenia | 264
procalcitonin value 1.15 ng/mL | 264
blood cultures grew R. mannitolilytica | 264
blood cultures grew R. pickettii | 264
susceptible to ciprofloxacin | 264
susceptible to trimethoprim-sulfamethoxazole | 264
fever persisted despite ciprofloxacin | 264
additional blood cultures positive for Candida parapsilosis | 456
additional blood cultures positive for R. pickettii | 456
additional blood cultures positive for R. mannitolilytica | 456
cultures of central venous catheter negative | 456
cultures of respiratory secretions negative | 456
cultures of urine negative | 456
cultures of rectal swab negative | 456
transthoracic echocardiogram negative for vegetations | 456
funduscopic examinations negative | 456
MRI showed thrombosis of internal carotid artery | 456
anticoagulant therapy with enoxaparin | 456
clearance of candidemia | 456
trimethoprim-sulfamethoxazole added | 600
blood cultures still positive for Ralstonia | 600
antibiotic treatment discontinued | 960
Ralstonia bacteraemia relapsed | 1008
treated with trimethoprim-sulfamethoxazole | 1008
treated with ciprofloxacin | 1008
cranioplasty surgery | 1248
developed fever | 1920
R. pickettii grown from blood cultures | 1920
ciprofloxacin administered | 1920
clinical improvement | 1920
transferred to rehabilitation centre | 1920
eight-week therapy course | 1920
no further relapse | 1920
breast implants | 0
thyroidectomy | 0
