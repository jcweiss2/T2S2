40 years old | 0
    woman | 0
    vomiting | -24
    diarrhea | -24
    loss of consciousness | -24
    common cold treatment | -24
    garenoxacin | -24
    hypothyroidism | -24
    febrile | 0
    shock | 0
    dopamine | 0
    noradrenaline | 0
    antibiotics | 0
    referral to Critical Care Center | 24
    body temperature 38.6°C | 0
    blood pressure 62/46 mmHg | 0
    heart rate 100–110 beats/min | 0
    respiratory rate 20 breaths/min | 0
    oxygen saturation 100% | 0
    Glasgow Coma Scale 15/15 | 0
    unremarkable physical examination | 0
    elevated white blood cell count | 0
    elevated C-reactive protein | 0
    elevated procalcitonin levels | 0
    sepsis-induced disseminated intravascular coagulation | 0
    elevated creatinine kinase | 0
    elevated creatinine kinase MB | 0
    elevated troponin T | 0
    sequential organ failure assessment score 8 | 0
    unremarkable chest radiography | 0
    unremarkable computed tomography | 0
    negative rapid antigen kit test for group A streptococcus | 0
    septic shock with unknown focus | 0
    meropenem | 0
    vancomycin | 0
    clindamycin | 0
    continuous renal replacement therapy | 0
    intravenous immunoglobulin | 0
    arginine vasopressin | 0
    hydrocortisone | 0
    dobutamine | 0
    pulse-induced contour cardiac output monitoring | 0
    intubation | 0
    mechanical ventilation | 0
    circulatory status not improved | 5
    MAP 40 mmHg | 5
    pulse contour cardiac index 1.34 L/min/m2 | 5
    administration of 2.3 L fluids | 5
    catecholamines | 5
    widespread ST elevation | 5
    ST depression | 5
    reduced LVEF 20% | 5
    diffuse hypokinesia | 5
    cardiogenic shock | 5
    coronary angiography no stenosis | 6
    Swan-Ganz catheter low cardiac output | 6
    IABP introduction | 6
    assist ratio 1:1 | 6
    stable circulatory status | 6
    HR 101 beats/min | 6
    MAP 84 mmHg | 6
    improved left ventricle motion | 6
    LVEF 40% | 6
    CRRT initiation | 9
    renal dysfunction | 9
    oliguria | 9
    reduced noradrenaline | 25
    reduced dobutamine | 25
    discontinuation of dobutamine | 36
    IABP assist ratio 1:2 | 40
    IABP discontinuation | 72
    vasoactive agents discontinuation | 72
    no IABP-related complications | 72
    fever resolved | 144
    CRRT discontinued | 168
    mechanical ventilation terminated | 264
    LVEF 54% | 168
    improvement in wall motion | 168
    inflammatory markers improved | 168
    inflammatory markers normal | 336
    discontinued antibiotics | 336
    returned to previous hospital | 528
    highly elevated anti-streptolysin O | 408
    anti-streptokinase detected | 408
    normal thyroid function | 1368
    <|eot_id|>
    