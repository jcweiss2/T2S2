33 years old | 0
male | 0
admitted to the hospital | 0
fever | -2160
diarrhea | -2160
anemia | -2160
liver dysfunction | -2160
elevated ferritin | -2160
unexplained anemia | -2160
splenomegaly | -2160
denies previous blood transfusion | 0
married | 0
2 children | 0
no family history of familial disease except for thalassemia in a sister | 0
provided written informed consent | 0
fever (>40°C) | -2160
received medical attention at the First Affiliated Hospital of Sun Yat-sen University | -2160
blood chemistry panel | -2160
hemoglobin (88 g/l) | -2160
ferritin (1,068.47 mg/l) | -2160
total bilirubin (392.4 mmol/l) | -2160
conjugated bilirubin (335.7 mmol/l) | -2160
γ-glutamyl transpeptidase (γ-GT; 150 U/l) | -2160
fibrinogen (1.53 g/l) | -2160
mechanical ventilation | -2153
respiratory failure | -2153
antibiotic treatment for suspected pneumonia and cholecystitis | -2153
diarrhea with watery stool | -2143
treatment with itraconazole and norvancomycin | -2143
colonoscopy | -2137
inflammatory colitis | -2137
immunohistochemical analysis of colon biopsy specimen identified CMV | -2137
treatment with ganciclovir | -2137
abdominal pain and bloating dissipated | -2127
body temperature returned to normal | -2127
diarrhea did not improve | -2127
immunohistochemical examination of the peripheral blood | -2121
no CMV | -2121
bone marrow aspiration | -2121
no hemophagocytosis | -2121
blood chemistry | -2121
improvement in total bilirubin (86.7 mmol/l) | -2121
conjugated bilirubin (43.9 mmol/l) | -2121
γ-GT (71 U/l) | -2121
fibrinogen (1.24 g/l) | -2121
requested discharge from the hospital | -2111
presented to us at the First Affiliated Hospital of Guangzhou University of Chinese Medicine | 0
body temperature was 41.0°C | 0
jaundice of the skin and sclera | 0
lower abdomen was distended | 0
no tenderness or rebound tenderness | 0
hepatomegaly and splenomegaly | 0
bedside chest X-ray | 0
no abnormality | 0
nutritional support | 0
blood chemistry analysis | 0
anemia (hemoglobin, 36 g/l) | 0
hyperbilirubinemia (total bilirubin, 234.9 mmol/l; conjugated bilirubin, 147.5 mmol/l) | 0
fever persisted (40°C) | 0
transferred to the intensive care unit | 240
CMV-immunoglobulin M testing | 240
negative result | 240
T lymphocyte count | 240
cluster of differentiation (CD)3+ (79.2.2%) | 240
CD4+ (38.2%) | 240
CD8+ (35.3%) | 240
T helper/suppressor cell ratio (1.08) | 240
hemoglobin was 39 g/l | 240
red blood cell count was 1.61×10^12/l | 240
leukocyte count was 2.67×10^9/l | 240
platelet count was 57×10^9/l | 240
ferritin was substantially elevated (7,931.21 mg/l) | 240
blood chemistry analysis | 240
total bilirubin value of 299.5 mmol/l | 240
conjugated bilirubin value of 215.7 mmol/l | 240
urinalysis | 240
occult blood (++) | 240
urinary bilirubin (++) | 240
10 erythrocytes/HPF | 240
abdominal computed tomography (CT) scan | 240
splenomegaly | 240
multiple gall bladder stones | 240
inflammatory changes in the gall bladder | 240
Wright-Giemsa staining | 240
bone marrow smears | 240
active hemophagocytosis | 240
phagocytosis of nucleated red blood cells and platelets | 240
whole-body positron emission tomography/CT scan | 240
no tumor mass | 240
peripheral blood and bone marrow aspiration sample specimens | 240
culture agar | 240
L. pseudomesenteroides | 240
identified using a VITEK 2 GP Test kit | 240
results from a stool culture for Clostridium difficile (C. difficile) was negative | 240
blood and bone marrow aspirate culture | 240
results came back positive on day 14 after admission for L. pseudomesenteroides | 336
drug sensitivity test | 336
vancomycin-resistant | 336
clindamycin-sensitive | 336
clindamycin (150 mg, taken orally every 12 h for 1 week) | 336
4 units of red blood cell suspension | 336
350 ml frozen plasma | 336
partial parenteral nutrition | 336
fever subsided rapidly (37.0°C) after 1 day of clindamycin therapy | 360
patient became afebrile after 7 days of clindamycin therapy | 504
repeat blood culture 10 days later identified L. pseudomesenteroides | 696
blood chemistry 5 days later | 696
improvement in hemoglobin (77 g/l) | 696
red blood cell count (3.05×10^12/l) | 696
platelet count (139×10^9/l) | 696
total (71.5 mmol/l) and conjugated bilirubin (45.2 mmol/l) | 696
body temperature returned to normal (36.5°C) | 696
volume of stool was reduced to 350 ml/day | 696
repeat blood culture 2 weeks later was negative for L. pseudomesenteroides | 1008
requested discharge due to financial concern | 1008
telephone follow-up 2 weeks later | 1128
continued treatment at Pengpai Memorial Hospital (Shanwei, China) | 1128
blood culture for L. pseudomesenteroides was negative | 1128
visited our hospital 8 months later | 4032
complete blood count test | 4032
continued to be anemic (hemoglobin at 89 g/l) | 4032
no other complaints | 4032