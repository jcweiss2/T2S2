13 years old | 0
female | 0
DiGeorge syndrome | 0
prior neonatal truncus arteriosus repair | 0
severe left pulmonary artery hypoplasia | 0
methicillin-sensitive staphylococcal bacteremia | -72
infective endocarditis | -72
septic pulmonary emboli | -72
bilateral pyelonephritis | -72
septic shock | -72
worsening respiratory failure | -24
pulmonary hemorrhage | -24
venovenous extracorporeal membrane oxygenation (V-V ECMO) | -24
acute hemorrhage | -144
right chest tube | -144
endotracheal tube | -144
computed tomography angiography | -144
patent conduit | -144
right ventricle | -144
pulmonary artery | -144
acute right hemothorax | -144
mycotic aneurysm | -144
medial basal segment | -144
right lower lobe pulmonary artery | -144
extravasation | -144
intercostal artery | -144
general anesthesia | -120
perfusionist team | -120
ECMO circuit | -120
left common femoral vein access | -120
micropuncture set | -120
9-French Flexor sheath | -120
inferior vena cava | -120
7-French APC catheter | -120
main pulmonary artery | -120
digital subtraction arteriography | -120
patent pulmonary artery conduit | -120
19-mm bilobed mycotic aneurysm | -120
guiding sheath | -120
right pulmonary artery | -120
5-French vertebral tip catheter | -120
AngioDynamics | -120
angled tip Glidewire | -120
Terumo | -120
branch vessel | -120
friable mycotic aneurysm | -120
embolization | -120
balloon occlusion technique | -120
ethylene-vinyl alcohol copolymer (EVOH) | -120
Onyx | -120
Scepter C Occlusion Balloon Catheter | -120
Microvention | -120
Synchro 0.014-inch wire | -120
Stryker Neurovascular | -120
Cadence Precision injector syringe | -120
dimethyl sulfoxide | -120
EVOH (Onyx 34) | -120
embolization of mycotic aneurysm | 0
pulmonary arteriography | 0
occlusion of mycotic aneurysm | 0
preserved flow | 0
normal lung parenchyma | 0
right femoral arterial access | 0
thoracic aortogram | 0
extravasation | 0
right intercostal artery | 0
coils | 0
Gelfoam | 0
total procedure time | 0
132 minutes | 0
pediatric intensive care unit | 24
stable condition | 24
hemorrhage | 24
right chest tube | 24
endotracheal tube | 24
resolved | 24
neurologic deterioration | 72
care withdrawn | 72
autopsy declined | 72