9 years old | 0
male | 0
idiopathic bone marrow aplasia | 0
admitted to pediatric ICU | 0
septic shock | 0
respiratory insufficiency | 0
mechanical ventilation | 0
cardiac monitoring | 0
severe neutropenia | 0
fever of unknown origin | 0
broad-spectrum antibiotic therapy | 0
antifungal therapy | 0
no clinical improvement | 0
circular erythematous lesions | -1080
necrotic center under cardiac monitoring electrodes | -1080
extensive necrosis | -1080 + 240
second biopsy | -1080 + 240
septate hyaline hyphae | -1080 + 240
Grocott staining | -1080 + 240
many septate hyphae with branches at acute angles | -1080 + 240
culture of material in Sabouraud dextrose agar plate | -1080 + 240
darker reverse coloration | -1080 + 240
microcultive in lamina technique | -1080 + 240
Aspergillus niger species | -1080 + 240
whole body computed tomography scan | -1080 + 240
no disseminated fungal infection | -1080 + 240
amphotericin B | 0
fluconazole | 0
voriconazole | -1080 + 240
no improvement | -1080 + 240
death | 2160
primary cutaneous aspergillosis | -1080 + 240
inoculation of Aspergillus species | -1080 
non-sterile cardiac monitoring electrodes | -1080 
use of non-sterile devices | -1080 
immunocompromised patient | 0 
infectious disease suspected | -1080 + 240 
biopsy and cultures performed | -1080 + 240 
pathogen identification | -1080 + 240 
sterile disposable devices recommended | -1080 + 240 
preventable risk of PCA | -1080 + 240 
importance of monitoring skin changes | -1080 + 240