79 years old| 0
female | 0
hypertension | 0
type 2 diabetes mellitus | 0
dyslipidemia | 0
hyperuricemia | 0
IgG/λ multiple myeloma | -1464
increased total serum proteins | -1464
increased γ-globulins | -1464
increased IgG heavy chains | -1464
increased free λ light chains | -1464
IgG/λ monoclonal gammopathy | -1464
hypocellular medullary aspirate | -1464
abnormal plasmocytes | -1464
anemia | -1464
lytic bone lesions | -1464
oral melphalan | -1464
prednisolone | -1464
ECOG Performance Status 1 | -1464
admitted to emergency department | 0
fatigue | 0
severe bone pain | 0
diarrhea | 0
hemodynamic instability | 0
oliguria | 0
oxygen requirement | 0
decreased breath sounds | 0
anemia | 0
leukocytosis | 0
neutrophilia | 0
thrombocytopenia | 0
elevated C-reactive protein | 0
elevated creatinine | 0
hypoalbuminemia | 0
type 1 respiratory insufficiency | 0
hyperlactacidemia |
