42 years old | 0
    multiparous | 0
    gestational age of 35 + 2 weeks | 0
    presented to the ER | 0
    altered mentation | 0
    seizures | 0
    high fever of 38.3 °C | 0
    nasopharyngeal COVID-19 PCR test positive | -48
    throat pain | -48
    endotracheal intubation | 0
    emergency call to obstetrics and gynecology department | 0
    mechanical ventilation | 0
    delivered a healthy baby by cesarean section two years ago | -17520
    no specific underlying diseases | 0
    no remarkable events during prenatal examinations | 0
    no history of drug abuse | 0
    no history of smoking | 0
    no history of drinking | 0
    no family history of genetic diseases | 0
    no family history of autoimmune diseases | 0
    no family history of thyroid diseases | 0
    generalized tonic-clonic seizure | 0
    drooling | 0
    continuous upper eyeball deviation | 0
    pupillary reflex prompt | 0
    pupillary reflex symmetric | 0
    pupillary reflex consensual | 0
    blood pressure of 121/71 mmHg | 0
    heart rate of 115 beats per minute | 0
    increased C-reactive protein | 0
    increased erythrocyte sedimentation rate |9| 0
    increased D-dimer | 0
    no proteinuria | 0
    normal urine protein-to-creatinine ratio | 0
    normal liver function test | 0
    normal serum electrolytes | 0
    normal blood glucose | 0
    normal blood urea nitrogen | 0
    normal creatinine | 0
    suppressed TSH | 0
    elevated free T4 | 0
    elevated total T3 | 0
    Burch-Wartofsky Point Scale score 65 | 0
    no acute intracranial hemorrhage | 0
    no focal parenchymal lesions | 0
    no visible causes of seizure | 0
    no focal neurological signs | 0
    no significant uterine contractions | 0
    fetal growth appropriate for gestational age | 0
    fetal heartbeat normal | 0
    fetal movements normal | 0
    initial diagnosis of eclampsia | 0
    maternal blood pressure normal | 0
    no fetal growth restriction | 0
    no thrombocytopenia | 0
    no kidney failure | 0
    no hepatic dysfunction | 0
    diagnosis of atypical eclampsia | 0
    final diagnosis of status epilepticus | 0
    final diagnosis of thyroid storm | 0
    final diagnosis of preexisting Graves’ disease | 0
    SARS-CoV-2 trigger for thyroid storm | 0
    treatment with labetalol | 0
    treatment with magnesium sulfate | 0
    treatment with midazolam | 0
    seizures persisted | 0
    consciousness not restored | 0
    cesarean section performed | 24
    newborn infant weight 2680 g | 24
    Apgar scores 8 at 1 min | 24
    Apgar scores 8 at 5 min | 24
    seizures continued post-cesarean | 24
    low-level sedation maintained | 24
    seizures decreased | 24
    consciousness restored | 24
    newborn's COVID-19 PCR test negative | 24
    newborn's thyroid function tests normal | 24
    no specific MRI findings | 24
    no specific electroencephalogram findings | 24
    TSH suppressed | 0
    free T4 elevated | 0
    total T3 elevated | 0
    TSH receptor antibody elevated | 0
    diffusely enlarged thyroid gland | 0
    round-shaped lobes | 0
    diffusely heterogeneous echotexture | 0
    coarse echotexture | 0
    isthmus nodule suspected malignant | 0
    fine-needle aspiration performed | 0
    cytology result papillary carcinoma | 0
    thyroidectomy scheduled | 0
    methimazole prescribed | 0
    methylprednisolone prescribed | 0
    propranolol prescribed | 0
    discharged ten days after cesarean | 240
    thyroid function tests near normal after one month | 720
    <|eot_id|>
    