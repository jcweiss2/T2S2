58 years old | 0
    male | 0
    admitted to the hospital | 0
    fecal occult blood | 0
    endoscopic mucosal resection (EMR) | -72
    electrocoagulation electro resection | -72
    cold resection | -72
    broad-based polyps | -72
    pedicled polyps | -72
    cecum polyps | -72
    ascending colon polyps | -72
    transverse colon polyps | -72
    descending colon polyps | -72
    sigmoid colon polyps | -72
    shock | -72
    dyspnea | -72
    sweating | -72
    blood pressure decreased | -72
    oxygen saturation decreased | -72
    heart rate increased | -72
    stable vital signs | 0
    normal coagulation function | 0
    colonoscopy | 96
    ulcerative foci | 96
    EMR of polyps | 96
    titanium clips placement | 96
    blood pressure decreased | 144
    heart rate increased | 144
    oxygen saturation dropped | 144
    mental irritability | 144
    gastrectomy | -8760
    gastric ulcers | -8760
    surgical treatment for oral cancer | -96
    fecal occult tests positive | -96
    painless colonoscopy | -96
    colon polyps | -96
    no adverse events | -96
    no family genetic history | 0
    blood gas analysis | -72
    pH 7.33 | -72
    partial pressure of carbon dioxide 37 mmHg | -72
    partial pressure of oxygen 211 mmHg | -72
    lactate levels 4.8 mmol/L | -72
    bicarbonate radical concentration 19.5 mmol/L | -72
    base excess -5.8 mmol/L | -72
    potassium ion concentration 2.9 mmol/L | -72
    PaO2/FiO2 221 mmHg | -72
    white blood cell count 3.29 × 10^9/L | -72
    neutrophil percentage 87.8% | -72
    platelet count 142 × 10^12/L | -72
    procalcitonin 1.66 ng/mL | -72
    interleukin-6 > 5000 pg/mL | -72
    prothrombin time 36.2 s | -72
    international normalized ratio 3.6 | -72
    prothrombin activity 21% | -72
    activated partial thromboplastin time 69.1 s | -72
    fibrinogen concentration < 0.6 g/L | -72
    fibrin degradation product > 360 μg/mL | -72
    D-dimer > 40 μg/mL | -72
    antithrombin III 69% | -72
    blood culture negative | -72
    blood gas analysis | 144
    pH 7.23 | 144
    partial pressure of carbon dioxide 33 mmHg | 144
    partial pressure of oxygen 149 mmHg | 144
    lactate level 7.1 mmol/L | 144
    bicarbonate radical concentration 13.8 mmol/L | 144
    base excess -12.7 mmol/L | 144
    potassium ion concentration 6.5 mmol/L | 144
    PaO2/FiO2 186 mmHg | 144
    white blood cell count 12.38 × 10^9/L | 144
    neutrophil percentage 86.4% | 144
    hemoglobin concentration 84 g/L | 144
    platelet count 192 × 10^12/L | 144
    procalcitonin 1.26 ng/mL | 144
    interleukin-6 > 5000 pg/mL | 144
    prothrombin time 36.5 s | 144
    international normalized ratio 3.64 | 144
    prothrombin activity 20% | 144
    activated partial thromboplastin time 62 s | 144
    fibrinogen concentration < 0.6 g/L | 144
    fibrin degradation product > 360 μg/mL | 144
    D-dimer > 40 μg/mL | 144
    antithrombin III 65% | 144
    thromboelastography abnormalities | 144
    white blood cell count 20.46 × 10^9/L | 168
    hemoglobin concentration 62 g/L | 168
    procalcitonin 5.72 ng/mL | 168
    platelet count normal | 168
    coagulation function normal | 168
    abdominal computed tomography | 168
    superior mesenteric artery CT angiography | 168
    no intestinal perforation | 168
    no lumbar lesion | 168
    no vascular damage | 168
    sepsis | 0
    septic shock | 0
    gastrointestinal bleeding | 168
    postpolypectomy syndrome | 0
    Moraxella osloensis infection | 168
    no abdominal pain | 0
    respiratory support | -72
    fluid resuscitation | -72
    oxygen treatment | -72
    transferred to ICU | -72
    regained consciousness | -72
    no abdominal pain | -72
    no abdominal distension | -72
    blood pressure recovery | -72
    heart rate 115 beats/min | -72
    respiratory rate 25 breaths/min | -72
    oxygen saturation 95% | -72
    temperature 38.9 °C | -72
    cefoxitin administration | -72
    plasma transfusion | -72
    fluid resuscitation | -72
    antiallergic therapy | 144
    vasoactive drugs | 144
    dark red bloody stools | 144
    cefoxitin administration | 144
    plasma infusion | 144
    cryoprecipitate infusion | 144
    red blood cells infusion | 144
    vital signs stable | 168
    gastrointestinal bleeding ceased | 168
    discharged | 192