4 years old | 0
female | 0
relapsed refractory pre-B cell ALL | 0
diagnosis of standard risk pre-B ALL | -199*24
blasts coexpressed CD19, CD22, CD58, CD10, CD38 | -199*24
cytogenetics revealed p53 deletion | -199*24
t(1;19) with a complex karyotype | -199*24
no CNS disease | -199*24
treated with National Mexican Protocol | -199*24
no evidence of morphologic or minimal residual disease via flow cytometry at end of induction chemotherapy | -199*24
relapsed 199 days after diagnosis | -199*24
failed reinduction chemotherapy | -199*24
failed two cycles of blinatumomab | -199*24
treated with reinduction therapy per ALL R3 | -199*24
did not achieve remission | -199*24
high burden of extramedullary disease in liver | -199*24
high burden of extramedullary disease in spleen | -199*24
high burden of extramedullary disease in kidneys | -199*24
high burden of extramedullary disease in lymph nodes | -199*24
chloroma to left orbit | -199*24
cranial nerve II palsy | -199*24
renal insufficiency | -199*24
requiring long-term electrolyte replacement | -199*24
poor response to therapy | -199*24
plans made for transfer of care for CAR T-cell therapy | -199*24
received bridging oral chemotherapy with 6-mercaptopurine | -199*24
received bridging oral chemotherapy with methotrexate | -199*24
treated for Staphylococcal epidermidis central catheter infection | -2*168
treated for septic shock with 10-day course of vancomycin | -2*168
received lymphoid depleting chemotherapy with fludarabine | -2*168
received lymphoid depleting chemotherapy with cyclophosphamide | -2*168
presented to emergency department on day 2 of lymphoid depleting therapy | -2*168
fever | -2*168
nausea | -2*168
headache | -2*168
fatigue | -2*168
initial resuscitation | -2*168
work-up | -2*168
initiation of broad-spectrum antibiotics | -2*168
admitted to hematology/oncology team | -2*168
transferred to PICU due to progressive septic shock with hypotension | 36
afebrile | 36
blood pressure 69/31 | 36
heart rate 165 beats per minute | 36
respiratory rate 56 breaths per minute | 36
oxygen saturation 100% on room air | 36
poor perfusion | 36
capillary refill time of 5 seconds | 36
pulses 3+ in bilateral radial arteries | 36
no murmur | 36
no gallop | 36
hypotension despite aggressive fluid resuscitation | 36
high doses of inotropes | 36
broad-spectrum antibiotics | 36
intubation for persistent shock | 36
contacted oncology team to discuss expected prognosis | 36
initiated on VA ECMO | 48
decannulated | 6*24
extubated | 10*24
blood culture positive for Escherichia coli | 36
suspected multidrug resistant | 36
mechanical ventilation | 36
initial echocardiogram revealed severe global hypokinesis of left ventricle | 36
ejection fraction 31% | 36
on vasoactive support including epinephrine | 36
on vasoactive support including norepinephrine | 36
on vasoactive support including vasopressin | 36
maximal Vasoactive-Inotropic Score of 98 | 36
ongoing shock state | 36
acute kidney injury | 36
severe oliguria | 36
total body fluid overload 18% | 36
lack of response to escalation of vasoactive support | 36
stress dose steroids | 36
bicarbonate infusion | 36
continuous renal replacement therapy initiated | 36
progression to multiple organ dysfunction | 36+8
ongoing shock (peak lactate 24 mmol/L) | 36+8
myocardial ischemia (troponin 2.03 nanogram/mL) | 36+8
renal dysfunction (three-fold rise in baseline serum creatinine 0.2–0.6) | 36+8
coagulopathy (prothrombin time 28.6 s, partial thromboplastin time 111.2 s, international normalized ratio 2.50) | 36+8
hepatobiliary dysfunction (aspartate aminotransferase 224 unit/L, total bilirubin 4.3 mg/dL, direct bilirubin 3.7 mg/dL) | 36+8
continued conversations between pediatric intensivist and oncologist | 36+8
ECMO candidacy and prognosis discussed | 36+8
family consented for venoarterial ECMO | 36+8
cannulated for venoarterial ECMO | 36+8
indwelling central catheter removed | 36+8
anticoagulation managed with systemic heparin | 36+8
CRRT via Prismaflex | 36+8
therapeutic plasma exchange (1.5× volume day 1 followed by 1× volume for 5 days) | 36+8
broad-spectrum antimicrobial therapy (meropenem, ceftazidime/avibactam, gentamicin, micafungin) | 36+8
weaned off vasoactive and inotropic support | 48
initiated on milrinone | 48
maintained good antegrade flow across aortic valve | 48
bacteremia cleared | 48
cardiac dysfunction improved | 48
repeat echo demonstrated low normal biventricular systolic function | 48+120
ejection fraction 51% during ECMO clamp trial | 48+120
CAR T-cell infusion (tisagenlecleucel) | 17*24
transferred to hematology/oncology service | 17*24
developed cytokine release syndrome | 17*24
requiring tocilizumab | 17*24
brief PICU readmission | 17*24
identified in remission 1 month later | 10*24
discharged | 10*24
diagnosis of standard risk pre-B ALL | -4776
blasts coexpressed CD19, CD22, CD58, CD10, CD38 | -4776
cytogenetics revealed p53 deletion | -4776
t(1;19) with a complex karyotype | -4776
no CNS disease | -4776
treated with National Mexican Protocol | -4776
no evidence of morphologic or minimal residual disease via flow cytometry at end of induction chemotherapy | -4776
relapsed 199 days after diagnosis | -4776
failed reinduction chemotherapy | -4776
failed two cycles of blinatumomab | -4776
treated with reinduction therapy per ALL R3 | -4776
did not achieve remission | -4776
high burden of extramedullary disease in liver | -4776
high burden of extramedullary disease in spleen | -4776
high burden of extramedullary disease in kidneys | -4776
high burden of extramedullary disease in lymph nodes | -4776
chloroma to left orbit | -4776
cranial nerve II palsy | -4776
renal insufficiency | -4776
requiring long-term electrolyte replacement | -4776
poor response to therapy | -4776
plans made for transfer of care for CAR T-cell therapy | -4776
received bridging oral chemotherapy with 6-mercaptopurine | -4776
received bridging oral chemotherapy with methotrexate | -4776
treated for Staphylococcal epidermidis central catheter infection | -336
treated for septic shock with 10-day course of vancomycin | -336
received lymphoid depleting chemotherapy with fludarabine | -336
received lymphoid depleting chemotherapy with cyclophosphamide | -336
presented to emergency department on day 2 of lymphoid depleting therapy | -336
fever | -336
nausea | -336
headache | -336
fatigue | -336
initial resuscitation | -336
work-up | -336
initiation of broad-spectrum antibiotics | -336
admitted to hematology/oncology team | -336
decannulated | 144
extubated | 240
progression to multiple organ dysfunction | 44
ongoing shock (peak lactate 24 mmol/L) | 44
myocardial ischemia (troponin 2.03 nanogram/mL) | 44
renal dysfunction (three-fold rise in baseline serum creatinine 0.2–0.6) | 44
coagulopathy (prothrombin time 28.6 s, partial thromboplastin time 111.2 s, international normalized ratio 2.50) | 44
hepatobiliary dysfunction (aspartate aminotransferase 224 unit/L, total bilirubin 4.3 mg/dL, direct bilirubin 3.7 mg/dL) | 44
continued conversations between pediatric intensivist and oncologist | 44
ECMO candidacy and prognosis discussed | 44
family consented for venoarterial ECMO | 44
cannulated for venoarterial ECMO | 44
indwelling central catheter removed | 44
anticoagulation managed with systemic heparin | 44
CRRT via Prismaflex | 44
therapeutic plasma exchange (1.5× volume day 1 followed by 1× volume for 5 days) | 44
broad-spectrum antimicrobial therapy (meropenem, ceftazidime/avibactam, gentamicin, micafungin) | 44
repeat echo demonstrated low normal biventricular systolic function | 168
ejection fraction 51% during ECMO clamp trial | 168
CAR T-cell infusion (tisagenlecleucel) | 408
transferred to hematology/oncology service | 408
developed cytokine release syndrome | 408
requiring tocilizumab | 408
brief PICU readmission | 408
identified in remission 1 month later | 240
discharged | 240
