54 years old | 0
male | 0
uncontrolled diabetes mellitus | 0
HbA1c of 13% | 0
admitted to the hospital | 0
right frontal headache | -120
vomiting | -120
normal complete blood count | 0
normal renal profile | 0
normal hepatic profile | 0
elevated glucose level | 0
negative blood culture | 0
negative HIV serology | 0
normal CD4 count | 0
brain CT scan | 0
circumferential mucosal thickening in the sphenoid sinuses | 0
right side | 0
mild scattered mucosal thickening in the other paranasal sinuses | 0
fluid opacification of the mastoid air cells | 0
fluid opacification of the middle ear cavities | 0
insulin | 0
Augmentin | 0
complained of sudden loss of vision in the right eye | 120
complained of jaw pain | 120
brain CT scan repeated | 120
progression of the inflammatory changes in the paranasal sinuses | 120
no acute brain insult | 120
suspected giant cell arteritis | 120
pulse intravenous methylprednisolone 1 gm daily | 120
temporal artery biopsy performed | 168
normal temporal artery biopsy | 168
corticosteroids discontinued | 168
symptoms worsened | 168
third CT scan brain | 168
progression of the sinusitis to the retropharyngeal abscess | 168
sinonasal biopsy obtained | 168
histopathological examination | 168
positive GMS stain for fungus | 168
mucormycosis | 168
treated with amphotericin B | 168
developed sepsis | 240
broad-spectrum antibiotics | 240
vancomycin | 240
meropenem | 240
chest CT scan | 240
abdominal CT scan | 240
mild bilateral pleural effusions | 240
mucosal edema involving the ascending colon | 240
no obstruction | 240
no significant lymphadenopathy | 240
developed melena | 336
developed streaks of blood | 336
hemoglobin drop from 83 to 75 g/L | 336
upper GI endoscopy | 336
sigmoidoscopy | 336
severe erythematous gastritis | 336
huge gastric ulcer | 336
necrotic-looking tissues | 336
non-bleeding visible vessel | 336
clipped | 336
multiple biopsies obtained | 336
pale mucosa | 336
ischemic changes 18–25 cm from the anal verge | 336
biopsies obtained | 336
severe acute chronic inflammation | 336
fibrinous exudate | 336
extensive ulceration | 336
fibrin microthrombi | 336
numerous fungal microorganisms | 336
single and clustered small (2–10 μm) narrow-based budding yeasts | 336
cryptococcus species | 336
refractory septic shock | 336
multiorgan failure | 336
passed away | 336