63 years old | 0
male | 0
admitted to the hospital | 0
right sided hemiparesis | -0.3
altered mental status | -0.3
confused | -0.3
aphasic | -0.3
right upper and lower extremity hemiparesis | -0.3
NIH stroke scale was 18 | 0
stroke alert | 0
non-contrast CT scan of the brain | 0
chronic opacification of left mastoid air cells | 0
fluid in mastoid air spaces bilaterally | 0
CT angiography of the head and neck | 0
tissue plasminogen activator (tPA) not given | 0
worsening encephalopathy | 2
intubated for airway protection | 2
fever 103 degrees Fahrenheit | 2
heart rate increased to 120 beats per minute | 2
newly dilated, non-reactive right pupil | 2
central nervous system infection | 2
uncal herniation | 2
stat repeat NCCT scan of the brain | 2
rapidly developing white matter edema | 2
lumbar puncture (LP) attempted | 2
empiric intravenous vancomycin, ceftriaxone, ampicillin and acyclovir administered | 2
white blood cell count of at 15,200/ μL | 2
lactic acid measurement of 3.2 mmol/L | 2
severe sepsis | 2
critical care medicine consulted | 2
admitted to the intensive care unit | 2
cerebrospinal fluid analysis | 4
gram-positive cocci in chains | 4
Streptococcus pneumoniae | 4
acute on chronic mastoiditis | 4
surgical intervention | 4
left sided myringotomy with tympanostomy tube placement | 8
cranial nerve palsy resolved | 8
ceftriaxone administered | 8
intravenous dexamethasone given | 8
follow up NCCT scan of the brain | 12
improvement of the previously identified extensive white matter edema | 12
weaned off of sedation | 96
neurologically stable for extubation | 96
encephalopathy resolved | 96
right sided motor weakness completely resolved | 96
transferred to the general medical floor | 96
diabetes mellitus 2 | -8760
bilateral mastoidectomies | -8760
progressive left ear pain | -72
discharged | 168