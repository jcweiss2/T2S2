3 years old | 0
    female | 0
    complex congenital heart disease | 0
    previous cardiac surgeries | 0
    admitted to the pediatric intensive care unit | 0
    shock | 0
    cardiopulmonary arrest | 0
    resuscitation | 0
    thrombosis in right ventricle-to-pulmonary artery conduit | 0
    severe hypoxic+ischemic encephalopathy | 0
    acute kidney injury | 0
    neurological rehabilitation | 0
    transition to home ventilation | 0
    dystonia | 0
    heart failure | 0
    endocarditis | 0
    pulmonary embolism | 0
    stem cell therapy investigated | 0
    metformin initiated | -408
    metformin dose increased | -144
    wide complex bradycardia | 0
    blood pressure 90/40 mmHg | 0
    respiratory rate 26 breaths per minute | 0
    temperature 37.2 °C | 0
    oxygen saturation 87% | 0
    prolonged capillary refill time | 0
    lethargic | 0
    severe lactic acidosis | 0
    hyperkalemia | 0
    hyperglycemia | 0
    hypotension | 0
    propranolol discontinued | 0
    dopamine infusion | 0
    norepinephrine infusion | 0
    higher ventilator support | 0
    clinical status improved | 3
    support therapies weaned | 3
    recurrence of serum lactate rise | 12
    recurrence of hyperkalemia | 12
    metformin discontinued | 12
    creatinine levels doubled | -120
    AKI resolved | 0
    metformin levels not collected | 0
    sepsis ruled out | 0
    rhabdomyolysis ruled out | 0
    blood cultures sterile | 0
    recovered rapidly | 12
    normal creatinine kinase levels | 0
    no new anti-infective agents | 0
    
</|end_header_id|>

3 years old | 0
female | 0
complex congenital heart disease | 0
previous cardiac surgeries | 0
admitted to the pediatric intensive care unit | 0
shock | 0
cardiopulmonary arrest | 0
resuscitation |?| 0
thrombosis in right ventricle-to-pulmonary artery conduit | 0
severe hypoxic-ischemic encephalopathy | 0
acute kidney injury | 0
neurological rehabilitation | 0
transition to home ventilation | 0
dystonia | 0
heart failure | 0
endocarditis | 0
pulmonary embolism | 0
stem cell therapy investigated | 0
metformin initiated | -408
metformin dose increased | -144
wide complex bradycardia | 0
blood pressure 90/40 mmHg | 0
respiratory rate 26 breaths per minute | 0
temperature 37.2 °C | 0
oxygen saturation 87% | 0
prolonged capillary refill time | 0
lethargic | 0
severe lactic acidosis | 0
hyperkalemia | 0
hyperglycemia | 0
hypotension | 0
propranolol discontinued | 0
dopamine infusion | 0
norepinephrine infusion | 0
higher ventilator support | 0
clinical status improved | 3
support therapies weaned | 3
recurrence of serum lactate rise | 12
recurrence of hyperkalemia | 12
metformin discontinued | 12
creatinine levels doubled | -120
AKI resolved | 0
metformin levels not collected | 0
sepsis ruled out | 0
rhabdomyolysis ruled out | 0
blood cultures sterile | 0
recovered rapidly | 12
normal creatinine kinase levels | 0
no new anti-infective agents | 0