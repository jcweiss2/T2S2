48 years old | 0
male | 0
admitted to the Emergency Department | 0
coronary artery disease | -672
chronic kidney disease | -672
chest pain | 0
shortness of breath | 0
stabilized in the ED | 0
transferred to the intermediate general ward | 0
drug optimization | 0
hemodialysis | 0
coronary angiography | 0
3-vessel CAD | 0
61% ejection fraction | 0
overweight | 0
history of CKD | 0
history of hemodialysis | 0
history of stroke | 0
history of angina | 0
history of diabetes | 0
history of dyslipidemia | 0
history of smoking | 0
scheduled for urgent CABG surgery | 0
preoperative screening | 0
no rapid testing | 0
anemia | 0
leukocytosis | 0
increased cardiac enzymes | 0
decreased pCO2 | 0
increased pO2 | 0
decreased HCO3 | 0
thorax X-ray showed cardiomegaly | 0
CABG surgery | 192
transferred to the Intensive Care Unit | 192
extubated | 212
transferred to the intermediate ward | 216
transferred to the ward | 240
complained of increased difficulty in breathing | 336
decreased saturation | 336
low PO2 | 336
fever | 336
transferred to the isolation ICU room | 336
reintubated | 336
tested for COVID-19 | 336
RT-PCR test | 336
positive for COVID-19 | 336
neutrophil-to-lymphocyte ratio | 360
consolidation of both lungs | 360
pneumonia | 360
hemodynamically unstable | 432
sepsis | 432
deterioration of urea and creatinine levels | 432
considered for continuous renal replacement therapy | 432
respiratory failure | 456
died | 528
respiratory distress | 528
COVID-19 infection | 528