60 years old | 0
female | 0
hepatitis C-related cirrhosis | -672
recurrent hepatic encephalopathies | -672
chronic portal vein thrombosis | -672
liver transplantation | 0
construction of an end-to-side anastomosis of the donor portal vein to the superior mesenteric vein | 0
end-to-end bile duct anastomosis | 0
massive venous bleeding from local varices | 0
iliac conduit construction | 0
recovered well after surgery | 0
normal liver graft function | 0
stenosis of the bile duct anastomosis | 2160
biliary leakage | 2160
elevated liver enzymes | 2160
pigtail placement | 2160
FCSCEMS insertion | 2268
persisting leakage | 2268
stent extraction | 2592
hepatitis C reinfection | 2592
recurrent stenosis of the biliary anastomosis | 2592
ERCP | 2592
balloon dilatations | 2592
pigtail placements | 2592
stent placements | 2592
biopsy-proven significant fibrosis | 8760
treatment with pegylated interferon and ribavirin | 8760
elective ERCP | 10296
recovery of 3 plastic double-pigtails | 10296
cholangiogram | 10296
large portobiliary fistula | 10296
slight hemobilia | 10296
placement of FCSEMS | 10296
prophylactic antibiotic treatment with ciprofloxacin | 10296
septic shock | 10344
admitted to the intensive care unit | 10344
hemodynamic support | 10344
empiric broad-spectrum antibiotic treatment | 10344
computed tomography | 10344
angiography | 10344
chronic obliteration of the iliac conduit | 10344
partial perfusion of the hepatic artery by gastroduodenal collaterals | 10344
anuric kidney failure | 10344
continuous venovenous hemofiltration | 10344
intermittent hemodialysis | 10344
recovered well | 10344
evaluation for liver re-transplantation | 10344
FCSEMS replacement | 10944
extraction of the lying FCSEMS | 10944
no evidence of persisting leakage | 10944
no relevant stenosis | 10944