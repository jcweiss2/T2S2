29 years old | 0
male | 0
admitted to the hospital | 0
intermittent fevers | -48
forehead headache | -48
consumed unpasteurized cooked beef | -48
type 2 diabetes mellitus | 0
fatty liver | 0
smoking | 0
drinking | 0
nuchal rigidity | 0
glucose high | 0
C-reactive protein high | 0
erythrocyte sedimentation rate high | 0
white blood cells normal | 0
red blood cells normal | 0
hemoglobin normal | 0
urea normal | 0
creatinine normal | 0
serum minerals normal | 0
autoimmune antibodies normal | 0
turbid cerebrospinal fluid | 0
leukocytes 2090/mm3 | 0
protein 233.85 mg/dL | 0
glucose 1.4 mmol/L | 0
pressure > 33 cmH2O | 0
Gram-positive rods | 0
L. monocytogenes | 192
ampicillin | 192
erythrocin | 192
meropenem | 192
penicillin | 192
sulfamethoxazole | 192
ceftriaxone | 0
meropenem | 48
fever | 48
sinus tachycardia | 48
tachypnea | 48
confusion | 48
bilateral horizontal nystagmus | 48
bilateral abducens nerve palsy | 48
dysarthria | 48
weakness of all four limbs | 48
transferred to ICU | 120
Glasgow Coma Scale score 12/15 | 120
Glasgow Coma Scale score 5/15 | 192
intubated and ventilated | 192
etimicin discontinued | 288
extraventricular drainage | 528
rehaemorrhagia of the lateral ventricle | 696
anisocoria | 696
died | 744
L. monocytogenes rhombencephalitis | 0
hydrocephalus | 336
intracranial hemorrhage | 336
abnormally high T2 flow attenuated inversion recovery signal | 96
prominent temporal horns with enlargement of the ventricles | 96
hemorrhage of the right pons | 336
gross hydrocephalus and hemorrhage | 336
significant dilatation of fourth ventricle | 528
no remission in lateral ventricles | 528
rehaemorrhagia of the lateral ventricle and a larger ventricular system | 696