13 years old | 0
male | 0
admitted to the hospital | 0
Joubert syndrome | -120 months
mitochondrial disease | -12 months
sepsis | -156 weeks
neonatal intensive care unit | -156 weeks
end-stage renal disease | -60 months
hemodialysis | -60 months
intracranial hemorrhage | -36 months
high blood pressure | -36 months
hyperkalemia-induced cardiac arrest | -24 months
cardiopulmonary resuscitation | -24 months
intensive care unit | -24 months
post-CPR care | -24 months
heart problems | -12 months
lung problems | -12 months
kidney problems | -12 months
hypotension | 0
norepinephrine infusion | 0
stuporous | 0
Glasgow coma scale score 11 | 0
percutaneous endoscopic gastrostomy tube | 0
mean blood pressure 90-106 mmHg | 0
heart rate 95-107 beats/min | 0
shallow breathing | 0
100% oxygen saturation | 0
pre-anesthetic assessment | 0
jaw small | 0
mouth slightly protruding | 0
short neck | 0
reduced cervical mobility | 0
airway management | 0
anesthesia induction | 0
oral airway | 0
stylets | 0
Macintosh direct laryngoscope | 0
video-laryngoscope | 0
fiberoptic bronchoscope | 0
supraglottic airway device | 0
endotracheal tube | 0
blood sugar 132 mg/dl | 0
noninvasive blood pressure | 0
electrocardiography | 0
pulse oximetry | 0
invasive blood pressure monitoring | 0
left radial artery cannulation | 0
train-of-four stimulation | 0
bispectral index monitoring | 0
propofol | 0
remifentanil | 0
rocuronium | 0
anesthesia started | 0
mask ventilation | 0
I-gel insertion | 0
I-gel removal | 0
tracheal intubation | 0
mechanical ventilation | 0
end-tidal carbon dioxide | 0
oxygen saturation | 0
operation lasted 45 min | 45
hemodynamics stable | 45
norepinephrine infusion 0.03-0.07 µg/kg/min | 45
TOF count 1-2 | 45
no additional injection of muscle relaxants | 45
no additional opioids | 45
spontaneous breathing returned | 45
BIS 73 | 45
TOF ratio 76% | 45
midazolam | 45
transferred to SICU | 45
ventilator applied | 45
synchronized intermittent mandatory ventilation mode | 45
FiO2 0.25 | 45
tidal volume 6 ml/kg | 45
respiratory rate 20 breaths/min | 45
pressure support 13 cmH2O | 45
Glasgow coma scale score 6 | 45
trachea extubated | 60
100% oxygen saturation | 60
venous blood gas analysis | 60
venous pH 7.30 | 60
PCO2 53 mmHg | 60
PO2 47 mmHg | 60
base excess 0.3 mmol/L | 60
SO2 78% | 60
glucose 130 mg/L | 60
lactate 0.3 mmol/L | 60