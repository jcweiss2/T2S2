65 years old | 0
female | 0
admitted to the hospital | 0
right flank pain | -168
fatigue | -168
diabetes mellitus | -8760
breast cancer | -87600
Glasgow Coma Scale: E4V5M6 | 0
blood pressure 77/55 mm Hg | 0
heart rate 120 beats/min | 0
temperature 36.2°C | 0
respiratory rate 42/min | 0
mildly distended abdomen | 0
right flank and costovertebral angle tenderness | 0
white bleed cell count 18.5x10^9/L | 0
hemoglobin 11.7 × 10^-1 g/L | 0
platelet 7.8×10^-5/L | 0
blood urea nitrogen 67.9 mg/dL | 0
creatinine 3.53 mg/dL | 0
sodium 124 mEq/L | 0
potassium 3.7 mEq/L | 0
chloride 84 mEq/L | 0
prothrombin time-international normalized ratio 1.29 | 0
blood glucose 543 mg/dL | 0
glycosylated hemoglobin A1c 12.1% | 0
metabolic acidosis | 0
pH 7.41 | 0
arterial oxygen pressure 101.6 mm Hg | 0
PaCO2 16.1 mm Hg | 0
bicarbonate 10.0 mEq/L | 0
base excess 12.1 mEq/L | 0
lactic acid 3.43 mmol/dL | 0
urinalysis showed white blood cell 3+ | 0
occult blood 3+ | 0
emphysematous changes in the right kidney | 0
right emphysematous pyelonephritis (EPN) class 3B | 0
admitted to the intensive care unit (ICU) | 0
meropenem administered | 0
vancomycin administered | 0
intravenous fluids administered | 0
vasopressors administered | 0
steroids administered | 0
intubated | 6
mechanical ventilation | 6
portable abdominal X-ray | 6
progression of emphysematous changes in the right kidney | 6
exploratory laparotomy | 6
swelling in Gerota’s fascia | 6
foul-smelling gas released | 6
renal parenchyma spongy and drained purulent material | 6
right nephrectomy | 6
copious irrigation | 6
abdomen closed | 6
Escherichia coli in blood culture | 24
Escherichia coli in urine culture | 24
Escherichia coli in purulent material culture | 24
antibiotics continued | 24
leukocytosis | 168
fever | 168
acute renal failure | 168
hemodialysis | 168
tracheostomy | 168
weaned from hemodialysis | 336
weaned from mechanical ventilation | 336
transferred to a rehabilitation hospital | 504