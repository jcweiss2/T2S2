60 years old | 0
female | 0
impaired consciousness | -72
atrial fibrillation | -672
dilated cardiomyopathy | -672
oral warfarin | -672
biventricular pacing implantable cardioverter defibrillator | -672
found lying at home | -1
transported to hospital | -1
arrival at hospital | 0
Japan Coma Scale score II-10 | 0
Glasgow Coma Scale score 14 | 0
no clear neurological deficits | 0
non-contrast head CT | 0
hemorrhage in third and fourth ventricles | 0
hemorrhage in bilateral lateral ventricles | 0
brain 3D-CTA | 0
spot enhancement on lateral wall of anterior horn of left lateral ventricle | 0
blood pressure control | 0
ventricular drainage not performed | 0
cerebral angiograph | 72
aneurysm at distal site of mLSA | 72
embolization | 72
endovascular treatment | 72
N-butyl-2-cyanoacrylate injection | 72
aneurysm embolization | 72
postoperative head CT | 96
no hemorrhagic complications | 96
no cerebral infarction | 96
sepsis triggered by pneumonia | 120
decrease in muscle strength | 120
disuse | 120
rehabilitation | 720
discharged | 720
modified Rankin Scale 1 | 720
intraventricular aneurysm | 0
distal medial lenticulostriate artery aneurysm | 0
primary intraventricular hemorrhage | 0
intracerebral hemorrhage | 0
subarachnoid hemorrhage | 0
hypertension | 0
arteriovenous malformation | 0
trauma | 0
Moyamoya disease | 0
cavernous malformation | 0
coagulation abnormalities | 0
spot sign | 0
intracerebral hematoma | 0
extravasation of contrast medium | 0
enlargement of hematoma | 0
bleeding in cerebral parenchyma | 0
primary vascular injury | 0
secondary vascular injury | 0
aneurysm regression | 0
spontaneous thrombosis | 0
transient aneurysm regression | 0
re-rupture | 0
idiopathic intraventricular aneurysms | 0
true aneurysm | 0
pseudoaneurysm | 0
pathological evaluation | 0
radical surgery | 0
trans-cortical approach | 0
trans-callosal approach | 0
cortical injury | 0
postoperative epilepsy | 0
endovascular treatment | 0
liquid embolic material | 0
coil embolization | 0
flow-directed catheter | 0
cerebral infarction | 0
apathy | 0
personality changes | 0
biventricular pacing implantable cardioverter defibrillator | 0
MRI evaluation | 0
postoperative CT | 0
proximal perforating artery embolization | 0
cerebral infarction risk | 0
embolization | 0
direct surgery | 0