83 years old | 0
male | 0
admitted to the hospital | 0
syncope | -24
fell to the ground | -24
leg ecchymosis | 0
anuric | 0
rhabdomyolysis-induced AKI | 0
sepsis | 0
acute prostatitis | 0
increased urea | 0
increased creatinine | 0
increased myoglobin | 0
increased CPK | 0
increased LDH | 0
increased CRP | 0
increased PCT | 0
increased total bilirubin | 0
increased direct bilirubin | 0
increased AST | 0
increased ALT | 0
increased PSA | 0
increased white blood cell count | 0
volume expansion | 0
diuretic treatment | 0
antibiotic treatment | 0
femoral central venous catheter placement | 0
HFR-Supra treatment | 0
myoglobin removal | 0
inflammatory status reduction | 0
fluid balance maintenance | 0
furosemide administration | 0
piperacillin/tazobactam administration | 0
meropenem administration | 0
HFR-Supra sessions | 0
myoglobin reduction | 120
CPK reduction | 120
LDH reduction | 120
CRP reduction | 120
PCT reduction | 120
femoral hemodialysis catheter removal | 144
right jugular central venous catheter placement | 144
on-line hemodiafiltration | 144
high-flux hemodialysis | 144
dialysis therapy prolongation | 144
urine output increase | 192
urea reduction | 504
creatinine reduction | 504
CRP reduction | 504
total bilirubin reduction | 504
AST reduction | 504
ALT reduction | 504
PSA reduction | 504
white blood cell count reduction | 504
discharge | 504
urea level at 6 months | 2160
creatinine level at 6 months | 2160
GFR at 6 months | 2160