18 years old|0
    male|0
    admitted to the emergency|0
    fever| -192
    abdominal discomfort| -192
    anorexia| -192
    persistent vomiting| -192
    decreased urine output| -24
    thrombocytopenia| -24
    leukopenia| -24
    elevated transaminases| -24
    admitted to the intensive care unit|0
    normal hemoglobin|0
    leukopenia|0
    thrombocytopenia|0
    deranged liver function tests|0
    deranged kidney function tests|0
    urea|0
    creatinine|0
    uric acid|0
    hemodialysis|0
    negative malaria tests|0
    negative IgM anti-HAV|0
    negative IgM anti-HEV|0
    negative HBsAg|0
    negative dengue serology|0
    proteinuria|0
    hematuria|0
    white blood cells in urine|0
    normal chest X-ray|0
    normal 2D-echocardiography|0
    hepatosplenomegaly|0
    splenic infarcts|0
    bulky distal body and tail of pancreas|0
    mild ascites|0
    raised amylase|0
    raised lipase|0
    negative autoimmune workup|0
    negative rickettsia tests|0
    negative post streptococcal glomerulonephritis tests|0
    negative Weil–Felix|0
    negative ASO titer|0
    negative COVID RT-PCR|0
    negative leptospiral serology|0
    negative urine culture|0
    myalgia|0
    leg pains|0
    elevated creatinine phosphokinase|0
    blood culture grew S. enterica serovar typhi|96
    acute hepatitis|0
    acute pancreatitis|0
    splenic infarcts|0
    acute renal failure|0
    lower gastrointestinal bleeding|120
    hemoglobin drop|120
    intravenous antibiotics|0
    blood transfusions|0
    hemodialysis|0
    afebrile|168
    no gastrointestinal bleed|168
    hemoglobin stabilized|168
    good urine output|168
    creatinine decreased|168
    discharged|168
    serial creatinine phosphokinase decline|168
    follow-up kidney function normal|312
    transaminases normal|312
    creatinine phosphokinase normal|312
    
    