54 years old | 0
African-American | 0
female | 0
admitted to the hospital | 0
fevers | -336
cough | -336
shortness of breath | -336
deep vein thrombosis | -3024
pulmonary embolism | -3024
anticoagulated with warfarin | -3024
oxygen saturation 99% | 0
blood pressure 100/70 mmHg | 0
heart rate 75 b.p.m. | 0
respiratory rate 30 breaths/min | 0
elevated D-dimer | 0
ferritin 683.2 ng/mL | 0
lactate dehydrogenase 929 U/L | 0
aspartate aminotransferase 190 U/L | 0
alanine aminotransferase 131 U/L | 0
decreased platelet count | 0
white blood cell count 3.9 | 0
absolute lymphocyte count 0.59 | 0
elevated probrain natriuretic peptide | 0
troponin elevation | 0
electrocardiogram showed right ventricular strain | 0
transthoracic echocardiogram showed dilated right ventricle | 0
McConnell’s sign | 0
computed tomography angiography showed bilateral pulmonary emboli | 0
respiratory failure | 0
intubated | 0
ARDS | 0
right ventricular thrombus | 24
azithromycin | 0
doxycycline | 24
hydroxychloroquine | 24
intravenous heparin | 24
enoxaparin | 336
catheter-directed thrombolysis discussed | 24
extubated | 336
transferred to step-down unit | 408
transferred to general medical floors | 408
discharged to inpatient rehabilitation unit | 456
right popliteal deep vein thrombosis | 408
D-dimer remained elevated | 456
therapeutic dose of enoxaparin | 456
SARS-CoV-2 positive | 96
COVID-19 PCR | 96
inpatient rehabilitation therapy | 456
hoarse voice | 336
improved daily | 408
follow-up with primary care physician | 456
follow-up with primary cardiologist | 456