46 years old | 0
    male | 0
    road traffic collision | -336
    erythematous changes over the trunk | -336
    chest to abdomen erythema | -336
    severe abnormalities of the extremities | -336
    bilateral lung contusions | -336
    mild hemothorax | -336
    right third to fifth rib fractures | -336
    liver laceration | -336
    minor active bleed | -336
    trans-arterial embolization of the right hepatic artery | -336
    admitted to ICU | 0
    sinus tachycardia | 0
    ventricular premature complex | 0
    elevated troponin-I | 0
    echocardiogram arranged | 0
    no cardiac wall abnormality | 0
    no pericardial effusion | 0
    pigtail chest catheter placed | 96
    subsequent echocardiogram | 96
    progression of left pleural effusion | 96
    no pleural effusion over the right costophrenic angle | 96
    dark red drainage fluid | 96
    CXR rechecked | 96
    improvement in hemithorax white-out | 96
    improvement in fluid amount | 96
    pigtail catheter size not revised | 96
    transferred to regular ward | 240
    chest pigtail catheter removed | 240
    shortness of breath | 288
    recurrent massive left pleural effusion | 288
    echo-guided pigtail insertion | 288
    minimal turbid fluid drained | 288
    culture positive for Staphylococcus aureus | 288
    symptoms temporarily improved | 288
    severe chest pain | 336
    worsening shortness of breath | 336
    frequent VPC | 336
    cardiomegaly observed | 336
    CT scan | 336
    severe purulent pericardial effusion | 336
    suspected purulent pericarditis | 336
    cardiac tamponade | 336
    pericardiectomy | 336
    debridement | 336
    purulent exudate removal | 336
    RA/SVC junction tear repair | 336
    penicillin beta-lactam antibiotic | 336
    oxacillin administered | 336
    gentamycin administered | 336
    dyspnea | 504
    desaturation | 504
    follow-up CT | 504
    bilateral lung pleural effusion | 504
    empyema | 504
    decortication surgery | 504
    multiple bilateral loculated effusions | 504
    exudates removed | 504
    intravenous antibiotics | 504
    discharged | 720
    