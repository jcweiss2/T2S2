76 years old | 0 | 0 
male | 0 | 0 
admitted to the hospital | 0 | 0 
pancreatic adenocarcinoma | -672 | 0 
metastasis to the liver | -672 | 0 
diastolic heart failure | -672 | 0 
atrial fibrillation | -672 | 0 
coronary artery disease | -672 | 0 
severe hyponatremia | 0 | 0 
sodium level of 116 mmol/L | 0 | 0 
x-ray findings consistent with pneumonia | 0 | 0 
broad-spectrum antibiotics | 0 | 24 
fluid for hyponatremia | 0 | 24 
transferred to the intensive care unit | 0 | 0 
jugular vein distention | 0 | 0 
lower extremity pitting edema | 0 | 0 
transthoracic echocardiogram | 0 | 0 
left ventricular cavity size normal | 0 | 0 
mildly reduced systolic function | 0 | 0 
septal flattening | 0 | 0 
left atrial enlargement | 0 | 0 
suspected MV vegetation | 0 | 0 
severe mitral regurgitation | 0 | 0 
tricuspid regurgitation | 0 | 0 
elevated RV systolic pressure | 0 | 0 
type 2 and type 3 pulmonary arterial hypertension | 0 | 0 
ill-defined thickening in the TV leaflets | 0 | 0 
afebrile | 0 | 0 
leukocytosis | 0 | 0 
recent urethral instrumentation | -24 | 0 
blood cultures obtained | 0 | 0 
infectious disease specialist consulted | 0 | 0 
transesophageal echocardiogram | 24 | 24 
normal left ventricular size and function | 24 | 24 
normal RV size and function | 24 | 24 
hypermobile interatrial septum | 24 | 24 
no left atrial or left atrial appendage thrombus | 24 | 24 
vegetations on the atrial aspect of MV leaflets | 24 | 24 
severe mitral regurgitation | 24 | 24 
systolic flow reversal in the pulmonary vein | 24 | 24 
vegetation on the TV leaflet | 24 | 24 
tricuspid regurgitation | 24 | 24 
RVSP 47 mm Hg | 24 | 24 
blood cultures negative | 24 | 48 
polymerase chain reaction testing negative | 24 | 48 
workup for antiphospholipid syndrome unremarkable | 24 | 48 
marantic endocarditis suspected | 24 | 48 
apixaban discontinued | -168 | 0 
low molecular weight heparin or unfractionated heparin recommended | 48 | 0 
computed tomography imaging of the head | 48 | 48 
infectious disease recommended discontinuation of broad-spectrum antibiotics | 48 | 48 
enoxaparin started | 72 | 0 
platelets recovered to above 50,000 109/L | 72 | 72 
expired | 168 | 168