3-year-old | 0
female | 0
intermittent fever | -144
drowsiness | -24
second child | 0
no family history of neurological disorders | 0
full-term cesarean section | 0
non-consanguineous marriage | 0
no birth complications | 0
nodding spasm | -17520
no treatment for nodding spasm | -17520
no intellectual developmental disorder | 0
no developmental language delay | 0
no history of liver disease | 0
no substance abuse | 0
intermittent seizures | -432
electroencephalogram spiked slow waves | -432
multi-spiked slow waves | -432
generalized spiked waves | -432
decreasing dominant rhythm in occipital region | -432
video-EEG myoclonic seizures | -432
no positive routine blood findings | -432
no positive liver function findings | -432
no positive kidney function findings | -432
no positive electrolyte test results | -432
no positive computed tomography scan of head | -432
epilepsy diagnosis | -432
myoclonia diagnosis | -432
sodium valproate treatment | -432
epilepsy well controlled | -432
discharged after previous admission | -432
continue sodium valproate | -432
routine blood tests | 0
liver function tests | 0
kidney function tests | 0
electrolyte tests | 0
MOF | 0
hemophagocytic syndrome | 0
jaundice | 0
drowsiness at admission | 0
anuria | 0
bilateral pupil size | 0
sensitivity to light reflex | 0
temperature 36.8 °C | 0
pulse rate 103 beats per minute | 0
respiratory rate 22 breaths per minute | 0
blood pressure 109/67 mmHg | 0
oxygen saturation 99% | 0
height 103 cm | 0
body weight 17 kg | 0
pharyngeal congestion | 0
low and dull cardiac sounds | 0
hepatomegaly | 0
no other abnormalities | 0
hemoglobin 77 g/L | 0
platelet 68×109/L | 0
troponin I elevated | 0
NT-proBNP elevated | 0
hyperbilirubinemia | 0
hypoalbuminemia | 0
serum creatinine elevated | 0
electrolyte disturbance | 0
PT increased | 0
APTT increased | 0
D-dimer increased | 0
fibrinogen decreased | 0
interleukin-2 receptor elevated | 0
serum ferritin elevated | 0
serum aminotransferases elevated | 0
lactate dehydrogenase elevated | 0
hyperlactatemia | 0
hyperammonemia | 0
no positive pathogen findings | 0
hepatomegaly on abdominal ultrasound | 0
thickening of gallbladder wall | 0
no positive cardiac ultrasound | 0
no positive kidney ultrasound | 0
acute liver failure | 0
grade 3 acute kidney injury | 0
disseminated intravascular coagulation | 0
meropenem treatment | 0
methylprednisolone treatment | 0
plasma exchange | 0
hemodialysis | 0
immunosupportive therapy | 0
component transfusion | 0
organ protection | 0
sodium valproate discontinued | 0
pulmonary hemorrhage | 36
respiratory failure | 36
mechanical ventilation | 36
genetic metabolic disease considered | 0
peripheral blood DNA extraction | 0
plasma exchange performed 4 times | 0
hemodialysis performed 5 times | 0
remained unconscious | 0
anuria persisted | 0
MOF uncorrected | 0
parents decided to forgo treatment | 0
patient died | 0
NEXMIF heterozygous variant | 0
other variants detected | 0
no mitochondrial abnormalities | 0
de novo variant in NEXMIF | 0
no pathogenic variants in parents | 0
