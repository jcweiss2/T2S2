23 years old | 0
woman | 0
admitted to Medical Intensive Care Unit | 0
organophosphorus poisoning | 0
mechanical ventilation | 0
ionotropic support | 0
left femoral artery catheter inserted | 0
fever | 168
tachycardia | 168
erythematous papules on the left lower limb | 216
white blood cell count 16,500/mm3 | 216
neutrophils 84% | 216
lymphocytes 12% | 216
monocytes 3% | 216
eosinophils 1% | 216
blood cultures sent | 216
intra-arterial catheter removed | 216
skin lesions biopsied | 216
skin lesions became blackish with necrotic areas | 240
blood cultures yielded Pseudomonas aeruginosa | 240
catheter tip cultures yielded Pseudomonas aeruginosa | 240
skin lesion cultures yielded Pseudomonas aeruginosa | 240
Pseudomonas aeruginosa sensitive to ceftazidime | 240
biopsy of the skin lesion revealed acute neutrophilic infiltration | 240
necrotic area | 240
treated with ceftazidime | 240
lesions resolved completely | 480
full recovery from organophosphorus poisoning | 480
discharged home | 480
ecthyma gangrenosum | 240