54 years old | 0
male | 0
admitted to the hospital | 0
shortness of breath | -168
multiple episodes of seizure | -168
right lung non-small cell lung cancer (squamous cell carcinoma) | 0
metastasis to brain | 0
superior vena caval syndrome (stage IV) | 0
started on tab phenytoin 300 mg at bedtime | 0
anti-edema measures with steroids (tab dexamethasone 8 mg 3 times daily during RT) | 0
tapered over 2 weeks post RT | 0
received palliative RT to the mediastinum and whole brain | 0
total dose of 20 Gray in 5 fractions over one week with Co-60 gamma rays | 0
two weeks post radiotherapy | 336
general condition improved | 336
received one cycle of palliative chemotherapy with paclitaxel-carboplatin combination | 336
three weeks after completing the RT | 504
presented with painful, erythematous lesions in the scalp | 504
lesions generalized | 504
afebrile | 504
pulse rate 98/min | 504
respiratory rate 28/min | 504
blood pressure 109/83 mm Hg | 504
features of mild dehydration | 504
erythematous, tender macules over the scalp, face, trunk, and limbs | 504
confluent epidermal detachment | 504
blistering involving almost 30% of his body surface area | 504
conjunctivitis | 504
hemorrhagic crusting on lips | 504
erosions over buccal and nasal mucosa | 504
erosions over the glans penis | 504
TEN caused by phenytoin | 504
hemogram normal | 504
biochemical parameters normal | 504
hyponatremia | 504
phenytoin immediately discontinued | 504
managed with intravenous fluid replacement | 504
electrolyte correction | 504
systemic antibiotics | 504
steroids (dexamethasone 16 mg/day tapered at 2 mg/day over one week) | 504
local skin care with antibiotic and antifungal dressings | 504
condition worsened | 504
died due to septicemia | 504
seventh day of hospital admission | 168
acute onset | 504
painful skin lesions | 504
fever >39°C (102.2°F) | 504
sore throat | 504
oral mucosal complications | 504
ocular mucosal complications | 504
rapidly spreading confluent and extensive epidermal detachment | 504
dehydration | 504
dyselectrolytemia | 504
systemic disease | 504
mortality 25-35% | 504
risk factors: age >40 years | 504
risk factors: malignancy | 504
risk factors: heart rate >120/min | 504
risk factors: initial percentage of epidermal detachment over 10% | 504
risk factors: serum urea >10 mmol/litre | 504
risk factors: serum glucose >14 mmol/litre | 504
risk factors: bicarbonate <20 mmol/litre | 504
aromatic anticonvulsants (phenytoin, phenobarbitone, carbamazapine) as high risk agents | 504
phenytoin use for seizure control | 504
phenytoin use for prophylactic use in brain metastasis | 504
risk of TEN 8.3 per 10,000 new users | 504
occurs within 8 weeks of drug use | 504
radiation alone not resulted in SJS-TEN syndrome | 504
concurrent use of whole brain RT and phenytoin induces cutaneous type IV hypersensitivity reactions | 504
erythema multiforme (EM) | 504
SJS | 504
TEN | 504
first case reported by Delattre et al | 504
EMPACT syndrome | 504
dusky macules in the RT portal | 504
spread to other regions | 504
eruptive disorder with systemic involvement | 504
immunologically mediated type IV hypersensitivity to phenytoin and metabolites | 504
augmented by concurrent use of RT | 504
lesions in non-cranial RT sites | 504
component of concurrent whole brain RT as trigger | 504
carboplatin based chemotherapy as potential trigger | 504
management in intensive care unit | 504
immediate cessation of phenytoin | 504
fluid replacement | 504
electrolyte replacement | 504
systemic steroids | 504
antibiotics | 504
local wound care | 504
high dose corticosteroids within 24-48 hours of TEN | 504
rapid tapering over 2 weeks | 504
increased mortality from sepsis | 504
gastrointestinal bleed | 504
delayed wound healing | 504
use of phenytoin avoided during RT | 504
replaced with sodium valproate, benzodiazepines, gabapentin, or topiramate | 504
complications anticipated and managed aggressively | 504
disclosure of no conflicts of interest | 504
funded by Sultan Qaboos University Hospital | 504
