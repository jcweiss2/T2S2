22 years old | 0
African American | 0
female | 0
admitted to the emergency room | 0
worsening respiratory distress | -336
drooping of eyelids | -336
systemic lupus erythematosus (SLE) | -3960
lupus nephritis | -3960
cyclophosphamide | -3960
mycophenolate | -3960
azathioprine | -672
prednisone | -672
hypothyroidism | 0
hypertension | 0
myasthenia gravis | 0
acute hypoxic respiratory failure | 0
endotracheal intubation | 0
mechanical ventilation | 0
febrile | 0
tachycardia | 0
decreased breath sounds | 0
pneumonia | 0
respiratory muscle weakness | 0
myasthenia crisis | 0
sepsis | 0
plasmapheresis | 0
steroids | 0
antimicrobial agents | 0
pyridostigmine | 24
increased bronchial secretions | 0
hypotensive | 192
oliguria | 192
acute renal failure | 192
acute tubular necrosis (ATN) | 192
abdominal tenderness | 216
abdominal computed tomography (CT) scan | 216
free air in the abdominal cavity | 216
emergent laparotomy | 216
peritonitis | 216
gastric cardia perforation | 216
worsening coagulation panel | 0
worsening liver function tests | 0
prothrombin time (PT) increased | 0
albumin level decreased | 0
bilirubin level stable | 0
alkaline phosphatase level stable | 0
aspartate aminotransferase (AST) level increased | 0
alanine aminotransferase (ALT) level increased | 0
AST level peaked | 240
ALT level peaked | 240
acute respiratory distress syndrome | 360
fatal cardiac arrest | 360
disseminated herpes | 0
herpetic hepatitis | 0
liver failure | 0
gastric perforation | 216
peritonitis | 216
pneumonia | 0
ARDS | 360
fulminant hepatic failure | 360
death | 360
acyclovir therapy | 0
liver transplantation | 0
lifelong acyclovir prophylaxis | 0