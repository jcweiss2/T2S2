63 years old | 0
African-American | 0
male | 0
presented | 0
food aversion | -96
subjective fevers | -96
chills | -96
chest pain | -96
abdominal pain | -96
remote history of tobacco use | -96
remote history of cocaine use | -96
no diabetes mellitus | 0
no medical illnesses | 0
not on prescription medications | 0
not on over-the-counter medications | 0
fever of 38.3°C | 0
hemodynamically stable | 0
poor dentition | 0
white cell count of 22.4 × 10^9/L | 0
aspartate aminotransferase of 93 units/L | 0
alanine aminotransferase of 110 units/L | 0
total bilirubin of 1.2 mg/dL | 0
computed tomography of chest | 0
computed tomography of abdomen | 0
computed tomography of pelvis | 0
multiple indeterminate hypoAattenuating lesions throughout liver | 0
abdominal sonogram | 0
multiple complex hypoechoic foci throughout liver | 0
magnetic resonance imaging of abdomen | 0
multiple cystic lesions with enhancing internal septations | 0
marked diffusion restriction | 0
largest lesion measured 4.5 cm × 4.1 cm × 3.8 cm | 0
empiric treatment with broad-spectrum antibiotics initiated | 0
immediate resolution of fever | 24
aspiration from one abscess cavity | 24
placement of three drainage catheters in right hepatic lobe | 24
drainage grew Fusobacterium nucleatum | 24
antibiotics narrowed based on culture and sensitivities | 24
liver aspirate testing for acid-fast organisms negative | 24
aerobic cultures negative | 24
fungal cultures negative | 24
stool cultures negative | 24
examination for ova negative | 24
examination for parasites negative | 24
examination for giardia negative | 24
examination for cryptosporidium negative | 24
examination for clostridium difficile negative | 24
examination for entamoeba negative | 24
blood cultures negative | 24
urine cultures negative | 24
testing for viral hepatitis negative | 24
testing for human immunodeficiency virus negative | 24
tumor markers for alpha-fetoprotein unremarkable | 24
cancer antigen 19-9 unremarkable | 24
carcinoembryonic antigen unremarkable | 24
trans-thoracic echocardiogram revealed no valvular vegetations | 24
colonoscopy | 24
two 4-8 mm adenomatous polyps in rectum | 24
mild diverticulosis in sigmoid colon | 24
no evidence of prior inflammation | 24
no evidence of current inflammation | 24
no evidence of infection | 24
panorex demonstrated multiple missing teeth | 24
lucency around root of left mandibular premolar | 24
likely periapical abscess | 24
output from hepatic drains continued to decrease | 336
drains removed | 336
affected teeth extracted | 336
antibiotics transitioned to oral route | 336
discharged home | 672
asymptomatic at 6 weeks post-hospitalization | 1008
liver enzymes trended down to normal levels | 1008
repeat cross-sectional imaging | 1008
significant interval decrease in rim enhancement | 1008
significant interval decrease in size of liver abscesses | 1008
treatment response | 1008
