17 years old | 0
    female | 0
    infective endocarditis | -72
    intravenous antibiotics | -72
    vegetations in mitral valve leaflet | -72
    Staphylococcus aureus | -72
    sudden deterioration of mental status | 0
    disoriented | 0
    dizzy | 0
    high-grade fever | 0
    intracranial abscess | 0
    mycotic aneurysm of the right cerebral hemisphere | 0
    no evidence of rupture of aneurysm | 0
    no significant mass effect | 0
    conservative treatment | 0
    neurosurgical consultation upon discharge | 0
    discharged | 0
    