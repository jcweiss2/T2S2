61 years old | 0
    male | 0
    presented with 2-month history of systemic erythema | -1440
    presented with 1.5-month history of oedema of the lower limbs | -1080
    administered allopurinol tablets two months ago | -1440
    developed systemic rash | -1440
    rash scattered throughout the body | -1440
    granular with dark red papules | -1440
    accompanied by scratches | -1440
    partial ulceration | -1440
    scabs | -1440
    denied cough | 0
    denied cold | 0
    denied fever | 0
    denied joint pain | 0
    denied diarrhea | 0
    denied urinary symptoms | 0
    elevated white blood cell count (32.3 × 109/L) | -1440
    91.6% neutrophils | -1440
    2.6% eosinophils | -1440
    high C-reactive protein (175 mg/L) | -1440
    high ALT (133 U/L) | -1440
    diagnosed with drug-induced dermatitis | -1440
    given 60 mg glucocorticoid once a day | -1440
    reduced by 8 mg every 5 days | -1440
    loratadine | -1440
    cetirizine | -1440
    rash disappeared | -1440
    discharged | -1440
    presented with oedema of both lower limbs | -1080
    particularly the right lower limb | -1080
    redness on the back of the foot | -1080
    local tenderness | -1080
    higher skin temperatures | -1080
    history of hypertension (5 years) | 0
    history of secondary diabetes (2 months) | 0
    blood pressure 129/86 mmHg | 0
    heart rate 124 beats/min | 0
    temperature 38.7 °C | 0
    respiration 17 breaths per minute | 0
    saturation 95% without oxygen | 0
    localized red-purplish discoloration on both lower limbs | 0
    clear chest | 0
    soft abdomen | 0
    no guarding | 0
    no rigidity | 0
    white blood cell count 13.2 × 109/L | 0
    neutrophilia 93% | 0
    hemoglobin 79 g/L | 0
    elevated CRP 302 mg/L | 0
    elevated procalcitonin 2.84 ng/mL | 0
    degraded albumin 24 g/L | 0
    serum creatinine 4.95 mg/dL | 0
    elevated B-type natriuretic peptide 1791.6 pg/mL | 0
    glycosylated haemoglobin 9.2% | 0
    metabolic acidosis (pH: 7.32; base excess: -6.0 mEq/L) | 0
    normal blood electrolyte | 0
    normal liver function | 0
    chest radiography unremarkable | 0
    other laboratory data unremarkable | 0
    ultrasonography showed oedema of the dorsum of the feet | 0
    suspected intermuscular abscess of the right calf | 0
    MRI revealed multiple muscle and subcutaneous soft tissue swelling | 0
    intermuscular abscesses observed | 0
    diagnosed with necrotizing fasciitis caused by Staphylococcus aureus | 0
    started on cefoperazone/sulbactam (2g every 8h) | 0
    started on caspofungin (50mg daily) | 0
    received serum albumin intravenously | 0
    received fluids intravenously | 0
    immunoglobulins administered | 0
    blood glucose monitored | 0
    insulin injected subcutaneously | 0
    ultrasound-guided abscess puncture and drainage performed | 24
    105 mL bloody purulent fluid drained | 24
    temperature dropped to 37.4 °C | 48
    white blood cell count 10.5 × 109/L | 48
    neutrophilia 88.9% | 48
    CRP 128.50 mg/L | 48
    Gram staining showed Gram-positive cocci | 24
    culture confirmed Staphylococcus aureus | 24
    blood culture confirmed Staphylococcus aureus | 24
    sputum culture negative | 24
    methicillin-resistant Staphylococcus aureus not isolated | 24
    linezolid intravenous injection | 24
    fever recurrence | 72
    second ultrasound showed abscess narrowed | 72
    drainage not smooth | 72
    little purulent fluid drained daily | 72
    MRI confirmed multiple abscesses | 72
    surgical debridement of necrotic tissue within 48h | 72
    necrotic tissue in deep fascia greyish | 72
    purulent fluid confirmed diagnosis | 72
    culture of necrotic tissues revealed Staphylococcus infection | 72
    postoperative vacuum sealing drainage (VSD) | 72
    negative pressure maintained 40-60 kPa | 72
    saline continuous irrigation | 72
    second debridement for unhealed right leg | 168
    sudden cough with 3 mL bloody sputum | 240
    shortness of breath | 240
    saturation 93% with 33% oxygen | 240
    wheezes in both lungs | 240
    echocardiography showed left ventricular enlargement | 240
    ejection fraction 57% | 240
    pericardial effusions | 240
    hemoglobin 67 g/L | 240
    elevated brain natriuretic peptide (>9000 ng/mL) | 240
    elevated lactate dehydrogenase | 240
    CT scan showed acute bilateral pulmonary oedema | 240
    pleural effusions at base of both lungs | 240
    multi-disciplinary treatment organized | 240
    non-invasive positive pressure ventilation | 240
    glucocorticoids for toxaemia | 240
    diuretics used | 240
    intravenous fluid input adjusted | 240
    immunoglobulin administered | 240
    thymosin administered | 240
    red blood cells infused | 240
    erythropoietin supplementation | 240
    repeated CT scans showed pulmonary oedema absorption | 312
    pleural fluid absorption | 312
    repeated debridement once a week | 384
    total of 6 debridements | 2688
    skin grafting performed on dorsum of right foot | 2688
    discharged after 4 months | 2880
    alive with well-controlled diabetes during follow-up | 2880
    
    <|eot_id|>
    61 years old | 0
male | 0
admitted to the hospital | 0
systemic erythema | -1440
oedema of the lower limbs | -1080
allopurinol administration | -1440
systemic rash | -1440
rash scattered throughout the body | -1440
granular dark red papules | -1440
scratches | -1440
partial ulceration | -1440
scabs | -1440
no cough | 0
no cold | 0
no fever | 0
no joint pain | 0
no diarrhea | 0
no urinary symptoms | 0
elevated white blood cell count (32.3 × 109/L) | -1440
neutrophils 91.6% | -1440
eosinophils 2.6% | -1440
high CRP (175 mg/L) | -1440
high ALT (133 U/L) | -1440
diagnosed with drug-induced dermatitis | -1440
glucocorticoid 60 mg daily | -1440
glucocorticoid reduced by 8 mg every 5 days | -1440
loratadine | -1440
cetirizine | -1440
rash disappearance | -1440
discharged | -1440
oedema of both lower limbs | -1080
right lower limb oedema | -1080
redness on back of foot | -1080
local tenderness | -1080
higher skin temperatures | -1080
hypertension (5 years) | 0
secondary diabetes (2 months) | 0
blood pressure 129/86 mmHg | 0
heart rate 124 beats/min | 0
temperature 38.7 °C | 0
respiration 17 breaths/min | 0
saturation 95% without oxygen | 0
red-purplish discoloration on lower limbs | 0
clear chest | 0
soft abdomen | 0
no guarding | 0
no rigidity | 0
white blood cell count 13.2 × 109/L | 0
neutrophilia 93% | 0
hemoglobin 79 g/L | 0
CRP 302 mg/L | 0
procalcitonin 2.84 ng/mL | 0
albumin 24 g/L | 0
serum creatinine 4.95 mg/dL | 0
B-type natriuretic peptide 1791.6 pg/mL | 0
glycosylated haemoglobin 9.2% | 0
metabolic acidosis | 0
normal electrolytes | 0
normal liver function | 0
unremarkable chest radiography | 0
unremarkable other labs | 0
ultrasound showed dorsum oedema | 0
suspected right calf abscess | 0
MRI soft tissue swelling | 0
intermuscular abscesses | 0
diagnosed with necrotizing fasciitis | 0
cefoperazone/sulbactam started | 0
caspofungin started | 0
serum albumin administered | 0
fluids administered | 0
immunoglobulins given | 0
blood glucose monitoring | 0
insulin therapy | 0
ultrasound-guided drainage | 24
105 mL purulent fluid drained | 24
temperature drop to 37.4 °C | 48
white blood cell count 10.5 × 109/L | 48
neutrophils 88.9% | 48
CRP 128.50 mg/L | 48
Gram-positive cocci | 24
Staphylococcus aureus culture | 24
blood culture positive | 24
sputum culture negative | 24
methicillin-resistant S. aureus negative | 24
linezolid started | 24
fever recurrence | 72
second ultrasound abscess narrowed | 72
drainage not smooth | 72
daily purulent fluid | 72
MRI confirmed abscesses | 72
surgical debridement | 72
greyish necrotic tissue | 72
purulent fluid presence | 72
Staphylococcus culture from tissue | 72
VSD applied | 72
negative pressure 40-60 kPa | 72
saline irrigation | 72
second debridement | 168
cough with bloody sputum | 240
shortness of breath | 240
saturation 93% on oxygen | 240
wheezes in lungs | 240
left ventricular enlargement | 240
ejection fraction 57% | 240
pericardial effusions | 240
hemoglobin 67 g/L | 240
elevated BNP | 240
elevated lactate dehydrogenase | 240
CT bilateral pulmonary oedema | 240
pleural effusions | 240
multi-disciplinary treatment | 240
non-invasive ventilation | 240
glucocorticoids for toxaemia | 240
diuretics used | 240
fluid input adjusted | 240
immunoglobulin boost | 240
thymosin administered | 240
red blood cell transfusion | 240
erythropoietin given | 240
CT showed oedema absorption | 312
pleural fluid absorption | 312
repeated debridements weekly | 384
total 6 debridements | 2688
skin grafting | 2688
discharged after 4 months | 2880
alive with controlled diabetes | 2880