84 years old| 0
male| 0
dementia| 0
fever| -96
upper respiratory infection| -96
decline in blood pressure| -24
decrease in SpO2| -24
loss of consciousness| -24
referred to hospital| -24
respiratory failure| 0
shock| 0
blood pressure 77/48 mmHg| 0
pulse rate 107 beats per minute| 0
SpO2 84% with oxygen administration| 0
respiratory rate 32 breaths per minute| 0
body temperature 38.3℃| 0
coarse crackles on bilateral lung fields| 0
altered consciousness JCS III-200| 0
Glasgow Coma Scale 3 (E1V1M1)| 0
chest radiograph diffuse consolidation| 0
CT scan diffuse consolidation| 0
leukocytosis 27,180 /μL| 0
neutrophilia 98%| 0
high C-reactive protein 19.30 mg/dL| 0
slight elevation of liver enzymes| 0
hypoproteinemia| 0
renal dysfunction| 0
high creatine kinase| 0
thrombocytopenia| 0
prolonged prothrombin time| 0
elevated fibrin degradation products| 0
disseminated intravascular coagulopathy (DIC)| 0
septic shock| 0
severe aspiration pneumonia| 0
APACHEII score 30| 0
SOFA score 15| 0
meropenem hydrate 1.5 g/day| 0
dopamine hydrochloride 3 μg/kg/min| 0
nafamostat mesylate 0.07 mg/kg/hr| 0
nasogastric feeding tube insertion| 48
enteral nutrition started| 72
polymeric formula 5 kcal/kg/day| 72
infusion dose increased| 72
fever 39.5℃| 192
persistent decrease in SpO2 <90%| 192
white blood cell count 39,020 /μL| 192
chest radiograph fresh infiltrations| 192
aspiration from gastric feed reflux| 192
enteral feeding discontinued| 192
nasojejunal tube insertion| 240
jejunal feeding| 240
gastric decompression| 240
enteral feeding recommenced| 240
feeding dose increased| 240
gastric drainage volume 50-450 mL/day| 240
no drainage of enteral feed| 240
no recurrence of high grade fever| 240
no persistent decrease in SpO2| 240
evaluation by dysphagia team| 528
oral intake not safe| 528
percutaneous endoscopic gastrostomy (PEG)| 528
upper gastrointestinal endoscopy| 528
postoperative clinical course uneventful| 720
transferred to rehabilitation ward| 720
swallowing therapy| 1032
discharge| 1032
dopamine hydrochloride discontinued| 72
nafamostat mesylate discontinued| 120
meropenem hydrate discontinued| 336
sulfamethoxazole administered| 336
penicillin-susceptible streptococcus pneumoniae isolated| 0
