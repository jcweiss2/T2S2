60 years old | 0
female | 0
diabetes mellitus | -672
fever | -72
pain in the throat | -72
skin rash | -72
high CRP | -72
high sedimentation rate | -72
antibiotics | -72
admitted to hospital | 0
high P-CRP | 0
high B-leukocytes | 0
intravenous antibiotic with cefotaxime | 0
low systolic blood pressure | 24
confusion | 24
intensive skin rash | 24
fever persisted | 24
admitted to intensive care unit | 24
high ferritin level | 24
Still's disease suspected | 24
high Protrombinkomplex International Normalized Ratio | 24
high activated partial thromboplastin time | 24
elevated fibrin D-dimers | 24
low fibrinogen | 24
high CRP | 24
high blood sedimentation rate | 24
anemia | 24
thrombocytopenia | 24
leukopenia | 24
high procalcitonin | 24
meropenem | 24
gensumycin | 24
fluconazole | 24
high triglyceride values | 48
high soluble CD25R | 48
HLH diagnosis confirmed | 48
bone-marrow biopsy | 48
no signs of lymphoma or other malignancies | 48
skin biopsy | 48
non-specific inflammation | 48
18F-FDG PET/CT scan | 72
symmetrical and bilateral uptakes in lymph nodes | 72
no antibodies against parvovirus B19 | 72
no antibodies against Human Immunodefficiency Virus | 72
no antibodies against HHV 6 and 8 | 72
no antibodies against influenza A and B | 72
no antibodies against adenovirus | 72
no antibodies against coronavirus | 72
no antibodies against Respiratory syncytial virus | 72
elevated IgG against HSV | 72
elevated IgG against Varicella Zoster Virus | 72
EBV load of 2,400 copies/mL | 72
steroid treatment started | 96
60 mg prednisolone | 96
16.5 mg dexamethasone | 96
duration of therapy 3 months and 17 days | 96
dose gradually decreased | 120
therapy discontinued | 744
good response to steroid therapy | 168
no treatment with etoposide or cyclosporine | 168
fever disappeared | 168
blood pressure improved | 168
general condition improved | 168
skin rash decreased | 168
hemoglobin increased | 168
platelets increased | 168
ferritin decreased | 168
intense fatigue | 240
admitted to rehabilitation unit | 240
improvement of general condition | 336
normalized plasma ferritin | 744
no signs of HLH activation | 744