53 years old | 0
    female | 0
    presented with dizziness | -168
    presented with worsening shortness of breath | -168
    presented with increasing chest pressure | -168
    urinary tract infection | -672
    culture positive for Abiotrophia defectiva | -672
    sulfamethoxazole-trimethoprim 800/160 mg twice per day for a week | -672
    intramuscular injection of ceftriaxone | -672
    oral ciprofloxacin 500 mg twice per day for 7 days | -672
    admitted to hospital | 0
    lethargic | 0
    temperature 36.7°C | 0
    blood pressure 104/88 mmHg | 0
    heart rate 175 beats per minute | 0
    respiratory rate 21 breaths per minute | 0
    oxygen saturation 98% on room air | 0
    chest radiography unremarkable | 0
    electrocardiogram showed atrial fibrillation | 0
    atrial fibrillation with rapid ventricular rate to 180 beats per minute | 0
    brain natriuretic peptide elevated 819 pg/mL | 0
    initial troponin I 0.1 ng/mL | 0
    repeat troponin I 0.34 ng/mL | 0
    heparin infusion started | 0
    diltiazem infusion started | 0
    improvement in heart rate control | 0
    lactic acidosis | 0
    acute kidney injury | 0
    creatinine 1.62 mg/dL | 0
    thrombocytopenia 29,000/mm3 | 0
    transthoracic echocardiogram showed thickened and restricted mitral valve | 0
    large vegetation 21 mm x 19 mm on posterior leaflet | 0
    partial flail | 0
    severe regurgitation | 0
    vegetation obstructing inflow into left ventricle | 0
    stenotic physiology | 0
    aortic valve thickened | 0
    perforation of non-coronary cusp | 0
    ejection fraction normal | 0
    right ventricular systolic pressure severely elevated 70-80 mmHg | 0
    evidence of right ventricular overload | 0
    empiric vancomycin started | 0
    piperacillin/tazobactam started | 0
    switched to ampicillin 2 g every 4 hours | 24
    gentamycin 3 mg/kg every 24 hours | 24
    blood cultures growing gram-positive bacilli | 24
    surgical intervention deferred | 24
    acute heart failure | 168
    required emergent intubation | 168
    mechanical ventilation | 168
    ampicillin switched to ampicillin/sulbactam 3 g every 6 hours | 168
    daptomycin 6 mg/kg | 168
    sudden onset septic embolization to left lower limb | 168
    critical ischemia | 168
    new splenic infarcts | 168
    left lower extremity thrombectomy | 168
    four-compartment fasciotomy | 168
    blood cultures continued to show no definitive pathogen | 168
    surgical replacement of mitral valve | 168
    surgical replacement of aortic valve | 168
    intraoperative transesophageal echocardiogram showed enlarged left atrium 5.7 cm | 168
    thrombi present in left atrial appendage | 168
    thrombi present in right atrial appendage | 168
    aortic valve thinned | 168
    severe aortic insufficiency | 168
    posterior leaflet eroded by vegetation | 168
    micro-abscesses in posterior annulus | 168
    nodular extension up the endocardium into left atrium | 168
    pulmonary artery pressures elevated | 168
    inhaled epoprostenol initiated | 168
    good effect from epoprostenol | 168
    weaned slowly | 168
    postoperative course uncomplicated | 336
    blood culture pathogen identification showed Abiotrophia defectiva | 336
    gram-positive bacilli (cereus/thuringiensis, magaterium, subtilis) | 336
    discharged from intensive care unit | 672
    broad spectrum antibiotics for 6 weeks | 672