21 years old | 0
female | 0
primigravida | 0
admitted to the hospital | 0
asthma | -672
depression | -672
anxiety | -672
presented to an outside hospital | -336
suspected streptococcal pharyngitis | -336
discharged on oral Amoxicillin | -336
completed Amoxicillin | -288
presented to the emergency department | -168
discharged home | -168
broke out in a rash | -84
presented to an OSH ED | -84
fever | -84
sore throat | -84
body aches | -84
dry cough | -84
rash | -84
initial vital signs | -84
physical exam | -84
labs | -84
peripheral blood smear | -84
CXR on admission | -84
given intravenous fluids | -84
IV antibiotics | -84
infectious workup | -84
met 3/4 Systemic Inflammatory Response Syndrome criteria | -72
transferred to our facility | -72
bronchoscopy | -72
CT thorax | -72
multifocal pneumonia | -72
high-flow nasal cannula | -72
antibiotic regimen | -72
oral acyclovir | -72
IV acyclovir | -72
persistent fevers | -48
tachycardia | -48
tachypnea | -48
dyspneic | -24
hypoxic | -24
repeat CXR | -24
bilateral pleural effusions | -24
CT chest with contrast | -24
bilateral airspace disease | -24
immunological workup | -24
positive Coombs test | -24
elevated LDH | -24
ANA positive | -24
anti-RNP | -24
anti-Smith | -24
complement C3 | -24
complement C4 | -24
skin biopsy | -24
interface dermatitis | -24
vacuolar with atrophic epidermis | -24
subtle foci of vascular damage | -24
leukocytoclastic vasculitis | -24
BAL confirmed suspicion of alveolar hemorrhage | -24
Candida albicans | -24
respiratory viral and bacterial panel | -24
treated with cyclophosphamide | 0
IV methylprednisolone | 0
plasmapheresis | 0
cyclophosphamide | 0
high fever | 24
hypotension | 24
tachycardia | 24
candidemia | 24
ophthalmology evaluation | 24
bilateral cotton wool spots | 24
retinopathy | 24
extubated | 48
cyclophosphamide IV | 48
acute abdominal pain | 72
lipase | 72
amylase | 72
alkaline phosphatase | 72
total protein | 72
total bilirubin | 72
albumin | 72
CT chest, abdomen, pelvis | 72
acute pancreatitis | 72
discharged | 240
hydroxychloroquine | 240
prednisone taper | 240
preterm premature rupture of membranes | 336
spontaneous labor | 336
magnesium sulfate | 336
vaginal delivery | 336
healthy baby | 336