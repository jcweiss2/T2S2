21 years old | 0
male | 0
admitted to the hospital | 0
Prader-Willi syndrome (PWS) | -40320
birth weight of 3.3 kg | -174240
bilateral undescended testicles | -174240
obesity at age 4 | -146496
hyperphagia at age 5 | -144168
diagnosed with PWS | -113040
recombinant growth hormone (rGH) treatment | -113040
methylphenidate treatment | -113040
tonsillectomy | -113040
gonadotropin-releasing hormone deficiency | -51840
growth hormone deficiency | -51840
diagnosed with DM | -51840
stopped rGH therapy | -51840
metformin treatment | -51840
body mass index (BMI) 50.87 kg/m² | -51840
glipizide treatment | -24960
long-acting insulin (glargine) treatment | -24960
advised positive pressure ventilation | -24960
poor compliance | -24960
normal ventricle size | -24960
normal systolic function | -24960
dyspnea | 0
loss of consciousness | 0
BMI 69.04 kg/m² | 0
blood pressure 96/25 mmHg | 0
body temperature 39°C | 0
heart rate 93 beats per minute | 0
respiratory rate 28 per minute | 0
oxygen saturation 63% | 0
weight gain of 40 kg in one week | -168
oliguria (<100 mL/day) | 0
abdominal distension | 0
periorbicular cyanosis | 0
respiratory distress | 0
skin ulcers | 0
macular rash | 0
cardiomegaly | 0
haziness in the right lung | 0
arterial blood gas pH 6.9 | 0
PCO2 147 | 0
PO2 72.1 | 0
HCO3 29.3 | 0
admitted to the ICU | 0
intubation | 0
SIMV | 0
hemoglobin 15 g/dL | 0
white blood cell 19,620/μL | 0
erythrocyte sedimentation rate 49 mm/hr | 0
C-reactive protein 2.37 mg/dL | 0
lactic acid 10.37 mmol/L | 0
albumin 3.8 g/dL | 0
AST 51 U/L | 0
ALT 59 U/L | 0
BUN 34.9 mg/dL | 0
creatinine 0.93 mg/dL | 0
fasting glucose 141 mg/dL | 0
HbA1c 8.2% | 0
TSH 2.576 uIU/mL | 0
free T4 1.01 ng/dL | 0
Troponin I 0.844 ng/mL | 0
CK-MB 3.73 ng/mL | 0
proBNP 1,904 pg/mL | 0
bilateral pleural effusion | 0
peribronchial opacity | 0
normal saline infusion | 0
noradrenalin infusion | 0
cefotaxime treatment | 0
midazolam treatment | 0
fentanyl treatment | 0
physiotherapy | 0
negative respiratory virus tests | 0
dilated RV cavity | 0
decreased RV systolic function | 0
pulmonary hypertension (RV pressure 52 mmHg) | 0
RHF | 0
cor pulmonale diagnosis | 0
furosemide infusion (3 mg/hr) | 0
negative I/O balance (-1,000–1,500 mL/day) | 0
caloric restriction (1,500 kcal/day) | 0
ICU bed with pressure-relieving mattress | 0
positioning changes every 2 hours | 0
clindamycin treatment | 0
wound dressing | 0
total parenteral nutrition | 168
ventilator mode changed to PC SIMV | 168
weight loss of 5.8 kg | 168
adjusted I/O balance (-1,500–2,000 mL/day) | 168
weight loss of 1.8 kg/day | 168
improved lung congestion | 168
enteral nutrition started | 336
enteral feeding increased to 1,500 mL/day | 672
fluids and electrolytes correction | 672
weight 150.6 kg (-35.1 kg) | 672
extubation | 672
high flow oxygen (50 L/min) | 672
FiO2 0.4 | 672
decreased high flow to 20 L/min | 672
BiPAP during sleep | 840
rehabilitation training | 840
skin ulcers healed | 840
transferred to general ward | 864
weight 133 kg (-52.7 kg) | 864
oral feeding (1,000 kcal/day) | 1008
discharged | 1176
weight at discharge 131.4 kg (-54.3 kg) | 1176
furosemide 0.3 mg/kg/day | 1176
spironolactone 0.19 mg/kg/day | 1176
metformin 15.2 mg/kg/day | 1176
insulin 0.83 IU/kg/day | 1176
outpatient clinic visits every 3 months | 1176
HbA1c maintained at 8%–9% | 1176
continuing BiPAP during sleep | 1176
no congestive hepatopathy | 1176
no proBNP elevation | 1176
