50 years old | 0
male | 0
fatigue | 0
mild splenomegaly | 0
pancytopenia | 0
poor reticulocyte response | 0
splenic marginal zone lymphoma | 0
splenic involvement | 0
bone marrow involvement | 0
remission after 6 cycles of chemo-immunotherapy | 0
relapse after 1 year | -8760
pancytopenia (relapse) | -8760
splenic involvement (relapse) | -8760
bone marrow involvement (relapse) | -8760
partial remission after second line chemo-immunotherapy | 0
surveyed for 2 years | 0
supportive treatment with intravenous immunoglobuline | 0
hypogammaglobulinemia | 0
second relapse | -14448
third line chemo-immunotherapy | -14448
hospitalized with febrile neutropenia | -14448
pneumonia | -14448
bilateral ground-glass areas on thorax CT | -14448
admitted to chest diseases clinic | -14448
broad-spectrum antibiotherapy | -14448
discharged on February 7, 2020 | 0
partial clinical response | 0
laboratory response | 0
radiological regression | 0
admitted to emergency room with respiratory symptoms | 0
thoracic CT findings compatible with COVID-19 | 0
PCR positive for COVID-19 | 0
serum Na: 129 mmol/L | 0
CRP: 3.76 mg/dL | 0
D-dimer: 17.1 mg/L | 0
albumin: 3.4 g/dL | 0
sputum culture negative | 0
blood culture negative | 0
urine culture negative | 0
hydroxychloroquine treatment | 0
oseltamivir treatment | 0
favipiravir treatment | 0
immune plasma therapy | 0
broad spectrum antibiotic treatments | 0
clinical condition partially improved | 0
PCR positivity continued for 2 months | 1440
hospitalized for 64 days | 1536
negative PCR result on day 60 | 1440
discharged from hospital | 1536
admitted to emergency room again with respiratory complaints and fever | 1536
consolidation on thoracic CT | 1536
ground-glass density on thoracic CT | 1536
PCR positive for COVID-19 (July 2020) | 1536
serum Na: 135 mmol/L | 1536
CRP: 12.7 mg/dL | 1536
D-Dimer: 0.64 mg/L | 1536
albumin: 3.2 g/dL | 1536
Klebsiella pneumoniae in sputum culture | 1536
broad spectrum antibiotic treatments (July 2020) | 1536
immune plasma therapy (July 2020) | 1536
PCR negative after 5 days | 1536
radiological regression | 1536
discharged on 16th day | 1536
continued IVIG treatment in pandemic ward | 1536
admitted to emergency room again with diarrhea and general condition disorder | 3840
bilateral ground-glass areas on CT (August 2020) | 3840
PCR positive for COVID-19 (August 2020) | 3840
serum Na: 130 mmol/L | 3840
CRP: 7.59 mg/dL | 3840
D-dimer: 0.52 mg/L | 3840
albumin: 2.3 g/dL | 3840
sputum culture negative (August 2020) | 3840
blood culture negative (August 2020) | 3840
urine culture negative (August 2020) | 3840
metronidazole treatment | 3840
favipiravir treatment (August 2020) | 3840
prednol 40 mg IV | 3840
continued IVIG treatment | 3840
diarrhea continued | 3840
COVID-19 PCR positive in stool | 3840
high fever (38.5°C) | 3840
lobar pneumonia on chest radiograph | 3840
septic condition | 3840
admitted to intensive care unit | 3840
supportive treatments in ICU | 3840
death | 4272
hypogammaglobulinemia (ongoing) | 0
Non-Hodgkin lymphoma | 0
immune plasma therapy (third hospitalization) | 3840
intermittent PCR negative periods | varies
total PCR positivity duration: 110 days | 2640
longest viral shedding reported | 2640
chronic COVID-19 consideration | 2640
negative PCR after immune plasma (July 2020) | 1536
positive PCR after negative result (July 2020) | 3840
isolation since April 12 | 0
no viral culture performed | 0
possible chronic COVID-19 in immunosuppressed | 2640
