35 years old | 0
female | 0
gravida 3 | 0
para 0 | 0
infertility | -672
adenomyosis | -672
IVF | -672
amnion cavity acrinol-induced labor | -1344
gonadotropin-releasing hormone agonist | -672
control ovulation stimulation | -642
HP-HMG | -642
oocyte retrieval | -630
embryo transfer | -627
vaginal administration progesterone | -627
triplet pregnancy | -597
monozygotic twin | -597
singleton | -597
ultrasound-guided selective pregnancy reduction | -592
fetal nuchal translucency | -483
abnormal forearms and wrist joints | -483
single umbilical artery | -483
hospitalized | -364
genetic testing | -364
artificial abortion | -364
umbilical cord blood sampling | -363
labor induction | -363
fever | -48
right upper quadrant tenderness | -48
antibiotic administration | -48
carboprost administration | -48
postpartum hemorrhage | -24
hypotension | -24
septic shock | -24
DIC | -24
hemorrhagic shock | -24
total abdominal hysterectomy | 0
endometritis | 0
uterus cellulitis | 0
antibiotic administration | 0
abdominal debridement | 24
suturing | 24
discharged | 384
Escherichia coli infection | -24
vaginal discharge sample culture | -24
uterine discharge sample culture | 0