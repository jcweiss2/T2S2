54 years old | 0
female | 0
Roux-en-Y procedure | -7920
exploratory laparotomy | -72
altered mental status | -72
confusion | -72
hallucinations | -72
chest pain | -72
blood pressure 119/78 mmHg | 0
pulse 85 beats per minute | 0
temperature 97.8 F° | 0
respiratory rate 18/minute | 0
SpO2 84% | 0
Glasgow Coma Scale 13/15 | 0
bilateral coarse crackles | 0
expiratory wheezes | 0
regular rate and rhythm | 0
normal S1 and S2 | 0
no murmurs or gallops | 0
normal sinus rhythm | 0
no ST or T wave changes | 0
present bowel sounds | 0
mild diffuse tenderness | 0
abdominal wound healing well | 0
white blood cell count 11.8×10^3/mm^3 | 0
total bilirubin 3.2 mg/dL | 0
AST 131 U/L | 0
ALT 178 U/L | 0
ALK phosphate 339 IU/L | 0
urinalysis negative for infections | 0
urine drug screen positive for opiates | 0
urine drug screen positive for benzodiazepines | 0
arterial blood gas pH 7.37 | 0
arterial blood gas PCO2 40.7 | 0
arterial blood gas PO2 56 | 0
arterial blood gas HCO3 23.3 | 0
multi-lobar pneumonia | 0
right fronto-parietal infarct | 0
left cerebellar infarct | 0
BiPAP | 0
blood cultures drawn | 0
IV antibiotics started | 0
Vancomycin | 0
Cefepime | 0
Metronidazole | 0
transferred to critical care unit | 0
severe acute hypoxic respiratory failure | 24
intubated | 24
trans-esophageal echocardiogram | 24
prominent Eustachian valve | 24
multiple vegetations | 24
diffuse hypokinesia | 24
left ventricle ejection fraction 30% | 24
patent foramen ovale | 24
blood cultures revealed Staphylococcus capitis | 24
bronchoalveolar lavage culture revealed Methicillin Resistant Staphylococcus Aureus | 24
extubated | 72
mental status improved | 72
left facial droop | 72
left upper extremity weakness | 72
repeat transthoracic echocardiogram | 168
ejection fraction 45-50% | 168
normal Eustachian valve | 168
repeat blood cultures negative | 96
discharged to skilled nursing facility | 336
IV Vancomycin | 336
IV Cefepime | 336
follow-up exam | 1008
transthoracic echocardiogram | 1008
prominent Eustachian valve | 1008
no vegetation | 1008
ejection fraction 55% | 1008