52 years old | 0
female | 0
bipolar disorder | -8760
lithium treatment | -8760
risperidone treatment | -8760
dry cough | -168
sweats | -168
feeling feverish | -168
upper respiratory tract infection | -168
diagnosis of upper respiratory tract infection | -168
treatment for upper respiratory tract infection | -168
admitted to hospital | 0
delirium | 0
pain in upper right abdominal quadrant | 0
fever | 0
tachycardia | 0
irregular heart rhythm | 0
blood pressure 149/87 mm Hg | 0
tenderness of upper right abdominal quadrant | 0
normal white blood cell count | 0
elevated CRP | 0
hyponatraemia | 0
corrected calcium | 0
potassium level | 0
acute kidney injury | 0
urine culture positive for Escherichia coli | 0
elevated serum lithium concentration | 0
atrial fibrillation | 0
wide QRS complex | 0
ST-segment elevation | 0
previous ECG showed sinus rhythm | -2592
previous ECG showed narrow QRS | -2592
abdominal CT scan | 0
diagnosis of pyelonephritis | 0
discharged | 168
lithium suspended | 0
normal saline infusion | 0
empirical intravenous ceftriaxone | 0
switched to oral ciprofloxacin | 48
blood cultures remained sterile | 48
rapid clinical improvement | 24
heart-rate at 100-110 bpm | 24
no rate or rhythm control for AF | 24
spontaneous cardioversion of AF | 24
ECG showed sinus rhythm | 48
ECG showed first-degree atrioventricular block | 48
ECG showed narrow QRS | 48
ST-segment elevation | 48
reduced lithium posology | 168
discharged | 168
follow-up visit | 4320
lithium level in therapeutic range | 4320
ECG showed Brugada type 1 pattern | 4320
lithium withdrawal | 4320
valproic acid replacement | 4320
ECG showed no Brugada pattern | 4752
genetic testing for SCN5A mutation | 4752
brother's baseline ECG | 4752
brother's ajmaline provocation test | 4752
brother's genetic testing | 4752
SCN5A mutation | 4752
no implantable cardioverter-defibrillator | 4752
clinical follow-up | 4752