57 years old | 0
female | 0
visited the trauma and emergency department | 0
falling on the same level | -24
sudden onset of weakness | -72
nausea | -72
vomiting | -72
diarrhea | -72
known smoker | 0
obese | 0
uncontrolled hypothyroidism | 0
leukocytosis | 0
lymphopenia | 0
thrombocytopenia | 0
deteriorated renal function | 0
hyperglycemic hyperosmolar nonketotic state | 0
blood urea elevated | 0
serum creatinine elevated | 0
glycosuria | 0
pyuria | 0
blood glucose elevated | 0
glycated hemoglobin elevated | 0
hyperglycemic hyperosmolar non-ketotic state | 0
arterial blood gases normal pH | 0
serum osmolarity elevated | 0
CRP elevated | 0
PCT elevated | 0
afebrile | 0
vital signs stable | 0
intravenous hydration | 0
insulin infusion pump | 0
sedated | 12
intubated | 12
deterioration of medical condition | 12
ceftriaxone | 12
clindamycin | 12
abdominal and pelvic CT scan | 12
gas within left kidney | 12
infiltration of septa in perirenal space | 12
intraosseous gas in L3 and L4 | 12
emphysema in epidural space | 12
emphysematous pyelonephritis | 12
emphysematous osteomyelitis of the spine | 12
Klebsiella pneumoniae in urine culture | 12
meropenem | 12
septic shock | 48
multiple organ dysfunction | 48
died | 48
