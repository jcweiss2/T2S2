71 years old | 0
male | 0
new-onset atrial fibrillation | -20160
hospital admission for atrial fibrillation catheter ablation | -20160
ostium secundum atrial septal defect | -20160
mitral regurgitation | -20160
atrial fibrillation catheter ablation (radiofrequency) | -20160
transcatheter ostium secundum atrial septal defect repair | -20160
hospital admission for atrial fibrillation recurrence | -20160
left atrial mass related to the atrial septal defect closure device | -20160
anticoagulant optimization: apixaban to acenocoumarol | -20160
persistent left atrial mass | -20160
surgical removal of the mass | -20160
conclusive diagnosis of left atrial myxoma | -20160
last follow-up | -20160
patient clinically stable | -20160
permanent atrial fibrillation | -20160
good echocardiographic surgical result | -20160
admitted for pulmonary vein ablation | 0
no chronic disease | 0
no past medical history | 0
transoesophageal echocardiography (TEE) showed osASD | 0
significant left-to-right shunt | 0
coronary angiography excluded significant disease | 0
underwent AF ablation | 0
osASD transcatheter closure | 0
discharged on apixaban | 0
hospitalized after AF recurrence | 0
undergo external electrical cardioversion | 0
physical examination unremarkable | 0
completely asymptomatic | 0
transthoracic echocardiography revealed LA mass | 0
moderate mitral regurgitation | 0
device-related thrombus hypothesized | 0
apixaban replaced with acenocoumarol | 0
TEE showed mass size unchanged | 0
mass attached to infero-posterior margin of left disc | 0
isoechoic aspect with irregular margins | 0
extreme mobility | 0
severe mitral regurgitation | 0
cardiovascular MRI showed T1 isointensity | 0
T1 fat-saturated isointensity | 0
heterogeneous T2 hyperintensity | 0
absent first-pass perfusion enhancement | 0
late contrast enhancement sequences difficult to assess | 0
coronary angiography showed neovascularization | 0
case discussed in multidisciplinary heart team | 0
cardiac surgery indicated | 0
LA mass had myxoid appearance | 0
attached between closure device discs | 0
en bloc resection of mass and closure device | 0
LA septum reconstructed using pericardial patch | 0
mitral valve replaced with bioprosthesis | 0
severe regurgitation due to bileaflet prolapse | 0
mass had gelatinous, friable surface | 0
irregular edges | 0
histopathological diagnosis of myxoma | 0
protracted time in intensive care unit | 0
pneumonia | 0
septic shock | 0
acute kidney injury | 0
discharged to inpatient rehabilitation facility | 0
1-year follow-up asymptomatic | 0
permanent AF | 0
TTE shows good surgical result | 0
no tumor recurrence | 0
