66 years old | 0
male | 0
admitted to the emergency department | 0
dyspnea | 0
chest pain | 0
body temperature of 38.6°C | 0
heart rate of 140 beats/min | 0
blood pressure of 75/36 mm Hg | 0
respiratory rate of 26 breaths/min | 0
oxygen saturation of 92% on room air | 0
respiratory distress | 0
accessory muscle use | 0
erythema over the sternum | 0
pitting edema in both lower extremities | 0
feet that were cool to touch | 0
rapid rate | 0
regular rhythm | 0
soft systolic murmur | 0
jugular venous distension | 0
pulsus paradoxus | 0
tachypnea | 0
clear to auscultation | 0
aortic stenosis | -504
surgical mechanical aortic valve replacement | -504
chronic obstructive pulmonary disease | 0
cirrhosis secondary to alcohol use | 0
hypertension | 0
hyperlipidemia | 0
septic shock from sternal wound infection | 0
endocarditis | 0
cardiogenic shock | 0
postoperative complications | 0
tamponade due to postpericardiotomy syndrome | 0
postsurgical bleed | 0
bacterial or viral pneumonia | 0
acute coronary syndrome | 0
pneumothorax | 0
pulmonary embolism | 0
acute heart failure exacerbation | 0
chronic obstructive pulmonary disease exacerbation | 0
emergency bedside echocardiography | 0
moderate to large pericardial effusion | 0
tamponade physiology | 0
emergent echocardiography-guided pericardiocentesis | 0
access to the pericardial fluid | 0
intrapericardial position confirmed | 0
bright red blood removed | 0
hemopericardium | 0
initial hemodynamic improvement | 0
transthoracic echocardiography | 0
significant decrease in the size of the pericardial effusion | 0
pericardial effusion could not be fully drained | 0
pericardial fluid reaccumulated | 10
pericardial drain left in place | 10
cardiac surgery consulted | 10
fresh frozen plasma administered | 10
vitamin K administered | 10
admitted to the cardiac intensive care unit | 10
vasopressor support initiated | 10
broad-spectrum antibiotics started | 10
blood and pericardial cultures drawn | 10
chest computed tomography without intravenous contrast | 24
mid to lower sternotomy wound dehiscence | 24
fractured sternal wire | 24
puncturing the anterior pericardium | 24
intubated | 24
surgical exploration | 24
laceration of the RV free wall | 24
RV free wall repaired | 24
pericardial effusion caused by bleeding from the RV injury | 24
bleeding stopped | 24
pericardiocentesis | 24
right ventricle re-expanded | 24
bleeding resumed | 24
hypotension | 24
signs of shock | 24
vasopressor support | 24
blood and pericardial cultures positive for Staphylococcus aureus | 48
sternal bone cultures grew S aureus | 48
infectious disease specialty expertise consulted | 48
antibiotic therapy guided | 48
hospital course complicated by ongoing shock | 48
progressive acute kidney and liver injury | 48
multiple vasopressor support | 48
sternal wound debridement | 72
purulent exudate from the sternal wound | 72
transesophageal echocardiography | 168
new small vegetation on the mitral valve | 168
endocarditis | 168
comfort care | 336
passed away | 336
autopsy | 336
RV free wall injury confirmed | 336
infective endocarditis of the mitral valve confirmed | 336