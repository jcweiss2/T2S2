77 years old | 0
male | 0
admitted to the hospital | 0
fall | -72
fever | -72
weakness | -72
COVID-19 | -72
pneumonia | -72
bilateral ground-glass opacities | -72
intubated | 0
transferred to ICU | 0
hypertension | -672
cerebral infarction | -672
favipiravir | 0
tocilizumab | 0
paroxysmal atrial fibrillation | 24
CHADS2 VASC score | 24
HAS-BLED | 24
heparin | 24
ART-123 | 24
anterior chest hematoma | 48
Hb level dropped | 48
multiple hematomas | 48
chest wall hematoma | 48
obturatorius internus muscle hematoma | 48
emergency TAE | 72
angiography | 72
digital subtraction angiography | 72
extravasation | 72
embolization | 72
gelatin sponge | 72
coil | 72
hemostasis | 72
discharged from ICU | 168
follow-up CT | 504
chest hematoma decreased | 504
transferred to another hospital | 504 
bruising of the chest wall subsided | 120 
respiratory condition improved | 120
extubated | 120 
new-onset paroxysmal atrial fibrillation | 24 
activated partial thromboplastin time | 0 
prothrombin time | 0 
D-dimer | 0 
CRP | 0 
white blood cell count | 0 
hemoglobin | 0 
platelet | 0 
blood pressure | 0 
heart rate | 0 
SpO2 | 0 
body temperature | 0 
routine reverse transcription polymerase chain reaction test | 0 
severe acute respiratory syndrome coronavirus 2 infection | 0 
CT showed typical signs of pneumonia | 0 
worsening of respiratory symptoms | -72 
maximum barrier precautions | 72 
vinyl | 72 
negative pressure | 72 
caps | 72 
masks | 72 
eye guards | 72 
sterile gowns | 72 
sterile gloves | 72 
double glove use | 72 
N95 respirator masks | 72 
right common femoral artery | 72 
left axillary artery | 72 
acromial branch of the left thoracoacromial artery | 72 
left lateral thoracic artery | 72 
subclavian artery | 72 
coagulopathy | -72 
cytokines storm | -72 
damage-associated molecular patterns | -72 
cell-death mechanisms | -72 
vascular endothelial damage | -72 
hypercoagulable state | -72 
anti-inflammatory properties | 24 
anti-thrombotic prophylaxis | 24 
therapeutic dose of heparin | 24 
bleeding complications | 48 
informed consent | 0 
publication of clinical details and images | 0 
institutional approval | 0 
conflicts of interest | 0 
anticoagulants | 0 
management of Af and COVID-19 | 0 
potential bleeding complications | 0 
patient harm | 0 
emergency transcatheter embolization | 72 
TAE | 72 
axillary arteries | 72 
multiple hematomas | 48 
massive chest wall hematoma | 48 
obturatorius internus muscle hematoma | 48 
elderly patient | 0 
COVID-19 patient | 0 
severe infection | -72 
bacterial and viral infections | -72 
sepsis-associated coagulopathy | -72 
SAC | -72 
recombinant human soluble thrombomodulin | 24 
rTM | 24 
coagulation disorder | -72 
D-dimer level | -72 
DD | -72 
American Society of Hematology | 24 
ASH | 24 
anti-thrombotic prophylaxis dose | 24 
therapeutic dose | 24 
bleeding complications | 48 
SCARLET trial | 504 
randomized, double-blind, placebo-controlled, multinational, multicenter, parallel-group Phase 3 study | 504 
prothrombin fragments 1.2 | 504 
thrombin-antithrombin complex | 504 
baseline coagulation biomarker levels | 504 
mortality | 504 
Levi et al | 504 
subgroups | 504 
T1/2 | 504 
half-life | 504 
heparin and ART-123 | 24 
elderly COVID-19 patients | 24 
traumatic injury | 24 
potential bleeding complications | 24 
NIH COVID-19 Treatment Guidelines | 504 
mechanical ventilation | 504 
advanced stage of the disease | 504 
benefits | 504 
indication and administration | 24 
ART-123 and heparin | 24 
patient harm | 24 
anticoagulants | 0 
Af and COVID-19 | 0 
monitoring | 0 
bleeding complications | 0 
patient harm | 0 
emergency TAE | 72 
branches of the axial arteries | 72 
massive chest wall hematoma | 48 
obturatorius internus muscle hematoma | 48 
COVID-19 patient | 0 
multiple hematomas | 48 
fall | -72 
heparin | 24 
ART-123 | 24 
elderly patient | 0 
COVID-19 | 0 
severe infection | -72 
coagulopathy | -72 
anticoagulants | 0 
Af | 24 
COVID-19 associated coagulopathy | 24 
hypercoagulable state | -72 
anti-thrombotic prophylaxis | 24 
therapeutic dose of heparin | 24 
bleeding complications | 48 
informed consent | 0 
publication of clinical details and images | 0 
institutional approval | 0 
conflicts of interest | 0 
anticoagulants | 0 
management of Af and COVID-19 | 0 
potential bleeding complications | 0 
patient harm | 0 
emergency transcatheter embolization | 72 
TAE | 72 
axillary arteries | 72 
multiple hematomas | 48 
massive chest wall hematoma | 48 
obturatorius internus muscle hematoma | 48 
elderly patient | 0 
COVID-19 patient | 0 
severe infection | -72 
bacterial and viral infections | -72 
sepsis-associated coagulopathy | -72 
SAC | -72 
recombinant human soluble thrombomodulin | 24 
rTM | 24 
coagulation disorder | -72 
D-dimer level | -72 
DD | -72 
American Society of Hematology | 24 
ASH | 24 
anti-thrombotic prophylaxis dose | 24 
therapeutic dose | 24 
bleeding complications | 48 
SCARLET trial | 504 
randomized, double-blind, placebo-controlled, multinational, multicenter, parallel-group Phase 3 study | 504 
prothrombin fragments 1.2 | 504 
thrombin-antithrombin complex | 504 
baseline coagulation biomarker levels | 504 
mortality | 504 
Levi et al | 504 
subgroups | 504 
T1/2 | 504 
half-life | 504 
heparin and ART-123 | 24 
elderly COVID-19 patients | 24 
traumatic injury | 24 
potential bleeding complications | 24 
NIH COVID-19 Treatment Guidelines | 504 
mechanical ventilation | 504 
advanced stage of the disease | 504 
benefits | 504 
indication and administration | 24 
ART-123 and heparin | 24 
patient harm | 24 
anticoagulants | 0 
Af and COVID-19 | 0 
monitoring | 0 
bleeding complications | 0 
patient harm | 0 
emergency TAE | 72 
branches of the axial arteries | 72 
massive chest wall hematoma | 48 
obturatorius internus muscle hematoma | 48 
COVID-19 patient | 0 
multiple hematomas | 48 
fall | -72 
heparin | 24 
ART-123 | 24 
elderly patient | 0 
COVID-19 | 0 
severe infection | -72 
coagulopathy | -72 
anticoagulants | 0 
Af | 24 
COVID-19 associated coagulopathy | 24 
hypercoagulable state | -72 
anti-thrombotic prophylaxis | 24 
therapeutic dose of heparin | 24 
bleeding complications | 48 
informed consent | 0 
publication of clinical details and images | 0 
institutional approval | 0 
conflicts of interest | 0 
anticoagulants | 0 
management of Af and COVID-19 | 0 
potential bleeding complications | 0 
patient harm | 0 
emergency transcatheter embolization | 72 
TAE | 72 
axillary arteries | 72 
multiple hematomas | 48 
massive chest wall hematoma | 48 
obturatorius internus muscle hematoma | 48 
elderly patient | 0 
COVID-19 patient | 0 
severe infection | -72 
bacterial and viral infections | -72 
sepsis-associated coagulopathy | -72 
SAC | -72 
recombinant human soluble thrombomodulin | 24 
rTM | 24 
coagulation disorder | -72 
D-dimer level | -72 
DD | -72 
American Society of Hematology | 24 
ASH | 24 
anti-thrombotic prophylaxis dose | 24 
therapeutic dose | 24 
bleeding complications | 48 
SCARLET trial | 504 
randomized, double-blind, placebo-controlled, multinational, multicenter, parallel-group Phase 3 study | 504 
prothrombin fragments 1.2 | 504 
thrombin-antithrombin complex | 504 
baseline coagulation biomarker levels | 504 
mortality | 504 
Levi et al | 504 
subgroups | 504 
T1/2 | 504 
half-life | 504 
heparin and ART-123 | 24 
elderly COVID-19 patients | 24 
traumatic injury | 24 
potential bleeding complications | 24 
NIH COVID-19 Treatment Guidelines | 504 
mechanical ventilation | 504 
advanced stage of the disease | 504 
benefits | 504 
indication and administration | 24 
ART-123 and heparin | 24 
patient harm | 24 
anticoagulants | 0 
Af and COVID-19 | 0 
monitoring | 0 
bleeding complications | 0 
patient harm | 0 
emergency TAE | 72 
branches of the axial arteries | 72 
massive chest wall hematoma | 48 
obturatorius internus muscle hematoma | 48 
COVID-19 patient | 0 
multiple hematomas | 48 
fall | -72 
heparin | 24 
ART-123 | 24 
elderly patient | 0 
COVID-19 | 0 
severe infection | -72 
coagulopathy | -72 
anticoagulants | 0 
Af | 24 
COVID-19 associated coagulopathy | 24 
hypercoagulable state | -72 
anti-thrombotic prophylaxis | 24 
therapeutic dose of heparin | 24 
bleeding complications | 48 
informed consent | 0 
publication of clinical details and images | 0 
institutional approval | 0 
conflicts of interest | 0 
anticoagulants | 0 
management of Af and COVID-19 | 0 
potential bleeding complications | 0 
patient harm | 0 
emergency transcatheter embolization | 72 
TAE | 72 
axillary arteries | 72 
multiple hematomas | 48 
massive chest wall hematoma | 48 
obturatorius internus muscle hematoma | 48 
elderly patient | 0 
COVID-19 patient | 0 
severe infection | -72 
bacterial and viral infections | -72 
sepsis-associated coagulopathy | -72 
SAC | -72 
recombinant human soluble thrombomodulin | 24 
rTM | 24 
coagulation disorder | -72 
D-dimer level | -72 
DD | -72 
American Society of Hematology | 24 
ASH | 24 
anti-thrombotic prophylaxis dose | 24 
therapeutic dose | 24 
bleeding complications | 48 
SCARLET trial | 504 
randomized, double-blind, placebo-controlled, multinational, multicenter, parallel-group Phase 3 study | 504 
prothrombin fragments 1.2 | 504 
thrombin-antithrombin complex | 504 
baseline coagulation biomarker levels | 504 
mortality | 504 
Levi et al | 504 
subgroups | 504 
T1/2 | 504 
half-life | 504 
heparin and ART-123 | 24 
elderly COVID-19 patients | 24 
traumatic injury | 24 
potential bleeding complications | 24 
NIH COVID-19 Treatment Guidelines | 504 
mechanical ventilation | 504 
advanced stage of the disease | 504 
benefits | 504 
indication and administration | 24 
ART-123 and heparin | 24 
patient harm | 24 
anticoagulants | 0 
Af and COVID-19 | 0 
monitoring | 0 
bleeding complications | 0 
patient harm | 0 
emergency TAE | 72 
branches of the axial arteries | 72 
massive chest wall hematoma | 48 
obturatorius internus muscle hematoma | 48 
COVID-19 patient | 0 
multiple hematomas | 48 
fall | -72 
heparin | 24 
ART-123 | 24 
elderly patient | 0 
COVID-19 | 0 
severe infection | -72 
coagulopathy | -72 
anticoagulants | 0 
Af | 24 
COVID-19 associated coagulopathy | 24 
hypercoagulable state | -72 
anti-thrombotic prophylaxis | 24 
therapeutic dose of heparin | 24 
bleeding complications | 48 
informed consent | 0 
publication of clinical details and images | 0 
institutional approval | 0 
conflicts of interest | 0 
anticoagulants | 0 
management of Af and COVID-19 | 0 
potential bleeding complications | 0 
patient harm | 0 
emergency transcatheter embolization | 72 
TAE | 72 
axillary arteries | 72 
multiple hematomas | 48 
massive chest wall hematoma | 48 
obturatorius internus muscle hematoma | 48 
elderly patient | 0 
COVID-19 patient | 0 
severe infection | -72 
bacterial and viral infections | -72 
sepsis-associated coagulopathy | -72 
SAC | -72 
recombinant human soluble thrombomodulin | 24 
rTM | 24 
coagulation disorder | -72 
D-dimer level | -72 
DD | -72 
American Society of Hematology | 24 
ASH | 24 
anti-thrombotic prophylaxis dose | 24 
therapeutic dose | 24 
bleeding complications | 48 
SCARLET trial | 504 
randomized, double-blind, placebo-controlled, multinational, multicenter, parallel-group Phase 3 study | 504 
prothrombin fragments 1.2 | 504 
thrombin-antithrombin complex | 504 
baseline coagulation biomarker levels | 504 
mortality | 504 
Levi et al | 504 
subgroups | 504 
T1/2 | 504 
half-life | 504 
heparin and ART-123 | 24 
elderly COVID-19 patients | 24 
traumatic injury | 24 
potential bleeding complications | 24 
NIH COVID-19 Treatment Guidelines | 504 
mechanical ventilation | 504 
advanced stage of the disease | 504 
benefits | 504 
indication and administration | 24 
ART-123 and heparin | 24 
patient harm | 24 
anticoagulants | 0 
Af and COVID-19 | 0 
monitoring | 0 
bleeding complications | 0 
patient harm | 0 
emergency TAE | 72 
branches of the axial arteries | 72 
massive chest wall hematoma | 48 
obturatorius internus muscle hematoma | 48 
COVID-19 patient | 0 
multiple hematomas | 48 
fall | -72 
heparin | 24 
ART-123 | 24 
elderly patient | 0 
COVID-19 | 0 
severe infection | -72 
coagulopathy | -72 
anticoagulants | 0 
Af | 24 
COVID-19 associated coagulopathy | 24 
hypercoagulable state | -72 
anti-thrombotic prophylaxis | 24 
therapeutic dose of heparin | 24 
bleeding complications | 48 
informed consent | 0 
publication of clinical details and images | 0 
institutional approval | 0 
conflicts of interest | 0 
anticoagulants | 0 
management of Af and COVID-19 | 0 
potential bleeding complications | 0 
patient harm | 0 
emergency transcatheter embolization | 72 
TAE | 72 
axillary arteries | 72 
multiple hematomas | 48 
massive chest wall hematoma | 48 
obturatorius internus muscle hematoma | 48 
elderly patient | 0 
COVID-19 patient | 0 
severe infection | -72 
bacterial and viral infections | -72 
sepsis-associated coagulopathy | -72 
SAC | -72 
recombinant human soluble thrombomodulin | 24 
rTM | 24 
coagulation disorder | -72 
D-dimer level | -72 
DD | -72 
American Society of Hematology | 24 
ASH | 24 
anti-thrombotic prophylaxis dose | 24 
therapeutic dose | 24 
bleeding complications | 48 
SCARLET trial | 504 
randomized, double-blind, placebo-controlled, multinational, multicenter, parallel-group Phase 3 study | 504 
prothrombin fragments 1.2 | 504 
thrombin-antithrombin complex | 504 
baseline coagulation biomarker levels | 504 
mortality | 504 
Levi et al | 504 
subgroups | 504 
T1/2 | 504 
half-life | 504 
heparin and ART-123 | 24 
elderly COVID-19 patients | 24 
traumatic injury | 24 
potential bleeding complications | 24 
NIH COVID-19 Treatment Guidelines | 504 
mechanical ventilation | 504 
advanced stage of the disease | 504 
benefits | 504 
indication and administration | 24 
ART-123 and heparin | 24 
patient harm | 24 
anticoagulants | 0 
Af and COVID-19 | 0 
monitoring | 0 
bleeding complications | 0 
patient harm | 0 
emergency TAE | 72 
branches of the axial arteries | 72 
massive chest wall hematoma | 48 
obturatorius internus muscle hematoma | 48 
COVID-19 patient | 0 
multiple hematomas | 48 
fall | -72 
heparin | 24 
ART-123 | 24 
elderly patient | 0 
COVID-19 | 0 
severe infection | -72 
coagulopathy | -72 
anticoagulants | 0 
Af | 24 
COVID-19 associated coagulopathy | 24 
hypercoagulable state | -72 
anti-thrombotic prophylaxis | 24 
therapeutic dose of heparin | 24 
bleeding complications | 48 
informed consent | 0 
publication of clinical details and images | 0 
institutional approval | 0 
conflicts of interest | 0 
anticoagulants | 0 
management of Af and COVID-19 | 0 
potential bleeding complications | 0 
patient harm | 0 
emergency transcatheter embolization | 72 
TAE | 72 
axillary arteries | 72 
multiple hematomas | 48 
massive chest wall hematoma | 48 
obturatorius internus muscle hematoma | 48 
elderly patient | 0 
COVID-19 patient | 0 
severe infection | -72 
bacterial and viral infections | -72 
sepsis-associated coagulopathy | -72 
SAC | -72 
recombinant human soluble thrombomodulin | 24 
rTM | 24 
coagulation disorder | -72 
D-dimer level | -72 
DD | -72 
American Society of Hematology | 24 
ASH | 24 
anti-thrombotic prophylaxis dose | 24 
therapeutic dose | 24 
bleeding complications | 48 
SCARLET trial | 504 
randomized, double-blind, placebo-controlled, multinational, multicenter, parallel-group Phase 3 study | 504 
prothrombin fragments 1.2 | 504 
thrombin-antithrombin complex | 504 
baseline coagulation biomarker levels | 504 
mortality | 504 
Levi et al | 504 
subgroups | 504 
T1/2 | 504 
half-life | 504 
heparin and ART-123 | 24 
elderly COVID-19 patients | 24 
traumatic injury | 24 
potential bleeding complications | 24 
NIH COVID-19 Treatment Guidelines | 504 
mechanical ventilation | 504 
advanced stage of the disease | 504 
benefits | 504 
indication and administration | 24 
ART-123 and heparin | 24 
patient harm | 24 
anticoagulants | 0 
Af and COVID-19 | 0 
monitoring | 0 
bleeding complications | 0 
patient harm | 0 
emergency TAE | 72 
branches of the axial arteries | 72 
massive chest wall hematoma | 48 
obturatorius internus muscle hematoma | 48 
COVID-19 patient | 0 
multiple hematomas | 48 
fall | -72 
heparin | 24 
ART-123 | 24 
elderly patient | 0 
COVID-19 | 0 
severe infection | -72 
coagulopathy | -72 
anticoagulants | 0 
Af | 24 
COVID-19 associated coagulopathy | 24 
hypercoagulable state | -72 
anti-thrombotic prophylaxis | 24 
therapeutic dose of heparin | 24 
bleeding complications | 48 
informed consent | 0 
publication of clinical details and images | 0 
institutional approval | 0 
conflicts of interest | 0 
anticoagulants | 0 
management of Af and COVID-19 | 0 
potential bleeding complications | 0 
patient harm | 0 
emergency transcatheter embolization | 72 
TAE | 72 
axillary arteries | 72 
multiple hematomas | 48 
massive chest wall hematoma | 48 
obturatorius internus muscle hematoma | 48 
elderly patient | 0 
COVID-19 patient | 0 
severe infection | -72 
bacterial and viral infections | -72 
sepsis-associated coagulopathy | -72 
SAC | -72 
recombinant human soluble thrombomodulin | 24 
rTM | 24 
coagulation disorder | -72 
D-dimer level | -72 
DD | -72 
American Society of Hematology | 24 
ASH | 24 
anti-thrombotic prophylaxis dose | 24 
therapeutic dose | 24 
bleeding complications | 48 
SCARLET trial | 504 
randomized, double-blind, placebo-controlled, multinational, multicenter, parallel-group Phase 3 study | 504 
prothrombin fragments 1.2 | 504 
thrombin-antithrombin complex | 504 
baseline coagulation biomarker levels | 504 
mortality | 504 
Levi et al | 504 
subgroups | 504 
T1/2 | 504 
half-life | 504 
heparin and ART-123 | 24 
elderly COVID-19 patients | 24 
traumatic injury | 24 
potential bleeding complications | 24 
NIH COVID-19 Treatment Guidelines | 504 
mechanical ventilation | 504 
advanced stage of the disease | 504 
benefits | 504 
indication and administration | 24 
ART-123 and heparin | 24 
patient harm | 24 
anticoagulants | 0 
Af and COVID-19 | 0 
monitoring | 0 
bleeding complications | 0 
patient harm | 0 
emergency TAE | 72 
branches of the axial arteries | 72 
massive chest wall hematoma | 48 
obturatorius internus muscle hematoma | 48 
COVID-19 patient | 0 
multiple hematomas | 48 
fall | -72 
heparin | 24 
ART-123 | 24 
elderly patient | 0 
COVID-19 | 0 
severe infection | -72 
coagulopathy | -72 
anticoagulants | 0 
Af | 24 
COVID-19 associated coagulopathy | 24 
hypercoagulable state | -72 
anti-thrombotic prophylaxis | 24 
therapeutic dose of heparin | 24 
bleeding complications | 48 
informed consent | 0 
publication of clinical details and images | 0 
institutional approval | 0 
conflicts of interest | 0 
anticoagulants | 0 
management of Af and COVID-19 | 0 
potential bleeding complications | 0 
patient harm | 0 
emergency transcatheter embolization | 72 
TAE | 72 
axillary arteries | 72 
multiple hematomas | 48 
massive chest wall hematoma | 48 
obturatorius internus muscle hematoma | 48 
elderly patient | 0 
COVID-19 patient | 0 
severe infection | -72 
bacterial and viral infections | -72 
sepsis-associated coagulopathy | -72 
SAC | -72 
recombinant human soluble thrombomodulin | 24 
rTM | 24 
coagulation disorder | -72 
D-dimer level | -72 
DD | -72 
American Society of Hematology | 24 
ASH | 24 
anti-thrombotic prophylaxis dose | 24 
therapeutic dose | 24 
bleeding complications | 48 
SCARLET trial | 504 
randomized, double-blind, placebo-controlled, multinational, multicenter, parallel-group Phase 3 study | 504 
prothrombin fragments 1.2 | 504 
thrombin-antithrombin complex | 504 
baseline coagulation biomarker levels | 504 
mortality | 504 
Levi et al | 504 
subgroups | 504 
T1/2 | 504 
half-life | 504 
heparin and ART-123 | 24 
elderly COVID-19 patients | 24 
traumatic injury | 24 
potential bleeding complications | 24 
NIH COVID-19 Treatment Guidelines | 504 
mechanical ventilation | 504 
advanced stage of the disease | 504 
benefits | 504 
indication and administration | 24 
ART-123 and heparin | 24 
patient harm | 24 
anticoagulants | 0 
Af and COVID-19 | 0 
monitoring | 0 
bleeding complications | 0 
patient harm | 0 
emergency TAE | 72 
branches of the axial arteries | 72 
massive chest wall hematoma | 48 
obturatorius internus muscle hematoma | 48 
COVID-19 patient | 0 
multiple hematomas | 48 
fall | -72 
heparin | 24 
ART-123 | 24 
elderly patient | 0 
COVID-19 | 0 
severe infection | -72 
coagulopathy | -72 
anticoagulants | 0 
Af | 24 
COVID-19 associated coagulopathy | 24 
hypercoagulable state | -72 
anti-thrombotic prophylaxis | 24 
therapeutic dose of heparin | 24 
bleeding complications | 48 
informed consent | 0 
publication of clinical details and images | 0 
institutional approval | 0 
conflicts of interest | 0 
anticoagulants | 0 
management of Af and COVID-19 | 0 
potential bleeding complications | 0 
patient harm | 0 
emergency transcatheter embolization | 72 
TAE | 72 
axillary arteries | 72 
multiple hematomas | 48 
massive chest wall hematoma | 48 
obturatorius internus muscle hematoma | 48 
elderly patient | 0 
COVID-19 patient | 0 
severe infection | -72 
bacterial and viral infections | -72 
sepsis-associated coagulopathy | -72 
SAC | -72 
recombinant human soluble thrombomodulin | 24 
rTM | 24 
coagulation disorder | -72 
D-dimer level | -72 
DD | -72 
American Society of Hematology | 24 
ASH | 24 
anti-thrombotic prophylaxis dose | 24 
therapeutic dose | 24 
bleeding complications | 48 
SCARLET trial | 504 
randomized, double-blind, placebo-controlled, multinational, multicenter, parallel-group Phase 3 study | 504 
prothrombin fragments 1.2 | 504 
thrombin-antithrombin complex | 504 
baseline coagulation biomarker levels | 504 
mortality | 504 
Levi et al | 504 
subgroups | 504 
T1/2 | 504 
half-life | 504 
heparin and ART-123 | 24 
elderly COVID-19 patients | 24 
traumatic injury | 24 
potential bleeding complications | 24 
NIH COVID-19 Treatment Guidelines | 504 
mechanical ventilation | 504 
advanced stage of the disease | 504 
benefits | 504 
indication and administration | 24 
ART-123 and heparin | 24 
patient harm | 24 
anticoagulants | 0 
Af and COVID-19 | 0 
monitoring | 0 
bleeding complications | 0 
patient harm | 0 
emergency TAE | 72 
branches of the axial arteries | 72 
massive chest wall hematoma | 48 
obturatorius internus muscle hematoma | 48 
COVID-19 patient | 0 
multiple hematomas | 48 
fall | -72 
heparin | 24 
ART-123 | 24 
elderly patient | 0 
COVID-19 | 0 
severe infection | -72 
coagulopathy | -72 
anticoagulants | 0 
Af | 24 
COVID-19 associated coagulopathy | 24 
hypercoagulable state | -72 
anti-thrombotic prophylaxis | 24 
therapeutic dose of heparin | 24 
bleeding complications | 48 
informed consent | 0 
publication of clinical details and images | 0 
institutional approval | 0 
conflicts of interest | 0 
anticoagulants | 0 
management of Af and COVID-19 | 0 
potential bleeding complications | 0 
patient harm | 0 
emergency transcatheter embolization | 72 
TAE | 72 
axillary arteries | 72 
multiple hematomas | 48 
massive chest wall hematoma | 48 
obturatorius internus muscle hematoma | 48 
elderly patient | 0 
COVID-19 patient | 0 
severe infection | -72 
bacterial and viral infections | -72 
sepsis-associated coagulopathy | -72 
SAC | -72 
recombinant human soluble thrombomodulin | 24 
rTM | 24 
coagulation disorder | -72 
D-dimer level | -72 
DD | -72 
American Society of Hematology | 24 
ASH | 24 
anti-thrombotic prophylaxis dose | 24 
therapeutic dose | 24 
bleeding complications | 48 
SCARLET trial | 504 
randomized, double-blind, placebo-controlled, multinational, multicenter, parallel-group Phase 3 study | 504 
prothrombin fragments 1.2 | 504 
thrombin-antithrombin complex | 504 
baseline coagulation biomarker levels | 504 
mortality | 504 
Levi et al | 504 
subgroups | 504 
T1/2 | 504 
half-life | 504 
heparin and ART-123 | 24 
elderly COVID-19 patients | 24 
traumatic injury | 24 
potential bleeding complications | 24 
NIH COVID-19 Treatment Guidelines | 504 
mechanical ventilation | 504 
advanced stage of the disease | 504 
benefits | 504 
indication and administration | 24 
ART-123 and heparin | 24 
patient harm | 24 
anticoagulants | 0 
Af and COVID-19 | 0 
monitoring | 0 
bleeding complications | 0 
patient harm | 0 
emergency TAE | 72 
branches of the axial arteries | 72 
massive chest wall hematoma | 48 
obturatorius internus muscle hematoma | 48 
COVID-19 patient | 0 
multiple hematomas | 48 
fall | -72 
heparin | 24 
ART-123 | 24 
elderly patient | 0 
COVID-19 | 0 
severe infection | -72 
coagulopathy | -72 
anticoagulants | 0 
Af | 24 
COVID-19 associated coagulopathy | 24 
hypercoagulable state | -72 
anti-thrombotic prophylaxis | 24 
therapeutic dose of heparin | 24 
bleeding complications | 48 
informed consent | 0 
publication of clinical details and images | 0 
institutional approval | 0 
conflicts of interest | 0 
anticoagulants | 0 
management of Af and COVID-19 | 0 
potential bleeding complications | 0 
patient harm | 0 
emergency transcatheter embolization | 72 
TAE | 72 
axillary arteries | 72 
multiple hematomas | 48 
massive chest wall hematoma | 48 
obturatorius internus muscle hematoma | 48 
elderly patient | 0 
COVID-19 patient | 0 
severe infection | -72 
bacterial and viral infections | -72 
sepsis-associated coagulopathy | -72 
SAC | -72 
recombinant human soluble thrombomodulin | 24 
rTM | 24 
coagulation disorder | -72 
D-dimer level | -72 
DD | -72 
American Society of Hematology | 24 
ASH | 24 
anti-thrombot