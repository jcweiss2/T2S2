53 years old | 0
male | 0
admitted to the hospital | 0
subjective fever | -72
chills | -72
diffuse myalgias | -72
productive cough | -72
diagnosed with pneumonia | -24
prescribed Levofloxacin | -24
discharged home | -24
returned to the hospital | 24
dyspnea | 24
nausea | 24
emesis | 24
syncope | 24
tachycardic | 24
normotensive | 24
tachypneic | 24
normal oxygen saturations | 24
temperature of 37.1 degrees Celsius | 24
elevated WBC count | 24
elevated troponin-t | 24
elevated creatine kinase | 24
elevated lactate | 24
sinus tachycardia with frequent PVCs | 24
suspected sepsis | 24
blood cultures drawn | 24
treated with IV fluids | 24
treated with Piperacillin-Tazobactam | 24
transferred to the tertiary care centre | 48
heart rate of 122 beats per minute | 48
blood pressure of 111/88 mmHg | 48
respiratory rate of 25 breaths per minute | 48
oxygen saturation of 99% | 48
temperature of 36.5 degrees Celsius | 48
bilateral pulmonary crackles | 48
normal heart sounds | 48
elevated jugular venous pressure | 48
mottled skin | 48
cool extremities | 48
capillary refill time of six seconds | 48
benign abdominal exam | 48
unremarkable chest radiograph | 48
CT pulmonary angiogram | 48
pulmonary edema | 48
elevated NT-proBNP | 48
consulted to Cardiology | 48
suspected decompensated heart failure | 48
urgent cardiac transthoracic echocardiography | 48
severe global hypokinesis of the left ventricle | 48
ejection fraction of 15-20% | 48
small pericardial effusion | 48
probable myocarditis | 48
treated with Colchicine | 72
treated with high-dose Aspirin | 72
troponin peaked at 3871 ng/L | 96
nasopharyngeal swab completed | 96
sent for influenza antigen testing | 96
started on empiric Oseltamivir | 96
nasopharyngeal swab returned positive for Influenza B | 192
increasing dyspnea | 192
shortness of breath | 192
increased oxygen requirements | 192
new right-sided airspace opacity | 192
Vancomycin added to Piperacillin-Tazobactam | 192
pain to his forearms bilaterally | 192
elevated CK | 192
right forearm increased in sensitivity and became firm | 192
compartment pressure of 60 mmHg | 192
underwent a bedside right forearm fasciotomy | 192
transferred to the Medical-Surgical Intensive Care Unit | 192
intubation | 192
heart rate of 111 beats per minute | 192
blood pressure of 86/57 mmHg | 192
MAP of 67 mmHg | 192
saturating 97% | 192
pressure support of 8 cmH20 | 192
fraction of inspired oxygen of 45% | 192
positive end expiratory pressure of 10 cmH20 | 192
respiratory rate of 19 breaths per minute | 192
temperature of 37.1 degrees Celsius | 192
diffuse bilateral crackles in the lungs | 192
normal heart sounds | 192
elevated jugular venous pressure | 192
3+ pitting edema to his sacrum | 192
mottled skin | 192
cool extremities | 192
Norepinephrine started | 192
Furosemide infusion initiated | 192
Norepinephrine discontinued | 120
repeat TTE demonstrated complete recovery of his ejection fraction | 168
Oseltamivir continued | 168
anaerobic and aerobic blood cultures returned negative for growth | 168
repeat NP PCR test sent for Influenza | 168
repeat NP PCR test returned positive for Influenza B | 240
became oliguric | 240
creatinine of 416 umol/L | 240
underwent continuous renal replacement therapy | 240
recovery of renal function | 288
successfully extubated | 288
transferred to home hospital for rehabilitation | 312
discharged to his place of residence | 384