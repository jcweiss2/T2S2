54 years old | 0
male | 0
type 2 diabetes mellitus | -672
admitted to the hospital | 0
acute abdominal pain | -48
fever | -48
blood pressure 82/45 mm Hg | 0
pulse rate 135/min | 0
abdomen distended | 0
abdomen generally tight | 0
no jaundice | 0
diabetic ketoacidosis | 0
elevated white blood cells | 0
high C-reactive protein | 0
normal liver function tests | 0
abdominal ultrasonography | 0
massive ascites | 0
gases filling the intestines | 0
abdominal computerized tomography scan | 0
free fluid | 0
gallbladder wall thickness increased | 0
resolved gallbladder distention | 0
no pneumoperitoneum | 0
no choledocholithiasis | 0
diagnostic paracentesis | 2
bile leakage | 2
ascites with dark yellow-green color | 2
initial resuscitation | 2
emergent exploratory laparotomy | 4
diffuse biliary peritonitis | 4
peritoneal lavage | 4
no duodenal perforation | 4
no gallbladder perforation | 4
cholecystectomy | 4
intraoperative cholangiography | 4
extravasation from posterior wall of medium portion of choledochus | 4
perforation repaired over T-tube | 4
peritoneal cavity drained with two Salem tubes | 4
postoperative course uneventful | 24
discharged on 15th postoperative day | 360
T-tube removed on 32 postoperative day | 768
normal cholangiogram | 768
no biliary leakage | 768
no pancreaticobiliary junction or distal stricture | 768
pathological examination of cholecystectomy | 768
ulcerous acalculous cholecystitis | 768
follow-up after 3 months | 2160
no recurrence of symptoms | 2160