32 years old | 0
woman | 0
no significant past medical history | 0
referred to a dermatologist | -72
Nicolau syndrome | -72
presented to the emergency department | 0
severe pain | 0
redness | 0
swelling involving left buttock | 0
surrounding back area | 0
intramuscular injection of methocarbamol | -72
symptoms onset | -72
symptoms progressively worsened over three days | -72 to -48
purpose of injection to alleviate musculoskeletal pain | -72
motor vehicle accident | -72
anxious | 0
severe distress | 0
left buttock discolored | 0
dusky appearance | 0
marked erythema | 0
edema | 0
affected area extended from left buttock | 0
involved entire gluteal region | 0
spread to adjacent back area | 0
necrotic tissue | 0
black and eschar-like | 0
hypotension | 0
tachycardia | 0
leukocytosis | 0
left shift | 0
inflammatory response | 0
normal renal function | 0
normal hepatic function | 0
imaging studies ultrasound | 0
computed tomography | 0
massive tissue necrosis | 0
impaired peripheral perfusion | 0
aggressive resuscitation efforts | 0
broad-spectrum antibiotic therapy | 0
condition deteriorated | 24
hemodynamic instability | 24
cardiac shock | 24
death | 144
autopsy | 144
external examination | 144
internal examination | 144
tissue samples collected | 144
histopathological analysis | 144
toxicological analysis | 144
liver mild fatty changes | 144
kidney acute tubular necrosis | 144
acute kidney injury | 144
brain tissue normal | 144
therapeutic levels of metacarbamol | 144
compromised circulation | 0
cardiac shock | 144
