20 years old | 0
female | 0
insulin-dependent diabetes mellitus | -720
pulmonary tuberculosis | -144
productive cough | -720
weight loss | -720
fever | -720
anti-tuberculous medicines | -144
CT scan showing multiple cavitatory lesions in the right lung | 0
sepsis | 0
hypotension | 0
multi-organ failure | 0
diabetic ketoacidosis | 0
insulin infusion | 0
hypoxia | 0
acidosis | 0
pulseless ventricular tachycardia | 0
revived after ACLS protocol | 0
intubated | 0
VATS | 0
evacuation of the abscess | 0
major air leak | 0
oxygen saturation down to 60% | 0
jet ventilation | 0
desaturate again | 0
ruptured lung abscess at the right upper lobe | 0
lung isolation | 0
double lumen tube | 0
tracheal lumen clamped | 0
left lung ventilated differentially |; 0
recruitment maneuver | 0
oxygen saturation rises to 92% | 0
right upper lobe lobectomy | 0
packed red blood cell transfused | 0
phenylephrine boluses | 0
chest drain | 0
endotracheal tube replaced | 0
bronchoscopy | 24
no residual defect | 24
