29 years old | 0
male | 0
admitted to the hospital | 0
muscle pain | -144
joint pain | -144
general weakness | -144
fever | -144
liver dysfunction | -144
elevated total bilirubin | -144
elevated serum glutamic oxaloacetic transaminase | -144
elevated serum glutamic pyruvate transaminase | -144
elevated gamma-glutamyl transferase | -144
elevated lactate dehydrogenase | -144
systemic inflammation | -144
elevated C-reactive protein | -144
elevated procalcitonin | -144
elevated leukocyte levels | -144
acute respiratory failure | 0
altered state of consciousness | 0
intubation | 0
mechanical ventilation | 0
FiO2 100% | 0
SpO2 88.7% | 0
hemodynamic instability | 0
norepinephrine | 0
vasopressin | 0
broad-spectrum empirical antimicrobial therapy | 0
meropenem | 0
azithromycin | 0
oseltamivir | 0
methylprednisolone | 0
stress ulcer prophylaxis | 0
thromboprophylaxis | 0
UFH | 0
continuous sedation | 0
muscle relaxation | 0
prone position | 0
chest CT | 0
massive bilateral pneumonia | 0
minimal pleural effusions | 0
bedside focus ultrasound | 0
acute renal failure | 144
CRRT | 144
CytoSorb | 168
norepinephrine requirements lowered | 168
norepinephrine discontinued | 192
septic episode | 240
second CytoSorb therapy | 240
ICU delirium | 240
antipsychotics | 240
percutaneous tracheostomy | 240
hemodynamic stability | 240
weaned off from ventilator | 240
transferred to general ward | 1152
transferred to rehabilitation clinic | 1200