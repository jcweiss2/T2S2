33 years old | 0
woman | 0
presented with nausea | -24
presented with vomiting | -24
presented with abdominal pain | -24
discharged | -36
hospitalized for recurrent pericarditis | -36
treated with colchicine 0.6 mg twice daily | -36
febrile (temperature 38.6°C) | 0
hypotensive (blood pressure 66/39 mm Hg) | 0
physical examination benign | 0
leukocytosis (51.2 × 10^9/l) | 0
elevated serum lactate (12 mmol/l) | 0
acute kidney injury (serum creatinine 2.0 mg/dl) |;0
acute transaminitis (alanine aminotransferase 2,148 IU/l) | 0
acute transaminitis (aspartate aminotransferase 4,577 IU/l) | 0
severe coagulopathy (international normalized ratio >15) | 0
serum troponin within normal limits | 0
comprehensive toxicology screen negative | 0
electrocardiography normal sinus rhythm without ST-T changes | 0
transthoracic echocardiogram normal biventricular function | 0
transthoracic echocardiogram no valvular disease | 0
transthoracic echocardiogram no pericardial effusion | 0
sepsis from intrabdominal source suspected | 0
fluid resuscitation | 0
started on broad-spectrum antibiotics | 0
administered vasopressor therapy | 0
severe multisystem organ failure developed | 24
intubated | 24
paralyzed | 24
treated with intravascular volume repletion | 24
escalating doses of intravenous vasopressors (epinephrine) | 24
escalating doses of intravenous vasopressors (norepinephrine) | 24
escalating doses of intravenous vasopressors (vasopressin) | 24
broad-spectrum antibiotics | 24
stress-dose steroids | 24
high-dose vitamin B12 for refractory shock | 24
hemodynamics consistent with distributive shock | 24
cardiac output 7.4 l/min | 24
pulmonary artery diastolic pressure 8 mm Hg | 24
systemic vascular resistance indexed 1,572 dynes/s/cm^5/m^2 | 24
hemodynamics changed to cardiogenic shock | 48
pulmonary artery diastolic pressure 24 mm Hg | 48
cardiac output 4.3 l/min | 48
systemic vascular resistance indexed 2,298 dynes/s/cm^5/m^2 | 48
troponin increased to 73.14 ng/ml | 48
electrocardiogram unchanged | 48
transesophageal echocardiogram revealed severe biventricular failure (LVEF 15%) | 48
intravenous milrinone added for inotropic support | 48
started on continuous renal replacement therapy | 48
anuric renal failure | 48
hypotensive despite negative blood culture results | 48
improving leukocytosis | 48
consideration of colchicine toxicity | 48
packed red blood cell transfusion initiated | 48
CO normalized | 72
troponin decreased | 72
multisystem organ failure improved | 72
white blood cell count continued to fall | 96
neutropenic | 96
repeat echocardiogram showed LVEF 50-55% | 144
weaned from vasopressors | 312
off CRRT | 312
extubated | 312
hair loss | 576
admitted to taking 60 tablets of colchicine | 240
elevated serum colchicine level (5.7 ng/ml) | 240
elevated whole blood colchicine level (17 ng/ml) | 240
serum colchicine level 5.3 ng/ml | 264
whole blood colchicine level 7.6 ng/ml | 264
spent 15 days in intensive care unit | 360
discharged after nearly 3-week hospital stay | 504
complete renal recovery | 504
complete hepatic recovery | 504
complete cardiac recovery | 504
outpatient rehabilitation | 504
no further sequelae | 504
