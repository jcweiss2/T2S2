37 years old | 0
male | 0
no significant medical history | 0
no recent international travel | 0
no known contact with anyone with COVID-19 | 0
fever | -72
headache | -72
unilateral, painful neck swelling | -72
transported in an EpiShuttle | 0
admitted to the hospital | 0
area of redness in the posterior palate | 0
tender, non-fluctuant swelling extending from the left mandibular angle towards the sternocleidomastoid muscle | 0
denied any cough | 0
denied neck stiffness | 0
denied pain on swallowing | 0
denied respiratory distress | 0
denied chest pain | 0
febrile at 41°C | 0
tachycardic at 115 beats per minute | 0
normotensive at 119/76 mm Hg | 0
mentally alert | 0
intermittently raised respiratory rate varying between 12 and 22 breaths per minute | 0
peripheral oxygen saturation of 100% on room air | 0
unremarkable systemic examination | 0
unremarkable auscultation of the heart | 0
unremarkable auscultation of the lungs | 0
sinus tachycardia | 0
moderately flattened T-waves | 0
unremarkable chest X-ray | 0
respiratory alkalosis | 0
elevated C reactive protein (CRP) of 230 mg/L | 0
elevated procalcitonin of 2.1 μg/L | 0
normal leucocytes at 7.1×109/L | 0
elevated troponin T (TnT) at 90 ng/L | 0
raised N-terminal pro-B-type natriuretic peptide (NT-proBNP) at 160 ng/L | 0
echocardiography showing good ventricular function | 0
no hypokinesia | 0
no significant valve pathology | 0
subcutaneous oedema on the left side | 0
multiple enlarged lymph nodes up to 2.0×2.7 cm in diameter | 0
deterioration of the left ventricular function with reduced systolic function of 40% | 48
CRP rose to 344 mg/L | 48
procalcitonin rose to 12.9 μg/L | 48
transferred to intensive care due to respiratory distress | 72
cellulitis on the neck suspected | 0
started on broad-spectrum antibiotics cefotaxime and clindamycin | 0
raised TnT | 0
raised NT-proBNP | 0
suspected cardiac involvement | 0
less likely myocardial infarction | 0
suggested myocarditis as differential diagnosis | 0
received acetylsalicylic acid 300 mg | 0
observed with telemetry | 0
planned CT angiogram | 0
planned cardiac MRI | 0
nasopharyngeal swab positive for SARS-CoV-2 | 0
respiratory distress | 72
saturating 94% on room air | 72
placed on 3 L/min of oxygen | 72
lactate of 3.2 mmol/L | 72
partial pressure of arterial oxygen (PaO2) of 6.3 | 72
oliguria | 72
hypotension (83/41 mm Hg) | 72
invasive haemodynamic monitoring instituted | 72
high-preload, hyperdynamic, vasodilated state | 72
received intravenous furosemide | 72
required low-dose norepinephrine infusion | 72
maintained a middle arterial pressure of >60 mm Hg | 72
normalised urine output | 72
continuous positive airway pressure | 72
oxygen (2 L/min) by nasal cannula | 72
oxygen saturation remained >93% | 72
bibasal consolidations | 72
TnT rose to 1959 ng/mL | 72
NT-proBNP rose to 11,169 ng/L | 72
cardiac MRI revealing diffuse myocardial oedema | 120
CT angiogram showed no coronary artery stenosis | 120
discharged | 264
readmitted with unilateral, right-sided peripheral facial nerve palsy | 336
unremarkable neurological examination | 336
unremarkable general clinical status | 336
normal cerebral CT scan | 336
elevated protein of 1.0 g/L | 336
elevated IgG of 0.14 g/L | 336
mild mononuclear pleocytosis at 7×106/L | 336
empirically treated with doxycycline | 336
discharged | 336
no anti-Borrelia antibodies detected | 336
borderline raised CXCL13 of 20.3 pg/mL | 336
negative PCR for neurotropic agents in spinal fluid | 336
high levels of anti-SARS-CoV-2 IgG antibodies in serum | 336
low levels of anti-SARS-CoV-2 IgG antibodies in spinal fluid | 336
antibody index 1.47 | 336
antiganglioside antibodies detected in serum | 336
cerebral MRI normal | 336
recovered completely from facial palsy | 336
decreased exercise tolerance | 336
no shortness of breath | 0
denies chest pain | 0
