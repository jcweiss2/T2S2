38 years old | 0
male | 0
accidental traumatic forearm amputation | -1
steel rope hit his arm | -1
tourniquet applied by paramedics | -1
tourniquet released | 0
decision for replantation | 0
broad spectrum antibiotic treatment | 0
replantation surgery | 0
multiple samples for microbiological testing | 0
arterial and venous anastomosis | 48
saphenous vein grafts | 48
Coldex skin substitute | 48
progressive swelling | 168
increasing skin necrosis | 168
venous congestion | 168
emergent re-exploration | 168
thrombosis of all blood vessels | 168
avital extensor and flexor muscles | 168
superficial fungal contamination | 168
amputation at the level of the proximal forearm | 168
systemic antifungal therapy (Amphotericin B) | 168
repeated surgical debridement | 192
multiple microbiologic and histologic probes | 192
polymicrobial infection | 192
Bacillus cereus complex | 192
Yersinia enterocolitica group | 192
Staphylococcus capitis | 192
Pseudomonas putida | 192
Aspergillus fumigatus | 192
Mucor circinelloides | 192
uncertainty about Mucor invasiveness | 192
antifungal therapy escalated to Isavuconazol | 360
antibiotic treatment to Tienam | 360
acute renal and multi-organ failure | 432
transfer to intensive care unit | 432
histologic confirmation of colonization | 504
treatment plan changed | 504
closure of the skin defect | 840
fasciocutaneous hatchet flap | 840
meshed skin graft | 840
graft healed | 945
transfer to rehabilitation center | 1008
follow-up without complications | 8760