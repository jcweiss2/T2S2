45 years old | 0
male | 0
admitted to the hospital | 0
fever | -48
chills | -48
productive cough | -48
runny nose | -48
headache | -48
temperature of 39.8°C | 0
heart rate of 115 beats/min | 0
blood pressure of 130/70 mmHg | 0
respiratory rate of 18/min | 0
throat was injected | 0
examination of his ears and oral cavity was unremarkable | 0
total white blood cell count was slightly raised | 0
WBC count 15.45 × 10^9/L | 0
chest radiograph was normal | 0
symptomatic treatment for presumed upper respiratory tract infection | 0
discharged from the A and E | 0
seizures | 6
status epilepticus | 6
heart rate of 173 bpm | 6
blood pressure measuring 94/57 mmHg | 6
cardiac auscultation was normal | 6
confused | 6
consciousness was impaired | 6
reflexes were preserved | 6
pupils were equal and reactive | 6
no papilledema | 6
WBC count increased to 31 × 10^9/L | 6
predominant neutrophils | 6
CRP levels were grossly elevated | 6
intubated | 6
noncontrast computed tomography of the brain | 6
subtle fullness in the right frontal region | 6
mild sulcal effacement | 6
paranasal sinuses showed a diffuse mucosal thickening | 6
lumbar puncture | 12
cerebrospinal fluid analysis revealed an infective picture | 12
Glasgow Coma Scale dropped from 10 to 7 | 12
contrast-enhanced magnetic resonance imaging of the brain | 14
large peripherally enhancing right frontotemporoparietal subdural collection | 14
smaller collections in the left frontal region | 14
severe mass effect in the right cerebral hemisphere | 14
midline shift | 14
fluid-filled paranasal sinuses showed mucosal hyperenhancement | 14
small bony defect in the posterior wall of the left frontal sinus | 14
adjacent meningeal enhancement | 14
right frontal parenchymal edema | 14
diagnosis of sinogenic meningoencephalitis with multiple SDEs | 14
antibiotic treatment started | 14
vancomycin | 14
ceftriaxone | 14
right decompressive craniectomy | 18
evacuation of SDE | 18
Frank pus was drained | 18
Streptococcus intermedius | 18
sensitive to multiple antibiotics | 18
functional endoscopic sinus surgery | 18
pus from the infected sinus had the same organism and antibiotic sensitivity | 18
postoperatively treated with intravenous antibiotics | 18
intravenous meropenem | 18
vancomycin | 18
intensive care unit for 5 days | 18
condition improved gradually | 24
GCS of 10 | 24
vital signs becoming normal | 24
extubated on his fourth postoperative day | 96
follow-up CT showed improvement of mass effect and cerebral edema | 120
discharged with good neurological status | 480
inflammatory markers demonstrated a gradual decline | 480
CRP was 51.4 mg/L | 480
no change in his personality or cognitive functions | 480
no motor or sensory deficits | 480
developed scar epilepsy | 720
follow-up CTs demonstrated a significant parenchymal loss and gliosis | 720
oral sodium valproate | 720
levetiracetam | 720