71 years old | 0
man | 0
productive cough | -168
fever | -168
transferred to emergency room | 0
endoscopic removal of fish bone | -168
admitted to local clinic | -168
symptoms suggestive of mediastinitis | -168
esophageal endoscopic examination | -168
no mucosal defect found | -168
conservative management with nothing by mouth | -168
antibiotics | -168
productive cough progressed | 0
fever progressed | 0
chest computed tomography (CT) performed | 0
CT scan showed wide esophageal perforation | 0
mediastinal abscess | 0
right pleural empyema | 0
arrival at our institution | 0
blood pressure steady | 0
tachypneic | 0
gastrografin esophagogram showed perforation in middle thoracic esophagus | 0
urgent intervention necessary | 0
aspiration pneumonia progressed in intensive care unit | 0
history of traumatic hemothorax | -infinity
pleural drainage for empyema in right chest | -infinity
calcified pleural lesions visible on CT scan | 0
decision to avoid thoracic incision | 0
no conventional thoracotomy | 0
no video-assisted thoracoscopic surgery | 0
posterior mediastinal drainage with Barovac PS400L | 48
incision on left side of neck | 48
drainage insufficient | 72
esophageal endoscopy performed | 72
multiple sites of wall injuries | 72
perforation 26-30 cm from incisor | 72
3-mm perforation 32 cm from incisor | 72
2.5-cm-deep laceration 35 cm from incisor | 72
insertion of 2 Levin tubes via esophageal endoscopy | 72
12-Fr tube inserted into mediastinum | 72
12-Fr tube inserted into stomach for gastric drainage | 72
Stenotrophomonas maltophilia identified | 72
antibiotic regimen adjusted | 72
continuous suction of 60-80 mm Hg for mediastinal and gastric drainage | 72
aggressive mediastinal and gastric drainage started | 72
patient's condition improved | 72
jejunostomy performed | 216
gastrostomy performed | 216
Levin tube removed | 216
continuous suction maintained for mediastinal drainage | 216
natural drainage started during jejunostomy and gastrostomy | 216
extubated | 264
moved to general ward | 432
suction turned off for mediastinal drainage | 456
natural drainage started | 456
amount of drainage sufficiently reduced | 456
microbiologic culture on 13th hospital day | 312
no pathologic microorganism other than normal flora | 312
multiple consecutive microbiologic cultures same | 312
remaining Levin tube removed | 600
follow-up endoscopic examination on 26th hospital day | 624
previous injury sites nearly healed | 624
0.5-cm defect 28 cm from incisor | 624
follow-up chest CT scan on 29th hospital day | 696
notable decrease in mediastinal abscess | 696
follow-up esophagogram on 39th hospital day | 936
no evidence of leakage | 936
oral diet started | 936
discharged | 1104
follow-up esophagogram and endoscopic examination 6 months after initial presentation | 4320
no abnormal findings | 4320
esophageal perforation | 0
mediastinal contamination | 0
sepsis control | 0
perforation closure | 0
contamination drainage | 0
Stenotrophomonas maltophilia infection | 72
aspiration pneumonia | 0
mediastinal abscess drainage | 48
gastric drainage | 72
postpyloric nutrition | 216
esophageal injury healed | 624
failed E-VAC attempt | 0
high perioperative risk | 0
less-invasive methods chosen | 0
internal drainage | 72
adjuvant procedures | 72
conflict of interest | 0
no complications reported | 1104
