68 years old | 0
male | 0
biological aortic valve replacement | -2520
severe aortic stenosis | -2520
right coronary artery disease | -2520
persistent atrial fibrillation | -2520
admitted to the hospital | 0
fever | -72
dyspnoea | -72
dysarthria | -72
MSSA endocarditis | -72
aortic bioprosthesis | -72
secondary haemorrhagic stroke | -72
septic embolus | -72
treatment with intravenous antibiotics | -72
discharged | -744
neurological rehabilitation | -744
recurrent wide QRS complex tachycardia | 0
synchronized electrical cardioversions | 0
intravenous adenosine | 0
emergent electrophysiology study | 6
atrioventricular nodal catheter ablation | 6
incessant junctional ectopic tachycardia (JET) | 6
temporary pacemaker insertion | 6
recurrent JET | 72
redo catheter ablation | 72
permanent pacemaker insertion | 168
pacemaker interrogation | 2160
pseudoaneurysm of the right sinus of Valsalva | 0
infective endocarditis of a bioprosthetic valve | 0
haemodynamic collapse | 0
atrioventricular block (AVB) | 0
long PR intervals | 0
2:1 AVB | 0
normal left ventricular ejection fraction | 0
aortic bioprosthesis without dysfunction | 0
dilation of the right sinus of Valsalva | 0
multiple recurrences of the same tachycardia | 12
repeated synchronized electrical cardioversion | 12
increasing need for vasopressor drugs | 12
temporary wire insertion | 12
ventriculoatrial (VA) dissociation | 12
overdrive pacing | 12
synchronized shocks | 12
amiodarone administration | 12
emergency catheter ablation | 12
atrioventricular node (AVN) ablation | 12
His potential not visible | 12
ablation catheter positioned anatomically | 12
tachycardia stopped | 12
temporary pacing | 12
arrhythmia recurred | 48
redo ablation | 48
permanent pacemaker implantation | 168
blood cultures remained negative | 168
patient remained afebrile | 168
ejection fraction 65-70% | 1440
patient capable of walking and climbing stairs | 1440