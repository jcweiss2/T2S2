25 years old | 0
man | 0
intravenous drug abuse | 0
fevers | 0
back pain | 0
abdominal pain | 0
bilateral LE swelling | 0
sinus tachycardia | 0
extensive bilateral ileofemoral acute-on-chronic deep vein thrombosis | 0
extensive bilateral femoropopliteal acute-on-chronic deep vein thrombosis | 0
venous duplex imaging | 0
leukocytosis | 0
methicillin-resistant Staphylococcus aureus bacteremia | 0
tenderness to palpation in the epigastrium | 0
locally palpable thrill | 0
anasarca | 0
phlegmasia alba dolens of the bilateral LEs | 0
infrarenal MAAA | 0
spontaneous decompression via erosion into the IVC | 0
giant aortocaval fistula | 0
diminished distal arterial flow | 0
cavernous transformation of the ileofemoral venous network | 0
symmetrically diminished ankle-brachial indexes | 0
dampened aortoiliac pulse-volume recordings | 0
no evidence of active vegetation on echocardiography | 0
significant acute cardiopulmonary overload | 0
sepsis | 0
significant arterialization of the venous system | 0
endovascular aneurysm repair | -24
hemodynamic stability achieved | 0
resolution of tachycardia | 0
phlegmasia improved | 72
leukocytosis resolved | 144
negative blood cultures | 168
afebrile for 1 week | 168
bilateral axillary unifemoral bypass grafts | 168
ligation of the aortic stump | 168
ligation of the IVC | 168
endograft explant | 192
recovery in the intensive care unit | 192
discharged home | 240
vancomycin administered through a peripherally inserted central catheter | 240
follow-up at 1 month | 720
follow-up at 3 months | 2160
smooth recovery | 2160
no complications | 2160
venous duplex imaging |'0
