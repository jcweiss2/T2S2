female | 0 | 0 | Factual
59 years old | 0 | 0 | Factual
liver cancer | -672 | 0 | Factual
transarterial embolization | -392 | -392 | Factual
sorafenib | -168 | -56 | Factual
dizziness | -56 | -56 | Factual
skin ulcers | -56 | -56 | Factual
radiation therapy | -14 | -14 | Factual
liver transplantation | 0 | 0 | Factual
hepatitis B | 0 | 0 | Factual
entecavir | 0 | 0 | Factual
HBV serology test | 0 | 0 | Factual
immunosuppressive drugs | 24 | 24 | Factual
steroids | 24 | 24 | Factual
tacrolimus | 24 | 24 | Factual
acute renal failure | 24 | 24 | Factual
hematoma | 24 | 24 | Factual
hepatitis B immunoglobulin | 24 | 24 | Factual
fever | 240 | 552 | Factual
rash | 408 | 552 | Factual
procalcitonin | 240 | 312 | Factual
blood cultures | 312 | 312 | Factual
cytomegalovirus | 312 | 312 | Factual
Epstein-Barr virus | 312 | 312 | Factual
sirolimus | 408 | 408 | Factual
mycophenolate mofetil | 408 | 408 | Factual
Acinetobacter baumannii | 432 | 432 | Factual
methicillin-resistant Staphylococcus aureus | 432 | 432 | Factual
erythematous macules | 456 | 456 | Factual
papules | 456 | 456 | Factual
bone marrow suppression | 456 | 456 | Factual
white blood cell count | 456 | 456 | Factual
platelet count | 456 | 456 | Factual
hemoglobin | 456 | 456 | Factual
gamma globulin | 456 | 456 | Factual
skin biopsy | 504 | 504 | Factual
FISH analysis | 504 | 504 | Factual
donor lymphocytes | 504 | 504 | Factual
immunoglobin M | 504 | 504 | Factual
septic shock | 552 | 552 | Factual
multiple organ dysfunction syndrome | 552 | 552 | Factual
death | 552 | 552 | Factual