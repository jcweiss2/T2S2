28 years old | 0\
male | 0\
attended a health center | -24\
fatigue | -24\
anosmia | -24\
dyspnea | -24\
SpO2 levels were 55% | -24\
nasal cannula oxygen therapy | -24\
SpO2 levels were 75% | -24\
hospitalized | -24\
evaluated at an emergency department | -24\
chest radiography | -24\
bilateral lung infiltrates | -24\
RT-PCR swab tested positive for SARS-CoV-2 infection | -24\
admitted in a COVID-19 infirmary unit | -24\
non-invasive ventilation support | -24\
intubation | -24\
invasive mechanical ventilation | -24\
ventral decubitus positioning | -24\
Escherichia coli and methicillin-sensitive Staphylococcus aureus were detected on sputum culture | -48\
superinfection | -48\
prescription of an 8-day regimen of amoxicillin | -48\
blood culture revealed methicillin-resistant Staphylococcus aureus | -48\
steady clinical improvement | -48\
extubated | -48\
discharged | -168\
retrosternal thoracalgia irradiating to the left upper limb | -168\
abduction and external rotation were limited due to pain complaints | -168\
soft tissue swelling of the shoulder and arm | -168\
fever | -168\
increased levels of C-reactive protein | -168\
admitted for further investigation and treatment planning | -168\
gentamicin was prescribed and administered | -168\
thoracic CT with intravenous contrast administration | -159\
scapulohumeral synovitis | -159\
multiple intra-muscular collections | -159\
bilateral shoulder magnetic resonance imaging (MRI) with intravenous contrast administration | -156\
infraspinatus fossa and subscapular fossa collections | -156\
capsular thickening and increased signal intensity post-gadolinium administration | -156\
septic arthritis and rotator cuff collections | -156\
myonecrosis | -156\
aspiration of the infraspinatus fossa collection | -156\
seropurulent fluid | -156\
anaerobic and aerobic bacteria were negative | -156\
physical rehabilitation exercises | -156\
transferred to another hospital | -144\
indication to continue physical therapy and rehabilitation exercises | -144