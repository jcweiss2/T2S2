37 years old | 0
male | 0
quadriplegia | -672
chronic hypoxic respiratory failure | -672
mechanical ventilation | -672
tracheostomy | -672
admitted to the intensive care unit | 0
pneumonia | 0
serum creatinine level 1.39 mg/dl | 0
chest imaging result suggestive of multifocal pneumonia | 0
acute respiratory distress syndrome | 48
septic shock | 48
vasopressor therapy | 48
worsening oxygen requirement | 48
test result for novel coronavirus SARS-CoV-2 negative | 48
serum creatinine level worsened to 3.3 mg/dl | 72
decline in urine output | 72
renal sonogram obtained | 72
fractional excretion of urea 25.6% | 72
intravascular volume depletion | 72
diuretics | 72
bolus of i.v. fluid administered | 72
nephrology consultation requested | 72
question about possible glomerulonephritis | 72
pulmonary-renal syndrome | 72
antinuclear antibody test result positive | 72
bronchoscopy equivocal for alveolar hemorrhage | 72
mechanical ventilation | 0
fraction of inspired oxygen 70% | 0
positive end-expiratory pressure 12 cm H2O | 0
blood pressure 96/53 mm Hg | 0
pulse rate 92 beats per minute | 0
oxygen saturation 90% | 0
bilateral lung crackles | 0
trace pitting pedal edema | 0
urine output approximately 350 ml in the past 24 hours | 0
urine microscopy results demonstrated muddy brown casts | 0
tubular injury | 0
no dysmorphic red blood cells | 0
elevated serum creatinine levels | 0
mild hypernatremia | 0
hyperkalemia | 0
serum bicarbonate 25 mmol/l | 0
bedside ultrasound performed | 0
lung ultrasound revealed bilateral diffuse B-line pattern | 0
irregular pleural line | 0
focused cardiac ultrasound revealed hyperdynamic left ventricular systolic function | 0
enlarged right ventricle | 0
interventricular septal flattening | 0
D-sign | 0
volume and/or pressure overload | 0
inferior vena cava plethoric | 0
IVC-estimated right atrial pressure unreliable | 0
hepatic and portal vein Doppler performed | 0
hepatic vein Doppler waveform revealed S-wave reversal | 0
severely elevated RAP level | 0
portal vein Doppler waveform pulsatile with intermittent flow reversal | 0
severe venous congestion | 0
continuous renal replacement therapy initiated | 0
anti–double-stranded DNA negative | 72
antiglomerular basement membrane negative | 72
antineutrophil cytoplasmic antibodies negative | 72
renal biopsy not considered | 72
POCUS parameters used to guide decongestive therapy | 72
documented fluid balance negative 6.6 l | 72
hepatic vein Doppler showed S-wave below the baseline | 72
portal vein pulsatility improved | 72
blood pressure 115/57 mm Hg | 72
no vasopressors | 72
ultrafiltration continued | 72
fluid balance negative 5.1 l | 120
hepatic vein Doppler similar to previous tracing | 120
portal vein waveform normalized | 120
urine output 150 ml in the previous 24 hours | 120
continuous renal replacement therapy discontinued | 120
plan to transition to intermittent hemodialysis | 120
portal vein waveform improved before hepatic | 120
patient made more urine overnight | 144
did not require hemodialysis | 144
fluid balance negative 2 l | 192
hepatic vein Doppler normalized | 192
portal vein remained normal | 192
resolved venous congestion | 192
IVC remained dilated | 192
lung ultrasound showed improvement | 192
D-sign on cardiac ultrasound disappeared | 192
left ventricle returned to its normal circular shape | 192
serum creatinine level 2.1 mg/dl | 192
eventually trended down to 0.6 mg/dl | 336