42 years old | 0
female | 0
multiparous | 0
admitted to the ER | 0
altered mentation | 0
seizures | 0
high fever | 0
tested positive for COVID-19 | -48
throat pain | -48
nasopharyngeal COVID-19 PCR test | 0
endotracheal intubation | 0
emergency call to the obstetrics and gynecology department | 0
critical illness | 0
mechanical ventilation | 0
previous delivery by cesarean section | -10080
no underlying diseases | 0
no remarkable events during prenatal examinations | 0
no history of drug abuse | 0
no smoking | 0
no drinking | 0
generalized tonic-clonic type seizure | 0
drooling | 0
upper eyeball deviation | 0
prompt pupillary reflex | 0
blood pressure 121/71 mmHg | 0
heart rate 115 beats per minute | 0
increased C-reactive protein | 0
erythrocyte sedimentation rate | 0
D-dimer | 0
no proteinuria | 0
normal liver function test | 0
normal serum electrolytes | 0
normal blood glucose | 0
normal blood urea nitrogen | 0
normal creatinine | 0
thyroid function test | 0
TSH < 0.01 mIU/L | 0
free T4 1.95 ng/dL | 0
total T3 183.9 ng/dL | 0
overt hyperthyroidism | 0
Burch-Wartofsky Point Scale 65 | 0
brain computed tomography | 0
no acute intracranial hemorrhage | 0
no focal parenchymal lesions | 0
no visible causes of seizure | 0
chest X-ray | 0
electrocardiogram | 0
ultrasonography | 0
fetal growth appropriate for gestational age | 0
fetal heartbeat and movements normal | 0
no significant uterine contractions | 0
initial diagnosis of eclampsia | 0
atypical eclampsia | 0
final diagnosis of status epilepticus | 0
final diagnosis of thyroid storm | 0
final diagnosis of Graves’ disease | 0
treatment with labetalol | 0
treatment with magnesium sulfate | 0
treatment with midazolam | 0
cesarean section | 24
newborn infant weighed 2680 g | 24
1 min and 5 min Apgar scores 8 and 8 | 24
low-level sedation with midazolam | 24
intensive care unit | 24
seizures decreased | 36
consciousness restored | 36
newborn's nasopharyngeal COVID-19 PCR test negative | 24
thyroid function tests normal | 24
magnetic resonance imaging | 48
electroencephalogram | 48
no specific findings | 48
referral to endocrinologist | 48
evaluation and treatment of hyperthyroidism | 48
TSH < 0.01 mIU/L | 48
free T4 1.86 ng/dL | 48
total T3 175.3 ng/dL | 48
TSH receptor antibody 2.44 IU/L | 48
thyroid ultrasonography | 48
diffusely enlarged thyroid gland | 48
papillary carcinoma | 48
thyroidectomy scheduled | 48
methimazole | 48
methylprednisolone | 48
propranolol | 48
discharged in a healthy condition | 240
thyroid function test results close to normal values | 720