85 years old | 0
male | 0
admitted to the hospital | 0
severe valvular and ischaemic-hypertensive cardiopathy | 0
slight chronic renal failure | 0
chronic venous leg ulcers | 0
plunged his legs in seawater | -336
fever | 12
pain on the distal left lower limb | 0
ulcer on the left lateral ankle | 0
fibrinous, greenish and smelly coating | 0
varicose veins | 0
stasis dermatitis | 0
lipodermatosclerosis | 0
elevated CRP | 0
leucocytosis | 0
ankle-brachial pressure index | 0
X-ray | 0
infection of the wound | 0
intravenous antibiotic therapy with amoxicillin and clavulanic acid | 0
cellulitis in the left leg | 12
hypotension | 12
acute renal failure | 12
septic shock | 12
antibiotic changed to parenteral imipenem | 12
intravenous catecholamines | 12
blood cultures showed growth of V. parahaemolyticus | 12
bacteriological smear of the wounds showed growth of V. parahaemolyticus | 12
bacteriological smear of the wounds showed growth of Pseudomonas aeruginosa | 12
bacteriological smear of the wounds showed growth of Morganella morganii | 12
bacteriological smear of the wounds showed growth of Streptococcus mitis | 12
bacteriological smear of the wounds showed growth of Enterococcus spp | 12
stopped treatment with imipenem | 72
started targeted combined antibiotic therapy with oral ciprofloxacin and doxycycline | 72
normalization of haemodynamics | 168
return to the patient's usual renal parameters | 168
chronic hepatitis B infection | 0
hepatic function was globally intact | 0
sonography of the abdomen showed a “cardiac liver” with portal hypertension | 0
local therapy of the chronic wounds | 0
daily curettage | 0
application of topic sulphonamide | 0
pressure bandage of the lower limbs | 0
application of negative pressure wound treatment | 0
stopped negative pressure wound treatment | 72
discharged from the hospital | 168
treated the patient regularly in our outpatient clinic | 168
satisfactory granulation of the wound ground | 672
application of a split-thickness skin graft to the left leg | 672
complete wound healing | 720