67 years old | 0
    male | 0
    aorto-bi, iliac graft replacement placement for abdominal aortic aneurysm (AAA) | -8760
    AAA repair | -8760
    paraplegia | -8760
    graft leaking | -8760
    embolization | -8760
    fever | 0
    lethargy | 0
    tachycardia | 0
    tachypnea | 0
    hypotension | 0
    minimally responsive | 0
    unable to maintain airway | 0
    minimal peri-umbilical tenderness with deep palpation | 0
    no peritoneal signs | 0
    emergent intubation | 0
    transferred to medical critical care unit | 0
    white blood cell count 17,000/μL | 0
    hemoglobin 9.6 g/dL | 0
    platelet count 300,000/μL | 0
    BUN 66 mg/dL | 0
    Cr 2.1 mg/dL | 0
    minimal elevation of troponin | 0
    normal level of electrolytes | 0
    diagnosis of severe sepsis | 0
    septic shock of unknown source | 0
    empirical treatment with vancomycin | 0
    empirical treatment with meropenem | 0
    urine cultures negative | 0
    respiratory culture negative | 0
    blood culture demonstrated Eggerthella lenta | 0
    blood culture demonstrated Escherichia coli ESBL | 0
    blood culture demonstrated Enterococcus faecalis | 0
    transesophageal echocardiogram revealed no vegetation | 0
    abdominal CT with contrast demonstrated inflammatory changes around aorto-bi-iliac graft | 0
    no aortoenteric fistula | 0
    Indium-111 WBC scan showed increased activity in mid to lower abdomen | 0
    vascular surgery evaluation | 0
    unstable condition | 0
    vascular interventions deferred | 0
    frail condition | 0
    conservative strategy | 0
    IV vancomycin 1 g daily | 0
    IV meropenem 1 g twice daily | 0
    seven days course | 168
    continued fever | 168
    unable to wean from mechanical ventilation | 168
    repeat blood culture grew Eggerthella lenta | 168
    repeat blood culture grew Escherichia coli ESBL | 168
    repeat blood culture grew Enterococcus faecalis | 168
    antibiotic regimen changed to tigecycline 50 mg twice daily | 168
    tigecycline administered for 14 days | 168
    two days after tigecycline | 192
    repeat blood cultures negative | 192
    completion of antibiotics course | 336
    stabilization of comorbidities | 336
    discharged home | 336
    long term antibiotic therapy | 336
    close control of inflammation markers | 336
    
    