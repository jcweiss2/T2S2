26 years old | 0
    female | 0
    presented to the emergency department | 0
    first injection of ChAdOx1 nCoV-19 vaccine | -336
    headache nonresponsive to anti-inflammatory drugs | -336
    right-sided weakness | 0
    visual disturbances | 0
    combined (estrogen-progestogen) contraceptives | -87600
    general examination normal | 0
    vital signs normal | 0
    neurological examination severe right-sided weakness | 0
    CT scan hyperdense rectus sinus | 0
    CT scan hyperdense vein of Galen | 0
    MRI venography multifocal venous thrombosis | 0
    bilateral occlusion of parietal cortical veins | 0
    straight sinus occlusion | 0
    vein of Galen occlusion | 0
    internal cerebral veins occlusion | 0
    inferior sagittal sinus occlusion | 0
    transverse sinuses partially involved | 0
    extensive venous infarction with hemorrhagic transformation | 0
    D-dimer raised 12,204 mg/L | 0
    platelet count 134x10^9/L | 0
    treated with fondaparinux 5 mg subcutaneously | 0
    admitted to intensive care unit | 0
    clinical condition deteriorated | 24
    decreased consciousness | 24
    right-sided hemiplegia | 24
    complete Balint syndrome | 24
    blood collection T0 April 13 | -48
    blood collection T1 April 15 | 0
    blood collection T2 April 20 | 120
    PT normal | 0
    aPTT normal | 0
    FV-Leiden mutation absent | 0
    G20210A-prothrombin mutation absent | 0
    antithrombin normal | 0
    protein C/S normal | 0
    lupus anticoagulant negative | 0
    antiphospholipid antibodies negative | 0
    aPF4-heparin IgG ELISA positive | 0
    platelet activation test positive | 0
    PF4–heparin antibodies inhibited by heparin | 0
    platelet thrombus formation impaired | 0
    AUC smaller | 0
    OT longer | 0
    hypercoagulability | 0
    short lag-time | 0
    increased thrombin-peak | 0
    short time-to-peak | 0
    increased ETP | 0
    increased ETP-TM ratio | 0
    FVIII increased 200 U/dL | 0
    PC normal 88 U/dL | 0
    FVIII/PC ratio increased 2.3 | 0
    IVIG 1 g/kg o.d. for 2 days | 24
    dexamethasone 40 mg/day for 4 days | 24
    fondaparinux replaced by argatroban | 24
    argatroban increased to 3 mg/kg/min | 24
    neurological conditions improved | 72
    awake | 72
    fully responsive to stimuli | 72
    progressive recovery of right upper-limb strength | 72
    partial optic ataxia | 72
    regression of apraxia | 72
    CT scan normal rectus sinus | 120
    CT scan normal vein of Galen | 120
    oedema in brain tissue | 120
    MRI venography restored venous flow rectus sinus | 120
    MRI venography restored venous flow vein of Galen | 120
    right internal cerebral vein still occluded | 120
    bilateral frontoparietal cortical veins still occluded | 120
    intraparenchymal venous infarction unchanged | 120
    platelet count increased 339x10^9/L | 120
    D-dimer decreased to normal levels | 120
    aPF4 reactivity reduced | 120
    patient serum no platelet activation | 120
    moderate disability | 1680
    no neuropsychological deficits | 1680
    walk unassisted for short distances | 1680
    sustained clonus | 1680
    spasticity in right leg | 1680
    right arm almost fully recovered | 1680
    fondaparinux replaced with oral vitamin K antagonist | 1680
    VITT | 0
    cerebral venous thrombosis | 0
    bi8hemispheric hemorrhage | 0
    successful treatment with argatroban | 0
    successful treatment with IVIG | 0
    successful treatment with corticosteroids | 0
    high-titer aPF4 | 0
    signs of platelet activation | 0
    platelet count decreased by approximately 50% | 0
    avoided heparin treatment | 0
    immune modulating therapy | 0
    reduction of aPF4 titer | 0
    reduction of D-dimer | 0
    antibodies to PF4 induced platelet activation | 0
    loss of serum activity in PAT | 0
    IVIG blockade of FCγ platelet receptors | 0
    antibody suppression | 0
    platelets’ ability to promote thrombus formation reduced | 0
    laboratory tests correlated with clinical course | 0
    early multidisciplinary therapeutic approach | 0
    resolution of the syndrome | 0
    