27 years old | 0
female | 0
admitted to the emergency department | 0
ingested delayed-release venlafaxine | -12
ingested large amount of alcohol | -12
hallucinations | 0
hyperreflexia | 0
mydriasis | 0
trismus | 0
opsoclonus | 0
myoclonus | 0
serotonergic syndrome | 0
sinus tachycardia | 0
prolonged corrected QT-interval (QTc) 513ms | 0
standard QRS width | 0
blood-alcohol level 2.32 ‰ | 0
glucose level 238 mg/dL | 0
negative drug screening tests | 0
received 2000 ml Sterofundin | 0
received 12 mg midazolam | 0
transferred to intensive care unit | 0
recurring severe hypoglycemia | 12
received 200 ml 20% glucose solution | 12
blood pressure declined | 12
severe chest wall rigidity | 12
hypoxemia | 12
invasive ventilation | 12
received 5 mg midazolam | 12
received 50 μg sufentanil | 12
received 50 mg rocuronium | 12
vasopressors needed | 12
noradrenaline up to 10 mg/h | 12
dobutamine up to 30 mg/h | 12
progressive lactic acidosis | 12
lactic acid 1.8 mmol/L | 12
lactic acid increased to 19.1 mmol/L | 17
severe left-ventricular dysfunction | 13
LVEF 10-15% | 13
global left-ventricular hypokinesia | 13
hemodynamic instability | 17
veno(arterial extracorporeal life support (ECLS) | 17
diffuse bleeding | 17
INR 3.6 | 17
PTT 62 s | 17
antithrombin III 28% | 17
fibrinogen 0.4 g/L | 17
GOT > 7000 U/I | 17
acute liver failure | 17
disseminated intravascular coagulation | 17
venlafaxine serum concentration > 720 μg/L | 17
acute kidney failure | 17
slow low-efficiency dialysis initiated | 17
dialysis continued for fifteen days | 17
systemic heparin used | 17
ECLS explantation | 168
regional calcium citrate anticoagulation | 168
continuous heparin 400 IE/h | 168
septic shock | 96
procalcitonin 11.6 mmols/L | 96
serum lactate 5.6 mmol/L | 96
increased noradrenaline | 96
increased fluid replacement | 96
pressure-controlled ventilation | 96
oxygen demand increased | 96
chest X-ray infiltrates | 96
ventilator-associated pneumonia | 96
meropenem initiated | 96
vancomycin initiated | 96
anisocoria | 96
distorted pupils | 96
cranial imaging normal | 96
pupil abnormalities resolved | 144
high doses midazolam 1.2 mg/kg/h | 144
high doses sufentanil 0.8 μg/kg/h | 144
LVEF 45% | 168
LVEF 55% | 504
ECLS weaned | 168
extubated | 336
pneumonia improved | 336
oriented | 336
no neurological damage | 336
lesion of N. peroneus | 336
transferred to general ward | 336
transferred to rehabilitation | 336
