60 years old | 0
male | 0
diagnosed with glomerulonephritis secondary to anti-neutrophil cytoplasmic antibody-positive microscopic polyangiitis | -720
elevated creatinine | -720
treated with intravenous methylprednisolone | -720
treated with oral cyclophosphamide | -720
renal function normalized | -720
discharged home | -720
prednisolone | -720
cyclophosphamide | -720
admitted to regional hospital | -336
nausea | -336
vomiting | -336
diarrhea | -336
intolerance of oral intake | -336
large volume watery diarrhea | -336
transfer to tertiary hospital intensive care unit | -336
hemofiltration for hypovolemic acute kidney injury | -336
cyclophosphamide reduced to 50 mg daily | -336
cyclophosphamide ceased | -336
received approximately one month of cyclophosphamide | -336
total cyclophosphamide dose 2.1 g | -336
empiric antimicrobial therapy commenced | -336
tazobactam | -336
piperacillin | -336
intravenous metronidazole | -336
ganciclovir | -336
secretory diarrhea | -336
no infective agents identified | -336
vasoactive intestinal polypeptide non-diagnostic | -336
chromogranin levels non-diagnostic | -336
diffuse mural thickening of small and large bowel | -336
denuded and erythematous mucosa in duodenum | -336
denuded and erythematous mucosa in sigmoid colon to terminal ileum | -336
rectum relatively spared | -336
full thickness mucosal ulceration | -336
inflammation throughout terminal ileum and large bowel | -336
no features of inflammatory bowel disease | -336
no vasculitis | -336
no viral inclusions | -336
diarrhea persisted | -336
maximal doses of antidiarrheals | -336
octreotide | -336
cholestyramine | -336
repeat imaging failed to reveal etiology | -336
stool specimens negative | -336
endoscopic evaluation negative | -336
histopathology negative | -336
regenerative mucosal changes | -336
viral PCR negative | -336
bacterial cultures negative | -336
fungal cultures negative | -336
required continuous intravenous therapy | -336
electrolyte replacements | -336
total parenteral nutrition | -336
severe hypoalbuminemia | -336
infliximab administered | -336
no clinical improvement | -336
no endoscopic improvement | -336
septic complications with Enterobacter | -336
Candida glabrata bacteremia | -336
returned to intensive care | -336
died from severe acute respiratory distress syndrome | -336
post-mortem examination showed hemorrhagic ulceration in small bowel | -336
minimal residual mucosa in small bowel | -336
similar changes in ascending and transverse colon | -336
retained mucosa in descending colon | -336
relative sparing of rectum | -336
no evidence of vasculitis | -336
no thromboemboli | -336
no infectious etiology identified | -336
herpes simplex virus-1 DNA detected | -336
Enterobacter faecium cultured | -336
Candida krusei cultured | -336
Pneumocystis jiroveci cultured | -336
metastatic pulmonary calcification | -336
diffuse alveolar damage | -336
Candida krusei cultured in bowel | -336
severe multifocal ulcerative enterocolitis | -336
hemorrhagic enterocolitis | -336
acute hypovolaemic renal failure | -336
metabolic acidosis | -336
sepsis with Enterobacter | -336
Candida septicemia | -336
alterations in intestinal microbiome | -336
excessive reactive oxygen species | -336
upregulation of pro-inflammatory cytokines | -336
hemorrhagic cystitis absent | -336
large volume fluid replacement | -336
electrolyte replacement | -336
parenteral nutrition | -336
intestinal transplantation contraindicated | -336
prophylactic antimicrobial therapy | -336
early supportive care | -336
cessation of cyclophosphamide | -336
fatal enteropathy | -336
persistent hypokalemia | -336
hypomagnesemia | -336
hypophosphatemia | -336
hypoalbuminemia | -336
raised inflammatory markers | -336
no infective agents cultured | -336
computed tomography of abdomen showing diffuse mural thickening | -336
endoscopic biopsy showing full thickness ulceration | -336
no granulomas | -336
treatment with prophylactic antibiotics | -336
antivirals | -336
antifungals | -336
anti-diarrhoeals | -336
intravenous fluids | -336
electrolytes | -336
glucocorticoids | -336
infliximab | -336
hemorrhagic colitis resolved after cessation of cyclophosphamide | -336
neutropenic enterocolitis | -336
profound neutropenia absent | -336
IV steroid unsuccessful | -336
tissue PCR negative | -336
cultures negative | -336
prolonged immunosuppression | -336
failure of mucosal regeneration | -336
mucosal necrosis | -336
mucosal regeneration on repeat biopsies | -336
no repopulation of mucosal epithelium | -336
complications with malnutrition | -336
empiric treatment for infections | -336
early suspicion of adverse event | -336
timely cessation of cyclophosphamide | -336
prevention of morbidity | -336
prevention of mortality | -336
case report highlights fatal enteropathy | -336
etiology unclear | -336
risk factors unclear | -336
treatment unclear | -336
prophylactic antimicrobial therapy consideration | -336
early supportive care consideration | -336
disseminated message to protect future adverse events | -336
exempt from Institutional Review Board | -336
informed consent waived | -336
peer-review started | -336
first decision | -336
article in press | -336
no conflicts of interest | -336
no funding disclosed | -336
manuscript source: Unsolicited manuscript | -336
specialty type: Gastroenterology and hepatology | -336
country of origin: Australia | -336
peer-review report classification Grade A | -336
Grade B | -336
Grade C | -336
Grade D | -336
Grade E | -336
conflict-of-interest statement | -336
institutional review board statement | -336
informed consent statement | -336
peer-review timeline | -336
PEER REVIEW PROCESS | -336
references | -336
figures | -336
tables | -336
author contributions | -336
acknowledgments | -336
authors’ affiliations | -336
abbreviations | -336
competing interests | -336
availability of data and materials | -336
ethical approval | -336
consent for publication | -336
copyright | -336
license | -336
open access | -336
correspondence | -336
supplementary material | -336
footnotes | -336
keywords | -336
