76 years old | 0
female | 0
admitted to the hospital | 0
generalized malaise | -168
shortness of breath | -168
lower extremity swelling | -168
subjective fever | -168
denies chest pain | -168
denies orthopnea | -168
denies paroxysmal nocturnal dyspnea | -168
blood pressure 79/54 mmHg | -168
oral temperature 38.3°C | -168
heart rate 55 beats/min | -168
crackles up to the mid-lung fields bilaterally | -168
irregularly irregular heart rhythm | -168
2+ pitting edema up to the knees | -168
atrial fibrillation on coumadin | -672
rheumatic heart disease | -672
congestive heart failure | -672
digoxin | -672
congestive heart failure exacerbation | 720
readmitted to the hospital | 720
history of atrial fibrillation | 0
history of rheumatic heart disease | 0
history of congestive heart failure | 0
history of digoxin | 0
history of congestive heart failure exacerbation | 720
positive blood cultures for Pasteurella multicoda | 0
ceftriaxone | 0
digoxin immune fab (Digibind) | 0
echocardiogram | 0
ejection fraction of 45% to 49% | 0
possible vegetation on the mitral valve | 0
severe eccentric mitral and tricuspid regurgitation | 0
transesophageal echocardiogram | 0
mitral valve vegetation measuring 1.2×0.7 cm | 0
severe biatrial enlargement | 0
left atrium volume 101.40 mL/m2 | 0
right atrium volume 233.80 mL/m2 | 0
previous echocardiogram was unobtainable | 0
head computed tomography | 0
chronic infarctions likely from septic emboli | 0
owned 4 cats | 0
cardiothoracic surgery team evaluated the patient | 0
multi-valve replacement surgery and biopsy of the vegetation | 0
conserved treatment | 0
discharged to a skilled nursing facility | 168
6-week course of ceftriaxone | 168
readmitted for congestive heart failure exacerbation | 720
hospice care | 720
Note: The time stamps are approximate and based on the text.