22 years old | 0  
    woman | 0  
    admitted to the emergency department | 0  
    swallowing difficulties | 0  
    throat pain | 0  
    local inflammation of the tonsils on the left side | 0  
    acute tonsillitis | 0  
    symptomatic therapy with ibuprofen | 0  
    discharged | 0  
    presented at ophthalmology outpatient department | 144  
    acute paresis of the abducens nerve | 144  
    partial paresis of the right oculomotor nerve | 144  
    general mydriasis of the right eye | 144  
    impairment in function of the musculus levator | 144  
    general impairment in motion of the right eye | 144  
    paresis of the right abducens nerve | 144  
    prism cover test showed +40 pdpt when looking to the right | 144  
    primary position at +20 pdpt when looking to the left +10 pdpt | 144  
    discrete paralysis of the abducens nerve on the left eye | 216  
    onset of exophthalmos on the right side | 216  
    documented by the Hertel Exophthalmometer | 216  
    no pathological signs in fundus and retina | 216  
    neurological investigation revealed general photophobia | 216  
    incomplete trismus | 216  
    discrete signs of meningism | 216  
    fever | 216  
    sepsis | 216  
    substantial inflammation | 216  
    leucocytosis of 16,000/µL | 216  
    15,000/µL neutrophils | 216  
    45% left shift | 216  
    C-reactive protein of 271 g/L | 216  
    activated coagulation | 216  
    profound thrombocytopenia (21,000/µL) | 216  
    international normalized ratio of 1.27 | 216  
    MRI investigation of the head | 216  
    marked thromboses at various locations including the cavernous sinus on both sides | 216  
    more pronounced on the right side | 216  
    thrombosis of the superior ophthalmic vein in the right eye | 216  
    small starting abscess in the right temporal lobe | 216  
    computed tomography of the neck | 216  
    abscess in the left tonsil with a maximum diameter of 6 mm | 216  
    partially occluding thrombus in the right internal jugular vein | 216  
    computed tomography of the lung | 216  
    multiple septic emboli | 216  
    starting abscesses | 216  
    diagnosis of Lemierre's syndrome | 216  
    high-dose intravenous antibiotic therapy with amoxicillin/clavulanic acid | 216  
    clindamycin | 216  
    two pairs of blood cultures | 216  
    anticoagulation therapy with 20,000 units of heparin | 216  
    anaerobic cultures positive for Gram-negative pleomorphic bacilli | 216  
    identified as Fusobacterium necrophorum | 216  
    minimal inhibitory concentrations of 0.094 to 0.004 mg/L | 216  
    highly susceptible to penicillin | 216  
    amoxicillin | 216  
    ceftriaxon | 216  
    metronidazole | 216  
    operative drainage of the left tonsillary abscess delayed by 5 days | 216  
    thrombocytopenia | 216  
    progressive brain abscess in the right temporal lobe | 216  
    switched to ceftriaxon and metronidazole | 216  
    mycotic aneurysm in the right internal carotid artery | 216  
    transferred to neurosurgical intensive care unit | 216  
    intensive anti-coagulation therapy with heparin | 216  
    thromboses in the IJV | 216  
    thromboses in the cavernous sinus | 216  
    thromboses in the ophthalmic vein | 216  
    cranial nerve palsy | 216  
    persisted during the first two weeks | 216  
    discharged from the hospital | 216  
    discrete residual sign of an abducens nerve paralysis on both sides | 216  
    emphasis on the right side | 216  
    oculomotor nerve paralysis on the right side had completely disappeared | 216  
    no other complications | 216  
    Lemierre's syndrome | 216  
    acute bacterial pharyngitis | 216  
    oropharyngeal infection | 216  
    ipsilateral thrombophlebitis | 216  
    thrombosis in the ipsilateral internal jugular vein | 216  
    infection in the lateral parapharyngeal cavity | 216  
    hematogenic or lymphogenic connection | 216  
    thrombosis in the IJV | 216  
    septic dissemination | 216  
    abscesses in the lung | 216  
    abscesses in the bone | 216  
    abscesses in the joints | 216  
    abscesses in the soft tissues | 216  
    abscesses in the brain | 216  
    abscesses in the eyes | 216  
    abscesses in the cardiovascular system | 216  
    paresis of the oculomotor and abducens nerve | 216  
    impairment of the sixth and twelfth cranial nerves | 216  
    clival syndrome | 216  
    isolated paresis of the sixth cranial nerve | 216  
    meningitis | 216  
    evaluation of the IJV thrombosis | 216  
    contrast-assisted computed tomography | 216  
    MRI | 216  
    ultrasound | 216  
    imaging investigation of the lung | 216  
    computed tomography | 216  
    septic emboli in the lung | 216  
    absence of clinical symptoms like cough or sputum | 216  
    MRI investigation of the brain | 216  
    timely identification of abscesses | 216  
    intracranial venous thromboses | 216  
    uncharacteristic symptoms | 216  
    paresis of the abducens and oculomotor nerves | 216  
    interdisciplinary basis | 216  
    minimize the delay until the establishment of the diagnosis | 216  
    institution of therapy | 216  
    avoid any catastrophic or lethal outcome | 216  
    primary ophthalmological symptoms | 216  
    conflict of interest | 216  
    drooping right eyelid | 216  
    exophthalmos on the right side | 216  
    thrombosis in the cavernous sinus | 216  
    thrombosis in the superior ophthalmic vein | 216  
    intra-axial brain abscess in the right temporal lobe | 216  
    worsened rapidly despite treatment with a broad-spectrum antibiotic | 216  
    tonsillary abscess on the left side | 216  
    maximum diameter of 1.3 cm | 216  
    numerous septic emboli in both lungs | 216  
    mycotic aneurysm in the right internal carotid artery | 216  
    adjacent to the previously thrombosed cavernous sinus | 216  
    