56 years old | 0
woman | 0
presented to the emergency department | 0
high-grade fever | -48
shortness of breath | -48
ill-appearing | 0
hypotensive | 0
tachycardic | 0
tachypneic | 0
mottled cold extremities | 0
chest radiogram | 0
CT scan | 0
multilobar pneumonia | 0
laboured breathing | 0
hypotension | 0
intubated | 0
transferred to the medical Intensive care unit | 0
fluid resuscitation | 0
required intravenous norepinephrine | 0
vasopressin | 0
dopamine | 0
haemodynamic support | 0
blood cultures obtained | 0
intravenous vancomycin | 0
ceftriaxone | 0
azithromycin | 0
prolonged prothrombin time | 0
prolonged partial thromboplastin time | 0
elevated fibrin degradation products | 0
disseminated intravascular coagulopathy (DIC) | 0
positive urine Streptococcus pneumonia antigen | 0
blood cultures grew Streptococcus pneumoniae | 0
diffuse petechial rash | 72
non-blanching purpuric ecchymotic skin lesions | 72
flaccid bullae | 72
extensive skin sloughing off | 72
skin biopsy | 72
non-inflammatory vascular occlusion | 72
skin necrosis | 72
purpura fulminans (PF) | 72
14-day course of broad-spectrum antibiotics | 0
heparin drip | 0
blood products | 0
inadequate response to therapies | 72
hyperbaric oxygen therapy instituted | 72
hyperbaric oxygen therapy stopped | 312
anuric renal failure | 72
required haemodialysis | 72
bedside incisional fasciotomy | 72
no evidence of muscle necrosis | 72
no compartment syndrome | 72
transferred to the burns unit | 72
75% skin loss | 72
prolonged hospital stay | 0
dismal prognosis | 0
lack of meaningful recovery | 0
shared decision to pursue comfort measures only | 0
