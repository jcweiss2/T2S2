83 years old | 0
male | 0
admitted to the hospital | 0
fall | -12
syncope | -12
lying on the floor throughout the night | -12
leg ecchymosis | 0
anuria | 0
rhabdomyolysis-induced AKI | 0
septic state | 0
acute prostatitis | -12
increased urea (140 mg/dL) | 0
increased creatinine (7.96 mg/dL) | 0
increased myoglobin (15,560 ng/mL) | 0
increased CPK (124,841 U/L) | 0
increased LDH (1,199 U/L) | 0
increased CRP (53.6 mg/dL) | 0
increased procalcitonin (505.3 ng/mL) | 0
increased total bilirubin (7.53 mg/dL) | 0
increased direct bilirubin (4.24 mg/dL) | 0
increased AST (749 U/L) | 0
increased ALT (410 U/L) | 0
increased PSA (662 ng/mL) | 0
increased white blood cell count (26,460 cells/µL) | 0
increased neutrophils (93%) | 0
sodium 137 mEq/L | 0
potassium 4.9 mEq/L | 0
calcium 8.7 mg/dL | 0
albumin 2.6 g/dL | 0
phosphate 4.1 mg/dL | 0
blood pressure 105/75 mm Hg | 0
heart rate 110 bpm | 0
body temperature 37.4°C | 0
no hydronephrosis | 0
empty bladder | 0
traces of blood in bladder catheter | 0
no previous renal impairment | -24
serum creatinine 0.8 mg/dL | -24
prostatic hypertrophy (prostate volume: 190 mL) | -24
PSA 9.9 ng/mL | -24
overactive bladder | -24
recurrent prostatitis | -24
no statins use | -24
volume expansion | 0
diuretic | 0
alpha-agonist | 0
antibiotic treatment | 0
furosemide 125 mg intravenous daily | 0
femoral central venous catheter placement | 0
HFR-Supra treatment | 0
ultrafiltration | 0
ultrafiltrate regeneration | 0
solute and volume removal | 0
myoglobin removal | 0
reduction of inflammatory status | 0
maintenance of fluid balance | 0
urine output 300 mL per 24 hours | 96
urine output 2,400 mL after 8 days | 168
furosemide tapered to 50 mg oral | 168
piperacillin/tazobactam | 0
meropenem | 24
E. coli resistant to piperacillin/tazobactam | 24
significant reduction in myoglobin (98.4%) | 144
significant reduction in CPK (99.8%) | 144
significant reduction in LDH (72%) | 144
significant reduction in CRP (81%) | 144
significant reduction in PCT (98%) | 144
blood flow 250 mL/min | 0
endogenous ultrafiltrate flow 14 L per session | 0
ultrafiltration rate according to clinical status | 0
enoxaparin 4,000 IU bolus | 0
normalization of myoglobin | 144
improved signs of systemic inflammation | 144
renal failure not recovered | 144
femoral catheter removed | 144
right jugular central venous catheter placed | 144
HDF sessions | 144
high-flux hemodialysis sessions | 144
dialysis no longer required | 504
urine output 2,300 mL per day | 504
serum urea 96 mg/dL | 504
serum creatinine 3.06 mg/dL | 504
CRP 3.2 mg/dL | 504
total bilirubin 0.81 mg/dL | 504
AST 27 IU/L | 504
ALT 25 IU/L | 504
PSA 61 ng/mL | 504
white blood cells 6,300 cells/µL | 504
hospitalization length 21 days | 504
urea 89 mg/dL | 3024
creatinine 2.41 mg/dL | 3024
GFR (CKD8-EPI) 24 mL/min | 3024
chronic kidney disease | 3024
maladaptive renal repair | 3024
