70 years old | 0\
male | 0\
farmer | 0\
admitted to the emergency department | 0\
high-grade fever | -120\
generalized body ache | -120\
headache | -120\
altered sensorium | -24\
joint pains | -120\
epigastric pain | -120\
inguinal lymphadenopathy | 0\
mild generalized rash | 0\
no eschar | 0\
hemodynamically stable | 0\
disoriented | 0\
no focal neurological deficit | 0\
no neck rigidity | 0\
acute febrile illness with undifferentiated fever | 0\
malaria | -120\
dengue | -120\
typhoid | -120\
leptospira | -120\
Scrub typhus antigen card | 0\
Scrub immunoglobulin M (IgM) | 0\
leukocytosis | 0\
mild hyperbilirubinemia | 0\
transaminitis | 0\
slightly raised international normalized ratio | 0\
negative for hepatitis B antigen | 0\
negative for hepatitis C antibody | 0\
mild fatty infiltration of the liver | 0\
tablet doxycycline 100 mg twice daily | 0\
defervescence | 48\
orientation improved | 48\
weakness of both lower limbs | 96\
weakness of both upper limbs | 96\
absent deep tendon reflexes | 96\
flexor plantar responses | 96\
bladder incontinence | 96\
no bowel incontinence | 96\
breathing difficulty | 96\
respiratory distress | 96\
intubated | 96\
mechanical ventilation | 96\
MRI of the brain | 96\
MRI of the cervical spine | 96\
nerve conduction velocity | 96\
motor sensory demyelinating polyneuropathy | 96\
intravenous immunoglobulin therapy | 96\
tablet rifampicin 600 mg twice daily | 96\
improvement in weakness | 120\
improvement in respiratory parameters | 120\
weaned off and extubated from the ventilator | 216\
oral feeding | 216\
aggressive limb and chest physiotherapy | 216\
shifted out from ICU | 216\
discharged from the hospital | 672\
full neurological recovery | 672