41 years old | 0
female | 0
history of untreated hypertension | -672
morbid obesity | -672
chronic back pain | -672
IVDU | -672
2 weeks of worsening low back pain | -336
diffuse abdominal pain | -336
lower extremity weakness | -336
anorexia | -336
fever | -336
chills | -336
shortness of breath | -336
dizziness | -336
constipation | -336
recent use of acetaminophen | -336
recent use of gabapentin | -336
recent use of hydrocodone | -336
recent use of methamphetamines | -336
recent use of marijuana | -336
admitted to the hospital | 0
blood pressure of 79/53 mmHg | 0
heart rate of 149 bpm | 0
lactic acid of 4.2 mg dl-1 | 0
WBC 37 500 ul-1 | 0
erythrocyte sedimentation rate 75 mm h-1 | 0
urine toxicology was positive for cannabis | 0
urine toxicology was positive for amphetamines | 0
midline tenderness of the lumbar spine | 0
3/5 strength in bilateral lower extremities | 0
bilateral shoulder warmth | 0
bilateral shoulder erythema | 0
bilateral shoulder tenderness | 0
limited range of motion | 0
multiple needle puncture sites on the antecubital fossas bilaterally | 0
puncture wounds on the right foot | 0
blood cultures were collected | 0
empirically started on vancomycin | 0
empirically started on metronidazole | 0
empirically started on aztreonam | 0
empirically started on IV fluids | 0
MRSA bacteraemia | 0
vancomycin with an MIC of 1 mg l-1 | 24
rifampin with MIC of ≤1 mg l-1 | 24
levofloxacin with MIC of ≤1 mg l-1 | 24
clindamycin with MIC of ≤0.5 mg l-1 | 24
daptomycin with MIC of ≤0.5 mg l-1 | 24
linezolid with MIC of 2 mg l-1 | 24
bilateral shoulder plain radiographs showed no abnormalities | 24
arthrocentesis of the AC joints showed WBC of 93 137 ul-1 | 24
arthrocentesis of the AC joints showed WBC of 32 043 ul-1 | 24
arthrocentesis of the AC joints grew MRSA | 24
surgical debridement of the shoulders | 48
intubated | 48
MRI of the lumbar spine showed L3-L5 osteomyelitis | 48
MRI of the lumbar spine showed facet septic arthritis | 48
MRI of the lumbar spine showed dorsal paraspinous myositis | 48
MRI of the lumbar spine showed L2-L5 epidural abscess | 48
MRI of the lumbar spine showed bilateral psoas myositis | 48
MRI of the lumbar spine showed bilateral psoas abscesses | 48
MRI of the bilateral shoulders after debridement showed septic arthritis of the AC joints | 48
MRI of the bilateral shoulders after debridement showed right distal trapezius abscess | 48
MRI of the bilateral shoulders after debridement showed left supraclavicular abscess | 48
MRI of the brain showed no acute intracranial processes | 48
TTE was negative for any valvular vegetations | 48
cardiology deferred acquiring a transoesophageal echocardiogram | 48
repeat surgical debridement of the shoulders | 72
neurosurgery evaluated the patient for possible debridement of the epidural abscess | 72
recommended medical management | 72
leukocytosis continued to rise | 72
peaked at 52 100 ul-1 | 72
trough levels of vancomycin were being monitored | 72
repeat blood cultures continued to be positive for MRSA | 72
antibiotics were escalated to daptomycin | 240
antibiotics were escalated to ceftaroline | 240
blood cultures ultimately became negative | 336
rifampin was added | 336
required critical care | 336
repeat MRI of the lumbar spine showed worsening epidural abscess | 432
neurosurgery took the patient for surgical drainage with drain placement | 432
intraoperative wound cultures were positive for MRSA | 432
intraoperative wound cultures were positive for Proteus mirabilis | 432
improved clinically | 432
all drains were removed | 432
discharged | 672
prescribed oral levofloxacin | 672
prescribed oral rifampin | 672