70 years old | 0
male | 0
jaundice | -1344
repeated vomiting | -1344
total serum bilirubin 5.7 mg/dl | 0
direct bilirubin 4.7 mg/dl | 0
INR 1.2 | 0
normal ALT | 0
normal AST | 0
normal serum electrolytes | 0
normal serum creatinine | 0
ultrasound abdomen | 0
hepatomegaly | 0
dilated intrahepatic biliary channels | 0
dilated extrahepatic biliary channels | 0
no cirrhosis of liver | 0
no portal hypertension | 0
hypo-echoic lesion in head of pancreas | 0
contrast enhanced computed tomography (CECT) scan | 0
soft tissue mass head of pancreas | 0
haziness of fat planes between mass and stomach | 0
free superior mesenteric artery | 0
free portal vein | 0
free superior mesenteric vein | 0
mildly dilated stomach | 0
enlarged supra-pancreatic lymph nodes | 0
enlarged peri-portal lymph nodes | 0
no distant metastasis | 0
cancer head of pancreas | 0
possibility of gastric wall invasion | 0
surgical intervention | 0
preoperative plan pancreaticoduodenectomy | 0
evaluated by cardiac physician | 0
evaluated by pulmonary physician | 0
evaluated by anesthesia physician | 0
found fit for surgery | 0
intraoperative finding similar to preoperative imaging | 0
dissection of supra-pancreatic lymph nodes | 0
common hepatic artery injured | 0
repair with Proline 8/0 | 0
intraoperative Doppler on hepatic artery | 0
normal flow hepatic artery | 0
RI 0.6 | 0
PSV 100 cm/s pre anastomotic | 0
PSV 125 cm/s post anastomotic | 0
SAT 71 ms | 0
pyloric preserving pancreaticoduodenectomy | 0
admitted to Intensive care | 0
postoperative day one | 24
stable | 24
Doppler on hepatic artery | 24
no detectable flow hepatic artery | 24
ALT 1278 U/L | 24
AST 973 U/L | 24
CECT | 24
completely thrombosed common hepatic artery | 24
no detected contrast beyond repair site | 24
intrahepatic small accessory left hepatic artery | 24
hardly detectable middle hepatic artery | 24
arising from left gastric artery | 24
decision to follow patient | 24
ALT starts to decrease | 48
AST starts to decrease | 48
bilirubin starts to decrease | 48
gradual improvement of liver function parameters | 48
shifted from ICU to ward | 72
Doppler on hepatic artery | 72
no flow in hepatic artery | 72
ALT 137 U/L | 240
AST 34 U/L | 240
total bilirubin 1.3 mg/dl | 240
discharged | 240
follow up two weeks later | 624
normalization of liver function tests | 624
non-detectable hepatic artery flow | 624
no significant complaint | 624
follow up six months later | 4320
normal lab parameters | 4320
CECT scan | 4320
completely thrombosed hepatic artery | 4320
small accessory left hepatic artery | 4320
hardly detectable middle hepatic artery | 4320
no liver infarction | 4320
no abscess | 4320
no biliary complications | 4320
