7 years old | 0
male | 0
admitted to the hospital | 0
fever | -72
coughing | -72
pain in the legs | -72
dysesthesia | -72
waddling gait | -72
sister had flu-like syndrome | -168
symptomatic treatment | -72
aggravations | -72
deterioration of general state | -72
abdominal pain | -72
food intolerance | -72
acute respiratory failure | -72
tachycardia | 0
normal blood pressure | 0
respiratory retraction | 0
abdominal breathing | 0
diffuse rhonchi | 0
severe hypoxemia | 0
noninvasive ventilation | 0
high-flow oxygen therapy | 0
chest X-ray showed interstitial pneumonia | 0
transferred to pediatric intensive care unit | 0
chest X-ray control showed right basal consolidation | 24
dribble on the way to hospital | -72
probable aspiration | -72
neurological deterioration | 48
agitation | 48
bilateral mydriasis | 48
intubation | 48
sedation | 48
mechanical ventilation | 48
neurological manifestations progressed | 72
bulbar and peripheral motor deficit | 72
upper limb weakness | 72
central involvement | 72
normal consciousness | 72
no spontaneous movements of arms and legs | 72
dysfunctions in cranial nerves | 72
facial diplegia | 72
bilateral ptosis | 72
mydriasis | 72
severe swallowing disorders | 72
absence of cough | 72
tetraparesia | 72
hyperreflexia | 72
areflexia | 96
dysautonomia | 72
vascular fillings | 72
Mycoplasma pneumonia | 0
Haemophilus influenza | 0
inflammatory signs | 0
increased C-reactive protein | 0
procalcitonin | 0
toxicology studies negative | 0
microbiological tests negative | 0
immune tests normal | 0
cerebrospinal fluid examinations normal | 48
antiganglioside and antigalactocerebroside antibodies negative | 48
cerebral tomography scan normal | 48
cerebromedullar magnetic resonances normal | 120
ultrasonography showed phrenic paresia | 504
electroencephalogram normal | 48
sensitive evoked potentials normal | 456
electromyogram showed axonal motor polyneuropathy | 192
intravenous immunoglobulin treatment | 120
second course of immunoglobulin | 432
recovery started | 504
mechanical ventilation necessary for 48 days | 0
tracheostomy performed | 696
enteral feeding for 18 weeks | 0
salt supplementation | 0
speech and oral intake improved | 504
intensive functional and psychotherapeutic rehabilitation | 504
patient left hospital after 11 weeks | 840
examination after 20 weeks showed proximal weakness | 1200
decreased upper limb deep tendon reflexes | 1200
walking was fluid | 1200
no breathing or swallowing troubles | 1200
electromyogram showed improvements | 1200
tracheostomy and gastrostomy removed after 5 months | 2160
last examination showed discrete hypotonia | 8760
fine motor skill difficulties | 8760
fatigability | 8760
intermittent hand tremors | 8760
deep tendon reflexes normal | 8760
electromyogram still improving | 8760