84 years old | 0
    male | 0
    admitted to the emergency department | 0
    febrile | -24
    encephalopathic | -24
    melanotic stool | -24
    cerebrovascular accident | -8760
    residual left hemiparesis | -8760
    gastrointestinal bleed | -8760
    hypertension | -8760
    hyperlipidemia | -8760
    gastroesophageal reflux disease | -8760
    diverticular disease | -8760
    depression | -8760
    benign prostatic hypertrophy | -8760
    chronic iron deficiency anemia | -8760
    immobility | -8760
    heart rate 92 | 0
    blood pressure 95/51 | 0
    obtunded | 0
    acute anemia | 0
    acute renal failure | 0
    procalcitonin 14 ng/mL | 0
    stool heme-positive | 0
    dry mucous membranes | 0
    non-tender abdomen | 0
    non-distended abdomen | 0
    no evidence of skin changes | 0
    no evidence of infection | 0
    volume resuscitation | 0
    broad spectrum antibiotics initiated | 0
    admitted to ICU | 0
    presumed gastrointestinal bleed | 0
    presumed sepsis of unknown etiology | 0
    elevated lactic acid | 0
    hypotension | 0
    gastroenterology consultation | 0
    endoscopy deferred | 24
    no continued evidence of active bleeding | 24
    laboratory values normalized | 24
    hemodynamics normalized | 24
    returned to baseline mental status | 24
    no history of weight loss | -8760
    no history of decreased appetite | -8760
    no recurrent melanotic stool | -8760
    no alterations in bowel habits | -8760
    right hip erythema | 24
    right hip induration | 24
    right hip pain | 24
    no crepitus | 24
    CT right hip concern for necrotizing soft tissue infection | 24
    gas involving right retroperitoneum | 24
    gas involving upper thigh | 24
    no evidence of abscess | 24
    general surgery consultation | 24
    necrotizing fasciitis consultation | 24
    operative intervention declined | 24
    clinical improvement with non-operative treatment | 32
    CT abdomen and pelvis | 56
    7.1 cm proximal right colon mass | 56
    invasion into retroperitoneum | 56
    gas tracking into adjacent soft tissues | 56
    concerning perforated malignancy | 56
    colorectal surgery consultation | 56
    tumor resection with debridement discussed | 56
    widespread soft tissue infection | 56
    palliative care elected | 56
    transitioned to hospice care | 56
    expired | 240
    <|eot_id|>
    