48 years old | 0
    female | 0
    presented for an elective outpatient ERCP | 0
    evaluation of sphincter of Oddi dysfunction | 0
    recent acute pancreatitis | 0
    episodic abdominal pain | 0
    common bile and pancreatic ducts cannulated | 0
    basal sphincter pressures measured | 0
    cholangiography | 0
    pancreatography | 0
    cystic duct cannulated | 0
    cholecystokinin infusion | 0
    bile aspirated | 0
    microlithiasis analysis | 0
    no immediate complications | 0
    mild post-procedure discomfort | 0
    admitted to the hospital | 0
    developed chest pain | 24
    blood work revealed white blood cell count of 14.5 × 1,000/μL | 24
    hematocrit 32.9% | 24
    aspartate aminotransferase (AST) 176 U/L | 24
    alanine aminotransferase (ALT) 32 U/L | 24
    total bilirubin 0.46 mg/dL | 24
    serum lipase 93 U/dL | 24
    serum troponin 2.3 ng/mL | 24
    cardiology evaluation requested | 24
    non-ST elevation myocardial infarction | 24
    treated medically | 24
    developed abdominal pain with peritoneal signs | 24
    AST 250 U/L | 24
    ALT 55 U/L | 24
    total bilirubin 3.34 mg/dL | 24
    direct bilirubin 2.85 mg/dL | 24
    lipase of 192 U/dL | 24
    computerized tomography (CT) scan of the abdomen | 24
    large amount of air within and around the gallbladder | 24
    extensive free air in lesser sac, retroperitoneum, intraperitoneal cavity, and bile duct | 24
    loculated area of air in posterior segment of the right hepatic lobe | 24
    presumptive diagnosis of emphysematous cholecystitis | 24
    suspicion of bowel perforation | 24
    started on broad spectrum antibiotics (ampicillin/sulbactam) | 24
    laparotomy performed | 48
    completely gangrenous gallbladder | 48
    no evidence of bowel perforation | 48
    cholecystectomy performed | 48
    no gallstones present | 48
    common bile duct (CBD) without any abnormalities | 48
    common hepatic duct (CHD) markedly inflamed with possible gangrene | 48
    histopathologic examination of the gallbladder revealed gangrenous cholecystitis | 48
    gram-positive rods invading the gallbladder wall | 48
    cultures from the gallbladder and blood grew Clostridium perfringens | 48
    discharged home | 336
    presented with abdominal pain and fever | 432
    abdominal CT scan | 432
    two large abscesses in liver | 432
    percutaneous drainage catheters placed | 432
    left lobe abscess drained bilious fluid | 432
    cholangiography via percutaneous drain | 432
    communication of left lobe abscess with left intrahepatic biliary system | 432
    extravasation of contrast in peribiliary area | 432
    disruption and necrosis of intrahepatic ducts | 432
    CHD and CBD demonstrated necrosis and infarction | 432
    intramural tracking of contrast | 432
    trans-hepatic 8F locking loop draining catheter placed | 432
    continued on antibiotics and supportive measures | 432
    CHD drain exchanged for internal external percutaneous drain | 504
    discharged home | 504
    presented to emergency room with worsening abdominal pain and fever | 672
    serum creatinine 3.5 mg/dL | 672
    leukocytosis of 20,000/μL | 672
    required treatment of septic shock | 672
    broad spectrum antibiotics | 672
    supportive measures | 672
    revision of biliary drain catheters | 672
    recurrent hospital admissions due to cholangitis | 2160
    recurring hepatic abscesses | 2160
    sepsis with Enterococcus, Pseudomonas, Klebsiella, and Candida | 2160
    severe hypotension | 2160
    renal failure | 2160
    respiratory failure | 2160
    managed by percutaneous drains, antibiotics, and supportive care | 2160
    ERCP done 15 months after index ERCP | 10800
    multiple strictures and beading in intraEand extraEhepatic biliary tree | 10800
    hepatic abscesses resolved | 10800
    biliary strictures required management | 10800
    placement and exchange of biliary stents every 3 months | 10800
    evidence of progressive sclerosing cholangitis | 10800
    developed end-stage liver disease | 10800
    underwent successful living donor liver transplantation | 21600
    explant histopathology revealed secondary biliary cirrhosis | 21600
    bile duct necrosis | 21600
    fungal hyphae | 21600
    bacterial organisms | 21600
    maintained normal hepatobiliary function | 21600
    feeling well in 3 years of follow-up after liver transplantation | 21600