4 years old | 0
intact male | 0
Golden retriever | 0
admitted to the hospital | 0
abdominal distention | -72
melena | -72
lethargy | -72
anorexia | -72
azotemia | -72
hypoalbuminemia | -72
hydroxyethyl starch administration | 0
increased plasma osmolality | 0
6% hydroxyethyl starch 130/0.4 solution | 0
10 ml/kg, IV, bolus | 0
increased creatinine level | 168
proteinuria | 168
deteriorating azotemia | 168
deteriorating proteinuria | 168
referred to the Veterinary Medical Teaching Hospital | 336
severe azotemia | 336
ascites | 336
gastrointestinal bleeding | 336
normothermic | 336
normal heart rate | 336
normal respiratory rate | 336
hypertensive | 336
ecchymosis | 336
distended abdomen | 336
microcytic non-regenerative anemia | 336
neutrophilia | 336
thrombocytopenia | 336
hypoalbuminemia | 336
hypoproteinemia | 336
hyperbilirubinemia | 336
increased alkaline phosphatase | 336
increased gamma glutamyl transferase activity | 336
increased fasting bile acid | 336
mild increased activated partial thromboplastin | 336
metabolic acidosis | 336
hyponatremia | 336
hyperkalemia | 336
hypocalcemia | 336
anuria | 336
euthanized | 360
necropsy | 360
multifocal nodules on the liver surface | 360
petechial-to-ecchymotic hemorrhages in the heart | 360
gastrointestinal bleeding | 360
degeneration of the kidney cortex | 360
multiple hepatic nodules surrounded by thick fibrous septa | 360
moderate multiple calcium depositions in the necrotic areas | 360
severe multiple linear renal tubular necrosis | 360
moderate glomerular injury | 360
osmotic nephrosis lesions | 360
acute kidney injury | 168
liver cirrhosis | 360
platelet dysfunction | 336
uremic toxin production | 336
decreased liver function | 360
insufficient removal of HES molecules | 360
accelerated renal function impairment | 360