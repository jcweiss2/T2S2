31 years old | 0 | 0 
female | 0 | 0 
non-smoking | 0 | 0 
Caucasian | 0 | 0 
no past medical history | 0 | 0 
admitted to the hospital | 0 | 0 
sudden-onset severe headache | -840 | -840 
left arm numbness | -840 | -840 
cranial computed tomography (CT) scan | -840 | -840 
grade 2 (Hunt and Hess scale) SAH | -840 | -840 
no prior history of head injury | 0 | 0 
uncomplicated pregnancy | 0 | 0 
uncomplicated vaginal delivery | 0 | 0 
digital subtraction angiography (DSA) | -720 | -720 
ruptured right middle cerebral artery aneurysm | -720 | -720 
percutaneous endovascular coil embolization | -720 | -720 
no permanent neurological deficits | -720 | 0 
fever | -504 | -504 
chills | -504 | -504 
constant abdominal pain | -504 | -504 
purulent uterine discharge | -504 | -504 
no urinary symptoms | -504 | -504 
no respiratory symptoms | -504 | -504 
blood culture | -504 | -504 
piperacillin/tazobactam | -504 | -480 
vancomycin | -504 | -480 
azithromycin | -504 | -480 
sepsis | -480 | -480 
septic shock | -480 | -480 
transferred to intensive care unit | -480 | -480 
body temperature 38.3 °C | -480 | -480 
invasive blood pressure 90/65 mmHg | -480 | -480 
heart rate 135/min | -480 | -480 
arterial oxygen saturation 82 % | -480 | -480 
mild disorientation | -480 | -480 
slower capillary refill | -480 | -480 
coarse rales | -480 | -480 
sequential organ failure assessment (SOFA) score 4 | -480 | -480 
hemoglobin 6.8 g/dL | -480 | -480 
d-dimers 4.58 μg/mL | -480 | -480 
C-reactive protein 322 mg/L | -480 | -480 
fibrinogen concentration 6.4 mL | -480 | -480 
E. coli sensitive to piperacillin/tazobactam | -480 | -480 
chest radiography | -480 | -480 
pulmonary nodules | -480 | -480 
CT of the thorax | -480 | -480 
transvaginal ultrasound | -480 | -480 
enlarged uterus | -480 | -480 
complete loss of zonal anatomy | -480 | -480 
abdominal magnetic resonance imaging (MRI) | -480 | -480 
heterogenous myometrial mass | -480 | -480 
splenic metastatic lesion | -480 | -480 
serum β-human chorionic gonadotrophin (β-hCG) 232,085 mUI/mL | -480 | -480 
suction evacuation and curettage | -480 | -480 
choriocarcinoma diagnosis | -480 | -480 
International Federation of Gynecology and Obstetrics (FIGO) modified WHO prognostic scoring system | -480 | -480 
total score 12 | -480 | -480 
high risk of developing resistance to single-drug chemotherapy | -480 | -480 
multiagent chemotherapy regimen | -480 | -480 
low-dose etoposide | -480 | -456 
cisplatin | -480 | -456 
EMA/CO regimen | -456 | -168 
etoposide | -456 | -168 
methotrexate | -456 | -168 
actinomycin D | -456 | -168 
cyclophosphamide | -456 | -168 
vincristine | -456 | -168 
β-hCG levels plateaued | -168 | -168 
restaging with MRI of the brain | -168 | -168 
18F-fluorodeoxyglucose (FDG) positron emission tomography (PET)/CT scan | -168 | -168 
decreased pulmonary nodules | -168 | -168 
decreased uterine mass | -168 | -168 
low standardized uptake value (SUV) | -168 | -168 
revised FIGO score 7 | -168 | -168 
EP/EMA regimen | -168 | 0 
normalization of β-hCG | 0 | 0 
grade 3 neutropenia | -336 | -336 
granulocyte colony stimulating factor (G-SCF) | -336 | -336 
dose reduction of etoposide | -336 | -336 
dose reduction of actinomycin D | -336 | -336 
grade 2 alopecia | -336 | 0 
grade 2 nausea | -336 | 0 
dexamethasone | -336 | 0 
ondansetron | -336 | 0 
grade 2 fatigue | -168 | 0 
male condoms | 0 | 720 
follow-up | 0 | 720 
alive 21 months post diagnosis | 720 | 720