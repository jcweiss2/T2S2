18 years old | 0
male | 0
morbidly obese | 0
diabetes | 0
end-stage renal disease | 0
hemodialysis | 0
peripheral vascular disease | 0
left below knee amputation | 0
right above knee amputation | 0
right extra anatomical axillobifemoral bypass graft | 0
presented to emergency department | 0
right-sided abdominal pain | -48
vomiting | -48
fever | -48
conscious | 0
alert | 0
oriented | 0
pale and sick | 0
temperature 37.8°C | 0
blood pressure 150/90 mmHq | 0
oxygen saturation 95% | 0
abdomen distended and tympanic | 0
right upper quadrant and right flank tenderness | 0
total leukocyte count 20 × 10^3 | 0
hemoglobin 10.7 gm% | 0
acidotic | 0
pH 7.33 | 0
end-stage renal disease | 0
chest X-ray showing gas under the right hemi-diaphragm | 0
perforated viscous | 0
CT scan with contrast | 0
right perinephric collection with extension into the right sub-phrenic region | 0
gas in the right collecting system and urinary bladder | 0
no gas in the renal parenchyma | 0
right atrial thrombus | 0
started on parenteral antibiotics | 0
admitted to intensive care unit | 0
percutaneous drainage | 0
failed percutaneous drainage | 0
trial of percutaneous drainage | -24
open drainage of a very thick, foul smelly, loculated perinephric and sub-phrenic collection | -24
epidural anesthesia and sedation | -24
very abnormal bladder mucosa with multiple cystic lesions with air “bubbles” | -24
ureteric Double J stent inserted in the right ureter | -24
urethral catheter to drain the bladder | -24
culture of the collection showed Klebsiella pneumonia extended-spectrum β-lactamase | -24
severe sepsis and multiple organ failure | -48
died | -48