Mayer-Rokitansky-Küster-Hauser syndrome | 0
primary amenorrhea | 0
sigmoid neovaginoplasty | -9 years
lower abdominal pain | 0
bilateral pelvic pain | 0
no routine irrigation or dilation of neovagina | 0
penetrative sexual intercourse every couple of weeks | 0
no intercourse in a few months | 0
CT imaging of the abdomen | 0
tubular, heterogenous, fluid-filled structure | 0
abdominal pain acutely worsened | 24
diaphoresis | 24
significant distress due to pain | 24
leukocytosis | 24
absolute neutrophils | 24
empiric intravenous piperacillin-tazobactam | 24
transfer to hospital | 24
hypotensive | 24
tachycardic | 24
afebrile | 24
tachypneic | 24
oxygen saturation | 24
IV fluid boluses | 24
antimicrobials changed to IV ceftriaxone, IV vancomycin, and IV metronidazole | 24
exploratory laparotomy | 24
cystoscopy | 24
vaginoscopy | 24
normal bladder and urethra | 24
obliterated introitus | 24
diffuse intra-abdominal spillage of mucus | 24
perforated sigmoid neovagina | 24
purulent fluid drained | 24
intrabdominal drains placed | 24
intubated | 24
mechanical ventilation | 24
septic shock | 24
vasopressor agents | 24
antimicrobials changed to IV cefepime, IV vancomycin, and IV metronidazole | 24
peritoneal culture growing gram-negative rods | 24
blood cultures negative | 24
peritoneal cultures finalized to Bacterioides thetaioaomicron, Bacterioides caccae, and Actinomyces species | 168
antimicrobials changed to IV piperacillin-tazobactam | 168
weaned off vasopressors | 192
extubated | 192
transferred to general floor | 288
Infectious Diseases team consulted | 288
discharged home | 360
abdominal wound vacuum | 360
IV piperacillin-tazobactam for four weeks | 360
readmitted with sepsis | 504
generalized malaise | 504
diffuse abdominal pain | 504
white blood count | 504
absolute neutrophil count | 504
d-dimer | 504
lactate | 504
CT of chest, abdomen and pelvis | 504
bilateral pleural effusions | 504
loculated left pleural effusion | 504
multiple new abdominal abscesses | 504
transcutaneous drainage catheter in pelvis | 504
open anterior midline wound with wound vacuum | 504
hypoxemia | 504
transferred to ICU | 504
IV piperacillin-tazobactam continued | 504
placement of right perihepatic drain | 504
aspiration of purulence | 504
unsuccessful drainage of peri-splenic collection | 504
blood cultures negative | 504
interventional radiology reconsulted | 504
drainage of right perinephric abscess | 504
drainage of perisplenic abscess | 504
broad-spectrum PCR sent | 504
antimicrobials narrowed to IV ampicillin-sulbactam | 768
discharged | 768
broad spectrum PCR positive for Gleimia europaea, Alistipes onderdonkil, Varibaculum timonense, and Jonquetella anthropi | 768
follow-up at adult infectious diseases clinic | 1056
improved clinically | 1056
repeat CT abdomen | 1056
transitioned to oral amoxicillin-clavulanate | 1056
complete resolution of abscesses | 1056