46 years old | 0
male | 0
kidney transplantation | -1044
Basiliximab | -1044
tacrolimus | -1044
mycophenolic acid | -1044
prednisone | -1044
creatinine level 1.13 mg/dL | -84
productive cough | -72
diarrhea | -72
amoxicillin/clavulanic acid therapy | -72
MPA dose reduction | -72
MPA dose reduction | -69
Azithromycin | -69
reverse transcription polymerase chain reaction assay | -66
SARS-CoV-2 RNA positive | -66
admitted to the hospital | -66
body temperature 38.8°C | -66
persistent cough | -66
persistent diarrhea | -66
ill-defined left basal opacity | -66
right infra-hilar reticulonodular interstitial pattern | -66
leukocytopenia | -66
thrombocytopenia | -66
hypokalemia | -66
elevated C-reactive protein | -66
elevated lactate dehydrogenase | -66
MPA withdrawn | -66
Tac dose reduction | -66
hydroxychloroquine | -66
respiratory status deterioration | -60
renal function deterioration | -60
transferred to ICU | -60
marked dyspnea | -60
peripheral blood oxygenation 93% | -60
marked signs of dehydration | -60
diarrheic stool passage | -60
elevated acute phase reactants | -60
hyperleukocytosis | -60
thrombocytopenia | -60
raised D-dimers | -60
hypokalemia | -60
hyponatremia | -60
sepsis biomarkers negative | -60
no signs of hydronephrosis | -60
normal Doppler graft parameters | -60
hematuria | -60
proteinuria | -60
leukocyturia | -60
erythrocytes/field | -60
leucocytes/field | -60
COVID-19 pneumonia | -60
bacterial pneumonia | -60
intubation | -58
high-flow nasal cannula oxygen therapy | -58
respiratory rate 40/min | -58
O2 saturation 89% | -58
PaO2/FiO2 117 | -58
noninvasive mechanical ventilation | -56
oxygen therapy | -56
complete remission of respiratory insufficiency | -56
stage 3 acute kidney injury | -56
creatinine levels peak | -49
oliguria | -48
polyuria | -46
severe hyponatremia | -46
methylprednisolone | -46
methylprednisolone i.v. pulse therapy | -44
Tac reintroduced | -42
Tac dose increase | -38
discharged home | -36
hydroxychloroquine | -66
lopinavir/ritonavir | -66
broad-spectrum prophylactic antibacterial therapy | -66
antifungal therapy | -66
meropenem | -66
linezolid | -66
trimethoprim/sulfamethoxazole | -66
caspofungin | -66
transferred to pneumology unit | -42
discharged home | -36
creatinine level return to baseline | -35
Tac plasma level within target level | -36
prophylactic anticoagulation | -60
enoxaparin | -60