22 years old | 0
female | 0
multiparous | 0
pregnant | 0
24 week gestation | 0
altered consciousness | -1
vomiting | -1
bleeding per vaginum | -1
history of PV manipulation | -24
pale | 0
dehydrated | 0
tender and distended abdomen | 0
blood pressure 80/46 mm Hg | 0
heart rate 130/min | 0
respiratory rate 35/min | 0
Glasgow coma score 8 | 0
no neck rigidity | 0
reflexes normal | 0
gangrenous bowel loops protruding out from vagina | 0
gas under the diaphragm | 0
prolonged PR interval | 0
wide QRS complex | 0
peaked T wave | 0
rehydrated with normal saline | 0
invasive positive pressure ventilation | 0
Ryle's tube | 0
Foley's catheterization | 0
central venous cannulation | 0
midazolam infusion | 0
fentanyl infusion | 0
severe anaemia | 0
deranged renal functions | 0
metabolic acidosis | 0
hyperkalaemia | 0
hyponatraemia | 0
nebulised with salbutamol | 0
dextrose-insulin infusion | 0
unsafe abortion | -24
uterine perforation | -24
bowel perforation | -24
fluid replacement | 0
blood transfusion | 0
BP returned to 116/62 mm Hg | 2
emergency laparotomy | 2
general anaesthesia | 2
sudden hypotension | 2
cardiac arrest | 2
external cardiac massage | 2
colloid bolus | 2
inj adrenaline | 2
dopamine infusion | 2
revived after 2 minutes | 4
ketamine infusion | 4
nitrous oxide-oxygen combination | 4
neuromuscular blockade | 4
atracurium | 4
dead foetus extracted | 4
uterine perforation | 4
gangrenous bowel loops | 4
resection anastomosis | 4
subtotal hysterectomy | 4
end-colostomy | 4
blood transfusion | 4
fluid transfusion | 4
surgery lasted for 4 hours | 4
shifted to ICU | 4
SIMV mode | 4
dopamine infusion tapered | 24
extubated | 48
discharged | 240
no major organ failure | 240
no neurological deficit | 240