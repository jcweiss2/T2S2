66 years old| 0
    female | 0
    smoker | 0
    referred to emergency department | 0
    hypotension | 0
    colonoscopy | -504
    removal of two serrated polyps | -504
    generalized weakness | -336
    fatigue | -336
    blood pressure 60/30 mm Hg | -336
    sent to ED | -336
    confused | 0
    lethargic | 0
    fever | -120
    temperature 98.1 °F | 0
    blood pressure 74/45 mm Hg | 0
    heart rate 99 beats/min | 0
    respiratory rate 18 breaths/min | 0
    conjunctivae pink | 0
    no jaundice | 0
    lungs clear | 0
    heart sounds audible | 0
    no murmurs | 0
    no rubs | 0
    no gallops | 0
    abdominal tenderness | 0
    bilateral costovertebral angle tenderness | 0
    bowel sounds present | 0
    WBC count 28,700/mm3 | 0
    left shift | 0
    hemoglobin 8.3 g/dL | 0
    normal liver function | 0
    normal renal function | 0
    IV normal saline bolus | 0
    blood pressure 105/60 mm Hg | 0
    blood cultures obtained | 0
    urine cultures obtained | 0
    ceftriaxone | 0
    possible pyelonephritis | 0
    transferred to ICU | 0
    CT abdomen with contrast | 0
    intraabdominal abscess | 0
    hepatic abscess | 0
    perihepatic abscess | 0
    right lower quadrant abscess | 0
    interventional radiology consulted | 0
    surgery consulted | 0
    intraabdominal drains placed | 0
    pus drained | 0
    ceftriaxone discontinued | 0
    meropenem | 0
    vancomycin | 0
    metronidazole | 0
    pus culture | 72
    Streptococcus constellatus | 72
    meropenem discontinued | 72
    vancomycin discontinued | 72
    ceftriaxone restarted | 72
    metronidazole continued | 72
    alertness improved | 72
    appetite improved | 72
    abdominal tenderness decreased | 72
    WBC count improved | 168
    fluid drained less than 10 cc | 168
    repeat CT abdomen | 168
    abscess decreased | 168
    residual liver abscess | 168
    three drains removed | 168
    last drain removed | 336
    PICC placed | 336
    antibiotics for 6 weeks | 336
    discharged | 348
    nursing home | 348
    CT abdomen resolution | 672
    <|eot_id|>
    