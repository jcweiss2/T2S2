58 years old | 0
female | 0
Caucasian | 0
British | 0
admitted to the hospital | 0
found unresponsive | 0
complained of headache | -24
attended the ED with symptoms suggesting a urinary tract infection | -72
given unspecified oral treatment | -72
discharged | -72
mid-stream urine sample obtained | -72
reported as positive for E. coli | -72
Glasgow Coma Score of 6/15 | 0
right-sided weakness | 0
facial droop | 0
afebrile | 0
no neck stiffness | 0
myoclonic jerks in both arms | 0
anxiety | 0
treated with sertraline | 0
smoked approximately thirty cigarettes per day | 0
alcohol intake of seven units per day | 0
no recent history of travel | 0
no recent history of trauma | 0
no recent history of surgery | 0
intubated in the ED | 0
transferred to the Intensive Care Unit | 0
initial working diagnosis was of stroke | 0
ceftriaxone 2 grams 12-hourly started | 0
aciclovir 640 miligrams 12-hourly started | 0
blood tests on admission | 0
White cell count 9.8 109/L | 0
Neutrophils 8.8 109/L | 0
Lymphocytes 0.2 109/L | 0
Platelets 62 109/L | 0
C-reactive protein 643mg/L | 0
Creatinine 232 μmol/L | 0
Urea 19.7mmol/L | 0
CT of the brain showed signs of a left-sided middle cerebral artery infarct | 0
no hydrocephalus | 0
MRI of the brain showed a right internal capsule acute infarct | 0
debris in the ventricles suggestive of ventriculitis | 0
blood cultures taken | 0
reported as having grown E. coli | 24
lumbar puncture performed | 0
cerebrospinal fluid results | 0
White cell count 15 680 106/L | 0
Polymorphs 95% | 0
Lymphocytes 5% | 0
Turbid | 0
Red blood cells 220 106/L | 0
Protein 4.26g/L | 0
Glucose 0.4mmol/L | 0
Serum glucose 7.0mmol/L | 0
CSF gram-stain analysis revealed gram-negative organisms | 0
culture results were later reported as Escherichia coli | 24
unenhanced CT brain seven days after admission confirmed a recent right internal capsule infarct | 168
repeat LP on day 11 post-admission | 264
marked improvement | 264
no further bacterial growth | 264
mechanical ventilation for twenty-seven days | 0
sedation hold | 648
neurological examination | 648
marked left-sided hemiparesis | 648
ceftriaxone continued at the same dose and frequency until day 25 of admission | 0
dose reduced to 2 grams daily | 600
aciclovir stopped | 0
Strongyloides serology reported negative | 0
human immunodeficiency virus serology reported negative | 0
Hepatitis B serology reported negative | 0
Hepatitis C serology reported negative | 0
renal tract ultrasound showed no evidence of hydronephrosis or collection | 0
transthoracic echocardiogram reported as normal | 0
MRI brain with contrast on day 27 of hospital admission | 648
persistent features of ventriclitis | 648
subacute infarct in the right internal capsule | 648
trapped occipital horn of the right lateral ventricle | 648
tracheostomy performed | 648
decannulated in ICU | 696
stepped-down to the Stroke ward | 696
intensive physiotherapy and neuro-rehabilitation | 696
MRI brain on day forty-one post-admission | 984
mild reduction of a ring-enhancing lesion in the right lateral ventricle | 984
persistent ventricular debris | 984
discharged to a rehabilitation facility | 1392
follow-up imaging at four months | 2928
significant regression of the findings previously noted | 2928