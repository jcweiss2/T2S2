12-year-old | 0
boy | 0
trauma to right ankle | -72
pain in right ankle | -72
swelling in right ankle | -72
cough | -120
fever | -120
febrile (38.5°C) | 0
tachycardia (125/min) | 0
respiratory rate (25/min) | 0
right ankle swelling | 0
redness | 0
local rise of temperature | 0
tenderness over lateral malleolus | 0
tenderness over lower third leg laterally | 0
restriction of ankle movements | 0
no neurovascular deficits | 0
normal plain X-ray | 0
hemoglobin 12.5 g/dL | 0
total count 21.28K/uL | 0
neutrophils 19.77K/uL | 0
lymphocytes 0.75K/uL | 0
CRP 360.1 mg/L | 0
ESR 60 mm/hr | 0
RA factor negative | 0
ASO titre 400 IU/ML | 0
sickling negative | 0
normal urine routine | 0
admitted for suspected cellulitis | 0
pediatric consultation for cough | 0
chest X-ray pneumonia | 0
IV cloxacillin started | 0
Staphylococcus aureus in blood culture | 72
general condition deteriorated | 72
elevated temperature | 72
tachycardia (140/min) | 72
respiratory rate 40/min | 72
SPO2 87% | 72
moderate swelling right leg | 72
tender calf | 72
positive Homan sign | 72
D-Dimer negative | 72
CT angiogram no pulmonary embolism | 72
right pleural effusion | 72
bilateral patchy pneumonia | 72
duplex scan popliteal vein thrombosis | 72
thrombophilia workup negative | 72
low molecular heparin treatment | 72
IV cloxacillin continued | 72
clinical improvement | 168
calf swelling reduced | 168
blood parameters normalized | 168
discharged on day 14 | 336
warfarin treatment | 336
repeat duplex scan normal | 504
no recurrence in 6 months | 2160
