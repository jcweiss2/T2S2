86 years old | 0
overweight (BMI = 29) | 0
woman | 0
presented to the emergency department | 0
severe abdominal pain | -24
nausea | -24
vomiting | -24
appendectomy | -73032
implantation of heart pacemaker | -8760
heart rate: 88/min | 0
blood pressure: 110/50 mmHg | 0
saturation: 98% in room air | 0
body temperature: 36.6°C | 0
signs of dehydration | 0
tenderness localized in the middle upper abdomen | 0
no signs of peritoneal irritation | 0
clearly audible peristalsis | 0
serum amylase elevated (1218 U/l) | 0
urinary amylase elevated (8100 U/l) | 0
serum lipase elevated (5850 U/l) | 0
glucose level elevated (175 mg/dl) | 0
no previous diabetes diagnosis | 0
no diabetes medications | 0
serum C-reactive protein level normal (2.1 mg/l) | 0
serum white blood cell count normal (9.57 × 10^9/l) | 0
marginal dilatation of the common bile duct (9 mm) | 0
intrahepatic bile ducts not dilated | 0
gallbladder described as thin-walled | 0
no intraluminal gallstones | 0
pancreas impossible to evaluate due to bowel gas | 0
no intraperitoneal free fluid | 0
no free gas detected during ultrasound | 0
admitted to the surgery department | 0
suspicion of acute pancreatitis | 0
strict diet | 0
intravenous hydration | 0
analgesic treatment | 0
persistent severe abdominal pain | 0
hypotension | 0
oliguria | 0
serum C-reactive protein level slightly elevated (48 mg/l) | 0
decreased serum white blood cell count (2.27 × 10^9/l) | 0
high percentage of neutrophils (77.7%) | 0
increased serum aspartate aminotransferase (59 U/l) | 0
increased serum alanine aminotransferase (53 U/l) | 0
amylase levels comparable to initial | 0
lipase levels comparable to initial | 0
deteriorating general condition | 0
computed tomography (CT) of the abdomen | 16
free gas in the peritoneal cavity | 16
free gas retroperitoneally around duodenum, pancreas, liver | 16
radiologist suggested perforated duodenal diverticulum | 16
decision for emergency surgery | 16
laparotomy | 16
perforation of the duodenum ruled out | 16
significantly enlarged gangrenous gallbladder | 16
free fluid of purulent character | 16
cholecystectomy performed | 16
peritoneal cavity lavage | 16
drainage | 16
retrospective analysis of CT images | 16
gas in the gallbladder wall | 16
gas within pancreatic parenchyma | 16
pneumobilia in the left hepatic lobe | 16
gas penetration into abdominal wall muscles | 16
final diagnosis: emphysematous cholecystitis | 16
gangrenous pancreatitis | 16
retroperitoneal gangrene | 16
transferred to the intensive care unit | 16
critical condition | 16
septic shock | 16
multiorgan failure | 16
increased procalcitonin (38.96 ng/ml) | 16
increased C-reactive protein (118.2 mg/l) | 16
increased D-dimer (2000.0 ng/ml) | 16
increased lactate dehydrogenase (1290 U/l) | 16
increased creatine phosphokinase (3787 U/l) | 16
increased myoglobin (> 12,000 ng/ml) | 16
increased troponin (0.018 ng/ml) | 16
decreased red blood cell count (3.44 × 10^12/l) | 16
decreased hemoglobin level (107.0 g/l) | 16
relaparotomy to exclude intraperitoneal bleeding | 16
cardiac arrest | 16
resuscitation | 16
death | 16
