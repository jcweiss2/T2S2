22 years old | 0
female | 0
presented to the outpatient clinic | 0
fever | 0
sore throat | 0
acute bacterial pharyngitis | 0
oral antibiotics | 0
no improvement | 0
persistent fever | -240
confusion | -240
dyspnea | -240
cyanosed | -240
basal crackles in both lungs | -240
anterior infrahyoid soft neck swelling | -240
emergently intubated | -240
admitted to ICU | -240
leukocytosis | -240
absolute neutrophilia | -240
mild increase in creatinine | -240
high blood sugar | -240
positive acetone in urine | -240
chest x-ray | -240
computed tomography (CT) chest | -240
wide mediastinum | -240
moderate bilateral pleural effusion | -240
adjacent subpleural atelectasis | -240
bilateral basal lung infiltrates | -240
mild pericardial effusion | -240
intercostal tubes inserted | -240
pleural fluid analysis | -240
exudate | -240
pH 7.1 | -240
high white blood cell count | -240
predominantly neutrophils | -240
initial cultures negative | -240
community acquired pneumonia | -240
secondary bilateral empyema | -240
diabetic ketoacidosis | -240
newly diagnosed diabetes mellitus | -240
septic shock | -240
acute kidney injury | -240
progressive edema in all limbs | -336
increase in anterior soft neck swelling | -336
managed with mechanical ventilation | -336
intravenous fluids | -336
insulin | -336
vasopressors | -336
broad spectrum antibiotics | -336
antifungals | -336
no improvement | -336
referred to King Khalid University Hospital | -336
clinical evaluation upon admission | -336
high fever | -336
hypotension | -336
tachycardia | -336
hypoxemia on mechanical ventilation | -336
bilateral intercostal chest tubes | -336
generalized edema | -336
anterior infrahyoid soft neck swelling | -336
repeated CT chest and neck | -336
high density fluid collection in prethyroid region | -336
extending down to sternoclavicular joint | -336
multiple small mediastinal lymph nodes | -336
pretracheal lymph nodes | -336
paratracheal lymph nodes | -336
prevascular lymph nodes | -336
ultrasound guided aspiration of prethyroid fluid | -336
frank pus | -336
thoracic surgery team consulted | -336
conservative management | -336
sputum culture revealed Pseudomonas aeruginosa | -336
Acinetobacter baumannii | -336
antibiotics adjusted | -336
fever persisted | -336
hypotension persisted | -336
deterioration in renal function | -336
renal replacement therapy | -336
neck and chest CT scan repeated | -336
multiloculated collection in neck | -336
extending down to sternum | -336
large loculated cystic lesion in anterior mediastinum | -336
increased pericardial effusion | -336
increased bilateral pleural effusion | -336
basal atelectasis | -336
bilateral consolidation | -336
surgical intervention | -336
cervical dissection | -336
debridement | -336
drainage of pus | -336
left thoracotomy | -336
drainage of mediastinal collection | -336
drainage of left pleural collection | -336
pleuropericardial window | -336
right thoracotomy | -384
debridement | -384
drainage of right pleural collection | -384
samples sent for cultures | -384
no bacterial growth | -384
histopathology revealed acute inflammatory process | -384
gradual improvement in hemodynamics | -384
conscious level improvement | -384
renal function improvement | -384
inflammatory markers improvement | -384
difficult weaning from mechanical ventilation | -384
generalized weakness | -384
tracheostomy postponed | -384
infection in anterior neck | -384
inflammation in anterior mediastinum | -384
high fever | -624
tachycardia | -624
hypotension | -624
requiring vasopressors | -624
repeat CT neck and chest | -624
interval reduction in collections | -624
loculated pleural effusion | -624
bilateral lateral loculated fluid collections | -624
beneath thoracotomy sites | -624
drained by CT guided aspiration | -624
critical illness polyneuropathy | -624
critical illness myopathy | -624
tracheo-esophageal fistula | -624
managed conservatively | -624
tracheostomy | -624
feeding gastrostomy | -624
weaning from mechanical ventilation achieved | -1968
transferred to general ward | -1968
stayed for 6 weeks | -1968
healing of tracheo-esophageal fistula | -1968
oral feeding resumed | -1968
tracheostomy removed | -1968
gastrostomy tubes removed | -1968
discharged from hospital | -1968
