38 years old | 0
    Afro-Brazilian woman | 0
    sickle cell disease (Hb SS) | 0
    acute painful vasoCocclusive crises | -960
    bone infarcts | -960
    skin ulcer of the lower limb | -960
    acute chest syndrome | -960
    autosplenectomy | -960
    jaundice | -2880
    choluria | -2880
    dyspnea on light exertion | -2880
    pain in the right upper abdominal quadrant | -2880
    pain in the lower limbs | -2880
    blood pressure 140 × 90 mm Hg | 0
    heart rate 81 beats per minute | 0
    respiratory rate 18 breaths per minute | 0
    temperature 36.7 °C | 0
    oxygen saturation 96% | 0
    respiratory sounds normal | 0
    painful enlarged liver | 0
    anemia (Hb: 6.7 g/dL; hematocrit: 21%) | 0
    cholestasis (total bilirubin: 16.01 mg/dL; direct bilirubin: 12.11 mg/dL) | 0
    slight elevation of liver enzymes (AST: 138 U/L; ALT: 46 U/L; ALP 445 U/L; GGT 437 mg/dL) | 0
    albumin levels at lower normal limit (3.4 g/dL) | 0
    INR at upper normal limit (1.37) | 0
    serology tests negative for hepatitis B and C, HIV, autoimmune conditions | 0
    positive IgG antibodies for cytomegalovirus | 0
    positive IgG antibodies for Epstein-Barr virus | 0
    alpha-fetoprotein within normal ranges | 0
    ceruloplasmin within normal ranges | 0
    iron metabolism markers slightly altered (iron: 174 μg/dL; transferrin saturation: 68%; total iron binding capacity: 256 μg/dL; ferritin: 575 ng/dL) | 0
    renal function preserved (creatinine: 0.53 mg/dL) | 0
    blood cultures negative | 0
    chest X-ray no change of pulmonary parenchyma | 0
    Hb S fraction 74% (one month before) | -720
    MRI showing enlarged liver with slightly irregular contours and heterogeneous parenchyma | 0
    MRI suggestive of chronic liver disease | 0
    small volume ascites | 0
    gallbladder typical at MRCP | 0
    choledocus duct typical at MRCP |3 0
    slight focal dilatation of biliary tree in right hepatic lobe | 0
    no biliary obstruction detected | 0
    intravenous fluids | 0
    analgesia | 0
    folate | 0
    supplementary oxygen therapy | 0
    received 900 mL packed red blood cells | 0
    hematocrit increased to 25% | 0
    exchange blood transfusion (EBT) | 0
    clinical improvement | 0
    Hb S fraction dropped to 14.3–20.4% | 0
    resolution of respiratory distress | 0
    resolution of lower limb pain | 0
    jaundice persisted | 0
    choluria persisted | 0
    slight abdominal pain persisted | 0
    acute respiratory distress | 312
    fever | 312
    hypoxemia | 312
    chest X-ray diffuse lung opacities | 312
    acute chest syndrome | 312
    transferred to ICU | 312
    mechanical ventilation | 312
    meropenem therapy initiated | 312
    mental confusion | 312
    isolated seizure | 312
    posterior reversible encephalopathy syndrome (PRES) | 312
    normal levels of ammonia | 312
    hepatic encephalopathy discarded | 312
    increasing levels of direct bilirubin | 312
    elevated INR | 312
    Hb S below 25% | 312
    renal function progressively deteriorated | 312
    creatinine 3.31 mg/dL (day of death) | 768
    blood cultures negative in ICU | 312
    airway secretion cultures negative in ICU | 312
    refractory shock | 768
    death | 768
  