69 years old | 0
male | 0
admitted to the hospital | 0
left lower abdomen pain | -336
intermittent fever | -8760
weight loss | -8760
paraumbilical tenderness | 0
left lower quadrant tenderness | 0
abdominal distension | 0
leucocytosis | 0
neutrophilia | 0
eosinophilia | 0
Haemoglobin of 126 g/L | 0
Platelets of 518 * 10^9/L | 0
C-reactive protein 262.48 mg/L | 0
faecal impaction | 0
nonspecific distribution of bowel gases | 0
no air under diaphragm | 0
no signs of bowel obstruction | 0
multifocal segmental wall thickening in the distal ascending, proximal transverse, and distal descending colon | 0
fluid collections suggesting concealed perforations | 0
severe diverticulitis | 0
Piperacillin/Tazobactam | 0
nothing by mouth | 0
symptoms worsened | 96
blood-stained stool | 96
recurrence of multifocal segmental wall thickening | 96
interval increase in size of surrounding collections | 96
severe diverticulitis versus aggressive infections like basidiobolomycosis and actinomycetes | 96
surgical intervention | 96
biopsy for bacterial, TB, fungal cultures | 96
histopathology | 96
liposomal amphotericin B | 96
Amoxicillin/Clavulanic acid | 96
tigecycline | 96
persistently febrile | 192
white blood cells increased to 31.7 * 10^9/L | 192
absolute eosinophils count increased to 3.58 * 10^9/L | 192
haemoglobin dropped to 10 g/dL | 192
redemonstration of circumferential wall thickening of the colon | 192
interval increase in size of fluid collection measuring approximately 7.9 × 9 cm | 192
interval increase in abdominopelvic ascites with surrounding inflammatory changes | 192
faecal peritonitis | 216
multiple colon perforation at sigmoid, transverse, and descending colon | 216
small bowel adhesion | 216
adhesions between small bowel and transverse colon | 216
Adhesolysis | 216
total colectomy | 216
end ileostomy created | 216
placement of two drains | 216
absolute eosinophils count dropped immediately after surgery | 216
haemoglobin dropped to 69.0 g/L | 216
inotropic support | 216
transfused several units of packed red blood cells | 216
minimal ventilator settings | 216
minimal respiratory secretions | 216
no collection found | 216
Pseudomonas aeruginosa | 216
carbapenem resistant Klebsiella variicola | 216
Bacteroides fragilis | 216
Candida glabrata | 216
extensive inflammation involving the full thickness of the colon tissue | 216
extended to the serosal surface | 216
mixed inflammatory cells | 216
sheets of eosinophils | 216
multiple foci of fungal microorganism | 216
thin walled, occasionally septated and surrounded by thick eosinophilic cuff splendore-Hoeppli phenomenon | 216
continuing liposomal amphotericin B 5 mg/kg IV once per day | 216
Itraconazole 200 mg orally twice per day | 216
modifying antibacterial agents | 216
condition deteriorated | 216
passed away due to refractory septic shock | 216
