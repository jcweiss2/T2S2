26 years old | 0
male | 0
admitted to the hospital | 0
rash | 0
pain | 0
edema | 0
cellulitis | 0
body temperature 38.2 | 0
heart rate 110 | 0
blood pressure 140/70 | 0
respiration rate 22 | 0
hypotonia | -8760
poor sucking | -8760
cryptorchidism | -8760
pneumonia | -8760
diagnosis of PWS | -8760
mental retardation | -6336
diabetes | -6336
obesity | -6336
hyperphagia | -6336
chronic renal failure | -1092
hemodialysis | -1092
amputation advised | -24
skin disinfection | -24
antibiotic treatment | -24
obstruction in arteriovenous fistula | -24
aneurysmectomy | -24
vessel ligation | -24
local anesthesia | -24
anxiety | -24
guardian in operating room | -24
dual lumen catheterization | -24
left brachiocephalic fistula surgery | -24
general anesthesia requested | -24
hemoglobin 7.5 | -1
hematocrit 22.8 | -1
glomerular filtration rate 11.65 | -1
sodium 131 | -1
potassium 6.6 | -1
glucose 112-354 | -1
pH 7.311 | -1
PaCO2 36.0 | -1
PaO2 70.9 | -1
HCO3- 17.8 | -1
SaO2 93.0 | -1
EKG normal | -1
pulmonary edema | -1
cardiomegaly | -1
height 150 | -1
weight 105 | -1
BMI 46.7 | -1
short neck | -1
short limbs | -1
sleep apnea | -1
mild sleep apnea | -1
Mallampatti class II | -1
oxygen treatment | -1
mental retardation | -1
simple communication | -1
H2 antagonist | -1
vital signs | 0
body temperature 37.5 | 0
heart rate 85 | 0
blood pressure 160/90 | 0
respiration rate 22 | 0
invasive arterial pressure measurement | 0
USG guided arterial catheterization | 0
SaO2 95 | 0
oxygen administration | 0
upper body elevation | 0
remifentanil | 0
propofol | 0
loss of consciousness | 0
SaO2 drop | 0
mask ventilation | 0
tidal volume 250 | 0
EtCO2 20-30 | 0
atracurium | 0
endotracheal intubation | 0
SaO2 77 | 0
Cormack and Lehane classification | 0
vocal cords small | 0
intubation failed | 0
SaO2 58 | 0
mask ventilation | 0
SaO2 82 | 0
endotracheal intubation | 0
SaO2 70 | 0
pressure control ventilation | 0
airway pressure 30 | 0
respiration rate 15 | 0
FiO2 50 | 0
tidal volume 400 | 0
EtCO2 42 | 0
SaO2 93 | 0
FiO2 70 | 0
positive end expiratory pressure | 0
dexamethasone | 0
sevoflurane | 0
remifentanil | 0
SaO2 93-98 | 0
Hb 8.8 | 1
K+ 5.4 | 1
glucose 77 | 1
dextrose | 1
insulin | 1
spontaneous breathing | 1
atracurium | 1
vital signs stable | 3
systolic blood pressure 100-115 | 3
diastolic blood pressure 45-60 | 3
heart rate 75-85 | 3
ABGA | 3
electrolytes | 3
glucose | 3
Hb 7.8 | 3
K+ 5.8 | 3
glucose 96 | 3
PaCO2 52.5 | 3
PaO2 110 | 3
dextrose | 3
spontaneous breathing | 3
tidal volume 300 | 3
vital capacity 800 | 3
extubation | 3
oxygen mask | 3
SaO2 88 | 3
expiratory wheezing | 3
inhalation therapy | 3
steroids | 3
β2 agonist | 3
recovery room | 3
oxygen | 3
upper body elevation | 3
SaO2 95 | 3
intensive care unit | 3
chest X-ray | 3
SaO2 90 | 24
oxygen treatment | 24
vital signs stable | 48
general ward | 48