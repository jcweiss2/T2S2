22 years old | 0
female | 0
admitted to the hospital | 0
fever | -72
shortness of breath | -72
feeling generally unwell | -72
chest X-ray demonstrated multiple opacities | -72
CT of the chest and abdomen | -72
multiple cavitations | -72
pulmonary embolism | -72
femoral thrombosis | -72
GPA confirmed | -72
warfarin | -72
rituximab | -72
methylprednisolone | -72
Immunoglobulins (IgG) | -72
fluconazole | -72
second infusion of rituximab | -72
third infusion of rituximab | -72
prophylactic co-trimoxazole | -72
angioedema | -72
rash | -72
90% total body surface area (TBSA) | -72
oral and ophthalmic mucosa involved | -72
fluconazole stopped | -72
co-trimoxazole stopped | -72
steroids increased | -72
suspicion of Stevens-Johnson syndrome (SJS) | -72
deterioration | -72
100% TBSA | -72
critical care team support | -72
TEN suspected | -72
TEN confirmed | -72
skin biopsy | -72
SCORTEN score of 3 | -72
mortality risk of 35.3% | -72
referred to specialist burns centre | -72
Piperacillin/Tazobactam (Tazocin) | 0
Vancomycin | 0
sputum and wound swab sensitivities | 0
prednisolone reduced to 40 mg daily | 168
good re-epithelisation of the skin | 240
discharged | 504
physiotherapy | 504