36 years old | 0
    male | 0
    butcher | 0
    history of smoking | 0
    history of cannabinoid consumption | 0
    presented to the emergency room | 0
    severe headache | -24
    fever | -24
    dysarthria | -24
    confusion | -24
    psychomotor agitation | -24
    Glasgow Coma Scale 13 | 0
    nuchal rigidity | 0
    respiratory distress | 0
    desaturation | 0
    diminished breath sounds bilaterally | 0
    Brudzinski's sign absent | 0
    Kernig's sign absent | 0
    Lasegue's sign absent | 0
    leukocytosis | 0
    neutrophilia | 0
    elevated C-reactive protein | 0
    thrombocytopenia | 0
    unremarkable renal function | 0
    unremarkable hepatic function | 0
    unremarkable ionogram | 0
    unremarkable serology tests | 0
    negative urine toxicology tests | 0
    cerebral computerized tomography | 0
    hydrocephalus in third ventricle | 0
    cerebrospinal fluid analysis | 0
    glucose 1mg/dL | 0
    protein 671 mg/dL | 0
    white blood cell count 104 cells/mm3 | 0
    Gram-positive diplococci | 0
    acute bacterial meningitis | 0
    ceftriaxone | 0
    vancomycin | 0
    acyclovir | 0
    dexamethasone | 0
    thiamine supplementation | 0
    tested positive for SARS-CoV-2 | 0
    sedated | 0
    mechanically ventilated | 0
    transferred to ICU | 0
    vasopressor support | 0
    intracranial pressure monitoring | 0
    intracranial hypertension | 0
    cerebrospinal fluid drainage | 0
    seizures | 24
    epileptiform discharges | 24
    levetiracetam | 24
    cerebrospinal fluid culture positive | 24
    Streptococcus suis II | 24
    susceptible to penicillin | 24
    susceptible to ceftriaxone | 24
    antibiotic therapy for 14 days | 24
    dexamethasone discontinued after 5 days | 0
    improvement in oxygenation | 168
    hemodynamic stability | 168
    sedation stopped | 168
    weaned from mechanical ventilation | 168
    no recurrence of seizures | 168
    no focal neurological deficits | 168
    discharged to district hospital | 168
    complete resolution of symptoms | 168
    no hearing loss | 0
    no COVID-19 symptoms | 0
    no asplenia | 0
    no diabetes mellitus | 0
    no alcoholism | 0
    no malignancy | 0
    no structural heart disease | 0
    occupational exposure | 0
    frequent contact with nasal and oral cavity | 0
    