74 years old | 0
female | 0
admitted to the hospital | 0
lethargy | -48
weakness | -48
diagnosed with DM | -504
history of hypertension | 0
history of hyperlipidemia | 0
small cell lung cancer | 0
metastatic to the brain | 0
gamma knife radiation therapy | -168
dexamethasone | -504
cerebral edema | -504
elevated blood glucose level | -168
follow-up appointment with oncologist | -168
left eyelid swelling | 0
erythema | 0
preseptal cellulitis | 0
ophthalmoplegia | 24
visual impairment | 24
mental status worsened | 24
difficulty following commands | 24
aggressive hydration | 0
i.v. fluids | 0
insulin | 0
septic shock | 24
broad-spectrum antibiotics | 24
vasopressors | 24
central venous catheter | 24
computed tomography scan | 24
left ocular proptosis | 24
invasive rhinomaxillary fungal disease | 24
amphotericin B | 120
surgical debridement | 120
magnetic resonance imaging | 120
invasive fungal disease | 120
left inferior frontal lobe | 120
multidisciplinary meeting | 120
healthcare agent declined further surgery | 120
orbital exenteration | 120
skull base surgery | 120
conservative medical management | 120
surgical pathology report | 144
invasive mucormycosis | 144
R. oryzae | 144
S. maltophilia | 144
blood cultures | 144
MSSA | 144
liposomal amphotericin B | 120
cefazolin | 144
levofloxacin | 144
herpetic lesion | 168
valacyclovir | 168
vasopressor support | 0
electrolyte abnormalities | 120
hypokalemia | 120
potassium supplementation | 168
spironolactone | 168
discharged | 600
lost to follow-up | 600
declined appointments | 600