17 years old | 0
    female | 0
    admitted to the hospital | 0
    acute onset of behavioral change | 0
    extreme politeness | 0
    obedience | 0
    pre-morbid gregarious personality | -672
    progression to excessive and irrelevant talks | -672
    features of disinhibition | -672
    frank psychotic features | -240
    verbal aggression | -240
    physical aggression | -240
    muttering to herself | -240
    marked delusional thoughts | -240
    tendency to run amok | -240
    diagnosis of acute functional psychosis | -240
    oleanzapine started | -240
    behavioral syndrome persisted | -240
    mild reduction of psychomotor activity | -240
    stiffness of whole body | -240
    akinesia | -240
    mutism | -240
    evaluated by neurologist and psychiatrist | -240
    MRI brain scattered T2 and FLAIR hyperintensities | -240
    CSF examination no cells | -240
    normal CSF protein | -240
    normal CSF glucose levels | -240
    negative CSF viral markers | -240
    negative VDRL test | -240
    negative gram stain | -240
    negative AFB stain | -240
    negative India ink | -240
    negative cryptococcal antigen | -240
    negative bacterial cultures | -240
    negative mycobacterial cultures | -240
    negative fungal cultures | -240
    EEG non-specific diffuse theta delta slowing | -240
    low grade fever | -240
    serum Creatinine Phosphokinase raised to 1800 U/dl | -240
    diagnosis of NMS due to oleanzapine | -240
    dantrolene started | -240
    hydration started | -240
    slight reduction of rigidity | -240
    no other improvement noticed | -240
    clinical worsening over next 2 weeks | 336
    increasing mental obtundation | 336
    persistent akinetic mute state | 336
    frequent bouts of tachypnea | 672
    tachycardia | 672
    hypotension | 672
    sweating | 672
    deterioration over next 48 hours | 720
    gasping for breath | 720
    oxygen desaturation | 720
    endotracheal intubation | 720
    mechanical ventilation | 720
    brought to our center | 720
    widely fluctuating heart rate | 720
    widely fluctuating blood pressure | 720
    stimulus-induced sinus tachycardia | 720
    tachypnea | 720
    diaphoresis | 720
    sedative infusion | 720
    provisional diagnosis of sepsis syndrome | 720
    bilateral aspiration pneumonia | 720
    received critical care | 720
    received medical support | 720
    re-evaluated by neurology team | 720
    possibility of immune encephalitis considered | 720
    MRI brain repeated | 720
    similar changes as before | 720
    normal infectious meningoencephalitis workup | 720
    CSF samples sent for anti-NMDA receptor antibody | 720
    CSF samples sent for anti-VGKC antibody | 720
    CSF samples sent for anti# 100 Days of Code - Log

### R1

**Day 1**: January 1, 2021

**Today's Progress**: I worked on the freecodecamp responsive web design course. I finished the cat image page. I started the balance sheet challenge. I set up a basic html structure and started working on the css.

**Thoughts:** I'm finally starting my 100 Days of Code challenge. It's day 1 and I'm excited. I know I can do this. It's been a long time since I started working on web development. I'm going to use the fcc responsive web design course as my main resource. I also have a few projects that I need to finish.

**Link to work:** [Cat Image Project](https://github.com/ShivanshuS/freecodecamp-projects/blob/main/responsive-web-design/cat-photo-app/readme.md)

**Day 2**: January 2, 2021

**Today's Progress**: I worked on the balance sheet project. I added the header and main sections. I set up the colors, borders, and fonts. I added the data classes and the data entries. I tried to match the design as much as possible.

**Thoughts:** Today was a bit challenging. I had to figure out how to use the different CSS properties to match the design. I'm still getting the hang of it, but I'm making progress. The balance sheet is starting to look like the example.

**Link to work:** [Balance Sheet Project](https://github.com/ShivanshuS/freecodecamp-projects/blob/main/responsive-web-design/balance-sheet/readme.md)

**Day 3**: January 3, 2021

**Today's Progress**: I continued working on the balance sheet. I added the data entries and adjusted the colors. I fixed some alignment issues. I also started working on the navigation bar challenge.

**Thoughts:** The balance sheet is almost complete. I just need to adjust a few more details. The navigation bar is another challenge, but I'm confident I can tackle it. I'm getting better at using CSS Flexbox and Grid.

**Link to work:** [Balance Sheet Project](https://github.com/ShivanshuS/freecodecamp-projects/blob/main/responsive-web-design/balance-sheet/readme.md)

**Day 4**: January 4, 2021

**Today's Progress**: I finished the balance sheet project. I made the final adjustments to the layout and colors. It now matches the example perfectly. I also started the navigation bar challenge. I set up the HTML structure and added some basic CSS.

**Thoughts:** Completing the balance sheet was a relief. It's a good feeling to see the project come together. The navigation bar is next. I need to make it responsive and styled properly.

**Link to work:** [Balance Sheet Project](https://github.com/ShivanshuS/freecodecamp-projects/blob/main/responsive-web-design/balance-sheet/readme.md)

**Day 5**: January 5, 2021

**Today's Progress**: Worked on the navigation bar. Added the logo, links, and search bar. Styled the elements using Flexbox. Made the navigation bar responsive with media queries.

**Thoughts:** The navigation bar is taking shape. I had to adjust the spacing between elements and make sure it looks good on mobile. Flexbox is really helpful for layouts. I'm starting to understand media queries better.

**Link to work:** [Navigation Bar Project](https://github.com/ShivanshuS/freecodecamp-projects/blob/main/responsive-web-design/navigation-bar/readme.md)

**Day 6**: January 6, 2021

**Today's Progress**: Finished the navigation bar project. Adjusted the media queries for different screen sizes. Tested the responsiveness. Also started the registration form challenge.

**Thoughts:** The navigation bar is responsive and looks good on all devices. Now onto the registration form. I need to create a form with proper validation and styling.

**Link to work:** [Navigation Bar Project](https://github.com/ShivanshuS/freecodecamp-projects/blob/main/responsive-web-design/navigation-bar/readme.md)

**Day 7**: January 7, 2021

**Today's Progress**: Started the registration form. Set up the HTML structure with form elements. Added basic CSS styling. Began working on form validation using HTML5 attributes.

**Thoughts:** Forms can be tricky, especially with validation. I'm using HTML5 validation to make it easier. The form is starting to take shape. Need to add more styling and ensure it's responsive.

**Link to work:** [Registration Form Project](https://github.com/ShivanshuS/freecodecamp-projects/blob/main/responsive-web-design/registration-form/readme.md)

**Day 8**: January 8, 2021

**Today's Progress**: Continued work on the registration form. Added more form fields, styled them, and improved the layout. Worked on the CSS for different input types.

**Thoughts:** The form is getting more complex. Styling each input type requires attention to detail. I'm making sure the form is user-friendly and accessible.

**Link to work:** [Registration Form Project](https://github.com/ShivanshuS/freecodecamp-projects/blob/main/responsive-web-design/registration-form/readme.md)

**Day 9**: January 9, 2021

**Today's Progress**: Finished the registration form. Added final touches to the styling and validation. Tested the form for responsiveness and accessibility.

**Thoughts:** The registration form is complete. It's responsive, accessible, and validates inputs properly. Next up is the product landing page.

**Link to work:** [Registration Form Project](https://github.com/ShivanshuS/freecodecamp-projects/blob/main/responsive-web-design/registration-form/readme.md)

**Day 10**: January 10, 2021

**Today's Progress**: Started the product landing page project. Created the header, navigation, and hero section. Added basic CSS for layout and styling.

**Thoughts:** The product landing page is a bigger project. It requires multiple sections and a responsive design. I'm starting with the header and hero section.

**Link to work:** [Product Landing Page Project](https://github.com/ShivanshuS/freecodecamp-projects/blob/main/responsive-web-design/product-landing-page/readme.md)

**Day 11**: January 11, 2021

**Today's Progress**: Worked on the product landing page. Added features section and pricing cards. Styled the sections using CSS Grid and Flexbox.

**Thoughts:** The features and pricing sections are important parts of the landing page. Using Grid and Flexbox helps create a clean layout. I need to make sure the design is consistent.

**Link to work:** [Product Landing Page Project](https://github.com/ShivanshuS/freecodecamp-projects/blob/main/responsive-web-design/product-landing-page/readme.md)

**Day 12**: January 12, 2021

**Today's Progress**: Continued working on the product landing page. Added the footer and contact section. Adjusted the CSS for responsiveness.

**Thoughts:** The footer and contact sections complete the landing page. I'm testing responsiveness on different devices to ensure it looks good everywhere.

**Link to work:** [Product Landing Page Project](https://github.com/ShivanshuS/freecodecamp-projects/blob/main/responsive-web-design/product-landing-page/readme.md)

**Day 13**: January 13, 2021

**Today's Progress**: Finished the product landing page. Made final adjustments to the CSS and tested all sections. Ensured the page is fully responsive.

**Thoughts:** The product landing page is complete. It's a comprehensive project that covers many aspects of responsive design. I'm proud of how it turned out.

**Link to work:** [Product Landing Page Project](https://github.com/ShivanshuS/freecodecamp-projects/blob/main/responsive-web-design/product-landing-page/readme.md)

**Day 14**: January 14, 2021

**Today's Progress**: Started the technical documentation page project. Created the sidebar navigation and main content sections. Added basic CSS for layout.

**Thoughts:** The technical documentation page requires a fixed sidebar and responsive content. I'm using CSS Grid to layout the page. It's a new challenge but manageable.

**Link to work:** [Technical Documentation Page Project](https://github.com/ShivanshuS/freecodecamp-projects/blob/main/responsive-web-design/technical-documentation-page/readme.md)

**Day 15**: January 15, 2021

**Today's Progress**: Continued working on the technical documentation page. Added content sections and styled them. Implemented smooth scrolling for navigation links.

**Thoughts:** Adding content to the documentation page is time-consuming. I need to ensure the information is accurate and well-presented. Smooth scrolling improves user experience.

**Link to work:** [Technical Documentation Page Project](https://github.com/ShivanshuS/freecodecamp-projects/blob/main/responsive-web-design/technical-documentation-page/readme.md)

**Day 16**: January 16, 2021

**Today's Progress**: Finished the technical documentation page. Adjusted the CSS for responsiveness and tested all links. Added media queries for mobile devices.

**Thoughts:** The documentation page is now complete. It's fully responsive and the navigation works smoothly. Next up is the tribute page.

**Link to work:** [Technical Documentation Page Project](https://github.com/ShivanshuS/freecodecamp-projects/blob/main/responsive-web-design/technical-documentation-page/readme.md)

**Day 17**: January 17, 2021

**Today's Progress**: Started the tribute page project. Researched the subject and gathered content. Created the HTML structure and added basic styling.

**Thoughts:** The tribute page needs to be informative and visually appealing. I'm starting with the structure and will add styling later. The content is key here.

**Link to work:** [Tribute Page Project](https://github.com/ShivanshuS/freecodecamp-projects/blob/main/responsive-web-design/tribute-page/readme.md)

**Day 18**: January 18, 2021

**Today's Progress**: Continued work on the tribute page. Added images, timelines, and quotes. Styled the sections using CSS.

**Thoughts:** Incorporating images and timelines makes the page more engaging. Styling each section to highlight important information is crucial.

**Link to work:** [Tribute Page Project](https://github.com/ShivanshuS/freecodecamp-projects/blob/main/responsive-web-design/tribute-page/readme.md)

**Day 19**: January 19, 2021

**Today's Progress**: Finished the tribute page. Added final touches to the content and styling. Tested responsiveness on different devices.

**Thoughts:** The tribute page is complete. It tells the story effectively and looks good on all devices. I'm happy with the outcome.

**Link to work:** [Tribute Page Project](https://github.com/ShivanshuS/freecodecamp-projects/blob/main/responsive-web-design/tribute-page/readme.md)

**Day 20**: January 20, 2021

**Today's Progress**: Started the survey form project. Created the form structure and added various input types. Began styling with CSS.

**Thoughts:** The survey form is another form project but with different requirements. I need to include various form elements and style them appropriately.

**Link to work:** [Survey Form Project](https://github.com/ShivanshuS/freecodecamp-projects/blob/main/responsive-web-design/survey-form/readme.md)

**Day 21**: January 21, 2021

**Today's Progress**: Continued work on the survey form. Added more form fields and improved the layout. Implemented CSS for better visual hierarchy.

**Thoughts:** The form is getting more detailed. Each field needs to be styled to ensure clarity and usability. I'm focusing on user experience here.

**Link to work:** [Survey Form Project](https://github.com/ShivanshuS/freecodecamp-projects/blob/main/responsive-web-design/survey-form/readme.md)

**Day 22**: January 22, 2021

**Today's Progress**: Finished the survey form. Added validation and tested all form elements. Ensured the form is responsive and accessible.

**Thoughts:** The survey form is now complete. It's user-friendly and accessible. All form elements work as expected. Next project is the quiz page.

**Link to work:** [Survey Form Project](https://github.com/ShivanshuS/freecodecamp-projects/blob/main/responsive-web-design/survey-form/readme.md)

**Day 23**: January 23, 2021

**Today's Progress**: Started the quiz page project. Created the HTML structure for questions and answers. Added basic CSS for styling.

**Thoughts:** The quiz page requires dynamic content but I'm building it statically for now. I'll add JavaScript later for interactivity.

**Link to work:** [Quiz Page Project](https://github.com/ShivanshuS/freecodecamp-projects/blob/main/responsive-web-design/quiz-page/readme.md)

**Day 24**: January 24, 2021

**Today's Progress**: Continued working on the quiz page. Added more questions and styled the sections. Implemented CSS transitions for interactivity.

**Thoughts:** Styling the quiz page to make it engaging is important. Transitions add a layer of interactivity without JavaScript. It's looking better.

**Link to work:** [Quiz Page Project](https://github.com/ShivanshuS/ffreecodecamp-projects/blob/main/responsive-web-design/quiz-page/readme.md)

**Day 25**: January 25, 2021

**Today's Progress**: Finished the quiz page. Added final styling and tested responsiveness. Ensured the layout is consistent across devices.

**Thoughts:** The quiz page is complete. It's static but styled well. Next, I'll move on to JavaScript projects.

**Link to work:** [Quiz Page Project](https://github.com/ShivanshuS/freecodecamp-projects/blob/main/responsive-web-design/quiz-page/readme.md)

**Day 26**: January 26, 2021

**Today's Progress**: Started JavaScript algorithms and data structures course on freeCodeCamp. Completed the first few exercises on variables and functions.

**Thoughts:** Switching to JavaScript to strengthen my programming skills. The basics are straightforward, but I need to practice more complex problems.

**Link to work:** [freeCodeCamp Profile](https://www.freecodecamp.org/shivanshu)

**Day 27**: January 27, 2021

**Today's Progress**: Continued with JavaScript exercises. Worked on arrays, loops, and conditional statements. Solved problems like sum and multiply arrays.

**Thoughts:** Arrays and loops are fundamental. Practicing these exercises helps in understanding how to manipulate data structures.

**Link to work:** [freeCodeCamp Profile](https://www.freecodecamp.org/shivanshu)

**Day 28**: January 28, 2021

**Today's Progress**: Worked on more JavaScript exercises. Explored object manipulation and higher-order functions. Solved problems using map, filter, and reduce.

**Thoughts:** Higher-order functions are powerful. They make code cleaner and more efficient. I'm starting to see the benefits of functional programming.

**Link to work:** [freeCodeCamp Profile](https://www.freecodecamp.org/shivanshu)

**Day 29**: January 29, 2021

**Today's Progress**: Started