66 years old | 0
male | 0
atrial fibrillation | 0
common atrial flutter | 0
radiofrequency pulmonary vein isolation | 0
wide defragmentation of the left atrium | 0
creation of a posterior box | 0
sinus rhythm restored | 0
external electric shock at 200 J | 0
general anesthesia | 0
3D intracardiac navigation | 0
transseptal approach | 0
transoesophageal echocardiography | 0
fluoroscopic guidance | 0
oesophageal temperature monitored | 0
discharged from the hospital | 24
anticoagulant treatment | 24
proton pump inhibitors | 24
referred to the emergency department | 336
dyspnoea at rest | 336
thoracic discomfort | 336
rapid atrial fibrillation | 336
significant signs of inflammation | 336
CRP > 200 mg/L | 336
hyperleukocytosis | 336
hemodynamically stable | 336
poor tolerance of the arrhythmia | 336
beta-blockers initiated | 336
digoxin initiated | 336
unsuccessful cardioversion attempt with amiodarone | 336
abundant heterogeneous pericardial effusion | 336
circumferential pericardial effusion | 336
systolic-diastolic notch on the left atrium | 336
significant respiratory variation of the transvalvular flow | 336
pericardiocentesis | 336
removal of 400 cc of cloudy, orange pericardial fluid | 336
numerous polynuclear cells | 336
purulent fluid | 336
pericardial drain left in place | 336
hemodynamic failure | 336
hypotension | 336
fever | 336
acute respiratory failure | 336
acute anuric renal failure | 336
hepatic failure | 336
hyperlactatemia (6 mmol/L) | 336
severe acute right ventricular dysfunction | 336
cardiogenic shock | 336
septic shock | 336
broad-spectrum antibiotic treatment (piperacillin–tazobactam and amikacin flash) | 336
inotropic support with dobutamine | 336
multiphase thoracic–abdominal–pelvic CT scan | 336
minimal hydroaeric pericardial effusion | 336
upper-route opacification using a 1:10 diluted oral water-soluble contrast medium | 336
discontinuity in the anterior oesophageal wall | 336
extraluminal contrast leakage | 336
stagnation in the posterior portion of the cardiac mass | 336
oesophageal–pericardial fistula | 336
endoscopic management | 336
fistulous orifice visualized 31 cm from the dental arches | 336
18-cm covered oesophageal prosthesis placed | 336
final control with injection of water-soluble contrast medium into the esophagus | 336
rapid extubation | 336
weaning from amines | 336
sudden alteration in neurological state | 408
Glasgow Coma Scale of 3 | 408
cerebral CT scan revealed several ischaemic strokes of gaseous origin | 408
diffuse intraparenchymal and subarachnoid air embolism | 408
supratentorial and subtentorial air embolism | 408
migration of the oesophageal prosthesis | 408
presence of air bubbles in the left ventricle | 408
presence of air bubbles in the left auricle | 408
fistula between the esophagus and the right superior pulmonary vein | 408
brain MRI confirmed multiple ischaemic lesions | 432
mesencephalic involvement | 432
diffuse supra-tentorial cerebral edema | 432
subfalcine herniation | 432
very poor neurological prognosis | 432
brain death declared | 432
