53 years old | 0
female | 0
admitted to the emergency department | 0
dyspnoea | 0
chest tightness | 0
dizziness | 0
palpitations | 0
nausea | 0
vomiting | 0
oral glucose tolerance test | -12
transient hypoglycaemia | -12
impaired fasting glucose | -672
borderline haemoglobin A1c | -672
hypertension | -672
dyslipidaemia | -672
secondary hyperparathyroidism | -672
simvastatin | -672
calcium carbonate | -672
cholecalciferol | -672
metoprolol | -672
losartan | -672
pale skin | 0
cool extremities | 0
weak radial pulses | 0
prolonged capillary refilling time | 0
respiratory rate 40 breaths per minute | 0
oxygen saturation 80% | 0
heart rate 114 bpm | 0
blood pressure 111/75 mmHg | 0
bilateral inspiratory crackles | 0
soft abdomen | 0
no tenderness | 0
no palpable mass | 0
no focal neurological deficits | 0
body temperature 37.7°C | 0
hypoxaemia | 0
metabolic acidosis | 0
hyperglycaemia | 0
elevated cardiac troponin T | 0
normal C-reactive protein | 0
leucocytosis | 0
acute kidney injury stage 1 | 0
sinus tachycardia | 0
hypokinesia | 0
left ventricular ejection fraction 15% | 0
pulmonary oedema | 0
normal coronary arteries | 0
takotsubo-type contraction pattern | 0
fever 38.5°C | 24
lactate increased | 24
urinary output decreased | 24
heart rate 122 bpm | 24
systolic blood pressure 85 mmHg | 24
cardiac index 2.1 L/min/m² | 24
mean pulmonary artery pressure 23 mmHg | 24
norepinephrine | 24
levosimendan | 24
non-invasive ventilatory support | 24
antipyretics | 24
anxiolytics | 24
cardiac index 3 L/min/m² | 24
LVEF 20-25% | 24
LVEF 40-45% | 48
weaned from norepinephrine | 48
continued levosimendan | 48
insulin therapy | 24
empiric antibiotics | 24
negative cultures | 48
cardiac MRI confirmed takotsubo cardiomyopathy | 168
elevated S-cortisol | 168
normal S-renin | 168
normal S.aldosterone | 168
normal S.TSH | 168
normal S.T3 | 168
normal S.T4 | 168
elevated metanephrine | 168
elevated normetanephrine | 168
elevated methoxytyramine | 168
elevated chromogranin A | 168
readmitted due to abnormal catecholamines | 408
adrenergic blockade instituted | 408
CT revealed phaeochromocytoma | 504
left adrenalectomy | 1440
adrenergic blockade stopped | 1440
discharged | 1536
follow-up visit | 2544
scheduled CT | 8760
scheduled catecholamine testing | 8760
scheduled follow-up visit | 8760
