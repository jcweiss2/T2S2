56 years old | 0
female | 0
ESRD | 0
admitted to the ER | 0
fever | -48
painful rash on the hands | -48
abnormal blood culture report | -48
growth of yeast | -48
shortness of breath | -336
cough | -336
non-bloody white sputum | -336
subjective fever | -336
chills | -336
hemodialysis | -672
arteriovenous graft | -672
hypertension | 0
diabetes mellitus | 0
obese | 0
febrile | 0
blood pressure 156/86 mmHg | 0
oxygen saturation 98% | 0
violaceous macular lesions | 0
basilar crackles | 0
hypertensive retinopathy | 0
fungal chorioretinitis | 0
leukocytosis | 0
WBC count 1.34 × 10^4/μL | 0
blood cultures positive for yeast | 0
fluid collection around the arteriovenous graft | 0
fine needle aspiration | 12
culture grew candida zeylanoides | 12
excision of infected arteriovenous graft | 24
temporary Shiley catheter | 24
transesophageal echocardiogram | 24
negative for vegetation | 24
chest CT | 24
peripheral nodular lesions | 24
infective emboli | 24
bronchoscopy | 48
bronchoalveolar lavage | 48
white exudate | 48
tissue cultures | 48
Candida zeylanoides | 48
VITEK 2 system | 48
negative test for serum precipitins to Aspergillus fumigatus | 48
negative test for serum precipitins to Aspergillus niger | 48
caspofungin | 48
fluconazole | 72
repeat blood cultures | 72
negative for fungal growth | 72
discharged from the hospital | 168
parenteral fluconazole | 168
completed antifungal therapy | 1008
followed with us in dialysis center | 1008