59 years old | 0
female | 0
presented to the emergency department | 0
progressive central abdominal pain | -336
distention | -336
laparoscopic adjustable band insertion | -96336
nausea | -336
vomiting | -336
denied dysphagia | -336
denied odynophagia | -336
denied change in bowel habit | -336
afebrile | 0
tachycardic | 0
diffuse abdominal tenderness | 0
guarding | 0
elevated white cell count | 0
elevated C-reactive protein | 0
hyperlactatemia | 0
distended air-filled stomach | 0
intragastric band erosion | 0
internalization of gastric band and distal connector tubing | 0
moderate free fluid | 0
ascites | 0
mesenteric inflammatory fat stranding | 0
portal vein thrombosis | 0
exploratory laparotomy | 0
ischemic small bowel segment | 0
resected small bowel segment | 0
blood clots extruding from mesenteric vascular arcade | 0
on-table OGD | 0
deformed shaped stomach | 0
gastric band eroded through stomach wall | 0
biofilm formed around band device | 0
sealing perforation | 0
device retrieved | 0
stomach closed in two layers | 0
abdominal drains inserted | 0
monitored in intensive care unit | 0
hepatic ultrasound | 0
thrombosed portal vein | 0
commenced on tinzaparin sodium | 0
gastroenterology input | 0
dietician input | 0
physiotherapy input | 0
hematology input | 0
barium meal | 504
normal gastric contours | 504
no filling defects | 504
no gastric outlet emptying | 504
discharged | 504
