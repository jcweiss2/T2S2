48 years old | 0
female | 0
Roux-en-Y gastric bypass | -6720
Crohn's disease | -6720
rheumatoid arthritis | -6720
atrial fibrillation | -6720
anticoagulation | -6720
septic ascending cholangitis | -120
laparoscopic cholecystectomy | -120
endoscopic retrograde cholangiopancreatography (ERCP) | -120
admitted to the intensive care unit | -120
acute tubular necrosis | -120
temporary dialysis | -120
atrial fibrillation with rapid ventricular response | -120
spontaneous rectus sheath hematoma | -120
intravenous heparin | -120
cessation of anticoagulation | -96
blood transfusions | -96
embolization of right inferior epigastric artery | -96
hematoma perforated the right lateral wall of her bladder | -96
gross hematuria | -96
pain | -96
leaking around her foley catheter | -96
hematoma induced bladder spasms | -96
persistent lower urinary tract symptoms | -672
urgency/frequency | -672
dysuria | -672
gross hematuria | -672
cystoscopy | -24
large friable right sided bladder mass | -24
biopsy | -24
necrotic debris | -24
rare reactive urothelium | -24
referred to our institution | 0
magnetic resonance urography (MRU) | 0
hematoma decreased in size | 0
perforating through the right lateral wall of her bladder | 0
transurethral resection (TUR) | 24
large, smooth, homogeneous bladder mass | 24
resection to the level of the bladder mucosa | 24
clot visualized extending through a defect in the bladder wall | 24
pathology of the resected tissue showed a hematoma | 24
negative for malignancy | 24
worsening symptoms of urgency | 168
terminal voiding pain | 168
repeat MRU | 168
further extrusion of the hematoma within the bladder lumen | 168
trial of an indwelling catheter | 168
repeat endoscopic resection | 168
possible open surgery with partial cystectomy | 168
repeat TUR | 336
large, organized hematoma protruding from a 4 cm bladder wall cavity | 336
extensive resection | 336
entering the right lateral wall cavity | 336
identifying and amputating the base of the hematoma stalk | 336
visualized completely healed epithelium | 336
complete resolution of her irritative voiding symptoms | 336
MRU confirmed all the hematoma had been evacuated | 504
bladder had a sacculation of the right lateral bladder wall | 504
residual area of hematoma measuring 3.7 cm | 504
episode of gross hematuria | 17520
associated with a UTI | 17520
CT urogram demonstrated thickening of the right lateral bladder | 17520
tethering to the pelvic sidewall | 17520
cystoscopy confirmed a persistent right lateral diverticulum | 17520
well healed epithelium | 17520