64 years old | 0
male | 0
diabetes | -672
hypertension | -672
insulin | -672
amlodipine | -672
admitted to the intensive care unit | 0
septic shock | 0
leukocyturia | 0
fever | 0
desaturation | 0
hypotension | 0
tachycardia | 0
elevated blood sugar | 0
inflammatory syndrome | 0
elevated white blood cells | 0
elevated C-reactive protein | 0
thrombocytopenia | 0
normal renal function | 0
abdomino-pelvic CT scan | 0
painful infiltration | 0
crepitus | 0
destroyed left kidney | 0
aerial collection | 0
fluid resuscitation | 0
vasoactive drugs | 0
noradrenaline | 0
glycemic control | 0
insulin infusion | 0
empirical antibiotic therapy | 0
imipenem | 0
ciprofloxacin | 0
clinical improvement | 72
transfer to urology department | 240
discharge | 312
Emphysematous pyelonephritis | 0
septic shock diagnosis | 0
renal infection | -672
necrotizing renal infection | -672
gas in renal parenchyma | 0
gas in urinary tract | 0
gas in perineal tissue | 0
Escherichia coli infection | 0
Klebsiella pneumoniae infection | 0
Proteus mirabilis infection | 0
gram-positive cocci infection | 0
anaerobic organisms infection | 0
excretory tract obstruction | -672
pregnancy | -672
renal transplantation | -672
abdominal CT scan | 0
prognostic classification | 0
therapeutic decision | 0
left kidney involvement | 0
right kidney involvement | 0
bilateral involvement | 0
surgical intervention | 0
conservative treatment | 0
aggressive resuscitation | 0
broad-spectrum antibiotics | 0
third or fourth-generation cephalosporins | 0
carbapenems | 0
combination therapy | 0
gentamicin | 0
antimicrobial treatment | 0
nephrectomy | 0 
CT scan diagnosis | 0 
early diagnosis | 0 
good resuscitation | 0 
blood sugar control | -672 
urinary tract infection treatment | -672 
written informed consent | -24 
publication of case report | 312 
accompanying images | 312 
ethical approval | -24 
funding resources | -24 
author contribution | -24 
conflicts of interest | -24 
research registration | -24 
data availability | -24 
provenance and peer review | -24 
sponsorships | -24 
competing interests | -24