63 years old | 0
male | 0
African-American | 0
admitted to the hospital | 0
food aversion | -96
fever | -96
chills | -96
chest pain | -96
abdominal pain | -96
remote history of tobacco use | -100000
remote history of cocaine use | -100000
no diabetes mellitus | 0
no other medical illnesses | 0
not on any prescription or over-the-counter medications | 0
poor dentition | 0
fever of 38.3°C | 0
hemodynamically stable | 0
white cell count of 22.4 × 10^9/L | 0
aspartate aminotransferase of 93 units/L | 0
alanine aminotransferase of 110 units/L | 0
total bilirubin of 1.2 mg/dL | 0
multiple indeterminate hypo-attenuating lesions throughout the liver | 0
multiple complex hypoechoic foci throughout the liver | 0
multiple cystic lesions with enhancing internal septations and marked diffusion restriction | 0
empiric treatment with broad-spectrum antibiotics | 0
resolution of fever | 24
aspiration from one of the abscess cavities | 24
placement of three drainage catheters in the right hepatic lobe | 24
drainage from the hepatic abscess grew Fusobacterium nucleatum | 24
antibiotics were narrowed based on culture and sensitivities | 24
liver aspirate testing for acid-fast organisms was negative | 24
liver aspirate testing for aerobic and fungal cultures was negative | 24
stool cultures were negative | 24
examination for ova, parasites, giardia, cryptosporidium, clostridium difficile and entamoeba was negative | 24
blood and urine cultures were negative | 24
testing for viral hepatitis was negative | 24
testing for human immunodeficiency virus was negative | 24
tumor markers for alpha-fetoprotein, cancer antigen 19-9 and carcinoembryonic antigen were unremarkable | 24
trans-thoracic echocardiogram revealed no evidence of valvular vegetations | 24
endoscopic evaluation by colonoscopy revealed two 4 - 8 mm adenomatous polyps in the rectum | 24
mild diverticulosis in the sigmoid colon | 24
no evidence of prior or current inflammation or infection | 24
panorex demonstrated multiple missing teeth and lucency around the root of a left mandibular premolar | 24
periapical abscess | 24
output from the hepatic drains continued to decrease | 168
drains were eventually removed | 168
affected teeth were extracted | 168
antibiotics were transitioned to an oral route | 168
discharged home | 672
asymptomatic at 6 weeks post-hospitalization follow-up | 1008
liver enzymes trended down to normal levels | 1008
repeat cross-sectional imaging demonstrated a significant interval decrease in rim enhancement and size of the known liver abscesses | 1008