85 years old| 0
    male | 0
    admitted to a local hospital | -1344
    trismus | -1344
    hypertonia | -1344
    leg injury | -1344
    C. tetani infection | -1344
    immunoglobulins | -1344
    tetanus vaccination | -1344
    metronidazole | -1344
    transferred to ICU | -1320
    tracheostomy | -1320
    mechanical ventilation | -1320
    vasoactive support | -1320
    respiratory failure | -1320
    seizures | -1320
    baclofen | -1320
    midazolam | -1320
    diazepam | -1320
    severely slow cerebral activity | -1320
    worsening respiratory function | -1320
    opacity on chest radiography | -1320
    peripheral leukocytosis | -1320
    ventilator-associated pneumonia (VAP) | -1320
    blood cultures | -1320
    tracheal secretion samples | -1320
    Klebsiella pneumoniae | -1320
    methicillin-sensitive Staphylococcus aureus (MSSA) | -1320
    piperacillin-tazobactam | -1320
    moved to geriatric unit | -1296
    coma | -1296
    spontaneous breathing | -1296
    supplemental oxygen | -1296
    antibiotic therapy switched to linezolid | -1296
    VAP exacerbation | -1296
    meropenem | -1296
    septic shock | -1296
    awoke gradually | -1296
    feeding tube removed | -1296
    cholestasis | -1296
    acute edematous pancreatitis | -1296
    postponed endoscopic treatment | -1296
    urinary tract infection | -1296
    multidrug-resistant organisms (MDROs) | -1296
    K. pneumoniae | -1296
    Acinetobacter baumannii | -1296
    Enterococcus faecalis | -1296
    colistin | -1296
    amoxicillin-clavulanate | -1296
    clinical condition improved | -1296
    eligible for rehabilitation | -1296
    MDRO isolation | 0
    tracheal supplemental oxygen | 0
    bladder catheter | 0
    pressure ulcers (right unstageable, left stage II, sacrum stage II, right elbow stage III) | 0
    sarcopenic | 0
    low handgrip strength (9.9 kg) | 0
    low appendicular skeletal mass (ASM, 16.9 kg) | 0
    rehabilitation | 0
    Clostridioides difficile infection | 24
    oral vancomycin | 24
    AF with third-degree atrioventricular block | 72
    heart rate 30 beats/min | 72
    transferred to cardiac ICU | 72
    single-chamber pacemaker implantation | 72
    hyperkinetic delirium | 72
    transferred back to hospital | 96
    Pseudomonas aeruginosa bloodstream infection | 96
    ceftazidime-avibactam | 96
    amikacin | 96
    SARS-CoV-2 positive | 96
    remdesivir | 96
    droplet isolation | 96
    recurrence of C. difficile | 108
    transferred to geriatric medicine unit | 108
    fidaxomicin | 108
    bloodstream infection due to Candida parapsilosis | 240
    fluconazole-resistant | 240
    MSSA | 240
    Candida tropicalis | 240
    intravenous catheter replaced | 240
    caspofungin | 240
    cefazolin | 240
    bloodstream infection caused by P. aeruginosa | 408
    piperacillin-tazobactam | 408
    aztreonam | 408
    ceftazidime-avibactam (antibiotic resistance) | 408
    cefepime | 480
    tracheostomy closure | 624
    nutritional supplementation | 624
    malnutrition | 624
    sarcopenia | 624
    intensive rehabilitation compromised | 624
    infectious complications | 624
    non-infectious complications | 624
    short physiotherapy sessions | 624
    discharged | 624
    postural transition with assistance | 624
    motor reconditioning | 624
    respiratory reconditioning | 624
    posture transition training | 624
    aided transfers | 624
    axial stability | 624
    balance improvement exercises | 624
    breath-movement coordination exercises | 624
    thoracic expansion | 624
    girdle opening exercises | 624
    inhalation-exhalation exercises | 624
    wheelchairs recommended | 624
    walkers recommended | 624
    mobility deficit | 624
    ENT follow-up | 624
    geriatric follow-up | 624
    rehab evaluations recommended | 624