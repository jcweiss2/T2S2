70 years old | 0
male | 0
admitted to the hospital | 0
chronic diarrhea | -240
confusion | -240
gout | -720
discharged on colchicine | -720
discharged on allopurinol | -720
discharged on prednisone taper | -720
diarrhea began | -720
denied abdominal pain | 0
denied hematochezia | 0
denied melena | 0
denied nausea | 0
denied vomiting | 0
denied fevers | 0
denied chills | 0
denied night sweats | 0
tremulous | 0
weak | 0
worsening fatigue | 0
2 falls | -168
required 2 L of oxygen | 0
sleep apnea | 0
continuous positive airway pressure | 0
heart failure | 0
furosemide | 0
non-alcoholic steatohepatitis | 0
liver transplant | -3600
hypertension | 0
coronary artery disease | 0
drug eluting stent placement | 0
gout | 0
60-pack-year smoking history | 0
quit smoking | -10560
denied alcohol use | 0
denied drug use | 0
family history of thyroid disease | 0
tachycardia | 0
lethargic | 0
oriented only to person | 0
intact cranial nerves | 0
normal motor examination | 0
normal sensory examination | 0
morbidly obese | 0
no thyroid enlargement | 0
no ophthalmopathy | 0
white blood cells 4.76 K/cumm | 0
hemoglobin 10.0 g/dL | 0
platelets 106 K/cumm | 0
sodium 134.0 mmol/L | 0
potassium 5.20 mmol/L | 0
BUN 74.0 mg/dL | 0
creatinine 3.3 mg/dL | 0
magnesium 1.7 mg/dL | 0
phosphorus 7.2 mg/dL | 0
INR 1.54 | 0
blood cultures negative | 0
respiratory bacterial culture negative | 0
gastrointestinal PCR negative | 0
herpes simplex virus PCR negative | 0
cytomegalovirus PCR negative | 0
chest x-ray negative | 0
urinalysis negative | 0
VRE cultures negative | 0
MRSA cultures negative | 0
CT head negative | 0
urine drug screen negative | 0
tacrolimus levels within goal range | 0
hemoglobin A1c 4.7 | 0
glucose level 286 mg/dL | 0
lithium level less than 0.1 mmol/L | 0
procalcitonin level 0.09 ng/mL | 0
TSH level 0.01 mIU/L | 0
Free T4 level 5.91 ng/dL | 0
Free T3 level 14.5 pg/mL | 0
thyrotoxicosis | 0
thyroid storm | 0
diffuse mild hypervascularity | 0
no masses or nodules | 0
anti-thyroglobulin antibody 2555.0 IU/mL | 0
Burch-Wartofsky score 50 | 0
propanol 40 mg every six hours | 0
methimazole 20 mg three times a day | 0
prednisone 60 mg daily | 0
transferred to ICU | 0
non-ST-elevation myocardial infarction | 24
right lower lobe pneumonia | 24
piperacillin-tazobactam | 24
thrombocytopenia | 24
thyroid storm treatment | 0
thyroid uptake scan | 216
thyroiditis | 216
globally decreased uptake | 216
no active nodules | 216
prednisone 40 mg daily | 504
Free T3 level 2.1 pg/mL | 2160
T4 level 0.82 ng/dL | 2160
TSH level 16.23 mIU/L | 2160
levothyroxine 50 mcg daily | 2160
euthyroid | 3024
Free T3 level 2.5 pg/mL | 3024
T4 level 1.17 ng/dL | 3024
TSH level 1.38 mIU/L | 3024