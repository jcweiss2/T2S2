73 years old | 0
female | 0
duodenal switch surgery | -6720
pancreatic head adenocarcinoma | 0
obstructive jaundice | 0
DBE-ERCP attempted | 0
DBE-ERCP unsuccessful | 0
inability to reach the papilla | 0
EUS-guided choledochoenterostomy not attempted | 0
percutaneous transhepatic biliary drainage | 0
PTBD internalized | 0
common bile duct metal stent | 0
osseous metastasis | 0
nonsurgical candidate | 0
cholangitis | 1920
septic shock | 1920
obstructed CBD stent | 1920
refused PTBD placement | 1920
EUS-guided CDE | 1920
linear echoendoscope passed | 1920
extrahepatic bile duct examined | 1920
extrahepatic bile duct measured | 1920
common wall between small bowel and CBD interrogated | 1920
extrahepatic bile duct punctured | 1920
bile aspirated | 1920
cholangiogram showed obstruction | 1920
EUS-guided CDE with LAMS | 1920
double pigtail stent placed | 1920
sepsis improved | 1944
transferred from ICU to medical floor | 1944
discharged home | 1968