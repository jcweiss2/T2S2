high-grade fever | -120
generalized body ache | -120
headache | -120
altered sensorium | -24
joint pains | -120
epigastric pain | -120
ingual lymphadenopathy | 0
mild generalized rash | 0
no eschar | 0
disoriented | 0
no focal neurological deficit | 0
no neck rigidity | 0
provisional diagnosis of acute febrile illness with undifferentiated fever | 0
workup to rule out tropical infections | 0
malaria negative | 0
dengue negative | 0
typhoid negative | 0
leptospira negative | 0
Scrub typhus antigen card positive | 0
Scrub immunoglobulin M positive | 0
blood and other body fluid cultures sterile | 0
leukocytosis | 0
mild hyperbilirubinemia | 0
transaminitis | 0
slightly raised international normalized ratio | 0
hepatitis B antigen negative | 0
hepatitis C antibody negative | 0
mild fatty infiltration of the liver | 0
tablet doxycycline 100 mg twice daily | 0
defervescence | 48
orientation improved | 48
weakness of both lower limbs | 96
weakness progressed to upper limbs | 96
absent deep tendon reflexes | 96
flexor plantar responses | 96
bladder incontinence | 96
no bowel incontinence | 96
breathing difficulty | 96
respiratory distress | 96
intubated | 96
mechanical ventilation | 96
MRI of the brain without abnormality | 96
MRI of the cervical spine without abnormality | 96
nerve conduction velocity showed motor sensory demyelinating polyneuropathy | 96
cerebrospinal fluid analysis | 96
intravenous immunoglobulin therapy | 96
tablet rifampicin 600 mg twice daily | 96
improvement in weakness | 144
improvement in respiratory parameters | 144
weaned off mechanical ventilation | 216
extubated | 216
oral feeding started | 216
aggressive limb and chest physiotherapy | 216
shifted out from ICU | 240
discharged from hospital | 336
full neurological recovery | 336