43 years old | 0
male | 0
admitted to the hospital | 0
hypertension | -8760
mild lacunar infarction | -8760
perindopril | -8760
aspirin | -8760
community-acquired pneumonia | -24
respiratory failure | -24
invasive ventilatory support | -24
consolidation over the right lower zone | -24
leukocytosis | -24
raised C-reactive protein levels | -24
mild hypoalbuminemia | -24
hyperglycemia | -24
co-amoxiclav | -24
septic shock | -18
triple inotropes support | -18
piperacillin/tazobactam | -18
improved condition | -168
extubation | -168
failed to maintain adequate oxygenation | -168
reintubation | -168
tracheostomy | -120
persistent respiratory failure | -120
investigated for myasthenia gravis | -120
anti-acetylcholine receptor antibody level | -120
nerve conduction study | -120
decremental responses | -120
characteristic decremental compound muscle action potential amplitude | -120
diagnosis of myasthenia gravis | -120
IV immunoglobulin | -120
pyridostigmine | -120
prednisolone | -120
azathioprine | -120
improved condition | -48
removed tracheostomy | 0
discharged | 0
oral azathioprine | 0
oral pyridostigmine | 0
contrast-enhanced computed tomography scan | 0
no evidence of thymoma | 0
followed up every 3 months | 0
responded well to medication | 24
no further myasthenic crises | 24