56 years old | 0
male | 0
pre-diabetes | 0
hyperlipidemia | 0
admitted to the hospital | 0
ST-elevation myocardial infarction | 0
transported to the catheterization lab | 0
primary percutaneous intervention (PCI) | 0
left anterior descending (LAD) artery occluded | 0
stent implemented | 0
thrombus aspiration | 0
no-reflow phenomenon | 0
hemodynamically unstable | 0
ventricular fibrillation (VF) | 0
pulseless electrical activity (PEA) | 0
CPR commenced | 0
LUCAS3 device used | 0
ECMO decision | 0
cannulation | 0
CPR discontinued | 15
PCI finished | 15
LAD flow restored | 15
three-vessel disease | 15
transported to the ICU | 15
mechanical ventilation weaned off | 24
neurological consequences absent | 24
lactate levels increased | 24
vasopressors administered | 24
inotropes administered | 24
cannula positions checked | 24
ECMO machine operating | 24
hemoglobin (Hgb) fell | 24
probable bleeding focus | 24
massive blood transfusion protocol | 48
lactate dropped | 48
Hgb raised | 48
abdominal compartment syndrome | 72
intraabdominal hypertension | 72
declining urine output | 72
creatinine increased | 72
vasopressors increased | 72
lactate increased | 72
Hgb unchanged | 72
abdominal CT scan | 96
hemoperitoneum | 96
liver laceration | 96
transported to the operating room | 96
left lobectomy of the liver | 96
extubated | 120
condition improved | 120
vasopressors reduced | 120
lactate normalized | 120
PRBC transfusions | 120
ejection fraction (EF) improved | 168
arrhythmias | 168
non-sustained VT | 168
ventricular fibrillation | 168
repeat defibrillations | 168
EF reduced | 192
LVAD implantation decision | 192
transferred to another hospital | 168
ECMO support | 168
spontaneous breathing | 168
hemodynamically stable | 168
awake and alert | 168
no neurological sequelae | 168
catastrophic multiorgan failure | 240
sepsis | 240
death | 240