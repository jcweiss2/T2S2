11 years old | 0
male | 0
admitted to the hospital | 0
fever | -96
nausea | -96
abdominal pain | -96
pneumonia | -61368
contact with COVID-19 | -1200
elevated C-reactive protein | 0
elevated procalcitonin | 0
normal whole blood cell count | 0
bowel wall thickening in terminal ileum | 0
multiple enlarged lymph nodes along ileocolic artery | 0
intravenous antibiotics | 0
diarrhea | 48
hypotension | 72
inotropic agents | 72
white blood cell count 5.82 × 103/µL | 72
segmented neutrophils 92.1% | 72
platelet count 100 × 103/µL | 72
elevated serum CRP 189.50 mg/L | 72
elevated procalcitonin 14.55 mcg/L | 72
elevated aspartate aminotransferase | 72
elevated alanine aminotransferase | 72
elevated pro-brain natriuretic peptide | 72
elevated prothrombin time | 72
elevated activated partial thromboplastin time | 72
elevated fibrinogen | 72
elevated D-dimer | 72
normal cardiac markers | 72
cardiomegaly | 96
hypoalbuminemia | 96
intravenous immunoglobulin (IVIG) | 96
conjunctival injection | 144
cracked lips | 144
strawberry tongue | 144
left main coronary artery dilatation | 144
left anterior descending artery not tapered | 144
right coronary artery dilatation | 144
aneurysmal changes | 144
mild pericardial effusion | 144
pleural effusion | 144
lung parenchymal consolidation | 144
high-dose aspirin | 144
fever subsided | 192
erythematous papular rash | 192
finger desquamation | 192
aspirin dose reduction | 192
desquamation of left wrist | 312
desquamation of perianal area | 312
normalized inflammation markers | 312
normalized coagulopathy | 312
resolved cardiomegaly | 312
resolved pleural effusion | 312
reduced enlarged lymph nodes | 312
reduced coronary artery dilatation | 312
negative PCR for pathogens | 312
negative PCR for SARS-CoV-2 | 312
positive SARS-CoV-2 IgG antibody | 312
negative SARS-CoV-2 IgM antibody | 312
discharge | 312
