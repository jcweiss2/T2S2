80 years old | 0
female | 0
admitted to the intensive care unit | 0
dyspnea | -96
lethargy | -96
chest tightness | -96
denied cough | -96
denied hemoptysis | -96
denied fever | -96
denied gastrointestinal symptoms | -96
denied recent sick contacts | -96
denied traveling | -96
end-stage renal disease (ESRD) | -6720
severe pulmonary hypertension | -6720
chronic obstructive pulmonary disease (COPD) | -6720
former smoker | -6720
15-pack year history of cigarette use | -6720
no anti-coagulants | 0
no amiodarone | 0
no chemotherapeutic agents | 0
no recent nitrofurantoin use | 0
acute respiratory distress | 0
tachypnea | 0
hypoxemia | 0
oxygen saturation of 89% on room air | 0
oxygen saturation of 95% on 2 liters of oxygen via nasal cannula | 0
afebrile | 0
temperature of 36.7°C | 0
blood pressure of 89/55 mmHg | 0
heart rate of 89 beats per minute | 0
lungs examination was normal | 0
awake and alert | 0
cardiac examination was normal | 0
abdomen examination was normal | 0
no petechiae | 0
no bruising | 0
no gingival bleeding | 0
no oozing from sites of intravenous access | 0
anemia | 0
hemoglobin level of 9.9 g/dL | 0
leukocytosis | 0
white blood cell count was 13.0×103 cells/μL | 0
left shift | 0
neutrophil count was 10.8×103 cells/μL | 0
serum lactate of 3.7 mmol/L | 0
arterial blood gas done on room air with a pH of 7.317 | 0
pCO2 of 57.7 mmHg | 0
pO2 of 40.2 mmHg | 0
coagulation profile reported an international normalized ratio (INR) of 1.1 | 0
prothrombin time (PT) of 13.5 seconds | 0
partial thromboplastin time (PTT) of 30.6 seconds | 0
urine and serum toxicology were negative | 0
chest x-ray showed retrocardiac infiltrates | 0
nasopharyngeal swabs, rapid testing was positive for influenza A | 0
clinical status of the patient deteriorated rapidly | 12
development of shock | 12
intubated | 12
mechanical ventilation | 12
pressors | 12
vancomycin | 12
piperacillin-tazobactam | 12
azithromycin | 12
oseltamivir | 12
chest computed tomography (CT) showed left lower and right upper lobe infiltrates | 24
right lower lobe nodule | 24
no evidence of a pulmonary embolus | 24
fiberoptic bronchoscopy performed on day 2 of admission | 48
airway erythema of the left and right bronchial trees | 48
BAL performed in the left lower lobe showed progressive bloody returns | 48
consistent with DAH | 48
BAL done in the right lower lobe also produced similar findings | 48
bronchoscopy and blood and urine cultures were negative | 48
BAL cytology 4 1513 cells/mm3 for WBCs | 48
54% were segmented neutrophils | 48
44% were lymphocytes | 48
111 250 million cells/mm3 of red blood cells | 48
autoimmune workup including antinuclear antibody, cytoplasmic and perinuclear antineutrophilic cytoplasmic autoantibodies, and rheumatoid factor were negative | 48
echocardiogram showed severe pulmonary hypertension | 48
pulmonary artery systolic pressure of 78 mmHg | 48
hypoxic | 48
arterial to inspired oxygen (PaO2/FiO2) ratio of 102 mmHg | 48
on a positive end expiratory pressure of 8 mmHg | 48
intravenous methylprednisolone 250 mg/day was started | 48
improvement in oxygenation by day 3 | 72
arterial to inspired PaO2/FiO2 ratio of 317 mmHg | 72
repeated fiberoptic bronchoscopy done 3 days following the first | 96
normal mucosa | 96
progressively clear returns on BAL performed in the left lower lobe | 96
respiratory conditions improved | 96
decreased oxygen requirement | 96
septic shock | 168
died 2 weeks after admission | 336