29 years old | 0
Asian | 0
woman | 0
gravida 1 | 0
para 0 | 0
27 weeks of gestation | 0
acute onset of exacerbation of respiratory distress | 0
fever (>38°C) | -216
nasal discharge | -216
coughing | -216
antibiotics | -168
orthopnoea | 0
exacerbation of respiratory distress (wet-warm) | 0
systolic murmur (3/6 grade) at the apex | 0
bilateral coarse crackles | 0
bilateral leg oedema | 0
hypothyreosis | 0
levothyroxine | 0
sinus tachycardia | 0
complete right branch bundle block | 0
massive pulmonary congestion | 0
elevated brain natriuretic peptide (564.5 pg/mL) | 0
elevated C-reactive protein (4.86 mg/dL) | 0
elevated white blood cell count (13,890/μL) | 0
severe mitral valve regurgitation | 0
prolapse of the anterior mitral leaflet | 0
mobile vegetations (1.5 cm and 2 cm) | 0
severe pulmonary hypertension (112 mmHg) | 0
LVEF 71% | 0
suspected infective endocarditis | 0
emergent interventions | 0
multi-disciplinary conference | 0
betamethasone injection | 0
caesarean section | 0
delivery of male infant (1,154 g) | 0
APGAR scores 1, 5, 6 | 0
uterine compression suture | 0
mitral valve replacement with biological valve | 0
mitral valve leaflets occupied by vegetations | 0
anterior mitral leaflet perforation | 0
post-operative ICU admission | 0
histopathological examination showing acute neutrophil-dominant inflammation | 0
intravenous ceftriaxone | 0
intravenous sulbactam/ampicillin | 0
reduced LVEF (41%) | 144
abnormal anterior wall motion | 144
occlusion of mid-left anterior descending artery | 336
occlusion of peripheral right coronary artery | 336
multiple asymptomatic cerebral infarctions | 360
beta-blocker | 336
angiotensin-converting enzyme inhibitor | 336
discharge | 696
neonate discharge | 2280
normal mitral valve function at follow-up | N/A
slightly decreased LVEF (43%) at follow-up | N/A
