80 years old | 0
    female | 0
    referred for surgical treatment of recurrent RCC | 0
    first endoscopic surgery 2 years prior | -17520
    cyst fenestration | -17520
    partial cyst wall resection | -17520
    pedicled nasoseptal flap technique | -17520
    no CSF fistula observed | -17520
    bilateral reduction in visual acuity | -17520
    bitemporal hemianopsia | -17520
    mild bifrontal headache for 1 year | -17520
    no pituitary dysfunction | -17520
    preoperative sellar CT | -17520
    preoperative sellar MRI | -17520
    cystic sellar lesion | -17520
    recovered from visual disturbances | -17520
    returned to daily activities | -17520
    recurrence of visual disturbance | -8760
    recurrence of bifrontal headaches | -8760
    neurologic examination | 0
    anisocoric pupils | 0
    fixed mydriasis in left eye | 0
    bitemporal hemianopsia | 0
    new endoscopic transnasal transsphenoidal surgery | 0
    gross total resection achieved | 0
    CSF leak observed during cyst dissection | 0
    nasoseptal flap resurface | 0
    no hypertensive episodes during procedure | 0
    postoperative sellar MRI confirmed total resection | 0
    reservoir sign | 0
    CSF leakage | 0
    conservative approach with head elevation | 0
    neuro check | 0
    stable until 3rd postoperative day | 72
    minimal CSF outflow | 72
    no surgical procedure performed | 72
    subtle paraparesis | 96
    paraplegia | 96
    dorsal spine MRI revealed T3-T4 intramedullary lesion | 96
    hyperintense on T2 | 96
    right side on axial plane | 96
    emergency thoracic laminectomy T2-T5 | 96
    SDAVF observed | 96
    intramedullary hematoma observed | 96
    feeder artery on right T3 dural sleeve identified | 96
    arterial supply interrupted | 96
    vessels draining entered dura as single arterialized vein | 96
    dilated tortuous spinal vein on dorsal surface | 96
    draining vein-like varix thrombosed | 96
    partially projected into cord | 96
    intradural dorsal fistula | 96
    Type I spinal arteriovenous fistula | 96
    shunting point coagulated and divided | 96
    intramedullary hematoma evacuated | 96
    hematomyelia caused by rupture of draining vein | 96
    neurogenic shock | 96
    high doses of norepinephrine | 96
    admitted to ICU | 96
    no CSF rhinorrhea observed | 96
    progressive worsening of neurogenic shock | 240
    septic shock due to pneumonia | 240
    high doses of vasoactive amines | 240
    mean arterial pressure 50-60 mmHg | 240
    hypoxic encephalopathy | 240
    brain death | 240
    brain CT showed diffuse white matter hypodensity | 240
    no hypertensive episodes | 240
    no corticosteroid therapy | 240
    patient consent obtained | 240
    ethical standards followed | 240
    <|eot_id|>
    