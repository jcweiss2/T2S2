malaise | -72
fever | -72
loss of appetite | -72
chills | -72
nausea | -72
cardiac arrest | 0
ventricular fibrillation | 0
defibrillation | 0
adrenaline administration | 0
coved-type ST elevation in V1 and V2 | 0
hypercalcemia | 0
hypotension | 2
septic shock | 2
tazobactam-piperacillin administration | 2
vasopressors administration | 2
extubation | 48
fever reoccurrence | 120
liver abscess | 120
meropenem administration | 120
vancomycin administration | 120
puncture drainage | 120
pilsicainide test | 720
implantable cardioverter defibrillator implantation | 720
discharge | 720
tumor resection | 720
ectopic parathyroid adenoma diagnosis | 720
multiple endocrine neoplasia type 1 diagnosis | 720
nonfunctional pituitary adenoma diagnosis | 720
nonfunctional adrenal tumor diagnosis | 720
J point elevation | -1728
early repolarization | -1728
high parathyroid hormone levels | 720
abnormal uptake in the anterior mediastinum | 720
tumors in the pituitary and adrenal glands | 720 
no shortness of breath | 0 
denies chest pain | 0