65 years old | 0
    female | 0
    presented to the hospital | 0
    nausea | -48
    vomiting | -48
    diarrhea | -48
    CIDP | -2160
    prednisone 40–60 mg daily | -2160
    emigrated from Guatemala | -175200
    visited Guatemala annually | -175200
    prednisone 60 mg daily | 0
    positive Strongyloides serology | 0
    titer 2.11 index value | 0
    peripheral eosinophilia | 0
    no prior anti-helminthic treatment | 0
    blood pressure 94/72 mmHg | 0
    heart rate 158 beats/min | 0
    respiratory rate 26 breaths/min | 0
    oxygen saturation 94% | 0
    temperature 37.0 °C | 0
    rigors | 0
    dry mucous membranes | 0
    clear lung fields | 0
    suprapubic tenderness | 0
    WBC count 22,000/mm³ | 0
    19% bands | 0
    0% eosinophils | 0
    urinalysis 22 WBC/hpf | 0
    IV fluids | 0
    ciprofloxacin | 0
    metronidazole | 0
    methylprednisolone 100 mg IV | 0
    admitted to ICU | 0
    piperacillin-tazobactam | 0
    methylprednisolone discontinued | 0
    prednisone 30 mg twice daily | 0
    Escherichia coli in blood culture | 0
    Escherichia coli in urine culture | 0
    stool studies negative for enteric pathogens | 0
    hemodynamic improvement | 48
    transferred to medical ward | 48
    progressive hypoxemia | 120
    bilateral pleural effusions | 120
    diffuse perihilar opacities | 120
    diffuse peripheral air space opacities | 120
    progressive bilateral infiltrates | 192
    blood in tracheobronchial tree | 192
    persistently hemorrhagic BAL fluid | 192
    intubated | 192
    transferred to ICU | 192
    WBC count 24,000/mm³ | 192
    7% bands | 192
    13% eosinophils | 192
    platelets 348,000/mm³ | 192
    prothrombin time 13.9 s | 192
    DAH | 192
    methylprednisolone 1 g daily | 192
    oral ivermectin 200 mcg/kg | 192
    Strongyloides stercoralis in BAL fluid | 216
    corticosteroids discontinued | 216
    subcutaneous ivermectin 200 mcg/kg | 216
    resolving hemorrhage on bronchoscopy | 216
    ANCA negative | 216
    anti-GBM negative | 216
    ANA negative | 216
    HIV negative | 216
    HTLV-1 negative | 216
    stool monitoring for Strongyloides clearance | 216
    improvement over 10 days | 432
    discharged | 432
    oral ivermectin therapy for 4 weeks | 432
    
    