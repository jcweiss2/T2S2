56 years old | 0
    woman | 0
    presented to the emergency department | 0
    abdominal pain | -120
    persistent abdominal pain for five days | -120
    long-standing smoker | -0
    no previously diagnosed chronic medical conditions | 0
    no recent exposure to sick contacts | 0
    upper respiratory tract infection two weeks previously | -336
    self-resolved upper respiratory tract infection | -336
    no recent history of travel | 0
    tachycardic (110-115 beats/min) | 0
    hypertensive (169/110 mmHg) | 0
    afebrile | 0
    soft but tender abdomen | 0
    white blood cell count 20×10^9/L | 0
    CT angiography of abdomen and pelvis | 0
    infrarenal aortic aneurysm | 0
    periaortic hematoma 6.4 cm × 10 cm | 0
    suggestive of rupture | 0
    mild atheromatous changes in renal arteries and visceral vessels | 0
    unremarkable intra-abdominal structures | 0
    relatively young age | 0
    female sex | 0
    small size and inflammatory appearance of ruptured aneurysm | 0
    suggestive of mycotic aneurysm | 0
    blood cultures drawn | 0
    initiated ciprofloxacin | 0
    initiated cefazolin | 0
    emergent open repair through midline transperitoneal approach | 0
    edematous retroperitoneum | 0
    adherent duodenum | 0
    significant inflammatory changes in aorta | 0
    extending distally into iliac arteries | 0
    periaortic fluid nonpurulent | 0
    Gram stain of periaortic fluid | 0
    moderate polymorphs with no organisms seen | 0
    in situ aorto-bi-iliac 12 mm × 7 mm Hemashield graft | 0
    transferred to ICU | 0
    postoperative care | 0
    continued ciprofloxacin | 0
    continued cefazolin | 0
    acute occlusion of the graft | 24
    second surgery | 24
    extensive thrombectomy of both limbs of the graft | 24
    left iliofemoral bypass | 24
    consistently poor flow | 24
    declining condition | 24
    increasing pressors | 24
    broadened antibiotics to meropenem | 24
    broadened antibiotics to vancomycin | 24
    broadened antibiotics to fluconazole | 24
    sepsis treatment | 24
    negative blood cultures at initial presentation | 0
    need for hemodialysis | 24
    renal failure | 24
    culture results from aneurysm sac reported four days after surgery | 96
    subtyping performed shortly thereafter | 96
    Haemophilus influenzae type B infection | 96
    CT scan 19 days into admission | 456
    free air under diaphragm | 456
    free air around graft | 456
    exploratory laparotomy | 456
    perforated colon | 456
    gross graft contamination with stool and pus | 456
    subtotal colectomy | 456
    end-ileostomy | 456
    graft heavily irrigated | 456
    bilateral axillofemoral grafts placed | 456
    8 mm ringed polytetrafluoroethylene | 456
    explantation of infected graft four days later | 528
    edematous and friable bowel | 528
    two inadvertent enterotomies | 528
    additional surgeries for enterotomy repair | 528
    nine separate operations in two months | 0
    tracheostomy in ICU | 0
    prolonged ventilation | 0
    new-onset lumbar plexopathy | 0
    ongoing medical care | 0
    physiotherapy support | 0
    recovery | 0
    discharged to floor from ICU on postoperative day 82 | 1968
    antibiotics discontinued on postoperative day 91 | 2184
    discharged to home hospital on postoperative day 120 | 2880
    