70 years old | 0
    male | 0
    admitted to the Intensive Care Unit (ICU) | 0
    acute respiratory distress | -72
    fever | -72
    cerebrovascular accident (hemorrhagic stroke) | -4320
    anticoagulation therapy | -4320
    acute pulmonary embolism | -4320
    implantation of a vena cava filter | -4320
    hospital-acquired pneumonia | 0
    severe sepsis | 0
    hemodynamic collapse | 0
    hypotension | 0
    cold sweating | 0
    hypoxia | 0
    absence of lung infiltration at chest X-ray | 0
    transthoracic echocardiography | 0
    massive tricuspid insufficiency | 0
    papillary muscle rupture | 0
    suspected endocardial vegetation | 0
    transesophageal echocardiography | 0
    leaflet rupture | 0
    reflective metallic structures trapping in valvular leaflets | 0
    pericardial effusion | 0
    chest-abdominal X-ray | 0
    presence of metallic elements in the right heart | 0
    absence of the cava filter in the cava district | 0
    open heart surgery | 0
    tricuspid valve insufficiency | 0
    presence of 800 ml of blood in the pericardium | 0
    migration of the cava filter fragments through the interventricular septum | 0
    migration of the cava filter fragments through the right ventricular apex | 0
    removal of the tricuspid valve | 0
    removal of vena cava filter fragments | 0
    implantation of a prosthetic tricuspid valve | 0
    successful recovery | 24
    