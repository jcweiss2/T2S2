41 years old | 0
male | 0
admitted to the hospital | 0
altered mental status | -120
fever | -120
diffuse myalgia | -120
flu-like symptoms | -120
fever | -120
muscle pain | -120
severe fatigue | -120
presyncopal event | -24
intubated | 0
mechanical ventilation | 0
protect airway | 0
no nausea | 0
no vomiting | 0
no diarrhea | 0
no skin rashes | 0
chronic hepatitis C infection | 0
IV drug use | 0
no allergies | 0
no medications | 0
smoking | 0
blood pressure 144/95 mmHg | -1
heart rate 130 beats/minute | -1
oral temperature 101.9°F | -1
respiratory rate 18 breaths/minute | -1
oxygen saturation 97% | -1
AMS | 0
toxic | 0
moderate distress | 0
normocephalic | 0
atraumatic head | 0
no palpable masses | 0
poor dentition | 0
no lymphadenopathy | 0
no jugular venous distention | 0
no carotid bruits | 0
tachycardia | 0
normal S1 and S2 | 0
no murmurs | 0
no thrills | 0
clear breath sounds | 0
symmetric breath sounds | 0
no crackles | 0
no wheezes | 0
no rhonchi | 0
soft abdomen | 0
nondistended abdomen | 0
non-tender abdomen | 0
normal bowel sounds | 0
no organomegaly | 0
good skin turgor | 0
mild cyanosis | 0
no rashes | 0
no lesions | 0
no lower-extremity edema | 0
3+ radial pulses | 0
3+ posterior tibial pulses | 0
3+ dorsalis pedis pulses | 0
Glasgow coma score 8 | 0
sinus tachycardia | 0
normal axis | 0
PR duration 138 milliseconds | 0
no ST or T wave abnormalities | 0
normal chest X-ray | 0
normal CT head scan | 0
white blood cell count 18 600/mm3 | 0
hemoglobin 14.1 g/dL | 0
platelet count 50 000/mm3 | 0
CRP 24.3 MG/DL | 0
lactic acid 3.1 mmol/L | 0
normal chemistry panel | 0
normal renal function | 0
normal liver function | 0
normal electrolytes | 0
blood cultures sent | 0
ceftriaxone 2 grams every 12 h | 0
vancomycin 1 gram every 12 h | 0
initial working diagnosis of meningitis | 0
lumbar puncture not done | 0
thrombocytopenia | 0
intensive care unit | 0
extubated | 24
encephalopathy improved | 24
mechanical ventilation weaning trials | 24
MSSA bacteremia | 0
no skin wounds | 0
no lacerations | 0
no oral lesions | 0
TTE performed | 24
normal TTE results | 24
normal ejection fraction | 24
no valvular heart disease | 24
no vegetations | 24
repeat blood cultures | 72
MSSA bacteremia | 72
new CT chest findings | 72
bilateral diffuse alveolar disease | 72
septic emboli | 72
bilateral pleural effusions | 72
worsening respiratory distress | 72
repeat TTE | 72
no vegetations | 72
TEE performed | 120
moderate mitral regurgitation | 120
30×30 mm vegetation | 120
A1/A2 scallop of the anterior mitral valve leaflet | 120
cardiothoracic surgery consulted | 120
mitral valve replacement | 120
surgery performed | 504
mitral valve deemed irreparable | 504
#31 pericardial tissue valve placed | 504
annular and endocardial debridement | 504
resection of the abscess | 504
blood cultures no growth | 168
IV antibiotics | 0
mental status improved | 600
clinical status improved | 600
discharged | 600