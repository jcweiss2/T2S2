52 years old | 0
caucasian | 0
male | 0
living in western Black Sea region of Turkey | 0
no known past medical history | 0
jaundice | -96
darkening of urine color | -96
fatigue | -96
dyspnea | -96
emergency room visit | 0
computed tomography of the chest | 0
tested for COVID-19 with PCR | 0
COVID-19 PCR test negative | 0
chest CT consistent with COVID-19 pneumonia | 0
tachycardia | 0
heart rate 150 beats per minute | 0
normal blood pressure | 0
respiratory rate 50 breaths per minute | 0
oxygen saturation 80% | 0
15 L of O2 support | 0
admitted to medical ICU | 0
admission laboratory results | 0
diagnostic workup | 0
toxoplasma serology | 0
rubella serology | 0
HSV serology | 0
EBV serology | 0
CMV serology | 0
HIV serology | 0
hantavirus serology | 0
Leptospira serology | 0
ANA | 0
ANCA | 0
anti-dsDNA | 0
haptoglobin | 0
IGG | 0
IGM | 0
IGA | 0
IGE | 0
direct coombs | 0
indirect coombs | 0
complements C3 | 0
complements C4 | 0
peripheral blood smear no schistocytes | 0
abdominal ultrasonography mild hepatomegaly | 0
high-flow nasal cannula | 0
acute hypoxemic respiratory failure | 0
empirical treatment with meropenem | 0
empirical treatment with doxycycline | 0
blood culture pending | 0
femoral central venous catheter insertion | 0
plasmapheresis initiated | 0
severe hyperbilirubinemia | 0
total serum bilirubin more than 13 mg/dL | 0
60 units of fresh frozen plasma used | 0
five sessions of plasmapheresis | 0
total bilirubin dropped to 19.6 mg/dL | 24
Leptospira real-time PCR positive | 96
leptospirosis diagnosis confirmed | 96
medical treatment continued with meropenem | 96
medical treatment continued with doxycycline | 96
significant clinical improvement | 96
stayed in medical ICU for eight days | 192
weaned off oxygen | 192
laboratory values improved | 192
chest X-ray improved | 192
transferred to infectious diseases ward | 192
discharged from hospital | 192
uneventful recovery | 192
no further complications | 192
| Event | Timestamp (hours) |
|-------|-------------------|
| 52 years old | 0 |
| caucasian | 0 |
| male |D0 |
| living in western Black Sea region of Turkey | 0 |
| no known past medical history | 0 |
| jaundice | -96 |
| darkening of urine color | -96 |
| fatigue | -96 |
| dyspnea | -96 |
| emergency room visit | 0 |
| computed tomography of the chest | 0 |
| tested for COVID-19 with PCR | 0 |
| COVID-19 PCR test negative | 0 |
| chest CT consistent with COVID-19 pneumonia | 0 |
| tachycardia | 0 |
| heart rate 150 beats per minute | 0 |
| normal blood pressure | 0 |
| respiratory rate 50 breaths per minute | 0 |
| oxygen saturation 80% | 0 |
| 15 L of O2 support | 0 |
| admitted to medical ICU | 0 |
| admission laboratory results | 0 |
| diagnostic workup | 0 |
| toxoplasma serology | 0 |
| rubella serology | 0 |
| HSV serology | 0 |
| EBV serology | 0 |
| CMV serology | 0 |
| HIV serology | 0 |
| hantavirus serology | 0 |
| Leptospira serology | 0 |
| ANA | 0 |
| ANCA | 0 |
| anti-dsDNA | 0 |
| haptoglobin | 0 |
| IGG | 0 |
| IGM | 0 |
| IGA | 0 |
| IGE | 0 |
| direct coombs | 0 |
| indirect coombs | 0 |
| complements C3 | 0 |
| complements C4 | 0 |
| peripheral blood smear no schistocytes | 0 |
| abdominal ultrasonography mild hepatomegaly | 0 |
| high-flow nasal cannula | 0 |
| acute hypoxemic respiratory failure | 0 |
| empirical treatment with meropenem | 0 |
| empirical treatment with doxycycline | 0 |
| blood culture pending | 0 |
| femoral central venous catheter insertion | 0 |
| plasmapheresis initiated | 0 |
| severe hyperbilirubinemia | 0 |
| total serum bilirubin more than 13 mg/dL | 0 |
| 60 units of fresh frozen plasma used | 0 |
| five sessions of plasmapheresis | 0 |
| total bilirubin dropped to 19.6 mg/dL | 24 |
| Leptospira real-time PCR positive | 96 |
| leptospirosis diagnosis confirmed | 96 |
| medical treatment continued with meropenem | 96 |
| medical treatment continued with doxycycline | 96 |
| significant clinical improvement | 96 |
| stayed in medical ICU for eight days | 192 |
| weaned off oxygen | 192 |
| laboratory values improved | 192 |
| chest X-ray improved | 192 |
| transferred to infectious diseases ward | 192 |
| discharged from hospital | 192 |
| uneventful recovery | 192 |
| no further complications | 192 |
