60 years old | 0
menopausal | 0
postmenopausal bleeding | 0
endovaginal ultrasound | -24
intracavitary image | -24
polyp | -24
hysteroscopy | -24
polyp resection | -24
endometrial biopsy | -24
abdominal pelvic pain | 48
tachycardia | 48
fever | 48
hypotension | 48
diffuse abdominal sensibility | 48
CT scan | 48
desaturation | 48
hypotension | 48
C-reactive protein 360 | 48
blood gases | 48
lactate 4 | 48
intubation | 48
Glasgow coma scale 12 | 48
desaturation | 48
intra-uterine collection | 48
hydroaeric level | 48
increased uterus size | 48
gynecological examination | 48
aspiration of collection | 48
fetid blood | 48
bacteriological samples | 48
blood cultures | 48
antibiotic therapy | 48
imipinem | 48
amikacine | 48
vasoactive drug | 48
noradrenaline | 48
death | 51
bacteriological sampling | 51
blood culture | 51
Escherichia coli | 51
septic shock | 48
hypertension | -120
amlodipine | -120 
menopause | -120*10 
two children | 0 
admitted to recovery room | 48 
discharged | -1