4.5 years old | 0
male | 0
admitted to hospital | 0
disseminated varicella infection | 0
sepsis | 0
secondary staphylococci infection | 0
loss of consciousness | 0
intubated | 0
mechanical ventilatory support | 0
history of chicken pox | -240
treated with antipyretics | -240
treated with antipruritic lotions | -240
no acyclovir treatment | -240
swelling on right forearm | -72
bluish discoloration on right forearm | -72
ulceration on right forearm | -48
high-grade fever | 0
hypotension | 0
severe dehydration | 0
hepatomegaly | 0
abnormal bilateral extensor plantar response | 0
excoriated papules | 0
serohemorrhagic crusts | 0
hemorrhagic necrotic crust | 0
deep ulceration | 0
elevated d-Dimer | 0
elevated fibrinogen | 0
prolonged activated partial thromboplastin time | 0
prolonged protrombine time | 0
elevated white blood cells | 0
thrombocytopenia | 0
elevated alanine aminotransferase | 0
elevated aspartate aminotransferase | 0
elevated creatine kinase | 24
elevated CK-MB | 24
elevated lactate dehydrogenase | 24
elevated sedimantation | 24
elevated C-reactive protein | 24
hematuria | 24
proteinuria | 24
VZV immunglobuline M positive | 0
TORCH panel negative | 0
hepatitis markers negative | 0
anti-HIV negative | 0
diagnosed with purpura fulminans | 0
diagnosed with hepatitis | 0
diagnosed with probable rhabdomyolysis | 0
treated with vancomycin | 0
treated with cefotaxime | 0
treated with acyclovir | 0
topical silver sulfadiazine cream | 0
died | 96