48 years old | 0
female | 0
Roux-en-Y gastric bypass | -18240
Crohn's disease | -18240
rheumatoid arthritis | -18240
atrial fibrillation | -18240
anticoagulation | -18240
septic ascending cholangitis | -72
laparoscopic cholecystectomy | -24
endoscopic retrograde cholangiopancreatography (ERCP) | -24
admitted to intensive care unit | 0
acute tubular necrosis | 0
temporary dialysis | 0
atrial fibrillation with rapid ventricular response | 0
spontaneous rectus sheath hematoma | 0
intravenous heparin | 0
cessation of anticoagulation | 24
blood transfusions | 24
embolization of right inferior epigastric artery | 24
hematoma perforated right lateral wall of bladder | 24
bladder injury not recognized | 24
gross hematuria | 24
pain | 24
leaking around Foley catheter | 24
hematoma induced bladder spasms | 24
persistent lower urinary tract symptoms | 2160
urgency | 2160
frequency | 2160
dysuria | 2160
gross hematuria | 2160
cystoscopy | 2160
large friable right sided bladder mass | 2160
biopsy | 2160
necrotic debris | 2160
rare reactive urothelium | 2160
referred to institution | 2160
Magnetic resonance urography (MRU) | 2160
hematoma decreased in size from 15cm to 10cm | 2160
perforating through right lateral wall of bladder | 2160
transurethral resection (TUR) | 2160
large, smooth, homogeneous bladder mass | 2160
resection to bladder mucosa | 2160
clot extending through bladder wall defect | 2160
bladder diverticulum | 2160
pathology negative for malignancy | 2160
worsening urgency | 3504
terminal voiding pain | 3504
repeat MRU | 3504
further extrusion of hematoma within bladder lumen | 3504
discussion of management options | 3504
repeat TUR | 3504
large organized hematoma protruding from 4 cm cavity | 3504
extensive resection | 3504
entering right lateral wall cavity | 3504
amputating base of hematoma stalk | 3504
visualized healed epithelium | 3504
complete resolution of irritative voiding symptoms | 3504
MRU 13 weeks after second TUR | 5688
hematoma evacuated | 5688
bladder sacculation | 5688
residual hematoma 3.7 cm | 5688
episode of gross hematuria | 14448
UTI | 14448
CT urogram | 14448
thickening right lateral bladder | 14448
tethering to pelvic sidewall | 14448
cystoscopy | 14448
persistent right lateral diverticulum | 14448
well healed epithelium | 14448
