36 years old | 0 | 0 
female | 0 | 0 
pregnant | 0 | 0 
admitted to the hospital | 0 | 0 
recurrent vomiting | -24 | 0 
epigastric pain | -24 | 0 
diagnosed with uterine fibroid | -224 | -168 
weight loss | -672 | 0 
using iron tablets | -672 | 0 
history of weight loss | -672 | 0 
no change in bowel habits | -672 | 0 
no hematemesis or rectal bleeding | -672 | 0 
no history of hematuria or passing stones | -672 | 0 
looked ill | 0 | 0 
markedly dehydrated | 0 | 0 
drowsy | 0 | 0 
blood pressure 126/76 mmHg | 0 | 0 
pulse rate 94 min–1 | 0 | 0 
respiratory rate 30 min–1 | 0 | 0 
temperature 36.6°C | 0 | 0 
no lymphadenopathy | 0 | 0 
no thyromegaly | 0 | 0 
no edema | 0 | 0 
uterus size of 40 weeks | 0 | 0 
tender epigastric area | 0 | 0 
drowsy and hypotonic | 0 | 0 
brisk deep tendon reflexes | 0 | 0 
no obvious focal neurological sign | 0 | 0 
planter reflexes were down-going | 0 | 0 
chest and cardiovascular systems were unremarkable | 0 | 0 
hemoglobin 8.7 g/dl | 0 | 0 
WBCs 7000 μl–1 | 0 | 0 
platelets 445 000 μl–1 | 0 | 0 
ESR 109 mm/h | 0 | 0 
toxic granulation of WBCs | 0 | 0 
BUN 4.4 mmol/l | 0 | 0 
creatinine 59 μmol/l | 0 | 0 
HCO3 22 mmol/l | 0 | 0 
Na 138 mmol/l | 0 | 0 
Ca 4.8 mmol/l | 0 | 0 
uric acid 508 μmol/l | 0 | 0 
lactic acid 1.2 mmol/l | 0 | 0 
phosphorous 0.8 mmol/l | 0 | 0 
HIV serology was negative | 0 | 0 
calcium at 14 weeks’ gestation was 2.43 mmol/l | -448 | -448 
ALT 4 u/l | 0 | 0 
AST 11 u/l | 0 | 0 
ALP 150 u/l | 0 | 0 
total protein 72 g/l | 0 | 0 
albumen 30 g/l | 0 | 0 
cholesterol 4.05 mmol/l | 0 | 0 
triglyceride 3.59 mmol/l | 0 | 0 
PTH 3 pg/ml | 0 | 0 
TSH 0.68 mIU/l | 0 | 0 
free thyroxin 16.6 pmol/l | 0 | 0 
cortisol 1849 nmol/l | 0 | 0 
vitamin D 15 ng/ml | 0 | 0 
given normal saline infusion | 0 | 24 
given intramuscular calcitonin | 0 | 24 
transferred to the medical intensive care unit | 24 | 24 
rupture membrane | 48 | 48 
urgent cesarean section | 48 | 48 
hypercalcemia | -24 | 48 
reduction in the urine output | 48 | 48 
rise in serum creatinine | 48 | 48 
nephrologist was consulted for urgent hemodialysis | 48 | 48 
hemodialysis | 72 | 72 
surgery was complicated by bleeding | 72 | 72 
hypotension | 72 | 72 
required blood transfusion | 72 | 72 
successful delivery of a baby girl | 72 | 72 
removal of uterine masses | 72 | 72 
histopathology report was consistent with leiomyoma with calcifications | 72 | 72 
no evidence of malignancy | 72 | 72 
septicemia | 96 | 96 
septic shock | 96 | 96 
required vasopressors | 96 | 96 
required broad-spectrum antibiotics | 96 | 96 
serum calcium 2.34 mmol/l | 96 | 96 
phosphorus 1.1 mmol/l | 96 | 96 
BUN 6.2 mmol/l | 96 | 96 
Cr 75 mmol/l | 96 | 96 
Na 143 mmol/l | 96 | 96 
K 4.2 mmol/l | 96 | 96 
HCO3 16 mEq/l | 96 | 96 
chloride 113 mEq/l | 96 | 96 
albumin 21 g/l | 96 | 96 
serum lactate 5.19 | 96 | 96 
serum PTH 155 pg/ml | 96 | 96 
serum amylase 88 u/l | 96 | 96 
serum lipase 73 u/l | 96 | 96 
Hb 5.8 g/dl | 96 | 96 
platelets 125 000 μl1 | 96 | 96 
CT scan of the chest and pelvis showed no evidence of mass lesion or organomegaly | 96 | 96 
MRI of the brain showed evidence of infarcts | 96 | 96 
MRA revealed evidence of vasospasm | 96 | 96 
diffuse ischemic changes secondary to hypoxic insult | 96 | 96 
condition began to improve | 120 | 120 
required extensive physiotherapy | 120 | 168 
discharged home | 168 | 168 
final diagnosis of humoral hypercalcemia associated with a uterine fibroid | 168 | 168 
serum calcium remained within the normal range | 168 | 504 
calcium level during pregnancy | -672 | 0 
calcium level after delivery | 0 | 168 
calcium level 6 months after delivery | 504 | 504