57 years old | 0
    woman | 0
    severe rheumatic mitral stenosis | -168
    severe aortic stenosis | -168
    severe tricuspid regurgitation | -168
    implantation of 25 mm mitral On-X valve | 0
    implantation of 19 mm aortic On-X valve | 0
    de Vega tricuspid annuloplasty | 0
    Maze procedure | 0
    cardiopulmonary bypass | 0
    aortic cross-clamp | 0
    chronic atrial fibrillation | -168
    hypertension | -168
    pacemaker placement for sick sinus syndrome | -168
    warfarin use | -168
    no history of bleeding | -168
    preoperative echocardiogram | -168
    preoperative right heart catheterization | -168
    severe pulmonary hypertension | -168
    pulmonary arterial systolic pressures of 75 mmHg | -168
    severe right ventricular dilatation | -168
    intubated | 0
    high infusion rates of inotropic agents | 0
    high infusion rates of vasopressor agents | 0
    epinephrine infusion | 0
    norepinephrine infusion | 0
    vasopressin infusion | 0
    milrinone infusion | 0
    severe hypocoagulable | 0
    thrombocytopenia | 0
    hypofibrinogenemia | 0
    elevated INR levels | 0
    started subcutaneous heparin 5000 IU every 12 h | 192
    deep vein thrombosis prophylaxis | 192
    no antiplatelet therapy | 0
    no therapeutic heparinization | 0
    precarious medical condition | 0
    removal of epicardial pacing wires | 216
    pericardial tamponade | 216
    emergent sternum opening | 216
    worsening pulmonary hypertension | 216
    severe right heart failure | 216
    biventricular failure | 216
    intra-aortic balloon pump placement | 216
    inhalational epoprostenol therapy | 216
    renal failure | 216
    continuous renal replacement therapy | 216
    consumptive thrombocytopenia | 216
    thrombocytopathia | 216
    disseminated intravascular coagulopathy (DIC) | 504
    desmopressin administration | 504
    cryoprecipitate transfusion | 504
    factor VII transfusion | 504
    DIC resolved | 504
    waxing and waning coagulopathy | 504
    waxing and waning thrombocytopenia | 504
    profuse life-threatening bleeding | 1008
    bleeding from respiratory tract | 1008
    bleeding from upper gastrointestinal tract | 1008
    bleeding from natural orifices | 1008
    attempts to initiate anticoagulation | 1008
    prophylactic heparin doses | 1008
    diagnostic bronchoscopy | 1008
    upper gastrointestinal endoscopy | 1008
    lower gastrointestinal endoscopy | 1008
    extensive arteriovenous malformations (AVMs) in respiratory tract | 1008
    extensive arteriovenous malformations (AVMs) in gastrointestinal tract | 1008
    lack of preoperative endoscopy | 1008
    AVMs not restricted to colon | 1008
    difficult definitive diagnosis of Heyde's syndrome | 1008
    possible acquired von Willebrand factor deficiency | 1008
    possible aortic valve patient-prosthetic mismatch | 1008
    no anticoagulation | 0
    frequent transthoracic echocardiograms | 0
    frequent transesophageal echocardiograms | 0
    no valve thrombi | 0
    discharged to long-term acute care facility | 3984
    aspirin use | 3984
    warfarin use | 3984
    subtherapeutic INR of 1.6 | 3984
    higher risk for bleeding | 3984
    no history of thromboembolism | 3984
    no further bleeding episodes | 3984
    died | 3984
    pulmonary aspiration | 3984
    sepsis | 3984
    