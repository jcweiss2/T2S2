33 years old | 0
male | 0
admitted to the hospital | 0
severe anemia | 0
unresponsive to hemotransfusions | 0
increasing doses of erythropoietin | 0
membranoproliferative glomerulonephritis | -1800
treated with steroids | -1800
treated with immunosuppressants | -1800
persistent proteinuria | -1800
microhematuria | -1800
renal biopsy | -1800
membranoproliferative glomerulonephritis with glomerular sclerosis | -1800
mesangiocapillary global proliferation | -1800
no fibrinoid necrosis | -1800
no vascular thrombosis | -1800
no extracapillary proliferation | -1800
Congo red staining for amyloid negative | -1800
immunofluorescence results showed tiny granular deposits | -1800
immunoglobulin G (IgG) positive | -1800
C3 positive | -1800
immunoglobulin A (IgA) negative | -1800
immunoglobulin M (IgM) negative | -1800
C1q negative | -1800
κ and λ light chains negative | -1800
modest accumulation of intravascular fibrinogen | -1800
treated with azathioprine | -1800
treated with mycophenolate | -1800
steroid therapy only | -1800
rapid reduction in proteinuria | -1800
disappearance of microhematuria | -1800
bilateral aseptic necrosis of the femoral head | -720
stopped steroids | -720
slow worsening renal function | -720
mean serum creatinine 2.5 mg/dL | -720
proteinuria 1.5-2 g/24 h | -720
anemia | -720
treated with darbepoetin alfa | -720
severe anemia | 0
hemoglobin 6 g/dL | 0
severe asthenia | 0
dyspnea | 0
hemotransfusion of 2 units of packed red blood cells | 0
colonoscopy | 0
gastroscopy | 0
no significant alterations | 0
peripheral smear | 0
no schistocytes | 0
direct Coombs test negative | 0
indirect Coombs test negative | 0
G6PDH normal | 0
haptoglobin reduced | 0
lactate dehydrogenase increased | 0
autoimmunity normal | 0
persistent slight reduction in C3 | 0
methylprednisolone | 72
azathioprine | 72
low-flow oxygen therapy | 72
anti-glomerular basement membrane (anti-GBM) antibodies negative | 72
C-ANCA negative | 72
P-ANCA negative | 72
transnasal endoscopy | 96
bleeding striae in the first tracheal rings | 96
bronchoscopy | 120
no lesions visible at tracheal level or in both bronchial trees | 120
bronchoalveolar lavage | 120
blood in bronchoalveolar lavage | 120
improvement in clinical picture | 168
improvement in test results | 168
fatigue reduced | 168
dyspnea reduced | 168
oxygen saturation improved | 168
no further transfusions | 168
peripheral oxygen saturation constantly maintained at around 98% | 168
rapid deterioration of renal function | 168
initial filtrate 17 mL/min | 168
reduced to 11 mL/min | 168
increase in blood urea | 168
increase in creatinine values | 168
increase in potassium | 168
increase in phosphorus concentrations | 168
peritoneal dialysis | 240
CT control chest | 480
considerable improvement | 480
spirometry and DLCO test improved | 480
immunosuppressive therapy reduced | 480
discharged | 480
hemoglobin level maintained | 720
average value 11 g/dL | 720
erythropoiesis-stimulating agent doses reduced | 720
automated peritoneal dialysis | 720
moderate mental and physical well-being | 720
no notable disorders | 720
anti-GBM antibodies negative again | 840