27 years old | 0
female | 0
hepatitis C | 0
current IVDU | 0
tricuspid valve replacement | 0
infective endocarditis | 0
surveillance blood cultures positive for methicillin-sensitive Staphylococcus aureus | 0
surveillance blood cultures positive for Candida parapsilosis | 0
gingival hemorrhage | 0
spontaneous bruising | 0
abdominal swelling | 0
supratherapeutic international normalized ratio >10 | 0
thrombocytopenia (12 × 109 μL) | 0
large pericardial effusion | 0
hepatosplenomegaly | 0
mild ascites | 0
nafcillin initiated | 0
amphotericin B initiated | 0
echocardiogram shows large mobile mass involving the tricuspid valve | 0
echocardiogram shows prolapse into the right atrium | 0
echocardiogram shows flail and dehisced tricuspid valve | 0
very large pericardial effusion (4.21 cm posteriorly and 3.73 cm anteriorly) | 0
elevated intrapericardial pressure causing diastolic compression of the right ventricle | 0
ultrasound-guided pericardiocentesis | 24
removal of 600 mL serous fluid | 24
residual moderate effusion | 24
no right ventricular diastolic collapse | 24
nafcillin switched to cefazolin | 24
continued amphotericin B | 24
blood cultures positive for Mycobacteria | 72
amphotericin B discontinued | 72
fluconazole initiated | 72
echocardiogram shows severe tricuspid valve thickening | 72
large vegetation pedunculated and mobile | 72
ruptured tricuspid valve chordae | 72
flail septal leaflet | 72
effusion measures 2.8 cm anteriorly and 3.8 cm posteriorly | 72
some evidence of right ventricular compression without collapse | 72
blood cultures positive for Candida parapsilosis | 168
clinical deterioration with tachycardia | 168
increased dyspnea | 168
abdominal distension | 168
lower extremity edema | 168
persistent fevers | 168
lactic acid elevation | 168
transferred to CICU | 168
echocardiogram shows severe torrential tricuspid regurgitation | 168
flail septal leaflet with echodensity | 168
vegetation attached to tricuspid leaflet no longer visualized | 168
embolization suspected | 168
cefazolin switched to liposomal amphotericin B | 168
fluconazole switched to amikacin | 168
fluconazole switched to imipenem | 168
fluconazole switched to azithromycin | 168
continued clinical deterioration requiring intubation | 192
pressors initiated | 192
severe metabolic acidosis (lactic acid 19, pH 7.27) | 216
signs of multiorgan failure | 216
emergent tricuspid valve replacement | 216
redo sternotomy | 216
tricuspid valve replaced with Biocor valve | 216
removal of embolized CorMatrix valve from right pulmonary artery | 216
blood cultures positive for Mycobacterium | 216
switched to micafungin | 216
continued amikacin | 216
continued imipenem | 216
continued azithromycin | 216
patient discharged home | 672
pulmonary embolism | -432
Coumadin initiated | -432
intravenous drug use | -2160
tricuspid valve endocarditis | -2160
bacteraemia (Candida and Staphylococcus aureus) | -2160
treated with vancomycin | -2160
treated with daptomycin | -2160
treated with linezolid | -2160
treated with cefepime | -2160
treated with micafungin | -2160
CorMatrix extracellular-based material tricuspid valve replacement | -2160
post-operative pulmonary embolism | -2160
Coumadin initiated | -2160
completed 6-week course of antibiotics | -2160
recurrent IVDU | -432
positive blood cultures for AFB | 720
TEE reveals new tricuspid valve vegetations | 720
treated with linezolid | 720
treated with imipenem | 720
lost to follow-up | 720
