liver cirrhosis | -72
hepatocellular carcinoma | -72
admission | 0
intravenous glycoppyrolate administration | 0
general anesthesia induction | 0
intubation | 0
mechanical ventilation | 0
stable vital signs | 0
hepatectomy with CUSA | 0
sudden decrease in arterial blood pressure | 1
tachycardia | 1
ST elevation on EKG | 1
resuscitation with colloid and catecholamines | 1
diagnosis of VAE and PAE | 1
intraoperative ultrasonography | 1
arterial blood gas analysis | 1
catecholamine administration | 1.17
restoration of end-tidal carbon dioxide | 1.5
norepinephrine infusion | 1.5
fluid resuscitation | 1.5
disappearance of air emboli from left heart | 2.17
completion of hepatectomy | 2.17
end of surgery | 5
intensive care unit admission | 5
mechanical ventilation | 5
norepinephrine infusion | 5
abnormal PT/PTT | 5
abnormal fibrinogen | 5
abnormal d-dimer | 5
abnormal antithrombin III | 5
abnormal CK-MB | 5
abnormal troponin-T | 5
ST elevation on EKG | 5
recovery of EKG findings | 24
trans-thoracic echocardiogram | 24
tapering out norepinephrine infusion | 24
unchanged mental status | 120
brain CT | 120
brain MRI | 120
multiple acute cerebral infarctions | 120
weaning to spontaneous ventilation | 264
extubation | 264
unstable vital signs | 360
intravenous administration of catecholamines | 360
panperitonitis | 360
cardiac arrest | 744
death | 744