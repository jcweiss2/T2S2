48 years old | 0
male | 0
chronic renal failure | 0
ischemic stroke | 0
insulin-dependent diabetes | 0
fever | -96
malaise | -96
oliguria | -96
haematuria | -96
nausea | -96
vomiting | -96
febrile | 0
blood pressure normal | 0
abdomen depressible | 0
painful prostate | 0
leukocytosis | 0
renal failure | 0
high C-reactive protein | 0
hyperglycemia | 0
acidosis | 0
positive acetonuria | 0
male urinary tract infection suspected | 0
diabetic ketoacidosis suspected | 0
emphysematous lesions in prostate | 0
emphysematous lesions in seminal vesicles | 0
normal kidneys | 0
no dilatation of excretory cavities | 0
empirical intravenous antibiotics administered | 0
cefotaxime | 0
ciprofloxacine | 0
suprapubic catheterization | 0
Enterobacter cloacae isolated | 0
imipeneme | 0
apyretic | 72
aggravation of biological inflammatory syndrome | 72
increase of white blood cells | 72
increase of CRP | 72
severe metabolic acidosis | 72
emergency hemodialysis | 72
prostatic hydroaeric collections | 72
trans-rectal aspiration | 72
purulent liquid | 72
same germ isolated | 72
generalized convulsive seizures | 96
regression of biological inflammatory syndrome | 96
white blood cells decreased | 96
CRP decreased | 96
correct metabolic balance | 96
chronic renal failure | 96
head CT scan normal | 96
seizures attributed to antibiotics | 96
antibiotics changed | 96
piperacillin | 96
flagyl | 96
worsening of patient's state of consciousness | 336
septic shock | 336
transfer to intensive care department | 336
orotracheal intubation | 336
norepinephrine | 336
multi-organ failure | 336
death | 336