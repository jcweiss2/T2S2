39 years old | 0
male | 0
admitted to the hospital | 0
arterial hypertension | -8760
atypical chest pain | 0
blood pressure 180/110 mm Hg | 0
heart rate of 74 beats per minute | 0
loud systolic murmur at the base of the heart | 0
no symptoms of heart failure | 0
ECG showed sinus rhythm 73 beats per minute | 0
left ventricle hypertrophy (LVH) | 0
negative T waves in II, III, aVF | 0
coronary angiography | 0
atherosclerotic lesions | 0
maximum luminal diameter stenosis was 30–40% in the right coronary artery (RCA) | 0
troponin I level was detectable but not significantly elevated | 0
D-dimer level was elevated | 0
BAV with degenerative changes and calcifications | 0
aortic stenosis with the mean pressure gradient of 45 mm Hg | 0
mild aortic regurgitation | 0
concentric left ventricle hypertrophy | 0
maximum wall thickness up to 1.7 cm | 0
normal left ventricle systolic function (LVEF 65%) | 0
ascending aorta diameter was 5.6 cm | 0
thoracic aortic aneurysm (TAA) | 0
chronic pancreatitis | 0
type C chronic viral hepatitis | 0
hyperlipidemia | 0
refused to undergo surgery | 0
pharmacological treatment | 0
β-blocker | 0
angiotensin-converting enzyme inhibitor (ACEI) | 0
diuretic | 0
atorvastatin | 0
acetylsalicylic acid (ASA) | 0
cerebrovascular event | -876
aphasia of sudden onset | -876
hospitalization in a Department of Neurology | -876
echocardiography | -876
ultrasonography of cervical arteries | -876
calcified but not dissected | -876
abrupt onset of chest pain | 1092
severe retrosternal pain | 1092
radiated to the left upper limb | 1092
blood pressure 163/98 mm Hg | 1092
blood pressure 135/93 mm Hg | 1092
heart rate of 65 beats per minute | 1092
ECG showed sinus rhythm 72/min | 1092
LVH features with negative T waves in II, III, aVF and V3–V6 | 1092
troponin I level was mildly elevated | 1092
D-dimer level was elevated | 1092
acute aortic dissection (AAD) | 1092
bedside transthoracic echocardiography (TTE) | 1092
dissection flap in the dilated ascending aorta | 1092
CT confirmed BAV and dilatation of the ascending aorta | 1092
aortic dissection with intimal tear | 1092
Bentall procedure | 1096
total aortic root replacement | 1096
St Jude Medical 29 mm conduit | 1096
aortic valve | 1096
aortic root | 1096
ascending aorta | 1096
re-implantation of the coronary arteries | 1096
Datascope 22 mm prosthesis | 1096
distal part of the ascending aorta | 1096
postoperative day 1 | 1097
extubated | 1097
postoperative day 4 | 1100
fever of 39°C | 1100
septic shock | 1100
multiorgan failure | 1100
mediastinum was drained | 1100
empiric wide-spectrum antibiotic therapy | 1100
died on the 8th postoperative day | 1104
cardiopulmonary insufficiency | 1104