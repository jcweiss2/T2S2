59 years old | 0
African American woman | 0
hypertension | 0
hyperlipidemia | 0
type 2 diabetes mellitus | 0
end-stage renal disease | 0
diabetes mellitus nephropathy | 0
admitted to the hospital | 0
altered mental status | -8
bizarre behavior | -8
slow irrational speech | -8
delusions | -8
abnormal movements | -8
more somnolent than usual | -8
headaches | -72
worsening dyspnea | -72
dialysis scheduled | -24
altered mental status (dialysis) | -24
agitation | -24
automatisms | -24
hand movements | -24
head movements | -24
orofacial movements | -24
hypertensive (BP 160/63 mmHg) | 0
restless | 0
stereotypical movement of head turning | 0
staring | 0
nonsensical involuntary movements | 0
oriented to person infrequently | 0
not oriented to time | 0
not oriented to place | 0
could not follow commands | 0
responded inappropriately | 0
incomprehensible sounds | 0
Glasgow Coma Scale (GCS) 8/15 | 0
no focal weakness | 0
no facial droop | 0
no signs of meningeal irritation | 0
bibasilar rales | 0
altered mental status secondary to metabolic vs toxic encephalopathy | 0
CT scan of the head unremarkable | 0
chest X-ray cardiomegaly | 0
bilateral infiltrates suspicious for pulmonary edema | 0
toxicology screen negative | 0
blood ethanol level <10 mg/dl | 0
sodium 145 mEq/L | 0
potassium 5.1 mEq/L | 0
chloride 102 mEq/L | 0
bicarbonate 21 mmol/l | 0
glucose 197 mg/dl | 0
alkaline phosphatase 102 U/L | 0
alanine aminotransferase 76 U/L | 0
aspartate aminotransferase 43 mg/dl | 0
calcium 9.8 mg/dl | 0
magnesium 2.3 mg/dl | 0
BUN elevated 45 mg/dl | 0
creatinine elevated 8.2 mg/dl | 0
white counts 7800 cell/mcl | 0
hemoglobin 12.7 g/dl | 0
platelets 123000 cells/mcl | 0
C-reactive protein elevated 4.99 mg/dl | 0
ferritin elevated 1581 ng/ml | 0
ANA unremarkable | 0
anti-double stranded DNA unremarkable | 0
ANCA unremarkable | 0
RF unremarkable | 0
troponin mildly elevated | 0
pro-brain natriuretic peptide mildly elevated | 0
ECG normal sinus rhythm | 0
premature ventricular complexes | 0
confused | 24
not obeying commands | 24
no purposeful movements | 24
GCS 7/15 | 24
BP 190-210/70(100 mmHg | 24
episodes of severe agitation | 24
BUN trended up 70 mg/dl | 24
creatinine trended up 11.0 mg/dl | 24
nasogastric tube placed | 24
hydralazine started | 24
labetalol started | 24
hemodialysis on day 2 | 24
hemodialysis sessions days 3-10 | 72
BUN ranged 17-63 mg/dl | 72
clonidine added | 72
BP ranged 160-210/65-120 mmHg | 72
episodes of hypotension | 72
antihypertensive medications withheld | 72
repeat CT scan unremarkable | 168
CSF white counts elevated | 168
CSF protein elevated | 168
oligoclonal band negative | 168
EEG epileptiform discharges | 240
intravenous levetiracetam 1 g | 240
levetiracetam 250 mg twice daily | 240
levetiracetam after hemodialysis | 240
more alert | 264
oriented | 264
following verbal commands | 264
GCS improved 13/15 | 264
lethargic | 312
febrile | 312
BP 188/110 mmHg | 312
white counts elevated 25000 cells/mcL | 312
neutrophilia | 312
chest X-ray atelectatic changes | 312
CSF cell count unremarkable | 312
CSF protein unremarkable | 312
CSF glucose unremarkable | 312
blood cultures obtained | 312
urine cultures obtained | 312
CSF cultures obtained | 312
CSF viral panel PCR obtained | 312
CSF encephalopathy markers obtained | 312
transferred to ICU | 312
meropenem commenced | 312
acyclovir commenced | 312
repeat EEG diffuse encephalopathy | 360
MRI brain PRES findings | 360
continuous cardiopulmonary monitoring | 360
labetalol continuous infusion | 360
BP control goal <150/90 mmHg | 360
CSF viral panel PCR negative | 360
autoimmune encephalopathy markers negative | 360
acyclovir discontinued | 360
meropenem continued | 360
cultures negative | 360
leukocytosis resolution | 360
completely alert | 480
oriented | 480
obeying commands | 480
GCS 15/15 | 480
BP <150/80 | 480
regular hemodialysis | 480
outpatient antihypertensive regimen | 480
repeat MRI increased hemorrhage and encephalomalacia | 480
discharged | 480
modified Rankin scale 4 | 480
neurologist follow-up | 1440
repeat MRI residual brain abnormalities | 1440
long-term levetiracetam | 1440
