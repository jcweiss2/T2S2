70 years old | 0
male | 0
emergency esophageal diversion | -720
injury to the cervical esophagus | -720
spinal surgery | -720
gastric pull-up procedure | -504
postoperative anastomotic leakage | -504
endoscopy | -504
esophageal stent | -504
local cervical infection | -504
sepsis | -504
arterial hypertonus | 0
non-active smoking status | 0
ischemic stroke | 0
incomplete senso-motoric hemiparesis | 0
thyroidectomy | 0
open prostatectomy | 0
prostate cancer | 0
malnutrition | 0
systemic inflammation | 0
jugular phlegmon | 0
cervical phlegmon | 0
hemoglobin level of 6.7 g/dL | 0
white blood cell count of 6400 cells/μL | 0
platelet count of 210 × 10^3/μL | 0
creatinine level of 0.76 mg/dL | 0
unremarkable liver and cholestasis parameters | 0
albumin level of 2.8 g/dL | 0
chest computed tomography scan | 0
endoscopy | 0
dislodged esophageal stent | 0
esophageal perforation | 0
infected cavity | 0
esophageal stenosis | 0
stent removal | 0
endoscopic vacuum therapy | 24
EsoSponge system | 24
jugular and cervical phlegmon resolved | 336
repeated endoscopic balloon dilatation | 336
subtotal esophageal resection | 720
reconstruction using a free-jejunal graft interposition | 720
CT angiography | 720
partial sternotomy | 720
laparotomy | 720
jejunal segment harvested | 720
left carotid artery and left jugular vein used as recipient vessels | 720
graft implanted in an isoperistaltic position | 720
cervical anastomosis performed in an end-to-end fashion | 720
upper mediastinal gastro-jejunostomy performed in a side-to-side fashion | 720
upper sternum resected | 720
soft tissue defect covered with a sternocleidomastoid muscle flap | 720
abdominal reconstruction achieved by an end-to-end jejunojejunostomy | 720
postoperative course uneventful | 720
oral alimentation reestablished | 720
daily speech therapy | 720
anastomotic healing confirmed radiologically and endoscopically | 720
patient transferred to a rehabilitation clinic | 720
discharged | 720