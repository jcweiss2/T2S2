57 years old|0
    woman|0
    visual disturbance|0
    diplopia|0
    headaches|0
    visited another hospital|-10320
    MRI showing osteolytic, irregular enhancing lesion occupying the clivus|-10320
    T1-weighted gadolinium-enhanced images|-10320
    TSS|-10320
    excisional biopsy consistent with chordoma with chondroid differentiation|-10320
    not totally removed|-10320
    presented with diplopia again|-8760
    MRI showing clival chordoma increased in size|-8760
    extended TSS|-8640
    tumor still remained|-8640
    postoperative CSF leakage not observed|-8640
    tumor increased again|-6720
    Gamma knife radiosurgery|-6720
    treatment dose 18.5 Gy at tumor margin|-6720
    proton beam radiotherapy|-3120
    treatment dose 6960 cGy in 29 fractions|-3120
    presented with unpleasant odor inside nasal cavity|-2760
    visited radiation-oncology department several times|-2760
    took antibiotic drugs|-2760
    took steroids|-2760
    symptoms did not resolve|-2760
    visited emergency medical team|0
    copious epistaxis|0
    odor inside nasal cavity|0
    systemic inflammatory response syndrome|0
    body temperature 38.2 degrees|0
    WBC 30040/mm3|0
    imaging study to identify cause of epistaxis|0
    brain CT scan|0
    comatose mental state|0
    low blood pressure due to septic shock|0
    cardiopulmonary resuscitation|0
    vital signs recovered|0
    subsequent CT did not reveal cause of comatose mental state|0
    further evaluations in intensive care unit|0
    CSF examination by lumbar puncture|0
    MRI without enhanced gadolinium|0
    exploration inside nasal cavity with nasal endoscope|0
    synthetic materials in reconstruction of sellar floor|0
    nasal septum defect due to necrosis|0
    pale and fibrotic mucous membrane due to radiotherapy|0
    scarring and narrowing of blood vessels|0
    disruption and necrosis of mucous membrane|0
    CSF rhinorrhea not observed|0
    Enterococcus avium identified on mucosal culture|0
    Escherichia coli identified on mucosal culture|0
    CSF examination revealed increased WBC count 11280 cells/mm3|0
    CSF examination revealed protein level 345 mg/dL|0
    CSF examination revealed glucose level 4 mg/dL|0
    Enterococcus avium identified on CSF culture|0
    Escherichia coli identified on CSF culture|0
    Enterococcus avium identified on blood culture|0
    Escherichia coli identified on blood culture|0
    diagnosed with bacterial meningitis|0
    administered antibiotic therapy|0
    expired|168
    MRI follow-up in May 2011|-6720
    MRI follow-up in December 2012|-3120
    presented with sinusitis in December 2010|-8640
    prolonged steroid therapy|-2760
    chronic sinusitis|-2760
    sellar floor reconstruction with synthetic materials|-8640
    fulminant sinusitis|-2760
    delayed wound healing|-2760
    nasal septum defect|0
    synthetic materials in sellar floor reconstruction|0
    sinusitis worsened and infected adjacent mucosal membranes|0
    delayed bacterial meningitis|168
    fatal meningitis|168
    