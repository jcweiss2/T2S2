55 years old| 0
    male| 0
    admitted to emergency department| 0
    dyspnea| -24
    fever| -168
    cough| -168
    whitish sputum| -168
    former smoker| -168
    history of 5-pack-year| -168
    no alcohol abuse history| 0
    no known history of pulmonary diseases| 0
    no underlying diseases| 0
    no diabetes| 0
    no medications| 0
    no herbal medicines| 0
    admitted to coronary care unit| -72
    atypical chest pain| -72
    normal coronary angiography| -72
    chest radiography| -72
    normal chest radiograph| -72
    chest computed tomography| -72
    diffuse bronchial wall thickening| -72
    no evidence of emphysema| -72
    flu-like symptoms| -168
    fever| -168
    cough| -168
    sore throat| -168
    myalgia| -168
    conservative medication| -168
    no antiviral agents| -168
    blood pressure 130/90 mm Hg| 0
    heart rate 113 beats/min| 0
    respiratory rate 26 breaths/min| 0
    body temperature 37.8℃| 0
    conscious| 0
    acute ill-looking appearance| 0
    normal conjunctiva| 0
    no palpable lymph nodes| 0
    bilateral expiratory wheezes| 0
    white blood cells 15,200/mm3| 0
    neutrophils 84.9%| 0
    lymphocytes 8.6%| 0
    eosinophils 0.5%| 0
    hemoglobin 16.0 g/dL| 0
    platelets 144,000/mm3| 0
    C-reactive protein 46.5 mg/L| 0
    normal liver function tests| 0
    normal renal function tests| 0
    negative serologic tests for autoantibodies| 0
    negative rheumatoid factor| 0
    negative HIV test| 0
    negative VDRL test| 0
    normal CD4 count| 0
    arterial blood gas analysis| 0
    pH 7.45| 0
    PaO2 81.8 mm Hg| 0
    PaCO2 38.5 mm Hg| 0
    rapid influenza diagnostic test negative| 0
    negative anti-mycoplasma antibody| 0
    negative Legionella urinary antigen| 0
    negative pneumococcus urinary antigen| 0
    negative sputum culture| 0
    negative blood culture| 0
    negative acid-fast bacilli stain| 0
    positive serum galactomannan assay| 48
    chest radiograph bilateral infiltrates| 0
    chest CT patchy consolidations| 0
    ground-glass opacities| 0
    centrilobular nodules| 0
    prescribed ceftriaxone| 0
    prescribed clarithromycin| 0
    suspected community-acquired pneumonia| 0
    suspected acute exacerbation of asthma| 0
    initiated methylprednisolone 62.5 mg/day| 48
    no history of asthma| 0
    switched to piperacillin/tazobactam| 96
    switched to levofloxacin| 96
    worsening leukocytosis| 96
    hypoxemia| 96
    developed respiratory failure| 96
    transferred to ICU| 96
    mechanically ventilated| 96
    fever subsided| 96
    C-reactive protein declined to 6.6 mg/L| 96
    chest radiographic improvement| 192
    negative gram stain| 96
    negative tracheal aspiration culture| 96
    clinical deterioration| 216
    high fever| 216
    worsening chest radiograph| 216
    bronchoscopy| 216
    yellow-whitish exudative pseudomembranes| 216
    airway narrowing| 216
    acute-angle branching hyphae observed| 216
    BAL culture Aspergillus species| 216
    positive repeat serum galactomannan| 216
    PCR positive for influenza B| 216
    diagnosed probable IPA| 216
    initiated voriconazole| 216
    progressive worsening| 336
    death| 336
    