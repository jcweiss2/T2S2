30 years old | 0
male | 0
admitted to the hospital | 0
paralysis of both legs | -336
skin getting darker | -336
pain and darkening of the scrotum and penis | -336
strained waist | -336
felt very weak | -335
loss of urge to urinate and defecate | -335
bedwetting | -335
no haematuria | -336
no cloudy urine | -336
local bluish on the both legs | 0
diminished circulation to the lower part of the body | 0
necrosis from the penis to the scrotum | 0
hyperaemia without pus or active bleeding | 0
FC 16 French was placed | 0
normal urine production | 0
systemic infections | 0
WBC reached 27.000 per mm | 0
acute limb ischemia | 0
penile necrosis | 0
aorta thoracoabdominal CT Scan with contrast | 24
dissection from the aortic arch to the abdominal aorta | 24
intimal tear at the level of the aortic arch | 24
thrombus in the false lumen of the abdominal aorta | 24
occlusion of the distal abdominal aorta | 24
collateralization in the common bilateral femoral artery | 24
Thoracic Endovascular Aortic Repair (TEVAR) | 48
open thrombectomy | 48
unconscious | 48
put on ventilator | 48
debridement and amputation | 96
debridement of the penis and scrotum | 96
amputation above the knee procedure | 96
urinary diversion with percutaneous cystostomy | 96
necrotic tissue from the glans penis, penile shaft, and scrotum was removed | 96
septic shock | 192
multiorgan dysfunction | 192
died | 192