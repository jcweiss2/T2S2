64 years old | 0
male | 0
admitted to the ICU | 0
Escherichia coli Gram-negative septic shock | 0
purulent peritonitis | 0
rectosigmoid junction adenocarcinoma | 0
slightly disoriented | 0
hypotensive | 0
blood pressure of 110/55 mmHg | 0
lactic acidosis | 0
elevated white blood cell count | 0
WBC of 22680/μL | 0
PCT of 10 ng/mL | 0
renal insufficiency | 0
elevated creatinine of 1.88 mg/dL | 0
hyperglycemia of 263 mg/dL | 0
lactic acidosis | 0
base excess of -8.1 mmol/L | 0
lactate of 2 mmol/L | 0
fluids resuscitation | 0
crystalloids | 0
albumin | 0
broad-spectrum antibiotics | 0
meropenem | 0
metronidazole | 0
insulin | 0
invasive monitoring | 0
Vigileo monitor | 0
emergency surgical intervention | 0
intestinal subocclusions | 0
sepsis | 0
rectosigmoid palliative resection | 0
peritoneal lavage | 0
drainage | 0
bacteriological samples | 0
intubated | 0
mechanically ventilated | 0
febrile | 24
persistent leukocytosis | 24
WBC of 20090 /μL | 24
elevated PCT levels | 24
septic encephalopathy | 24
GCS of 10 points | 24
vasoactive support | 24
noradrenaline | 24
cardiac output of 7.3 L/min | 24
cardiac index of 3.1 L/min/m2 | 24
systemic vascular resistance index of 1897 dyn*s/cm5*m2 | 24
SOFA score of 10 points | 24
APACHE II score of 23 points | 24
blood cultures | 24
urine cultures | 24
vancomycin | 24
fluconazole | 24
extracorporeal endotoxin adsorption treatment | 24
Alteco LPS Adsorber | 24
double lumen 12Fr catheter | 24
unfractionated heparin | 24
haemofiltration | 24
blood flow rate of 150 ml/min | 24
duration of treatment of 120 minutes | 24
improvement in hemodynamic status | 48
reduction in noradrenaline infusion rate | 48
increase in MAP | 48
increase in CI | 48
reduction in PCT levels | 48
reduction in lactate levels | 48
decrease in SOFA score | 48
postoperative complication | 168
localised peritonitis | 168
ischemic bowel perforation | 168
death | 192
multiple organ failures | 192