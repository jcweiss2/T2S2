\boxed{70 years old| 0
male | 0
farmer | 0
admitted to the emergency department | 0
high-grade fever | -120
generalized body ache | -120
headache | -120
altered sensorium | -24
joint pains | -120
epigastric pain | -120
no other comorbidities | 0
no history of drug addiction | 0
no history of intoxication | 0
inguinal lymphadenopathy | 0
mild generalized rash | 0
no eschar | 0
hemodynamically stable | 0
disoriented | 0
no focal neurological deficit | 0
no neck rigidity | 0
provisional diagnosis of acute febrile illness | 0
workup for tropical infections | 0
negative for malaria | 0
negative for dengue | 0
negative for typhoid | 0
negative for leptospira | 0
positive scrub typhus antigen card | 0
positive scrub IgM | 0
sterile blood and body fluid cultures | 0
leukocytosis | 0
mild hyperbilirubinemia | 0
transaminitis | 0
slightly raised INR | 0
negative viral markers for hepatitis B | 0
negative viral markers for hepatitis C | 0
mild fatty infiltration of the liver | 0
treated with doxycycline | 0
defervescence | 48
improved orientation | 48
weakness of lower limbs | 96
weakness progressed to upper limbs | 120
absent deep tendon reflexes | 120
flexor plantar responses | 120
bladder incontinence | 120
no bowel incontinence | 120
shifted to ICU | 120
breathing difficulty | 120
respiratory distress | 120
intubated | 120
mechanical ventilation | 120
MRI brain without abnormality | 120
MRI cervical spine without abnormality | 120
NCV showed demyelinating polyneuropathy | 120
diagnosis of GBS | 120
CSF analysis | 120
started on IV immunoglobulin therapy | 120
added rifampicin for meningoencephalitis | 120
improvement in limb weakness | 168
improvement in respiratory parameters | 168
weaned off ventilator | 168
extubated | 168
oral feeding started | 168
aggressive limb and chest physiotherapy | 168
shifted out from ICU | 168
discharged from hospital | 672
full neurological recovery | 672
follow-up in outpatient department | 672
no functional disability | 672}