18 years old| 0
male | 0
admitted to the hospital | 0
fever | -72
rash | -72
acne |  -672
minocycline |  -672
increased WBC count | 0
eosinophilia| 0
systemic involvement| 0
diffuse erythematous or maculopapular eruption| 0
pruritis | 0
DRESS syndrome | 0
fever persisted | 0
rash persisted | 0
discharged | 24
Separate conjunctive phrases into its component events and assign them the same timestamp (for example, the separation of 'fever and rash' into 2 events: 'fever' and 'rash')  If the event has duration, assign the event time as the start of the time interval. Attempt to use the text span without modifications except 'history of' where applicable. Include all patient events, even if they appear in the discussion; do not omit any events; include termination/discontinuation events; include the pertinent negative findings, like 'no shortness of breath' and 'denies chest pain'.  Show the events and timestamps in rows, each row has two columns: one column for the event, the other column for the timestamp.  The time is a numeric value in hour unit. The two columns are separated by a pipe '|' as a bar-separated file. Skip the title of the table. Reply with the table only. Create a table from the following case:
<|eot_id|><|start_header_id|>user<|end_header_id|>
<|eot_id|><|start_header_id|>assistant<|end_header_id|>
73 years old | 0
myocardial infarction | -744
percutaneous coronary intervention | -744
stent insertion | -744
chills | -72
anorexia | -72
nausea | -72
diarrhea | -72
oxygen saturation 85% at room air | -72
HRCT chest showing ground-glass opacity | -72
admitted to COVID-19 ward | 0
therapeutic regimen for COVID-19 | 0
Tamiflu (Oseltamivir) | 0
hydroxychloroquine | 0
KALETRA (lopinavir/ritonavir) | 0
levofloxacin | 0
linezolid | 0
RT-PCR positive for COVID-19 | 0
breathing became harder | 24
oxygen saturation 94% with nasal cannula | 24
