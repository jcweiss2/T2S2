44 years old | 0  
    female | 0  
    hypothyroidism | 0  
    major depressive disorder | 0  
    electroconvulsive therapy | 0  
    intermittent headache | -48  
    progressive memory loss | -48  
    MRI showing enhancing lesion in right temporal lobe | -72  
    craniotomy with gross total resection | -24  
    WHO Grade III anaplastic astrocytoma diagnosis | -24  
    immunohistochemical stain positive for mutant IDH-1 | -24  
    widespread loss of ATRX | -24  
    strong p53 reactivity | -24  
    Ki-67 of 50% | -24  
    fluorescence in-situ hybridization showing loss of 19q | -24  
    polysomy of chromosome 1 | -24  
    initial CBC: Hgb 11.9 g/dL | -24  
    initial CBC: WBC 6.9 × 103/μL | -24  
    initial CBC: ANC 1.5 × 103/μL | -24  
    initial CBC: ALC 1.4 × 103/μL | -24  
    initial CBC: PLT 370 × 103/μL | -24  
    Karnofsky performance status 90% | 0  
    radiation therapy (5940 cGy in 33 fractions) | 0  
    temozolomide 75 mg/m2 | 0  
    grade-1 skin toxicity | 0  
    gastritis | 0  
    topical steroid cream | 0  
    ranitidine | 0  
    levetiracetam 500 mg daily | 0  
    levetiracetam discontinued after third cycle | 72  
    lymphopenia | 72  
    thrombocytopenia | 72  
    ALC 0.2 × 103/μL | 72  
    PLT 109 × 103/μL | 72  
    adjuvant temozolomide 150 mg/m2 for 6 cycles | 72  
    atovaquone started | 72  
    low CD4+ T-cell count | 72  
    allergy to sulfa drugs | 72  
    CBC prior to adjuvant TMZ: Hgb 9.3 | 72  
    CBC prior to adjuvant TMZ: WBC 3.2 | 72  
    CBC prior to adjuvant TMZ: PLT 248 | 72  
    CBC prior to adjuvant TMZ: ANC 2.4 | 72  
    CBC prior to adjuvant TMZ: ALC 0.2 | 72  
    neutropenia at 1 month follow-up | 432  
    WBC 1 | 432  
    ANC 0.6 | 432  
    ALC 0.1 | 432  
    Hgb 11.3 | 432  
    PLT 134 | 432  
    weekly CBC showing rapid decrease in WBC and PLT | 432  
    WBC 0.6 | 432  
    Hgb 9.3 | 432  
    PLT 11 | 432  
    emergency department presentation | 576  
    dyspnea | 576  
    rash | 576  
    paronychia | 576  
    severe pancytopenia | 576  
    WBC 0.1 | 576  
    ANC 0 | 576  
    ALC 0 | 576  
    Hgb 7.1 | 576  
    PLT 16 | 576  
    platelet transfusions | 576  
    red blood cell transfusions | 576  
    cefuroxime course | 576  
    fluconazole course | 576  
    cellulitis | 576  
    atovaquone discontinued | 576  
    bone marrow biopsy showing hypocellular marrow | 576  
    HIV negative | 576  
    HBV negative | 576  
    HCV negative | 576  
    EBV negative | 576  
    CMV negative | 576  
    parvovirus negative | 576  
    B12 204 pmol/L | 576  
    B12 supplementation | 576  
    neutropenic fever | 1296  
    septic shock | 1296  
    Bartholin gland abscess | 1296  
    rectovaginal fistula | 1296  
    WBC 0.00 | 1296  
    Hgb 7.3 | 1296  
    PLT 11 | 1296  
    abscess drainage | 1296  
    broad-spectrum antibiotics | 1296  
    Enterococcus VRE bacteremia | 1296  
    repeat bone marrow biopsy showing pan-hypoplasia | 1296  
    aplastic anemia diagnosis | 1296  
    granulocyte monocyte-colony stimulating factor | 1296  
    eltrombopag | 1296  
    cord blood stem cell transplantation | 1296  
    fludarabine conditioning | 1296  
    melphalan conditioning | 1296  
    lung abscesses | 1296  
    pyelonephritis | 1296  
    acute hypoxic respiratory failure | 1296  
    ICU transfer | 1296  
    death due to septic shock | 1296  
    multiple organ failure | 1296  

