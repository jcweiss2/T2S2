83 years old | 0
man | 0
brought to the emergency facility | 0
dislodgment of gastrostomy feeding tube | -24
underwent gastrostomy | -6480
swallowing disorder acquired after acute ischemic stroke | -6480
Stamm's technique | -6480
stoma was stenotic | -6480
dilated | -6480
new tube inserted through original orifice | -6480
discharged | -6480
experienced abdominal pain | -24
experienced vomiting | -24
returned to the hospital | -24
ill-looking patient | 0
dehydrated | 0
hypotension | 0
tachycardia | 0
abdomen distended | 0
abdomen diffusely tender | 0
left hypochondrium and flank tenderness | 0
abdominal computed tomography | 0
iodine contrast medium infusion through gastrostomy tube | 0
cavity formed by peritoneal blockade filled by gas and fluid | 0
exploratory laparotomy | 0
significant amount of lumpy liquid in peritoneal cavity | 0
peritoneal adhesions between loops and abdominal wall | 0
false path at gastrostomy site | 0
purulent collection adjacent to stomach | 0
another gastrostomy performed | 0
stomach sutured to abdominal wall | 0
peritoneal cavity lavage with saline | 0
abdomen drained | 0
referred to intensive care unit | 0
evisceration requiring re-operation | 0
multiple organ failure | 0
died | 1032
peritonitis | 0
septicemia | 0
death | 1032
1. Patient is 83 years old | 0
2. Male | 0
3. Brought to emergency facility (admission) | 0
4. Dislodgment of gastrostomy tube | -24 (day before admission)
5. Gastrostomy (Stamm's technique) 9 months ago | -6480
6. Swallowing disorder after acute ischemic stroke | -6480
7. Stoma was stenotic | timestamp? This happened 9 months ago? No, the stoma became stenotic after the initial gastrostomy. But in the case report, when he presented with the dislodged tube, the stoma was stenotic, so during the initial admission (0), they dilated it. So the stoma being stenotic is at 0.
