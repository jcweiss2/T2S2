30 years old | 0
female | 0
IVDU | -672
admitted to the hospital | 0
bacterial pneumonia | 0
IE suspected | 0
septic pulmonary emboli | 0
transesophageal echocardiography (TEE) performed | 0
IE confirmed | 0
ravaged TV with fenestrations | 0
wide-open tricuspid regurgitation | 0
flail segments | 0
multiple mobile TV vegetations | 0
left ventricular ejection fraction preserved | 0
multidisciplinary management | 0
cardiology consultation | 0
cardiac surgery consultation | 0
infectious disease consultation | 0
tricuspid valvulectomy decision | 0
blood and valve cultures confirmed methicillin-susceptible S aureus | 0
refractory hypoxemia | 2
partial pressure of oxygen 60 mm Hg | 2
mechanical ventilation | 2
chest radiography showed no evidence of hemopneumothorax | 2
chest radiography showed no evidence of pulmonary edema | 2
chest radiography showed no evidence of lung consolidation | 2
aggressive diuresis | 2
inhaled epoprostenol initiated | 2
neuromuscular blockade initiated | 2
prone position | 2
VV ECMO cannulation | 4
ECMO support initiated | 4
adequate oxygenation | 4
ECMO specialty transport team sent | 4
patient transferred | 6
VV ECMO support continued | 6
transthoracic echocardiography performed | 12
TEE performed | 12
ventricularization of the right heart | 12
wide-open systolic regurgitant flow | 12
right ventricle dilated | 12
interatrial septum bowing | 12
VV ECMO cannulas correctly positioned | 12
return cannula positioned at the junction of the right atrium and superior vena cava | 12
outflow jet directed into the right atrium | 12
drainage cannula positioned at the junction of the right atrium and inferior vena cava | 12
reversal of hepatic vein flow | 12
severe tricuspid regurgitation | 12
patent foramen ovale (PFO) found | 12
significant right-to-left flow | 12
PFO closure decision | 24
TV replacement decision | 24
patient taken to the operating room | 24
PFO closure performed | 24
TV replacement performed | 24
31-mm St. Jude Epic porcine bioprosthetic valve used | 24
intraoperative TEE performed | 24
no residual tricuspid regurgitation | 24
no residual right-to-left shunt | 24
patient deccannulated from ECMO | 24
patient extubated | 24
IV antibiotic therapy initiated | 24
addiction specialist treatment initiated | 24
patient remained in the hospital for 19 days | 24
patient left the hospital against medical advice | 432
lost to follow-up | 432