18 years old| 0
male | 0
admitted to the hospital | 0
fever | -72
rash | -72
acne |  -672
minocycline |  -672
increased WBC count | 0
eosinophilia| 0
systemic involvement| 0
diffuse erythematous or maculopapular eruption| 0
pruritis |* 0
DRESS syndrome | 0
fever persisted | 0
rash persisted | 0
discharged | 24
Separate conjunctive phrases into its component events and assign them the same timestamp (for example, the separation of 'fever and rash' into 2 events: 'fever' and 'rash')  If the event has duration, assign the event time as the start of the time interval. Attempt to use the text span without modifications except 'history of' where applicable. Include all patient events, even if they appear in the discussion; do not omit any events; include termination/discontinuation events; include the pertinent negative findings, like 'no shortness of breath' and 'denies chest pain'.  Show the events and timestamps in rows, each row has two columns: one column for the event, the other column for the timestamp.  The time is a numeric value in hour unit. The two columns are separated by a pipe '|' as a bar-separated file. Skip the title of the table. Reply with the table only. Create a table from the following case:
<|eot_id|><|start_header_id|>user<|end_header_id|>
<|eot_id|><|start_header_id|>assistant<|end_header_id|>
65 years old | 0
hypertension | 0
COPD | 0
Parkinson's disease | 0
irregular treatment | 0
irregular follow-up | 0
progressive worsening of respiratory distress | -168
productive cough | -168
hypercapnic respiratory failure | 0
altered sensorium | 0
leukocytosis | 0
infective exacerbation of COPD | 0
intubated | 0
invasive mechanical ventilation | 0
ventilator-associated pneumonia | 216
Acinetobacter baumanii | 216
cefoperazone/sulbactam | 216
colistin | 216
significant fall in procalcitonin levels | 216
spontaneous breath trial failed | 216
worsening respiratory acidosis | 216
desaturation | 216
hypotension | 216
hypovolemic hypotension | 216
fluid responsive | 216
persistent polyuria | 216
hypokalemia | 216
hyponatremia | 216
hypocalcemia | 216
hypomagnesaemia | 216
excess renal loss of electrolytes | 216
high fractional excretion of sodium | 216
high transtubular potassium gradient | 216
concomitant polyuria | 216
parenteral correction of electrolytes | 216
recurrence of electrolyte abnormalities | 216
difficult weaning | 216
stopping colistin | 216
parameters started to reverse | 360
extubated | 384
grade III bed sores | 384
infected bed sores | 384
Klebsiella spp. | 384
restarted colistin | 648
electrolyte abnormalities recurred | 648
polyuria recurred | 648
hypovolemic hypotension recurred | 648
supraventricular tachycardia | 648
adenosine reversion | 648
low serum magnesium | 648
magnesium replacement | 648
no recurrence of SVT | 648
10 day colistin course | 648
repeated electrolyte corrections | 648
volume replacements | 648
discharged | 1008
resolution of abnormalities | 1008
Bartter syndrome diagnosis | 0
metabolic alkalosis | 0
hypokalemia | 0
normal blood pressure | 0
surreptitious vomiting excluded | 0
diuretic use excluded | 0
hyperaldosteronism excluded | 0
hypovolemic hypotension | 0
polyuria | 0
Bartter-like syndrome | 0
difficult weaning | 0
colistin use | 0
<|begin_of_text|><|start_header_id|>system<|end_header_id|>
pruritis | 0
hypotension |
