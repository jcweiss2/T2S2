14 years old | 0
female | 0
admitted to the hospital | 0
upper left teeth pain | -168
bulging of the maxillary region | -168
odontological assistance | -168
prescribed cephalexin | -168
cephalexin treatment | -168
behavioral alterations | -24
auditory hallucination | -24
sleep disturbances | -24
aggression | -24
frontal headache | -24
headache | -336
vomiting | 0
alternating periods of agitation | 0
aggressiveness | 0
somnolence | 0
mental confusion | 0
paranasal sinuses and brain computed tomography (CT) scan | 0
right maxillary and frontal sinuses opacification | 0
frontal sinus osseous erosion | 0
subdural empyema | 0
cerebral edema | 0
inflammatory alterations | 0
admission day laboratory work-up | 0
Hemoglobin | 0
Monocytes | 0
Hematocrit | 0
Platelets | 0
Leukocytes | 0
Urea | 0
Bands | 0
Creatinin | 0
CRP | 0
Lymphocyte | 0
Blood Culture | 0
referred to the pediatric intensive care unit | 0
empirically started on ceftriaxone | 0
levofloxacin | 0
vancomycin | 0
acyclovir | 0
meningoencephalitis | 0
cardiopulmonary arrest | 0
resuscitation maneuvers | 0
Glasgow Coma Scale (GCS) | 0
new CT scan | 0
diffuse cerebral edema | 0
brain herniation | 0
left internal jugular vein thrombosis | 0
died | 48
cerebrospinal fluid (CSF) analysis | 48
Appearance | 48
Protein | 48
WBC count | 48
Glucose | 48
Erythrocytes | 48
Lactate | 48
Neutrophils | 48
Lymphocytes | 48
Monocytes | 48
CSF culture | 48
autopsy | 48
craniotomy | 48
meningeal purulent exudate | 48
frontal bone erosion | 48
acute inflammation | 48
neutrophils | 48
acute osteomyelitis | 48
neuronal and glial necrosis | 48
diffuse encephalic ischemia | 48
left internal jugular vein thrombosis | 48
thrombophlebitis | 48
pneumonia | 48
alveolar edema | 48
liver | 48
spleen | 48
heart | 48
lymph nodes | 48
bone marrow | 48
sepsis | 48
acute tubular necrosis | 48
subdural empyema | 0
Lemierre syndrome | 0 
Fusobacterium necrophorum | 0 
septic embolization | 0 
odontogenic sinusitis | 0 
pulpitis | 0 
dental involvement | 0 
neurosurgical source of infection | 0 
contiguity | 0 
neurological sequelae | 0 
motor deficits | 0 
dysphagia | 0 
seizures | 0 
biphasic headache | 0 
orbital cellulitis | 0 
broad-spectrum antibiotics | 0 
surgery | 0 
craniotomy with drainage | 0 
third generation cephalosporin | 0 
vancomycin | 0 
metronidazole | 0 
CT scan | 0 
intracranial complications | 0 
ABS | 0 
acute rhinosinusitis | 0 
sinusitis | 0 
URI | 0 
upper respiratory infections | 0 
viral infections | 0 
bacterial infections | 0 
acute otitis media | 0 
ABS complications | 0 
local tissue | 0 
orbit | 0 
intracranial involvement | 0 
prognosis | 0 
neurological sequelae | 0 
mortality | 0 
developed countries | 0 
undeveloped countries | 0 
case series | 0 
Streptococcus spp | 0 
Streptococcus milleri | 0 
Fusobacterium necrophorum | 0 
Staphylococcus ssp | 0 
anaerobes | 0 
polymicrobial cultures | 0 
culture-negative secretions | 0 
toothache | -168 
odontogenic infection | -168 
maxillary sinusitis | -168 
frontal sinusitis | -168 
neurological signs | 0 
altered mental status | 0 
seizures | 0 
focal deficits | 0 
vomiting | 0 
swelling of the forehead | 0 
fever | 0 
rhinorrhea | 0 
nasal obstructions | 0 
URI symptoms | 0 
headache | -336 
fever | -24 
altered sensorium | -24 
Glasgow Coma Scale | 0 
CT scan | 0 
imaging exam | 0 
laboratory work-up | 0 
C-reactive protein | 0 
neutrophilia | 0 
shift to the left | 0 
Streptococcus spp | 0 
Fusobacterium necrophorum | 0 
Staphylococcus ssp | 0 
anaerobes | 0 
polymicrobial cultures | 0 
culture-negative secretions | 0 
intracranial complications | 0 
ABS | 0 
subdural empyema | 0 
extradural empyema | 0 
brain abscess | 0 
meningitis | 0 
cavernous sinus thrombophlebitis | 0 
sphenoid osteomyelitis | 0 
teenagers | 0 
males | 0 
headache | -336 
neurological signs | 0 
altered mental status | 0 
seizures | 0 
focal deficits | 0 
vomiting | 0 
swelling of the forehead | 0 
fever | 0 
rhinorrhea | 0 
nasal obstructions | 0 
URI symptoms | 0 
Glasgow Coma Scale | 0 
CT scan | 0 
laboratory work-up | 0 
C-reactive protein | 0 
neutrophilia | 0 
shift to the left | 0 
Streptococcus spp | 0 
Fusobacterium necrophorum | 0 
Staphylococcus ssp | 0 
anaerobes | 0 
polymicrobial cultures | 0 
culture-negative secretions | 0 
Lemierre syndrome | 0 
thrombophlebitis | 0 
septic embolization | 0 
lung | 0 
Fusobacterium necrophorum | 0 
neurological involvement | 0 
septic embolization | 0 
jugular thrombophlebitis | 0 
atypical Lemierre syndrome | 0 
bone perforation | 0 
contiguity | 0 
mastoid involvement | 0 
septic embolization | 0 
diffuse pneumonia | 0 
septic embolization | 0 
jugular-vein-infected thrombosis | 0 
Lemierre syndrome | 0 
Fusobacterium necrophorum | 0 
special culture media | 0 
laboratory techniques | 0 
negative results | 0 
intracranial complications | 0 
ABS | 0 
dangerous consequences | 0 
neurological sequelae | 0 
death | 0 
altered neurological findings | 0 
biphasic headache | 0 
failure of a former treatment | 0 
orbital cellulitis | 0 
CT scan | 0 
advanced stage of the disease | 0 
hospital | 0 
treatment | 0 
broad-spectrum antibiotics | 0 
surgery | 0 
craniotomy with drainage | 0 
third generation cephalosporin | 0 
vancomycin | 0 
metronidazole | 0 
CT scan | 0 
intracranial complications | 0 
ABS | 0 
acute rhinosinusitis | 0 
sinusitis | 0 
URI | 0 
upper respiratory infections | 0 
viral infections | 0 
bacterial infections | 0 
acute otitis media | 0 
ABS complications | 0 
local tissue | 0 
orbit | 0 
intracranial involvement | 0 
prognosis | 0 
neurological sequelae | 0 
mortality | 0 
developed countries | 0 
undeveloped countries | 0 
case series | 0 
Streptococcus spp | 0 
Streptococcus milleri | 0 
Fusobacterium necrophorum | 0 
Staphylococcus ssp | 0 
anaerobes | 0 
polymicrobial cultures | 0 
culture-negative secretions | 0 
subdural empyema | 0 
Lemierre syndrome | 0 
Fusobacterium necrophorum | 0 
septic embolization | 0 
lung | 0 
Fusobacterium necrophorum | 0 
neurological involvement | 0 
septic embolization | 0 
jugular thrombophlebitis | 0 
atypical Lemierre syndrome | 0 
bone perforation | 0 
contiguity | 0 
mastoid involvement | 0 
septic embolization | 0 
diffuse pneumonia | 0 
septic embolization | 0 
jugular-vein-infected thrombosis | 0 
Lemierre syndrome | 0 
Fusobacterium necrophorum | 0 
special culture media | 0 
laboratory techniques | 0 
negative results | 0 
intracranial complications | 0 
ABS | 0 
dangerous consequences | 0 
neurological sequelae | 0 
death | 0 
altered neurological findings | 0 
biphasic headache | 0 
failure of a former treatment | 0 
orbital cellulitis | 0 
CT scan | 0 
advanced stage of the disease | 0 
hospital | 0 
treatment | 0 
broad-spectrum antibiotics | 0 
surgery | 0 
craniotomy with drainage | 0 
third generation cephalosporin | 0 
vancomycin | 0 
metronidazole | 0 
CT scan | 0 
intracranial complications | 0 
ABS | 0 
acute rhinosinusitis | 0 
sinusitis | 0 
URI | 0 
upper respiratory infections | 0 
viral infections | 0 
bacterial infections | 0 
acute otitis media | 0 
ABS complications | 0 
local tissue | 0 
orbit | 0 
intracranial involvement | 0 
prognosis | 0 
neurological sequelae | 0 
mortality | 0 
developed countries | 0 
undeveloped countries | 0 
case series | 0 
Streptococcus spp | 0 
Streptococcus milleri | 0 
Fusobacterium necrophorum | 0 
Staphylococcus ssp | 0 
anaerobes | 0 
polymicrobial cultures | 0 
culture-negative secretions | 0 
subdural empyema | 0 
Lemierre syndrome | 0 
Fusobacterium necrophorum | 0 
septic embolization | 0 
lung | 0 
Fusobacterium necrophorum | 0 
neurological involvement | 0 
septic embolization | 0 
jugular thrombophlebitis | 0 
atypical Lemierre syndrome | 0 
bone perforation | 0 
contiguity | 0 
mastoid involvement | 0 
septic embolization | 0 
diffuse pneumonia | 0 
septic embolization | 0 
jugular-vein-infected thrombosis | 0 
Lemierre syndrome | 0 
Fusobacterium necrophorum | 0 
special culture media | 0 
laboratory techniques | 0 
negative results | 0 
intracranial complications | 0 
ABS | 0 
dangerous consequences | 0 
neurological sequelae | 0 
death | 0 
altered neurological findings | 0 
biphasic headache | 0 
failure of a former treatment | 0 
orbital cellulitis | 0 
CT scan | 0 
advanced stage of the disease | 0 
hospital | 0 
treatment | 0 
broad-spectrum antibiotics | 0 
surgery | 0 
craniotomy with drainage | 0 
third generation cephalosporin | 0 
vancomycin | 0 
metronidazole | 0 
CT scan | 0 
intracranial complications | 0 
ABS | 0 
acute rhinosinusitis | 0 
sinusitis | 0 
URI | 0 
upper respiratory infections | 0 
viral infections | 0 
bacterial infections | 0 
acute otitis media | 0 
ABS complications | 0 
local tissue | 0 
orbit | 0 
intracranial involvement | 0 
prognosis | 0 
neurological sequelae | 0 
mortality | 0 
developed countries | 0 
undeveloped countries | 0 
case series | 0 
Streptococcus spp | 0 
Streptococcus milleri | 0 
Fusobacterium necrophorum | 0 
Staphylococcus ssp | 0 
anaerobes | 0 
polymicrobial cultures | 0 
culture-negative secretions | 0 
subdural empyema | 0 
Lemierre syndrome | 0 
Fusobacterium necrophorum | 0 
septic embolization | 0 
lung | 0 
Fusobacterium necrophorum | 0 
neurological involvement | 0 
septic embolization | 0 
jugular thrombophlebitis | 0 
atypical Lemierre syndrome | 0 
bone perforation | 0 
contiguity | 0 
mastoid involvement | 0 
septic embolization | 0 
diffuse pneumonia | 0 
septic embolization | 0 
jugular-vein-infected thrombosis | 0 
Lemierre syndrome | 0 
Fusobacterium necrophorum | 0 
special culture media | 0 
laboratory techniques | 0 
negative results | 0 
intracranial complications | 0 
ABS | 0 
dangerous consequences | 0 
neurological sequelae | 0 
death | 0 
altered neurological findings | 0 
biphasic headache | 0 
failure of a former treatment | 0 
orbital cellulitis | 0 
CT scan | 0 
advanced stage of the disease | 0 
hospital | 0 
treatment | 0 
broad-spectrum antibiotics | 0 
surgery | 0 
craniotomy with drainage | 0 
third generation cephalosporin | 0 
vancomycin | 0 
metronidazole | 0 
CT scan | 0 
intracranial complications | 0 
ABS | 0 
acute rhinosinusitis | 0 
sinusitis | 0 
URI | 0 
upper respiratory infections | 0 
viral infections | 0 
bacterial infections | 0 
acute otitis media | 0 
ABS complications | 0 
local tissue | 0 
orbit | 0 
intracranial involvement | 0 
prognosis | 0 
neurological sequelae | 0 
mortality | 0 
developed countries | 0 
undeveloped countries | 0 
case series | 0 
Streptococcus spp | 0 
Streptococcus milleri | 0 
Fusobacterium necrophorum | 0 
Staphylococcus ssp | 0 
anaerobes | 0 
polymicrobial cultures | 0 
culture-negative secretions | 0 
subdural empyema | 0 
Lemierre syndrome | 0 
Fusobacterium necrophorum | 0 
septic embolization | 0 
lung | 0 
Fusobacterium necrophorum | 0 
neurological involvement | 0 
septic embolization | 0 
jugular thrombophlebitis | 0 
atypical Lemierre syndrome | 0 
bone perforation | 0 
contiguity | 0 
mastoid involvement | 0 
septic embolization | 0 
diffuse pneumonia | 0 
septic embolization | 0 
jugular-vein-infected thrombosis | 0 
Lemierre syndrome | 0 
Fusobacterium necrophorum | 0 
special culture media | 0 
laboratory techniques | 0 
negative results | 0 
intracranial complications | 0 
ABS | 0 
dangerous consequences | 0 
neurological sequelae | 0 
death | 0 
altered neurological findings | 0 
biphasic headache | 0 
failure of a former treatment | 0 
orbital cellulitis | 0 
CT scan | 0 
advanced stage of the disease | 0 
hospital | 0 
treatment | 0 
broad-spectrum antibiotics | 0 
surgery | 0 
craniotomy with drainage | 0 
third generation cephalosporin | 0 
vancomycin | 0 
metronidazole | 0 
CT scan | 0 
intracranial complications | 0 
ABS | 0 
acute rhinosinusitis | 0 
sinusitis | 0 
URI | 0 
upper respiratory infections | 0 
viral infections | 0 
bacterial infections | 0 
acute otitis media | 0 
ABS complications | 0 
local tissue | 0 
orbit | 0 
intracranial involvement | 0 
prognosis | 0 
neurological sequelae | 0 
mortality | 0 
developed countries | 0 
undeveloped countries | 0 
case series | 0 
Streptococcus spp | 0 
Streptococcus milleri | 0 
Fusobacterium necrophorum | 0 
Staphylococcus ssp | 0 
anaerobes | 0 
polymicrobial cultures | 0 
culture-negative secretions | 0 
subdural empyema | 0 
Lemierre syndrome | 0 
Fusobacterium necrophorum | 0 
septic embolization | 0 
lung | 0 
Fusobacterium necrophorum | 0 
neurological involvement | 0 
septic embolization | 0 
jugular thrombophlebitis | 0 
atypical Lemierre syndrome | 0 
bone perforation | 0 
contiguity | 0 
mastoid involvement | 0 
septic embolization | 0 
diffuse pneumonia | 0 
septic embolization | 0 
jugular-vein-infected thrombosis | 0 
Lemierre syndrome | 0 
Fusobacterium necrophorum | 0 
special culture media | 0 
laboratory techniques | 0 
negative results | 0 
intracranial complications | 0 
ABS | 0 
dangerous consequences | 0 
neurological sequelae | 0 
death | 0 
altered neurological findings | 0 
biphasic headache | 0 
failure of a former treatment | 0 
orbital cellulitis | 0 
CT scan | 0 
advanced stage of the disease | 0 
hospital | 0 
treatment | 0 
broad-spectrum antibiotics | 0 
surgery | 0 
craniotomy with drainage | 0 
third generation cephalosporin | 0 
vancomycin | 0 
metronidazole | 0 
CT scan | 0 
intracranial complications | 0 
ABS | 0 
acute rhinosinusitis | 0 
sinusitis | 0 
URI | 0 
upper respiratory infections | 0 
viral infections | 0 
bacterial infections | 0 
acute otitis media | 0 
ABS complications | 0 
local tissue | 0 
orbit | 0 
intracranial involvement | 0 
prognosis | 0 
neurological sequelae | 0 
mortality | 0 
developed countries | 0 
undeveloped countries | 0 
case series | 0 
Streptococcus spp | 0 
Streptococcus milleri | 0 
Fusobacterium necrophorum | 0 
Staphylococcus ssp | 0 
anaerobes | 0 
polymicrobial cultures | 0 
culture-negative secretions | 0 
subdural empyema | 0 
Lemierre syndrome | 0 
Fusobacterium necrophorum | 0 
septic embolization | 0 
lung | 0 
Fusobacterium necrophorum | 0 
neurological involvement | 0 
septic embolization | 0 
jugular thrombophlebitis | 0 
atypical Lemierre syndrome | 0 
bone perforation | 0 
contiguity | 0 
mastoid involvement | 0 
septic embolization | 0 
diffuse pneumonia | 0 
septic embolization | 0 
jugular-vein-infected thrombosis | 0 
Lemierre syndrome | 0 
Fusobacterium necrophorum | 0 
special culture media | 0 
laboratory techniques | 0 
negative results | 0 
intracranial complications | 0 
ABS | 0 
dangerous consequences | 0 
neurological sequelae | 0 
death | 0 
altered neurological findings | 0 
biphasic headache | 0 
failure of a former treatment | 0 
orbital cellulitis | 0 
CT scan | 0 
advanced stage of the disease | 0 
hospital | 0 
treatment | 0 
broad-spectrum antibiotics | 0 
surgery | 0 
craniotomy with drainage | 0 
third generation cephalosporin | 0 
vancomycin | 0 
metronidazole | 0 
CT scan | 0 
intracranial complications | 0 
ABS | 0 
acute rhinosinusitis | 0 
sinusitis | 0 
URI | 0 
upper respiratory infections | 0 
viral infections | 0 
bacterial infections | 0 
acute otitis media | 0 
ABS complications | 0 
local tissue | 0 
orbit | 0 
intracranial involvement | 0 
prognosis | 0 
neurological sequelae | 0 
mortality | 0 
developed countries | 0 
undeveloped countries | 0 
case series | 0 
Streptococcus spp | 0 
Streptococcus milleri | 0 
Fusobacterium necrophorum | 0 
Staphylococcus ssp | 0 
anaerobes | 0 
polymicrobial cultures | 0 
culture-negative secretions | 0 
subdural empyema | 0 
Lemierre syndrome | 0 
Fusobacterium necrophorum | 0 
septic embolization | 0 
lung | 0 
Fusobacterium necrophorum | 0 
neurological involvement | 0 
septic embolization | 0 
jugular thrombophlebitis | 0 
atypical Lemierre syndrome | 0 
bone perforation | 0 
contiguity | 0 
mastoid involvement | 0 
septic embolization | 0 
diffuse pneumonia | 0 
septic embolization | 0 
jugular-vein-infected thrombosis | 0 
Lemierre syndrome | 0 
Fusobacterium necrophorum | 0 
special culture media | 0 
laboratory techniques | 0 
negative results | 0 
intracranial complications | 0 
ABS | 0 
dangerous consequences | 0 
neurological sequelae | 0 
death | 0 
altered neurological findings | 0 
biphasic headache | 0 
failure of a former treatment | 0 
orbital cellulitis | 0 
CT scan | 0 
advanced stage of the disease | 0 
hospital | 0 
treatment | 0 
broad-spectrum antibiotics | 0 
surgery | 0 
craniotomy with drainage | 0 
third generation cephalosporin | 0 
vancomycin | 0 
metronidazole | 0 
CT scan | 0 
intracranial complications | 0 
ABS | 0 
acute rhinosinusitis | 0 
sinusitis | 0 
URI | 0 
upper respiratory infections | 0 
viral infections | 0 
bacterial infections | 0 
acute otitis media | 0 
ABS complications | 0 
local tissue | 0 
orbit | 0 
intracranial involvement | 0 
prognosis | 0 
neurological sequelae | 0 
mortality | 0 
developed countries | 0 
undeveloped countries | 0 
case series | 0 
Streptococcus spp | 0 
Streptococcus milleri | 0 
Fusobacterium necrophorum | 0 
Staphylococcus ssp | 0 
anaerobes | 0 
polymicrobial cultures | 0 
culture-negative secretions | 0 
subdural empyema | 0 
Lemierre syndrome | 0 
Fusobacterium necrophorum | 0 
septic embolization | 0 
lung | 0 
Fusobacterium necrophorum | 0 
neurological involvement | 0 
septic embolization | 0 
jugular thrombophlebitis | 0 
atypical Lemierre syndrome | 0 
bone perforation | 0 
contiguity | 0 
mastoid involvement | 0 
septic embolization | 0 
diffuse pneumonia | 0 
septic embolization | 0 
jugular-vein-infected thrombosis | 0 
Lemierre syndrome | 0 
Fusobacterium necrophorum | 0 
special culture media | 0 
laboratory techniques | 0 
negative results | 0 
intracranial complications | 0 
ABS | 0 
dangerous consequences | 0 
neurological sequelae | 0 
death | 0 
altered neurological findings | 0 
biphasic headache | 0 
failure of a former treatment | 0 
orbital cellulitis | 0 
CT scan | 0 
advanced stage of the disease | 0 
hospital | 0 
treatment | 0 
broad-spectrum antibiotics | 0 
surgery | 0 
craniotomy with drainage | 0 
third generation cephalosporin | 0 
vancomycin | 0 
metronidazole | 0 
CT scan | 0 
intracranial complications | 0 
ABS | 0 
acute rhinosinusitis | 0 
sinusitis | 0 
URI | 0 
upper respiratory infections | 0 
viral infections | 0 
bacterial infections | 0 
acute otitis media | 0 
ABS complications | 0 
local tissue | 0 
orbit | 0 
intracranial involvement | 0 
prognosis | 0 
neurological sequelae | 0 
mortality | 0 
developed countries | 0 
undeveloped countries | 0 
case series | 0 
Streptococcus spp | 0 
Streptococcus milleri | 0 
Fusobacterium necrophorum | 0 
Staphylococcus ssp | 0 
anaerobes | 0 
polymicrobial cultures | 0 
culture-negative secretions | 0 
subdural empyema | 0 
Lemierre syndrome | 0 
Fusobacterium necrophorum | 0 
septic embolization | 0 
lung | 0 
Fusobacterium necrophorum | 0 
neurological involvement | 0 
septic embolization | 0 
jugular thrombophlebitis | 0 
atypical Lemierre syndrome | 0 
bone perforation | 0 
contiguity | 0 
mastoid involvement | 0 
septic embolization | 0 
diffuse pneumonia | 0 
septic embolization | 0 
jugular-vein-infected thrombosis | 0 
Lemierre syndrome | 0 
Fusobacterium necrophorum | 0 
special culture media | 0 
laboratory techniques | 0 
negative results | 0 
intracranial complications | 0 
ABS | 0 
dangerous consequences | 0 
neurological sequelae | 0 
death | 0 
altered neurological findings | 0 
biphasic headache | 0 
failure of a former treatment | 0 
orbital cellulitis | 0 
CT scan | 0 
advanced stage of the disease | 0 
hospital | 0 
treatment | 0 
broad-spectrum antibiotics | 0 
surgery | 0 
craniotomy with drainage | 0 
third generation cephalosporin | 0 
vancomycin | 0 
metronidazole | 0 
CT scan | 0 
intracranial complications | 0 
ABS | 0 
acute rhinosinusitis | 0 
sinusitis | 0 
URI | 0 
upper respiratory infections | 0 
viral infections | 0 
bacterial infections | 0 
acute otitis media | 0 
ABS complications | 0 
local tissue | 0 
orbit | 0 
intracranial involvement | 0 
prognosis | 0 
neurological sequelae | 0 
mortality | 0 
developed countries | 0 
undeveloped countries | 0 
case series | 0 
Streptococcus spp | 0 
Streptococcus milleri | 0 
Fusobacterium necrophorum | 0 
Staphylococcus ssp | 0 
anaerobes | 0 
polymicrobial cultures | 0 
culture-negative secretions | 0 
subdural empyema | 0 
Lemierre syndrome | 0 
Fusobacterium necrophorum | 0 
septic embolization | 0 
lung | 0 
Fusobacterium necrophorum | 0 
neurological involvement | 0 
septic embolization | 0 
jugular thrombophlebitis | 0 
atypical Lemierre syndrome | 0 
bone perforation | 0 
contiguity | 0 
mastoid involvement | 0 
septic embolization | 0 
diffuse pneumonia | 0 
septic embolization | 0 
jugular-vein-infected thrombosis | 0 
Lemierre syndrome | 0 
Fusobacterium necrophorum | 0 
special culture media | 0 
laboratory techniques | 0 
negative results | 0 
intracranial complications | 0 
ABS | 0 
dangerous consequences | 0 
neurological sequelae | 0 
death | 0 
altered neurological findings | 0 
biphasic headache | 0 
failure of a former treatment | 0 
orbital cellulitis | 0 
CT scan | 0 
advanced stage of the disease | 0 
hospital | 0 
treatment | 0 
broad-spectrum antibiotics | 0 
surgery | 0 
craniotomy with drainage | 0 
third generation cephalosporin | 0 
vancomycin | 0 
metronidazole | 0 
CT scan | 0 
intracranial complications | 0 
ABS | 0 
acute rhinosinusitis | 0 
sinusitis | 0 
URI | 0 
upper respiratory infections | 0 
viral infections | 0 
bacterial infections | 0 
acute otitis media | 0 
ABS complications | 0 
local tissue | 0 
orbit | 0 
intracranial involvement | 0 
prognosis | 0 
neurological sequelae | 0 
mortality | 0 
developed countries | 0 
undeveloped countries | 0 
case series | 0 
Streptococcus spp | 0 
Streptococcus milleri | 0 
Fusobacterium necrophorum | 0 
Staphylococcus ssp | 0 
anaerobes | 0 
polymicrobial cultures | 0 
culture-negative secretions | 0 
subdural empyema | 0 
Lemierre syndrome | 0 
Fusobacterium necrophorum | 0 
septic embolization | 0 
lung | 0 
Fusobacterium necrophorum | 0 
neurological involvement | 0 
septic embolization | 0 
jugular thrombophlebitis | 0 
atypical Lemierre syndrome | 0 
bone perforation | 0 
contiguity | 0 
mastoid involvement | 0 
septic embolization | 0 
diffuse pneumonia | 0 
septic embolization | 0 
jugular-vein-infected thrombosis | 0 
Lemierre syndrome | 0 
Fusobacterium necrophorum | 0 
special culture media | 0 
laboratory techniques | 0 
negative results | 0 
intracranial complications | 0 
ABS | 0 
dangerous consequences | 0 
neurological sequelae | 0 
death | 0 
altered neurological findings | 0 
biphasic headache | 0 
failure of a former treatment | 0 
orbital cellulitis | 0 
CT scan | 0 
advanced stage of the disease | 0 
hospital | 0 
treatment | 0 
broad-spectrum antibiotics | 0 
surgery | 0 
craniotomy with drainage | 0 
third generation cephalosporin | 0 
vancomycin | 0 
metronidazole | 0 
CT scan | 0 
intracranial complications | 0 
ABS | 0 
acute rhinosinusitis | 0 
sinusitis | 0 
URI | 0 
upper respiratory infections | 0 
viral infections | 0 
bacterial infections | 0 
acute otitis media | 0 
ABS complications | 0 
local tissue | 0 
orbit | 0 
intracranial involvement | 0 
prognosis | 0 
neurological sequelae | 0 
mortality | 0 
developed countries | 0 
undeveloped countries | 0 
case series | 0 
Streptococcus spp | 0 
Streptococcus milleri | 0 
Fusobacterium necrophorum | 0 
Staphylococcus ssp | 0 
