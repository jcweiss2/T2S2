40 years old | 0
male | 0
admitted to hospital | 0
hemiplegia of the right limb | -1
coma | -2
cerebral hemorrhage in the left basal ganglia region | 0
craniotomy | 0
hematoma removal | 0
decompression | 0
bone flap removal | 0
subdural effusion | 72
CSF leakage | 552
high body temperature | 552
lumbar puncture | 552
cloudy CSF | 552
elevated CSF protein | 552
elevated white blood cells in CSF | 552
decreased CSF glucose | 552
subcutaneous drainage | 560
drainage tube fixed | 560
subcutaneous effusion decreased | 576
body temperature normal | 576
subcutaneous drainage tube removed | 576
intracranial infection | 576
lumbar cistern catheter drainage | 600
CSF culture and drug sensitivity results | 600
carbapenem-resistant Klebsiella pneumoniae | 600
amikacin intravenous injection | 608
gentamicin intrathecal injection | 608
co-trimoxazole oral | 608
body temperature controlled | 624
CSF white blood cells decreased | 624
CSF glucose normal | 624
CSF protein normal | 624
lumbar cistern blocked | 648
tube removed | 648
head CT normal | 672
hydrocephalus | 720
infection controlled | 720
consciousness regained | 720
discharged to rehabilitation hospital | 720