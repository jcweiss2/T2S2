54 years old | 0
    man | 0
    admitted to a local hospital | 0
    discomfort in the hepatic region | 0
    cirrhosis | -8760
    hypersplenism | -8760
    portal hypertension | -8760
    multiple nodules at S4 and S5 in the liver | -24
    hepatocellular carcinoma | -24
    interventional surgery | -24
    multiple early stage lung tumors | -24
    referred to our hospital for surgery | -24
    significant decrease in platelets | -48
    significant decrease in fibrin | -48
    treated with thrombopoietin | -48
    treated with cryoprecipitate | -48
    white blood cell count 6.07×109/L | 0
    hemoglobin 124 g/L | 0
    platelet count 297×109/L | 0
    total bilirubin 29.3 µmol/L | 0
    direct bilirubin 11.8 µmol/L | 0
    total serum protein 59.5 g/L | 0
    albumin 32.7 g/L | 0
    prothrombin time 15.40 s | 0
    partial thromboplastin activation time 33.90 s | 0
    carcinoembryonic antigen 4.89 ng/mL | 0
    carbohydrate antigen 199 269.10 U/mL | 0
    carbohydrate antigen 724 7.19 U/mL | 0
    cytokeratin 19 fragment 6.30 ng/mL | 0
    hepatitis B virus DNA <5.00E+02 IU/mL | 0
    Child-Pugh classification grade B | 0
    Child-Pugh score of 8 points | 0
    hybrid ground glass density nodules in the posterior segment of the left upper lung | -24
    hybrid ground glass density nodules in the anterior segment of the right upper lobe | -24
    no evidence of lymph node metastases | -24
    no evidence of distant metastases | -24
    preoperative diagnosis lung cancer: clinical T1 N0 M0 stage IA | -24
    performed left superior segmentectomy | 0
    performed right superior wedge resection | 0
    rapid operative pathological diagnosis indicated adenocarcinomas on both sides | 0
    amount of bleeding 200 mL | 0
    length of operation 3 hours and 10 minutes | 0
    no blood transfusions | 0
    invasive adenocarcinoma on the left | 0
    well-differentiated adenocarcinoma on the right | 0
    negative margins | 0
    no evidence of metastasis in the lymph nodes | 0
    left thoracic duct effused 1,200 mL sanguineous drainage | 6
    increased heart rate | 6
    hypotension | 6
    plasma transfused | 6
    red blood cells transfused | 6
    platelets transfused | 6
    cryoprecipitate transfused | 6
    atrial fibrillation | 24
    dyspnea | 24
    acute respiratory distress syndrome | 24
    diffused alveolar hemorrhage | 24
    stale blood clots in the phlegm | 24
    violent coughing | 24
    white blood cell count 13.2×109/L | 48
    hemoglobin 66 g/L | 48
    platelet count 123×109/L | 48
    prothrombin time 15.80 s | 48
    partial thromboplastin activation time 35.40 s | 48
    fibrinogen 1.45 g/L | 48
    total bilirubin 33.7 µmol/L | 48
    direct bilirubin 15.3 µmol/L | 48
    total serum protein 50.1 g/L | 48
    albumin 33.3 g/L | 48
    postoperative CT scan patchy infiltrates scattered throughout both lungs | 96
    noninvasive ventilator-assisted ventilation | 96
    pulse oxygen saturation dropped to 85% | 96
    sanguineous drainage from the left thoracic duct | 96
    plasma transfused | 96
    red blood cells transfused | 96
    heart failure | 96
    pulmonary edema | 96
    standard heart failure treatments | 96
    low-dose steroids | 96
    left thoracic duct drainage gradually diminished | 168
    oxygenation improved | 168
    partial pressure of oxygen improved | 168
    sputum culture showed Klebsiella pneumoniae | 240
    sputum culture showed Candida albicans | 240
    meropenem employed | 240
    voriconazole employed | 240
    chest CT reexamination fewer patchy infiltrates | 312
    repeated sputum culture Candida albicans | 336
    voriconazole per os advised | 336
    discharged from the hospital | 384
    no evidence of recurrent disease at 3-month follow-up | 2160
    