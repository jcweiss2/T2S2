44 years old | 0
female | 0
admitted to the emergency department | 0
left groin and inner thigh redness | -72
left groin and inner thigh pain | -72
left groin and inner thigh swelling | -72
fever | -72
chills | -72
vomiting | -72
treated with intravenous vancomycin | -24
discharged from urgent care | -24
presented to the ED | 0
afebrile | 0
normotensive | 0
tachycardia | 0
mild tachypnea | 0
left inner thigh and groin induration | 0
morbidly obese | 0
lactate 3.5 mmol/L | 0
WBC 18.2 × 103 per mm3 | 0
hemoglobin 12.3 g/dL | 0
sodium 136 mmol/dL | 0
glucose 225 mg/dL | 0
creatinine 1.8 mg/dL | 0
LRINEC score of 6 | 0
bedside ultrasound performed | 0
subcutaneous thickening | 0
air | 0
fascial fluid | 0
started on intravenous vancomycin and piperacillin/tazobactam | 0
surgery consulted | 0
operative debridement | 0
excision of 15 cm × 23 cm of tissue | 0
extensive washout | 0
admitted to the surgical intensive care unit | 0
septic shock | 0
requiring vasopressors | 0
ventilator dependence | 0
repeat washouts with minor debridements | 24
lactate normalization | 72
down-trending WBC to 13.5 × 103 per mm3 | 72
extubated | 120
transferred to a step-down unit | 120
plastic surgery consulted | 120
evaluated for possible skin graft | 120
deemed to be a poor graft candidate | 216
wound vacuum-assisted closure (V.A.C.) device placed | 216
transferred to the plastic surgery service | 216
discharged home with a wound V.A.C. | 672
received a skin graft | 672