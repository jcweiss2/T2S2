43 years old | 0 | 0 
female | 0 | 0 
admitted to the hospital | 0 | 0 
difficult-to-manage bronchial asthma | -192 | 0 
hospitalized in the last 8 months on 10 occasions for acute exacerbations | -192 | 0 
asthmatic crisis | -192 | 0 
dry cough | -24 | 0 
progressive dyspnea | -24 | 0 
psychomotor agitation | -24 | 0 
audible wheezing | -24 | 0 
salbutamol | -24 | 0 
ipratropium bromide | -24 | 0 
diaphoretic | 0 | 0 
tachycardic | 0 | 0 
dyspneic | 0 | 0 
supraclavicular retractions | 0 | 0 
Glasgow coma scale 12/15 | 0 | 0 
arterial blood gases analysis | 0 | 0 
respiratory acidosis | 0 | 0 
hypoxemia | 0 | 0 
invasive ventilatory support | 0 | 0 
midazolam | 0 | 48 
propofol | 0 | 48 
hydrocortisone | 0 | 192 
magnesium sulfate | 0 | 192 
antibiotics | 0 | 192 
piperacillin tazobactam | 0 | 192 
clarithromycin | 0 | 192 
neuromuscular blocking agents | 48 | 96 
cisatracurium | 48 | 96 
improvement in ABG | 96 | 96 
ventilatory weaning | 96 | 96 
dual sedation suspended | 96 | 96 
NMB suspended | 96 | 96 
light sedation with dexmedetomidine | 96 | 240 
GCS 15/15 | 144 | 144 
weakness of the neck flexor muscles | 144 | 240 
facial paresis | 144 | 240 
quadriplegia | 144 | 240 
flaccid hyporeflexia | 144 | 240 
preserved sensitivity | 144 | 240 
brain MRI | 144 | 144 
cervical MRI | 144 | 144 
cerebrospinal fluid study | 144 | 144 
MRC score 37 points | 144 | 144 
electromyography | 144 | 144 
denervation | 144 | 240 
irritability | 144 | 240 
myopathic pattern | 144 | 240 
polyneuropathic compromise | 144 | 240 
axonal pattern | 144 | 240 
physiotherapy | 240 | 720 
comprehensive rehabilitation | 240 | 720 
ventilator withdrawn | 240 | 240 
MRC score 55 points | 720 | 720 
normal ABG control | 720 | 720 
symptomatic resolution | 720 | 720 
discharged | 720 | 720