63 years old | 0
male | 0
white | 0
peripheral vascular disease | -8760
claudication | -8760
hypertension | -8760
diabetes mellitus type-2 | -8760
chronic low back pain | -8760
dyspepsia | 0
melanic stools | -72
ibuprofen | -4320
sinus tachycardia | 0
hypotension | 0
left lower extremity weakness | 0
pallor | 0
pulselessness | 0
diffuse skin pallor | 0
severe anemia | 0
leukocytosis | 0
lactic acidosis | 0
acute renal failure | 0
hyponatremia | 0
hypokalemia | 0
positive occult blood | 0
positive blood cultures | 0
pantoprazole | 0
packed red blood cells | 0
crystalloid | 0
gastroenterology consultation | 0
vancomycin | 0
piperacillin/tazobactam | 0
CT angiogram | 0
EGD | 0
multiple bleeding duodenal ulcers | 0
cauterization | 0
epinephrine | 0
abdominal pain | 8
distension | 8
diaphoresis | 8
tachypnea | 8
fever | 8
hypertension | 8
tachycardia | 8
respiratory distress | 8
abdominal guarding | 8
rebound tenderness | 8
diffuse abdominal tenderness | 8
intubation | 8
general surgery consultation | 8
CT scan | 8
pneumo-peritoneum | 8
duodenal perforation | 8
norepinephrine | 9
vasopressin | 9
non-operative management | 9
strict bowel rest | 9
intravenous antibiotics | 9
intravenous fluconazole | 9
enteric antifungal coverage | 9
renal function deterioration | 120
oliguria | 120
acute tubular necrosis | 120
compartment syndrome | 120
extubation | 168
re-intubation | 180
hemodialysis | 192
left lower extremity necrosis | 360
palliative care | 360
death | 456