37 years old | 0
male | 0
quadriplegia | 0
chronic hypoxic respiratory failure | 0
mechanical ventilation | 0
tracheostomy | 0
admitted to the intensive care unit | 0
pneumonia | 0
serum creatinine level at presentation 1.39 mg/dl | 0
chest imaging suggestive of multifocal pneumonia | 0
acute respiratory distress syndrome | 0
septic shock | 0
vasopressor therapy | 0
worsening oxygen requirement | 0
SARS-CoV-2 negative | 0
serum creatinine level worsened to 3.3 mg/dl | 0
decline in urine output | 0
renal sonogram excluded obstructive uropathy | 0
fractional excretion of urea 25.6% | 0
prerenal etiology | 0
intravascular volume depletion | 0
diuretics treatment | 0
increased extravascular lung water | 0
i.v. fluid bolus administered | 0
nephrology consultation requested | 0
glomerulonephritis considered | 0
pulmonary-renal syndrome considered | 0
antinuclear antibody positive 1:160 | 0
bronchoscopy equivocal for alveolar hemorrhage | 0
fraction of inspired oxygen 70% | 0
positive end-expiratory pressure 12 cm H2O | 0
blood pressure 96/53 mm Hg | 0
pulse rate 92 bpm | 0
oxygen saturation 90% | 0
bilateral lung crackles | 0
trace pitting pedal edema | 0
urine output 350 ml/24h | 0
urine microscopy with muddy brown casts | 0
tubular injury | 0
no dysmorphic red blood cells | 0
hemodynamic injury | 0
serum sodium 146 mmol/l | 0
hyperkalemia 5.9 mmol/l | 0
serum bicarbonate 25 mmol/l | 0
dehydration | 0
overdiuresis | 0
administer fluids | 0
bedside ultrasound performed | 0
lung ultrasound bilateral diffuse B-line pattern | 0
irregular pleural line | 0
focused cardiac ultrasound hyperdynamic left ventricular systolic function | 0
enlarged right ventricle | 0
interventricular septal flattening | 0
D-shaped left ventricle | 0
volume overload | 0
pressure overload | 0
decreased cardiac output | 0
low blood pressure | 0
IVC plethoric | 0
IVC-estimated RAP unreliable | 0
hepatic vein Doppler S-wave reversal | 0
diastolic D pattern | 0
elevated RAP level | 0
portal vein Doppler pulsatile with flow reversal | 0
severe venous congestion | 0
severely elevated extravascular lung water | 0
right ventricular enlargement | 0
severe systemic venous congestion | 0
continuous renal replacement therapy initiated | 0
anti-double-stranded DNA negative | 24
antiglomerular basement membrane negative | 24
antineutrophil cytoplasmic antibodies negative | 24
renal biopsy not considered | 24
documented fluid balance negative 6.6 l | 72
hepatic vein Doppler S < D | 72
portal vein pulsatility improved | 72
blood pressure 115/57 mm Hg | 72
ultrafiltration continued | 72
fluid balance negative 5.1 l | 120
hepatic vein Doppler S < D | 120
portal vein waveform normalized | 120
urine output 150 ml/24h | 120
discontinued continuous renal replacement therapy | 120
plan for intermittent hemodialysis | 120
urine output 600 ml | 168
hemodialysis not required | 168
fluid balance negative 2 l | 192
hepatic vein Doppler S > D | 192
portal vein Doppler normal | 192
IVC dilated | 192
lung ultrasound improved | 192
increased lung water not resolved | 192
D-sign resolved | 192
left ventricle normal circular shape | 192
serum creatinine 2.1 mg/dl | 192
serum creatinine trended down to 0.6 mg/dl | 240
