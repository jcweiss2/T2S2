22 years old | 0
female | 0
admitted to the outpatient clinic | -240
fever | -240
sore throat | -240
treated as acute bacterial pharyngitis | -240
oral antibiotics | -240
no improvement | -240
persistent fever | -240
confusion | -240
dyspnea | -240
brought to the emergency room | 0
cyanosed | 0
basal crackles | 0
small anterior infrahyoid soft neck swelling | 0
emergently intubated | 0
admitted to ICU | 0
leukocytosis | 0
absolute neutrophilia | 0
mild increase in creatinine | 0
high blood sugar | 0
positive acetone in urine | 0
Chest x-ray | 0
computed tomography (CT) chest | 0
wide mediastinum | 0
moderate bilateral pleural effusion | 0
adjacent sub pleural atelectasis | 0
bilateral basal lung infiltrates | 0
mild pericardial effusion | 0
no signs of pulmonary embolism | 0
intercostal tubes inserted | 0
pleural fluid analysis | 0
exudate | 0
pH of 7.1 | 0
high white blood cell count | 0
predominantly neutrophils | 0
diagnosed as community acquired pneumonia | 0
secondary bilateral empyema | 0
diabetic ketoacidosis | 0
newly diagnosed diabetes mellitus | 0
septic shock | 0
acute kidney injury | 0
complicated by | 0
mechanical ventilation | 0
intravenous fluids | 0
insulin | 0
vasopressors | 0
broad spectrum antibiotics | 0
antifungals | 0
progressive edema | 24
increase in the size of the anterior soft neck swelling | 24
referred to King Khalid University Hospital (KKUH) | 336
clinical evaluation | 336
high fever | 336
hypotension | 336
tachycardia | 336
hypoxemia | 336
mechanical ventilation | 336
bilateral intercostal chest tubes | 336
generalized edema | 336
anterior infrahyoid soft neck swelling | 336
repeated CT chest and neck | 336
high density fluid collection | 336
prethyroid region | 336
extending down to the sternoclavicular joint | 336
multiple small mediastinal | 336
pretracheal | 336
paratracheal | 336
prevascular lymph nodes | 336
ultrasound guided aspiration | 336
frank pus | 336
thoracic surgery team consulted | 336
conservative management | 336
sputum culture | 336
Pseudomonas aeruginosa | 336
Acinetobacter baumannii | 336
antibiotics adjusted | 336
fever persisted | 336
hypotension persisted | 336
further deterioration in renal function | 336
renal replacement therapy | 336
neck and chest CT scan repeated | 336
multi loculated collection | 336
middle part of the neck | 336
extending down to the sternum | 336
larger and more defined | 336
large well defined loculated cystic lesion | 336
anterior mediastinum | 336
pericardial effusion increased | 336
bilateral pleural effusion increased | 336
basal atelectasis | 336
bilateral consolidation | 336
surgical intervention | 360
cervical dissection | 360
debridement | 360
drainage of pus | 360
left thoracotomy | 360
debridement | 360
drainage of mediastinal | 360
left pleural collection | 360
pleuropericardial window | 360
right thoracotomy | 384
debridement | 384
drainage of right pleural collection | 384
samples sent for bacterial | 384
fungal | 384
mycobacterial stains | 384
cultures | 384
no bacterial growth | 384
histopathology | 384
acute inflammatory process | 384
gradual improvement | 384
hemodynamics | 384
conscious level | 384
renal functions | 384
inflammatory markers | 384
weaning from mechanical ventilation | 384
difficult | 384
generalized weakness | 384
tracheostomy postponed | 384
infection and inflammation subsided | 384
anterior neck | 384
anterior mediastinum | 384
high fever | 480
tachycardia | 480
hypotension | 480
vasopressors | 480
repeat CT neck and chest | 480
interval reduction | 480
size of previously noted collections | 480
loculated pleural effusion | 480
interval development | 480
bilateral lateral loculated fluid collections | 480
beneath the thoracotomy sites | 480
CT guided aspiration | 480
ICU course complicated | 480
critical illness polyneuropathy | 480
myopathy | 480
tracheo-esophageal fistula | 480
conservatively managed | 480
tracheostomy | 480
feeding gastrostomy | 480
successful weaning | 744
mechanical ventilation | 744
transferred to general ward | 744
healing of tracheo-esophageal fistula | 840
oral feeding resumed | 840
tracheostomy tube removed | 840
gastrostomy tube removed | 840
discharged from hospital | 840