65 years old | 0
male | 0
hypertension | 0
admitted to the hospital | 0
subarachnoid hemorrhage | 0
external ventricular drain | 0
coiling | 0
septic shock | -192
C. difficile toxin positive | -192
leukocytosis | -192
creatinine level of 1.86 mg/dL | -192
vancomycin liquid 125 mg | -192
IV metronidazole 500 mg | -192
fidaxomicin 200 mg | -128
worsening sepsis | -128
no improvement in diarrhea | -128
abdominal pain | -96
distension | -96
acute hypoxemic respiratory failure | -96
mechanical ventilation | -96
diffuse severe bowel wall thickening | -96
toxic megacolon | -96
extensive pseudomembranes | -96
laparoscopic loop ileostomy | -96
colonic lavage | -96
vancomycin irrigation | -96
persistent diarrhea | 0
fever | 0
leukocytosis | 0
gastroenterology team consulted | 0
antibiotics held | 0
polyethylene glycol preparation | 0
FMT | 0
donor stool administered | 0
clinical condition improved | 72
resolution of leukocytosis | 72
resolution of diarrhea | 72
transferred to general medical floor | 120
discharged to rehabilitation facility | 240
repeat colonoscopy | 4320
resolution of CDI | 4320
reversal of ileostomy | 4320