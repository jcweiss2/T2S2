47 years old | 0
    woman | 0
    headache | -48
    blurred vision | -48
    referred to the department | 0
    CT scan of the skull | -48
    large mass arising from the sella | -48
    eroding the bony structures | -48
    invading the nasal cavity | -48
    admitted | 0
    Glasgow coma scale (GCS) 15 | 0
    afebrile | 0
    neurological examination showed no alterations | 0
    visual field intact | 0
    body mass index (BMI) 28.2 | 0
    medical history included mild psoriasis | 0
    gastroesophageal reflux disease (GERD) | 0
    cholelithiasis | 0
    no relevant infections except in her infancy | 0
    no previous surgeries | 0
    no routine medications | 0
    mother of two children | 0
    regular menses | 0
    blood pressure within normal limits | 0
    heart rate within normal limits | 0
    blood test showed microcromic microcytic anemia | 0
    reticulocytosis | 0
    hemoglobin (Hb) 8.6g/dL | 0
    hematocrit (HCT) 27.8% | 0
    mean cell volume (MCV) 64.5 | 0
    mean corpuscular hemoglobin (MCH) 20 pg | 0
    mean corpuscular hemoglobin concentration (MCHC) 30.9 g/dL | 0
    red blood cell distribution width (RDW) 20.2% | 0
    leucocytes count within normal limits | 0
    inflammatory indexes within normal limits | 0
    hormone blood concentrations normal except slight decrease in TSH | 0
    slight decrease in FSH | 0
    β-17-estradiol 35.8 pg/mL | 0
    urine osmolality normal | 0
    enhanced MRI | 0
    solid-cystic lesion arising from the sella turcica | 0
    abutting both cavernous sinuses | 0
    wrapping both carotid siphons | 0
    diagnosed with large pituitary adenoma with mixed solid/cystic consistence | 0
    scheduled for surgery the same week | 0
    headache treated with pain medications | 0
    no vision problems | 0
    headache suddenly worsened | 24
    rapidly developed gaze palsy | 24
    rapidly developed nuchal rigidity | 24
    GCS fell from 15 to 6 | 24
    emergency CT showed no parenchymal infarction | 24
    emergency CT showed no extra-axial bleeding | 24
    emergency CT showed no fluid collection | 24
    emergency CT showed no ischemia | 24
    urgent craniotomy performed | 24
    right frontotemporal approach | 24
    dura mater opened | 24
    brain swelling | 24
    dense pus covering the brain surface | 24
    purulent material found within the tumor located in the sella | 24
    drained purulent material | 24
    taken to the ICU | 24
    did not recover | 72
    died | 96
    pathological analysis confirmed nonfunctioning pituitary adenoma | 24
    chronic inflammation | 24
    necrosis | 24
    cultures of intraoperative material negative | 24
    