12 years old | 0
female | 0
cerebral palsy | 0
admitted to Intensive Care Unit | 0
decreased level of consciousness | 0
sepsis | 0
respiratory distress | 0
gastrointestinal bleeding | 0
hypoglycemia | 0
noninvasive ventilation | 0
wide spectrum antibiotics | 0
hypertonic glucose | 0
pancytopenia | 0
Klebsiella pneumoniae | 0
white worms escaped from right nose | 240
nasal myiasis | 240
L. sericata | 240
Ivermectin | 240
no other worm detected | 552
