32 years old | 0
male | 0
admitted to the hospital | 0
complaint of cough | -96
complaint of sputum | -96
complaint of dyspnea | -96
5-year history of classic pyoderma gangrenosum | -12000
received methylprednisolone pulses | -168
oral prednisolone | -672
cyclosporine | -672
surgical wound therapy | -672
respiratory rate of 30 breaths/min | 0
temperature of 39°C | 0
heart rate of 150 beats/min | 0
oxygen saturation below 90% | 0
large and deeply diffuse necrotic skin lesions | 0
skin lesions on the upper limbs | 0
skin lesions on the chest and back | 0
White blood cell count was 9.8 × 10^9/l | 0
differential of 79% neutrophils | 0
differential of 22% lymphocytes | 0
differential of 3% monocytes | 0
differential of 1% eosinophil | 0
Platelets were 25 × 10^9/L | 0
no vegetation in transthoracic echocardiogram | 0
computed tomography scan of the lungs | 0
multiple 1-2 cm nodules in various stages | 0
feeding vessels sign | 0
cavitations in some of them | 0
halo sign | 0
area of low attenuation surrounding a nodular lesion | 0
air-crescent signs | 0
small size left pleural effusion | 0
respiratory failure | 48
intubated and mechanically ventilated | 48
bronchoscopy | 48
bronchoalveolar lavage specimen | 48
diagnosis of probable invasive pulmonary aspergillosis | 48
direct microscopy examination of endobronchial washing | 48
direct microscopy examination of BAL samples | 48
acute branching septate hyphae | 48
aspergillosis | 48
culture of the samples revealed Aspergillus flavus | 48
diagnosis of cutaneous fusariosis | 48
Fusarium proliferatum isolated from skin lesion biopsy | 48
polymerase chain reaction assays | 48
fungal internal transcribed spacer region of rRNA gene | 48
voriconazole administration | 48
antimicrobial drugs administration | 48
linezolid administration | 48
meropenem administration | 48
ciprofloxacin administration | 48
treatment failed | 240
patient expired | 288