73 years old | 0
    man | 0
    presented with epigastric pain | 0
    nausea | 0
    hematemesis | -2
    smoker | 0
    pacemaker | 0
    arteriovenous (AV) block (II degree) | 0
    pale skin | 0
    blood pressure 155/70 mm Hg | 0
    heart rate 85 beats/min | 0
    capillary oxygen saturation of 92% | 0
    abdomen diffusively tender | 0
    abdomen distended | 0
    no clear rigidity | 0
    hemoglobin 90 mg/dL | 0
    white blood count 16×10^9/L | 0
    C-reactive protein 122 mg/L | 0
    abdominal radiography revealed soft tissue shadow | 0
    lamellar gas in gastric wall | 0
    CT showed thickened stomach wall | 0
    gas in intramural venous branches | 0
    gas in intrahepatic portal vein branches | 0
    gastroscopy showed no tumor | 0
    stomach necrosis in distal corpus | 0
    urgent surgery indicated | 0
    ischemic stomach body | 0
    necrotic areas along greater curvature | 0
    partial gastrectomy | 0
    Roux en esophago-jejunal anastomosis | 0
    postoperative course uneventful | 168
    discharged on 7th postoperative day | 168
    free of symptoms | 8760
    unremarkable gastroscopy findings | 8760
    ischemic transmural necrosis in greater curvature | 0
    edematous and inflamed smaller curvature | 0
    no sign of ulcer | 0
    no tumor | 0
    no mucosal laceration | 0
    polymicrobial infection (Klebsiella pneumoniae, Pseudomonas aeruginosa, Bacteroides fragilis) | 0
    emphysematous gastritis diagnosis | 0
    epigastric pain and nausea of 6 hours duration | -6
    hematemesis for the past 2 hours | -2