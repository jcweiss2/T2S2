70 years old | 0
male | 0
farmer | 0
presented to the emergency department | 0
high-grade fever | -120
generalized body ache | -120
headache | -120
altered sensorium | -120
joint pains | -120
epigastric pain | -120
inguinal lymphadenopathy | -120
mild generalized rash | -120
no eschar | -120
hemodynamically stable | -120
disoriented | -120
no focal neurological deficit | -120
no neck rigidity | -120
acute febrile illness with undifferentiated fever | -120
malaria | -120
dengue | -120
typhoid | -120
leptospira | -120
negative | -120
scrub typhus antigen card positive | 0
scrub immunoglobulin M (IgM) positive | 0
scrub typhus | 0
leukocytosis | 0
mild hyperbilirubinemia | 0
transaminitis | 0
sterile blood and other body fluid cultures | 0
doxycycline 100 mg twice daily | 0
defervescence | 2
improved orientation | 2
weakness of both lower limbs | 4
progressed to upper limbs | 4
bladder incontinence | 4
absent deep tendon reflexes | 4
flexor plantar responses | 4
intubated and put on mechanical ventilation | 4
MRI of the brain | 4
MRI of the cervical spine | 4
nerve conduction velocity (NCV) | 4
motor sensory demyelinating polyneuropathy | 4
cerebrospinal fluid (CSF) analysis | 4
albuminocytologic dissociation | 4
intravenous immunoglobulin therapy | 4
tablet rifampicin 600 mg twice daily | 4
improved weakness of all four limbs | 8
improved respiratory parameters | 8
weaned off and extubated from the ventilator | 8
oral feeding | 8
aggressive limb and chest physiotherapy | 8
shifted out from ICU | 8
discharged from the hospital | 28
full neurological recovery | 28