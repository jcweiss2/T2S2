39 years old | 0
male | 0
admitted to the Emergency Department | 0
hematemesis | 0
hemorrhagic shock | 0
arterial hypertension | -672
autoimmune thyroiditis | -672
type 2 diabetes mellitus | -672
diabetic neuropathy | -672
retinopathy | -672
nephropathy | -672
stage 3 chronic renal failure | -672
non-steroidal anti-inflammatory drugs | -168
neuropathic lower limbs pain | -168
resuscitation | 0
esophagogastroduodenoscopy | 0
huge clot in the stomach | 0
active bleeding | 0
cardiac arrest | 0
cardiopulmonary resuscitation | 0
hemodynamic stability | 0
proton pump inhibitors | 0
abdominal Doppler ultrasonography | 0
no sign of liver disease | 0
normal flow into the vena porta | 0
abdominal meteorism | 0
celio-mesenteric arteriography | 12
no arterial blush | 12
gastrointestinal hemorrhage | 24
transfused with packed red blood cells | 24
transfused with plasma | 24
abdominal contrast-enhanced computed tomography | 48
severe atrophy of the whole pancreas | 48
chronic pancreatitis | 48
thrombosis of the splenic vein | 48
splenomegaly | 48
cavernomatous transformation of the splenic hilum | 48
gastric fundus varices | 72
recent bleeding | 72
splenectomy | 96
splenic artery embolization | 24
laparoscopic splenectomy | 96
intraoperative hemorrhage | 96
splenic artery | 96
gastroepiploic vein | 96
short gastric vessels | 96
endoscopic vascular stapler | 96
minimal blood losses | 96
no intraoperative complications | 96
spleen extracted | 96
postoperative course | 96
discharged | 120
alive | 8760
no further episode of gastric bleeding | 8760