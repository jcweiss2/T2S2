45 years old | 0
male | 0
right-handed | 0
HIV | -672
CD4+ T-cell count of 556 | 0
admitted to the hospital | 0
horizontal diplopia | -24
weakness of left face | -24
weakness of right arm | -24
weakness of right leg | -24
hemiparesis alternans | -24
MRI | 0
FLAIR signal hyperintensity | 0
diffusion weighted imaging (DWI) restriction | 0
acute ischemic stroke | 0
Millard-Gubler syndrome | 0
extra-axial, curvilinear, high-signal abnormality | 0
subarachnoid space | 0
MRA | 0
cardiac telemetry | 0
sinus tachycardia | 0
transthoracic echocardiography | 0
transesophageal echocardiography | 0
normal ejection fraction | 0
normal valves | 0
normal chambers | 0
no clot | 0
no vegetation | 0
no patent foramen ovale | 0
no septal defect | 0
hypercoagulable serum panel | 0
anticardiolipin antibodies | 0
lupus anticoagulant | 0
protein C and S levels | 0
anti-thrombin III | 0
fibrinogen | 0
factor VIII | 0
prothrombin 20210 | 0
homocystine | 0
lipoprotein (a) | 0
sickle cell screen | 0
severe headache | 24
meningismus | 24
stupor | 24
lumbar puncture | 24
opening pressure of 230 mm H2O | 24
250 red blood cells | 24
75 white blood cells | 24
glucose of 80 | 24
protein of 54 | 24
opportunistic infections | 24
Cryptococcus | 24
tuberculosis | 24
syphilis | 24
acid-fast bacilli test | 24
PPD | 24
chest X-rays | 24
RPR | 24
VDRL | 24
FTA-ABS | 24
polymerase chain reaction (PCR) | 24
Herpes simplex virus 1 | 24
Herpes simplex virus 2 | 24
cytomegalovirus | 24
varicella-zoster virus (VZV) | 24
seeping, pustular furuncles | 24
MRSA | 24
blood cultures | 24
intravenous vancomycin | 24
second MRI | 48
extension of intra-axial FLAIR signal hyperintensities | 48
diffusion restriction | 48
bilateral pons | 48
left cerebellum | 48
new cerebral infarctions | 48
exacerbating cerebral infarctions | 48
subarachnoid space DWI restriction | 48
increasing in size | 48
expanding more curvilinearly | 48
left posterior fossa | 48
communicating hydrocephalus | 48
effacement of the fourth ventricle | 48
dilation of the lateral and third ventricles | 48
CSF trans-exudation | 48
another lumbar puncture | 48
4 red blood cells | 48
112 white blood cells | 48
glucose of 130 | 48
protein of 2,126 | 48
high-dose, broad-spectrum antibiotics | 48
vancomycin | 48
ceftriaxone | 48
ampicillin | 48
aggressive intravenous fluids | 48
pressor agents | 48
ventriculostomy | 48
supportive care measures | 48
comatose | 72
third MRI | 72
marked diffusion restriction | 72
hyperintense FLAIR signals | 72
brainstem parenchyma | 72
entire pons | 72
medulla | 72
left cerebellum | 72
repeat MRA | 72
irregularity and narrowing | 72
vertebro-basilar circulation | 72
lack of flow-related enhancement | 72
left vertebral artery | 72
posterior cerebral arteries | 72
expired | 96
autopsy | 96
brain weighed 1,212 g | 96
basilar artery | 96
posterior cerebral arteries | 96
cerebellar arteries | 96
mostly patent | 96
variable arteritis | 96
thick lymphoplasmocytic infiltration | 96
partial large-vessel occlusion | 96
subtotal small-vessel occlusion | 96
fibrointimal proliferation | 96
basilar meninges | 96
thickened | 96
white purulent material | 96
inferior brainstem | 96
left cerebellum | 96
recent non-hemorrhagic infarcts | 96
inflammation | 96
vasculitis | 96
cervical spinal cord leptomeninges | 96
moderate dilatation | 96
lateral and third ventricles | 96
aqueduct | 96
moderate compression | 96
fourth ventricle | 96
Gram and GMS stains | 96
copious Gram-Positive cocci | 96
chains | 96
macrophage infiltrates | 96
capillary proliferation | 96
post-mortem microscopy | 96