18 years old | 0
male | 0
type 1 diabetic | 0
hypertensive | 0
amlodipine | 0
inguinal hernia | -20
admitted to the emergency room | 0
abdominal pain | 0
ketoacidosis decompensation | 0
uremic syndrome | 0
conscious | 0
hemodynamically stable | 0
dyspneic | 0
febrile | 0
39.6°C | 0
right lumbar tenderness | 0
oliguric | 0
diuresis at 300 ml/24h | 0
altered renal function | 0
creatinine at 92 mg/l | 0
urea at 3.1 g/l | 0
K+ at 6.9 mmol/l | 0
Na+ at 123 mmol/l | 0
blood sugar at 6.5 g/l | 0
alkaline reserves at 8 mEq/l | 0
infectious syndrome | 0
CRP at 418 mg/l | 0
white blood cells at 26000/ml | 0
hemoglobin at 12.3 g/dl | 0
leucocyturia 320,000 | 0
hematuria at 120,000 | 0
emphysematous pyelonephritis | 0
renal abscess | 0
ruptured in the intraperitoneal cavity | 0
moderate abundance of pneumoperitoneum | 0
dialysis sessions | 0
insulin therapy | 0
antibiotic therapy | 0
ceftriaxone | 0
metronidazole | 0
surgical drainage of abscesses | 0
rise of a right double J stent | 0
evolution was favorable | 0
apyrexia | 2
chronic renal failure | 10
normal diuresis | 10
creatinine plateau of 20 mg/l | 10
oral antibiotics | 10
abdominopelvic CT | 10
clear regression of the bubbles of air | 34
double J catheter was removed | 42
abdominal pain persisted | -5.8
febrile low back pain | -5.8
septic shock | -5.8
Pseudomonas Aeruginosa | -5.8
Escherichia coli | -5.8
Klebsiella pneumonia | -5.8
Enterococcus | -5.8
Proteus mirabilis | -5.8
Type I EPN | -5.8
Type II EPN | -5.8
Class 1 EPN | -5.8
Class 2 EPN | -5.8
Class 3A EPN | -5.8
Class 3B EPN | -5.8
Class 4 EPN | -5.8
untreated EPN | -5.8
surgical treatment | -5.8
medical treatment | -5.8
uncontrolled diabetes | -5.8
upper excretory tract obstruction | -5.8