54 years old | 0
    male | 0
    admitted to the hospital | 0
    24-hour history of nausea | -24
    nausea | -24
    vomiting | -24
    diarrhea | -24
    abdominal pain | -24
    denied ingestion of fish | 0
    denied ingestion of contaminated food | 0
    denied ingestion of contaminated water | 0
    generalized skin flushing | 0
    blood pressure 60/39 mmHg | 0
    heart rate 131/min | 0
    temperature 37.8°C | 0
    aggressive fluid resuscitation initiated | 0
    intravenous ciprofloxacin initiated | 0
    intravenous metronidazole initiated | 0
    white blood count 18.9 × 10^9/L | 0
    neutrophils 17.63 × 10^9/L | 0
    hemoglobin 162 g/L |7 0
    platelets 120 × 10^9/L | 0
    creatinine 445 μmol/L | 0
    estimated GFR 12 mL/min | 0
    venous blood gas pH 7.29 | 0
    metabolic acidosis | 0
    non-injected CT scan showing thickened terminal ileum | 0
    non-injected CT scan showing distended appendix (13 mm) | 0
    non-injected CT scan showing mild stranding of surrounding fat | 0
    hemodynamic instability | 0
    suspected intra-abdominal source | 0
    surgical exploration | 0
    turbid fluid retrieved from RLQ sent for Gram stain and culture | 0
    1 cm necrotic zone at base of appendix | 0
    no significant signs of appendicular inflammation | 0
    no significant signs of ileal inflammation | 0
    appendectomy performed | 0
    peritoneal lavage performed | 0
    intraoperative short colonoscopy performed | 0
    colonoscopy normal | 0
    transesophageal echocardiography performed | 0
    echocardiography normal | 0
    admitted to ICU | 0
    vasopressors support for 2 days | 0
    developed disseminated intravascular coagulation (DIC) | 48
    empirical intravenous ciprofloxacin and metronidazole for 7 days | 168
    oral amoxicillin/clavulanic acid for 7 days | 168
    flushing syndrome persisted for 6 days | 144
    left ICU after 6 days | 144
    recovered uneventfully | 240
    discharged on postoperative Day 10 | 240
    blood analysis with MALDI-TOF MS | 0
    RLQ fluid analysis with MALDI-TOF MS | 0
    presence of R. ornithinolytica | 0
    multisensitive to ciprofloxacin | 0
    multisensitive to amoxicillin/clavulanic | 0
    pathological analysis showing acute inflammation of appendicular muscularis | 0
    no inflammation of mucosa | 0
    no perforation | 0
    periappendicular inflammation of fatty tissue | 0
    no bronchospasm | 0
    no oral swelling | 0
    no respiratory distress | 0
    unexplained cutaneous flushing | 0
    R. ornithinolytica septic shock | 0
    appendicitis | 0
    severe acute kidney failure | 0
    