Event|Timestamp (hours)
trismus and hypertonia|-336
injured leg|-336
treatment with immunoglobulins, tetanus vaccination, and metronidazole|-336
transferred to ICU|-336
tracheostomy|-336
mechanical ventilation|-336
vasoactive support|-336
treated with baclofen, midazolam, and diazepam|-336
severely slow cerebral activity|-336
opacity on chest radiography|-336
peripheral leukocytosis|-336
tracheal secretions tested positive for Klebsiella pneumoniae and MSSA|-336
antibiotic therapy with piperacillin-tazobactam|-336
moved to geriatric unit|-336
coma|-336
breathed spontaneously on 4 L/min of supplemental oxygen|-336
antibiotic therapy switched to linezolid|-336
combined treatment with meropenem|-336
awoke|-336
feeding tube removed|-336
developed cholestasis|-336
acute edematous pancreatitis|-336
urinary tract infection|-336
treated with colistin and amoxicillin-clavulanate|-336
clinical condition improved|-336
placed in MDRO isolation|0
required tracheal supplemental oxygen (1 L/min)|0
bladder catheter|0
developed pressure ulcers|0
sarcopenic|0
low handgrip strength|0
appendicular skeletal mass (ASM)|0
underwent rehabilitation|0
Clostridioides difficile infection|0
oral vancomycin prescribed|0
AF with a third-degree atrioventricular block|0
transferred to cardiac ICU|0
single-chamber pacemaker implantation|0
hyperkinetic delirium|0
transferred to hospital|0
Pseudomonas aeruginosa bloodstream infection|0
treated with ceftazidime-avibactam and amikacin|0
tested positive for SARS-CoV-2|0
treated with remdesivir|0
second recurrence of C. difficile|0
transferred to geriatric medicine unit|0
treated with fidaxomicin|0
bloodstream infection due to Candida parapsilosis, MSSA, and Candida tropicalis|0
infected catheter replaced|0
treated with caspofungin and cefazolin|0
bloodstream infection caused by P. aeruginosa|0
antibiotic treatment with piperacillin-tazobactam|0
shifted to aztreonam and ceftazidime-avibactam|0
shifted to cefepime|0
tracheostomy closure|0
nutritional supplementation prescribed|0
intensive rehabilitation compromised|0
short physiotherapy sessions|0
able to perform postural transition with assistance|0
motor and respiratory reconditioning continued|0
posture transition training and aided transfers|0
axial stability and balance improvement exercises|0
breath-movement coordination exercises|0
thoracic expansion and girdle opening exercises|0
inhalation-exhalation exercises|0
wheelchairs and walkers recommended|0
rehabilitation, ENT, and geriatric follow-up evaluations recommended|0