68 years old | 0
    man | 0
    admitted to the hospital | 0
    right forearm bite | -24
    superficial right forearm bite | -24
    swollen right forearm | -24
    cyanotic right forearm | -24
    general discomfort | -4
    injury lesion not washed | -24
    injury lesion not disinfected | -24
    swelling distal right upper extremity | -8
    pain distal right upper extremity | -8
    diagnosed with gout arthritis | -8
    nonsteroidal anti-inflammatory treatment | -8
    gradual worsening swelling | -8
    gradual worsening pain | -8
    purpura around wound | -8
    purpura right hand | -8
    weakness | -8
    palpitation | -8
    cold sweats | -8
    acute pain | 0
    shock | 0
    hypotension | 0
    rapid pulse | 0
    cold sweats | 0
    flaky plaques right upper limb | 0
    swelling right upper limb | 0
    weak iliac artery pulsation | 0
    dopamine administered | 0
    laboratory examinations conducted | 0
    imaging examinations conducted | 0
    multidisciplinary medical treatment organized | 0
    swelling continued expansion | 0
    ecchymosis continued expansion | 0
    crepitus subcutaneous soft tissue | 0
    gas bubbles subcutaneous tissue | 0
    edema subcutaneous tissue | 0
    anti-infection treatment administered | 0
    limb lesions continued expansion | 0
    deterioration of consciousness | 0
    white blood cell count 4.85 × 10⁹/L | 0
    hemoglobin 70 g/L | 0
    platelet count 36 × 10⁹/L | 0
    C-reactive protein 68.35 mg/L | 0
    procalcitonin 48.960 ng/mL | 0
    normal blood coagulation | 0
    gas in soft tissue right hand | 0
    gas in soft tissue right forearm | 0
    Gram-negative bacilli in bite wound | 0
    gas gangrene-like infection | 0
    open amputation performed | 0
    fish mouth incision | 0
    proximal to lesion | 0
    vascular nerves disconnected | 0
    blood vessels ligated | 0
    humerus bone cut | 0
    stump trimmed | 0
    proximal muscles responded to electrotome | 0
    muscle sutured to bone end | 0
    wound not sutured | 0
    sterile wound dressing applied | 0
    ICU isolation treatment | 0
    endotracheal intubation | 0
    malodorous gas escaped | 0
    necrotic lesions | 0
    dark purple lesions | 0
    dissolved tissues | 0
    penicillin administered | 0
    meropenem administered | 0
    clindamycin administered | 0
    vasoactive drugs administered | 0
    intermittent fever | 24
    fever 40°C | 24
    elevated infection index | 24
    elevated procalcitonin | 24
    elevated C-reactive protein | 24
    decreased infection index | 72
    decreased procalcitonin | 72
    decreased C-reactive protein | 72
    low hemoglobin | 0
    low platelet count | 0
    Aeromonas hydrophila cultured | 72
    necrotic tissue | 0
    inflammatory cell infiltration | 0
    original granulocytes 16.5% | 72
    original naive mononuclear cells 21.0% | 72
    mild myeloid hyperplasia | 72
    decreased megakaryocytes | 72
    interstitial edema | 72
    megakaryocyte reduction | 72
    AML diagnosis | 72
    MDS revised to AML | 72
    wound dressing replaced daily | 0
    foul odor stump tissue | 72
    exudate stump tissue | 72
    muscle tissue necrosis | 72
    ecchymoses around wound | 72
    stump trimmed | 168
    necrotic tissue removed | 168
    6 cm humerus removed | 168
    wound sutured layer by layer | 168
    vacuum sponge applied | 168
    vacuum sponge removed | 240
    foul odor after first surgery | 72
    exudate after first surgery | 72
    muscle necrosis after first surgery | 72
    ecchymoses after first surgery | 72
    vital signs recovered | 264
    hemoglobin recovered | 264
    platelet count recovered | 264
    extubated | 264
    spontaneous breathing resumed | 264
    clear consciousness | 264
    wound healed | 264
    discharged | 264
    AML chemotherapy refused | 264
    died from blood system disease | 17520
    