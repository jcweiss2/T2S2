25 years old | 0\
female | 0\
admitted to the hospital | 0\
severe pain | -24\
shortness of breath | -24\
worsening pain | -24\
tachypneic | -24\
oxygen saturation 56% | -24\
tachycardia | -24\
pulse 121 bpm | -24\
afebrile 36°C | -24\
hypotensive | -24\
blood pressure 56/30 mmHg | -24\
noradrenaline infusion | -24\
IV heparin 5000 units | -24\
IV amoxicillin-clavulanate | -24\
electively intubated | 0\
metabolic acidosis | 0\
lactic acidosis | 0\
respiratory distress | 0\
grossly swollen right thigh | 0\
extensive blistering ecchymotic patches | 0\
necrotizing fasciitis | 0\
septicemic shock | 0\
acute kidney injury | 0\
rhabdomyolysis | 0\
coagulopathy | 0\
thrombocytopenia | 0\
ischemic hepatitis | 0\
IV meropenem | 0\
IV clindamycin | 0\
IV vancomycin | 0\
high vaginal swab | 0\
CT pulmonary angiography | 0\
bedside echocardiography | 0\
intravenous immunoglobulin | 0\
continuous veno-venous hemofiltration | 0\
critical condition | 0\
required 4 inotropes | 0\
skin lesion spread | 24\
bluish discoloration | 24\
blistering | 24\
Gram positive cocci in chains | 24\
S. pyogenes | 24\
multidisciplinary discussion | 144\
IV clindamycin | 144\
IV crystalline penicillin G | 144\
CVVH | 144\
succumbed to death | 168\
septic shock | 168\
tissue necrosis | 168\
toxic shock syndrome | 168