74 years old | 0
female | 0
admitted to the emergency department | -24
dizziness | -24
emphysematous chronic obstructive pulmonary disease | -24
smoking habit | -24
severe chronic ischemic heart disease | -24
hypercholesterolemia | -24
hypoxemic respiratory failure | -24
SpO2 82% | -24
respiratory frequency 24/min | -24
oxygen therapy with Venturi mask started | -24
electrocardiogram negative for ischemia | -24
body temperature 37.6°C | -24
lymphopenia | -24
C-reactive protein increase | -24
chest HRCT performed | -24
centrilobular emphysema | -24
ground glass opacity areas at ventral segment of superior right lobe | -24
ground glass opacity areas at lateral segment of middle right lobe | -24
tested for Coronavirus-19 | -24
positive real-time polymerase chain reaction | -24
admitted to the medicine department | 0
therapy with hydroxychloroquine started | 0
therapy with azithromycin started | 0
deteriorated | 168
admitted to the intensive care unit | 168
admitted to Covid-19 Sub8ICU | 168
noninvasive mechanical ventilation started | 168
intubation not indicated | 168
received 8 mg/kg tocilizumab | 168
methylprednisolone 1 mg/kg started | 168
enoxaparin 100 U/kg 2 times a day started | 168
respiratory failure improved | 216
HRCT repeated | 480
regression of ground glass opacities | 480
arterial blood gasses showed improvement of hypoxemia | 480
arterial oxygen partial pressure/fraction of inspired oxygen ratio 176 mm Hg | 480
discontinuation of noninvasive mechanical ventilation | 480
high flow oxygen required | 480
clinical conditions deteriorated | 528
increasing respiratory frequency | 528
worsening of hypoxemia | 528
new chest HRCT performed | 528
increasing basal nonspecific ground glass opacities | 528
sign of loss of volume | 528
traction bronchiectasis | 528
gram-positive sepsis | 528
treated with linezolid | 528
respiratory conditions worsened | 528
noninvasive mechanical ventilation started again | 528
arterial blood gasses showed very severe hypoxemic respiratory failure | 1320
arterial oxygen partial pressure/fraction of inspired oxygen ratio less than 40 mm Hg | 1320
last chest HRCT performed | 1320
radiological progression of pulmonary fibrosis at inferior lobes | 1320
global architecture distortion | 1320
died | 1440
severe hypoxemic respiratory failure | 1440
