male | 0 | 0 
premature birth | -672 | -672 
emergency cesarean delivery | -672 | -672 
abruptio placenta | -672 | -672 
birth weight 1090g | -672 | -672 
Apgar 4 and 8 | -672 | -672 
respiratory distress | -672 | 0 
respiratory rate 65 breaths per min | -672 | 0 
chest retraction | -672 | 0 
CPAP machine | -672 | 168 
positive end expiratory pressures | -672 | 168 
inspired oxygen 30% | -672 | 168 
cloudy eyes | 0 | 0 
ectropion | 0 | 0 
dry ichthyotic skin | 0 | 0 
undescended testicles | 0 | 0 
height 75th percentile | 0 | 0 
weight 25th percentile | 0 | 0 
head circumference 25th percentile | 0 | 0 
temperature 36.2°C | 0 | 0 
heart rate 167 beats per min | 0 | 0 
normal neurological examination | 0 | 0 
normal breath sounds | 0 | 0 
no organomegaly | 0 | 0 
normal blood count | 0 | 0 
normal electrolytes | 0 | 0 
normal liver function | 0 | 0 
respiratory distress syndrome | 0 | 168 
ground-glass opacity | 0 | 168 
minor respiratory acidosis | 0 | 168 
surfactant dosage | 0 | 168 
trophic feeding | 72 | 168 
bowel movement | 12 | 12 
abdominal distension | 144 | 144 
tachycardia | 144 | 144 
tachypnea | 144 | 144 
thrombocytopenia | 144 | 144 
neutropenia | 144 | 144 
elevated C-reactive protein | 144 | 144 
meropenem and vancomycin | 144 | 216 
stopped trophic feeding | 144 | 144 
restarted feeding | 216 | 216 
high-flow oxygen treatment | 168 | 1008 
relapses of unexplained apnea | 504 | 1008 
septic examination negative | 504 | 1008 
normal brain MRI | 504 | 504 
nasogastric tube | 504 | 1008 
conjugated hyperbilirubinemia | 504 | 1008 
neonatal cholestasis workup | 504 | 1008 
normal echocardiogram | 504 | 504 
normal eye test | 504 | 504 
craniosynostosis | 504 | 504 
hepatosplenomegaly not seen | 504 | 504 
no biliary atresia | 504 | 504 
normal-appearing gallbladder | 504 | 504 
no intrahepatic or extrahepatic biliary tree dilatation | 504 | 504 
declining albumin level | 504 | 1008 
elevated bilirubin | 504 | 1008 
elevated AST and ALT | 504 | 1008 
multiple albumin infusions | 504 | 1008 
ursodeoxycholic acid treatment | 504 | 1008 
infectious etiology investigation | 504 | 1008 
negative results | 504 | 1008 
normal TSH, T3, T4, and cortisol levels | 504 | 504 
negative metabolic disorders | 504 | 504 
caffeine treatment | 504 | 1008 
hemoglobin optimization | 504 | 1008 
phenobarbitone treatment | 504 | 1008 
severe cyanosis | 912 | 912 
apnea | 912 | 912 
bradycardia | 912 | 912 
cardio-respiratory resuscitation | 912 | 912 
intubation | 912 | 912 
mechanical breathing | 912 | 912 
epinephrine | 912 | 912 
septic shock | 912 | 1008 
multiorgan failure | 912 | 1008 
disseminated intravascular coagulation | 912 | 1008 
acute renal damage | 912 | 1008 
capillary leak syndrome | 912 | 1008 
inotropic support | 912 | 1008 
high-frequency oscillating ventilation | 912 | 1008 
continuous inhaled nitric oxide treatment | 912 | 1008 
death | 1008 | 1008 
whole-exome sequencing | 1008 | 1008 
NOTCH2 gene mutation | 1008 | 1008 
pathogenic heterozygous variant c.1076c>T (Ser359Phe) | 1008 | 1008 
ALGS2 diagnosis | 1008 | 1008 
genetic counseling | 1008 | 1008