57 years old | 0
    male | 0
    hypertension | 0
    presented to the emergency room | 0
    fever | -216
    chills | -216
    shortness of breath | -216
    malaise | -216
    poor appetite | -216
    oxygen saturation of 64% | 0
    bilateral crackles | 0
    leukocyte count within normal range | 0
    elevated procalcitonin | 0
    SARS-CoV-2 positive | 0
    sputum Gram stain 10–25 WBCs/LPF | 0
    methicillin susceptible Staphylococcus aureus | 0
    oropharyngeal microbiota | 0
    bilateral patchy airspace disease | 0
    increased interstitial opacities | 0
    severe COVID-19 disease | 0
    oral dexamethasone | 0
    intravenous remdesivir | 0
    oxygen support via non-rebreather mask | 0
    intravenous azithromycin | 0
    intravenous ceftriaxone | 0
    persistent hypoxia | 0
    inability to wean from non-rebreather mask | 0
    steroids continued beyond day 10 | 216
    clinical condition worsened | 336
    cyanotic | 336
    dyspneic | 336
    endotracheal intubation | 336
    progression of infiltrates | 336
    vancomycin initiated | 336
    meropenem initiated | 336
    oral dexamethasone changed to intravenous methylprednisolone | 336
    worsening renal function | 336
    continuous renal replacement therapy | 336
    periods of hypotension | 336
    diarrhea | 792
    Candida colitis | 792
    nystatin administered | 792
    hypoxia | 864
    hypotension | 864
    methylprednisolone changed to hydrocortisone | 864
    midodrine added | 864
    blood cultures revealed yeast | 864
    micafungin administered | 864
    antibiotics discontinued | 864
    Cryptococcus neoformans identified | 864
    lumbar puncture performed | 864
    opening pressure 28 cm H2O | 864
    cerebrospinal fluid 185 WBCs/μL | 864
    65,000 RBCs/μL | 864
    positive India ink | 864
    Cryptococcus neoformans culture confirmed | 864
    cerebrospinal fluid cryptococcal antigen positive | 864
    HIV negative | 864
    micafungin discontinued | 864
    liposomal amphotericin B administered | 864
    flucytosine administered | 864
    repeated lumbar punctures | 936
    opening pressures less than 20 cm H2O | 936
    new skin nodules | 960
    disseminated cryptococcal infection | 960
    died | 1008
    hypotensive episode | 1008
    