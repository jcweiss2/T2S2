23 years old | 0
male | 0
normal karyotype pre-B acute lymphoblastic leukemia | -672
FLAM protocol chemotherapy | -672
cyclophosphamide | 0
cytarabine | 0
pegaspargase | 0
fever | 48
abdominal pain | 48
diarrhea | 48
piperacillin/tazobactam | 48
fluconazole | 48
nifuroxazide | 48
temperature returned to normal | 72
symptoms receded | 72
condition improved | 72
fever | 168
abdominal pain | 168
diarrhea | 168
granulocytopenia | 168
WBC 0.1–0.0 G/l | 168
meropenem | 168
metronidazole | 168
itraconazole | 168
G-CSF | 168
filgrastim | 168
temperature returned to normal | 216
abdominal pain subsided | 216
nifuroxazide continued | 216
G-CSF continued | 216
agranulocytosis | 216
asymptomatic | 240
second cycle of chemotherapy | 432
fever | 434
abdominal pain | 434
diarrhea | 434
Candida albicans | 434
ketoconazole | 434
piperacillin/tazobactam | 434
vancomycin | 434
G-CSF | 434
Enterobacter cloacae | 434
improvement of general condition | 434
reduction of abdominal pain | 434
fever | 522
vomiting | 522
acute pain in right epigastrium | 522
abdominal ultrasound | 522
acalculous gallbladder | 522
wall thickening | 522
pericholecystic fluid | 522
acalculous cholecystitis | 522
broad spectrum antibiotic regimen | 522
G-CSF | 522
intravenous fluids | 522
fasting | 522
condition deteriorated | 528
renal failure | 528
liver failure | 528
life-saving surgery | 528
laparoscopic cholecystectomy | 528
platelet concentrate transfused | 528
platelet count increased | 528
histopathological evidence | 528
lymphocyte infiltration | 528
hyperemia | 528
no neutrophil infiltrations | 528
no leukemia cells | 528
no bacteria | 528
no fungal cells | 528
bile culture | 528
no micro-organisms | 528
intensive care ward | 528
broad spectrum antibiotic regimen | 528
G-CSF | 528
erythrocyte concentrate transfused | 528
PC transfused | 528
fever | 552
lower peripheral blood pressure | 552
atelectatic-inflammatory changes | 552
imipenem/cilastatin sodium | 552
vancomycin | 552
metronidazole | 552
teicoplanin | 552
ketoconazole | 552
ciprofloxacin hydrochloride | 552
co-trimoxazole | 552
therapy effective | 552
condition improved | 552
no abdominal symptoms | 576
abdominal pain | 576
diarrhea | 576
permitted to eat | 600
light diet | 600
well tolerated | 600
improvement in peripheral blood | 612
G-CSF discontinued | 612
antibiotic therapy discontinued | 614
transferred to Department of Hematology | 648
discharged from hospital | 816