28 years old | 0
female | 0
admitted to the hospital | 0
twin pregnancy | 0
Sheehan syndrome | 0
hypothyroidism | -17280
equivocal serum cortisol levels | -17280
pituitary apoplexy | -17280
tablet hydrocortisone | -17280
tablet thyroxine | -17280
intrauterine insemination | -17280
diamniotic monochorionic twins | 0
gestational diabetes mellitus | -168
elective lower segment cesarean section | 0
multiple metabolic derangements | 0
intrauterine growth retardation | 0
nil per oral | -8
tablet thyroxine | -8
tablet ranitidine | -8
tablet metoclopramide | -8
fasting blood sugar | 0
withheld insulin | 0
injection hydrocortisone | 0
hydrocortisone infusion | 0
subarachnoid block | 0
general anesthesia backup | 0
invasive blood pressure monitoring | 0
arterial cannula placement | 0
supplemental oxygen | 0
hyperbaric bupivacaine | 0
fentanyl | 0
left lateral tilt | 0
T4 block level | 0
lower segment cesarean section | 0
hemostasis | 0
hypotension episodes | 6
phenylephrine bolus | 6
live male babies | 0
APGAR scores | 0
neonatal intensive care unit | 0
oxytocin infusion | 0
intraoperative blood loss | 0
normal ABG | 0
normal blood sugar levels | 0
T10 block regression | 120
high dependency unit | 48
injection paracetamol | 48
uneventful postoperative period | 168
pyrexia | -17520
pyonephritis | -17520
severe hyperglycemia | -17520
metabolic acidosis | -17520
acute kidney injury | -17520
septicemic shock | -17520
bilateral pleural effusion | -17520
respiratory distress | -17520
loss of fetus | -17520
drainage of pus | -17520
broad-spectrum antibiotics | -17520
hemodialysis | -17520
difficulty conceiving | -17280
anemia | 0
postpartum hemorrhage | 0
sepsis | -17520
hypotension | -17520
delayed awakening | 0
residual neuromuscular blockade | 0
postoperative mechanical ventilation | 0
hypotension requiring inotropes | 0
delayed emergence from anesthesia | 0
perioperative stress management | 0
steroid management | 0
postoperative gastrointestinal complications | 0
neuropsychiatric complications | 0
electrolyte disturbances | 0
coagulation disturbances | 0
core body temperature decrease | 0
reduced anesthetic drug requirement | 0
successful anesthetic management | 0
