65 years old | 0
female | 0
admitted to the hospital | 0
stage IIIA lung cancer | -648
smoking history | -648
hypertension | -648
hypothyroidism | -648
dyslipidemia | -648
spiculated suprahilar RUL nodule | -648
lung-RADS 4X | -648
PET/CT scan | -648
bronchoscopy | -648
NSCLC | -648
adenocarcinoma | -648
lymph node sampling | -648
surgical resection | -648
carboplatin | -567
paclitaxel | -567
radiation therapy | -567
CT scan | -567
adjuvant immunotherapy | -567
durvalumab | -567
pneumonitis | -567
steroid taper | -567
staging chest CT | -567
abdominal pain | -24
pancreatic head lesion | -24
abdominal and pelvic CT scan | -24
epigastric pain | -12
constipation | -12
loss of appetite | -12
weight loss | -12
endoscopic ultra-sound-guided biopsy | 0
pancreatic mass | 0
tumor cells | 0
CK7 | 0
TTF-1 | 0
Napsin-A | 0
CDX-2 | 0
KOC | 0
synaptophysin | 0
Smad-4 | 0
PET/CT scan | 12
brain MRI scan | 12
palliative radiation therapy | 24
carboplatin | 24
pemetrexed | 24
chemotherapy | 24
electrolyte derangements | 48
acute anemia | 48
hemoglobin nadir | 48
transfusion | 48
CT scan | 48
left lower lobe nodule | 48
staging PET/CT scan | 72
dyspnea | 96
cough | 96
generalized weakness | 96
rapid response | 96
oxygen supplementation | 96
bilevel-positive airway pressure | 96
broad-spectrum antibiotics | 96
vancomycin | 96
azithromycin | 96
cefepime | 96
altered mentation | 102
worsening hypoxemia | 102
vasopressor support | 102
palliative medicine team | 102
inpatient hospice care | 108
death | 108