50 years old | 0
    man | 0
    admitted to the emergency department | 0
    high spiking fever | 0
    disorientation | 0
    antiphospholipid syndrome | -2160
    deep vein thrombosis | -2160
    ischemic stroke | -2160
    warfarin | -2160
    prosthetic tissue aortic valve replacement | -2160
    aortic stenosis | -2160
    admitted to another hospital | -2160
    brainstem hemorrhage | -2160
    nosocomial pneumonia | -2160
    severe renal failure | -2160
    hemodialysis | -2160
    permacath | -2160
    anticoagulant therapy switched to enoxaparin | -2160
    permacath retained | -2160
    permacath removal not attended | -2160
    temperature of 39°C | 0
    blood pressure of 80/50 mmHg | 0
    pulse of 128 beats per minute | 0
    oxygen saturation of 88% | 0
    disorientation | 0
    no obvious foci of infection | 0
    leukocytosis of 20,000 per cubic millimeter | 0
    hemoglobin concentration of 12 g/dL | 0
    platelets count of 550,000 per cubic millimeter | 0
    blood urea nitrogen slightly elevated | 0
    creatinine levels slightly elevated | 0
    chest x-ray normal | 0
    microscopic hematuria | 0
    blood culture drawn | 0
    urine culture drawn | 0
    permacath extracted | 0
    vancomycin | 0
    piperacillin-tazobactam | 0
    amikacin |9 0
    vasopressors | 0
    admitted to intensive care unit | 0
    blood cultures grew MRSA susceptible to vancomycin | 24
    MRSA susceptible to daptomycin | 24
    MRSA susceptible to rifampin | 24
    MRSA susceptible to TMP/SMX | 24
    permacath tip cultures yielded MRSA | 24
    transthoracic echocardiogram normal | 24
    condition stabilized | 48
    transferred to medical ward | 48
    treated with vancomycin | 48
    treated with rifampin | 48
    fever persisted | 48
    blood cultures grew MRSA | 48
    MRSA susceptible to vancomycin | 48
    MRSA resistant to rifampin | 48
    antimicrobial therapy switched to vancomycin plus piperacillin-tazobactam | 48
    TEE showed thrombus in SVC | 144
    whole body CT scan normal | 144
    antimicrobial therapy switched to daptomycin plus oxacillin | 144
    bacteremic with MRSA | 144
    MRSA non-susceptible to daptomycin | 144
    MRSA resistant to vancomycin | 144
    daptomycin dose increased to 12 mg/kg | 168
    TMP/SMX added | 168
    MRSA bacteremia cleared | 216
    enoxaparin continued | 216
    therapeutic anti Xa levels | 216
    serial blood cultures sterile | 216
    cardiac arrest | 288
    asystole | 288
    died | 288
    MRSA genotype sequence type 5 | 0
    MRSA spa type t002 | 0
    septic thrombus formation | 0
    SVC thrombosis | 0
    MRSA bacteremia persisted | 0
    asymptomatic | 0
    hemodynamically stable | 0
    anticoagulation | 0
    thrombus dislodgement | 288
    massive pulmonary embolus | 288
    no SVC syndrome | 0
    no signs of SVC syndrome | 0
    autopsy refused | 288
    <|eot_id|>
    