72 years old | 0
male | 0
admitted to the hospital | 0
shortness of breath | -72
intermittent chest pain | -72
altered level of consciousness | 0
respiratory distress | 0
heart rate of 122 beats/min | 0
blood pressure of 86/46 mm Hg | 0
respiratory rate of 43 breaths/min | 0
oxygen saturations of 78% on room air | 0
temperature of 37.8°C | 0
sinus tachycardia | 0
thready central and peripheral pulses | 0
elevated jugular venous pressure | 0
S1 and S2 were present | 0
absence of murmurs or extra heart sounds | 0
extremities were mottled and cool | 0
bilateral peripheral edema | 0
breath sounds were diminished at the lung bases | 0
diffuse crepitations bilaterally | 0
abdominal examination was unremarkable | 0
hypertension | -672
dyslipidemia | -672
type 2 diabetes mellitus | -672
oral anti-hyperglycemic medications | -672
40 pack-year smoking history | -672
atypical chest discomfort | -1344
myocardial perfusion imaging | -1344
mild ischemia in the left anterior descending artery | -1344
medical therapy | -1344
coronary angiogram scheduled | -1344
severe interstitial pulmonary edema | 0
inferolateral ST-segment elevation | 0
white blood cell count 8.4 × 10^9/L | 0
hemoglobin 104 g/L | 0
whole blood lactate 4.0 mmol/L | 0
creatinine kinase 1,178 μ/L | 0
high sensitivity troponin T 3,482 ng/L | 0
Killip IV inferolateral ST-segment elevation myocardial infarction | 0
intubated for hypoxemic respiratory failure | 0
emergency coronary angiogram | 0
culprit lesion in the proximal to mid LAD | 0
revascularized with 2 drug-eluding stents | 0
chronic total occlusion of the mid right coronary artery | 0
collaterals from the LAD and left circumflex | 0
intra-aortic balloon pump | 0
transferred to the cardiac intensive care unit | 0
severe left ventricular dysfunction | 0
ejection fraction estimated at 20% | 0
akinesis of the mid to distal anterior, apex, inferior, and lateral walls | 0
absence of left ventricular thrombus | 0
hemodynamically significant valvular disease | 0
pericardial effusion | 0
abnormalities of the myocardium | 0
shock state persisted | 0
requirements of the intra-aortic balloon pump | 0
multiple vasoactive and inotropic medications | 0
norepinephrine | 0
vasopressin | 0
phenylephrine | 0
dobutamine | 0
oliguric renal failure | 0
continuous renal replacement therapy | 0
borderline fevers | 0
broad spectrum antimicrobial therapy | 0
piperacillin/tazobactam | 0
vancomycin | 0
blood cultures returned positive | 12
gram-negative bacilli | 12
Enterobacter cloacae | 12
antimicrobial therapy escalated to meropenem | 12
mixed distributive/septic and cardiogenic shock | 0
recurrent ischemia secondary to stent complication | 0
evolving mechanical complication of acute coronary syndrome | 0
ventricular free wall rupture | 0
ventricular septal rupture | 0
papillary muscle rupture | 0
acute mitral regurgitation | 0
abrupt pulseless electrical activity cardiac arrest | 48
large circumferential pericardial effusion | 48
emergency pericardiocentesis | 48
pericardial effusion relentlessly reaccumulated | 48
refractory cardiac tamponade | 48
mechanical circulatory support | 48
uncontrolled septicemia | 48
multiorgan dysfunction | 48
baseline frailty | 48
prohibitive surgical risk | 48
resuscitation efforts were ultimately unsuccessful | 48
cause of death suspected to be secondary to left ventricular FWR | 48
large transmural myocardial infarction | 48
extensive necrosis | 48
extensive multiple myocardial abscesses | 48
gram-negative rods | 48
left ventricular FWR of the mid inferior wall | 48
hemopericardium | 48
severe acute pyelonephritis of the left kidney | 48
source of infection | 48
late presenting Killip IV inferolateral ST-segment elevation myocardial infarction | 0
septic shock with E cloacae bacteremia | 0
acute pyelonephritis | 0
left ventricular FWR at the site of a septic myocardial abscess | 48
discharged | -1