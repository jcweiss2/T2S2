69 years old | 0
    male | 0
    admitted to medical intensive care unit | 0
    cough | -72
    sputum | -72
    fever | 0
    drowsy mental status | 0
    traumatic intracranial hemorrhage | -5088
    epidural hemorrhage | -5088
    subdural hemorrhage | -5088
    accidental fall | -5088
    right craniectomy | -5088
    ventriculoperitoneal shunt placement | -5088
    posttraumatic hydrocephalus | -5088
    intensive rehabilitation treatment | -2688
    able to communicate with others | -2688
    walk with walker | -2688
    feed himself | -2688
    drowsy after ingesting antipsychotic medication | -168
    aggressive behaviors | -168
    aspiration event | -168
    respiratory symptoms | -168
    deteriorating mental status | -168
    chest radiography | 0
    focal infiltrate at left lower lung field | 0
    chest computed tomography | 0
    consolidation with air bronchogram at left lower lobe posterior basal segment | 0
    suspected aspirated materials at left upper lobe bronchus | 0
    suspected aspirated materials at left lower lobe segmental bronchus | 0
    appearance of food particles in esophagus | 0
    aspiration-induced pneumonia | 0
    brain CT scan | 0
    previously inserted ventriculoperitoneal shunt | 0
    focal encephalomalacic changes in right frontal lobe | 0
    mental change due to pneumonia-induced sepsis | 0
    PaO2 43.9 mm Hg | 0
    SaO2 79.4% | 0
    respiratory rate 24 breaths/minute | 0
    comfortable respiration | 0
    high-flow nasal oxygen therapy with FiO2 0.5 | 0
    flow 50 L/minute | 0
    flow increased to 60 L/minute | 0
    FiO2 decreased to 0.4 | 0
    SpO2 93-97% | 0
    respiratory rate 22-26 breaths/minute | 0
    repeated sudden desaturation | 24
    endotracheal intubation | 24
    mechanical ventilation | 24
    desaturation due to airway secretion | 24
    attempted weaning from mechanical ventilation | 48
    unable to effectively expectorate airway secretions | 48
    volume of secretions decreased | 48
    alert mental status | 48
    extubated | 48
    HFNC to prevent postextubation respiratory failure | 48
    HFNC FiO2 0.4 | 48
    HFNC flow 50 L/minute | 48
    SpO2 93!100% | 48
    transferred to general ward | 72
    HFNC flow changed to 40 L/minute | 72
    mentation became drowsy | 100
    stupor | 100
    brain CT scan | 100
    pneumocephalus | 100
    midline shifting | 100
    near-collapse of left ventricle | 100
    Mount Fuji sign | 100
    tension pneumocephalus | 100
    HFNC stopped | 100
    changed to simple nasal cannula | 100
    follow-up brain CT scan | 112
    pneumocephalus slightly decreased | 112
    facial bone CT scan | 112
    skull base fractures at right frontal and ethmoidal sinuses | 112
    mental status improved from stupor to drowsy | 112
    follow-up brain CT | 184
    pneumocephalus markedly decreased | 184
    midline shifting improved | 184
    left ventricle structure improved | 184
    pneumocephalus nearly resolved | 480
    difficulties in expectorating airway secretions | 480
    tracheostomy | 480
    mental status improved | 480
    sudden decline in mental status | 960
    stupor | 960
    intracranial infection | 960
    craniotomy for drainage | 960
    mental status did not fully recover | 960
    death | 960