9 years old | 0
male | 0
neutered | 0
domestic shorthair | 0
admitted to the hospital | 0
weakness | -72
suspected signs of lower urinary tract disease | -72
severe cardiovascular collapse | -1
referred to tertiary referral hospital | -1
obtunded | 0
prolonged capillary refill time | 0
bradycardia | 0
hypothermia | 0
weak femoral pulses | 0
blood pressure too low to detect | 0
intravenous bolus of lactated Ringer’s solution | 0
fluid rate of 29 ml/h | 0
point-of-care ultrasound of the thorax and abdomen | 0
moderate volume of free abdominal fluid | 0
no evidence of pleural/pericardial effusion or B-lines | 0
atrial standstill with idioventricular escape rhythms | 0
jugular venous sample obtained | 0
minimum database and blood gas analysis | 0
severe metabolic acidosis | 0
hyperkalemia | 0
presumptive diagnosis of uroabdomen | 0
abdominocentesis | 0
serosanguinous fluid | 0
fluid analysis consistent with uroabdomen | 0
cytological analysis of the fluid | 0
intracellular bacteria | 0
concern of urosepsis | 0
ceftazidime added to treatments | 0
7F × 13 cm triple-lumen central venous line placed | 2
percutaneously using a modified Seldinger technique | 2
local block to the abdominal wall | 2
urinary catheter placed | 2
connected to a closed urine collection system | 2
moderate degree of difficulty in passing the urinary catheter | 2
concern for urethral obstruction | 2
IV administration of a 10 ml/kg bolus of lactated Ringer’s solution | 2
monitoring of arterial blood pressure, heart rate and capillary refill time | 2
systolic blood pressure increased to 110 mmHg | 4
heart rate increased to 180 beats/min | 4
capillary refill time decreased to <2 s | 4
ECG rhythm changed to a sinus rhythm | 4
external heat support provided | 4
cat’s temperature returned to normal | 4
pain management initiated with injectable tramadol | 4
peritoneal dialysis performed | 8
peritoneal dialysis solution created | 8
initial dialysate volume of exchange | 8
dialysate infusion | 8
dwell time | 8
fluid removal by gravity | 8
treatment repeated every 2 h for the first 12 h | 8
volume of dialysate infusion increased | 8
blood gas analysis revealed improvement in electrolyte and pH values | 8
no complications observed with increased volume of dialysate infusion | 8
cat appeared brighter and more responsive | 8
diagnostic abdominal ultrasound performed | 18
evidence of large volume of gravity-dependent sediment in the urinary bladder | 18
suspected rupture at the dorsal aspect of the urinary bladder | 18
fever | 18
clindamycin added to antibiotic protocol | 18
cat remained stable | 18
recheck bloodwork showed significant improvement of azotemia, glucose and lactate | 36
peritoneal drainage/dialysis catheter removed | 36
retrograde contrast cystography performed | 36
evidence of urinary bladder rupture | 36
exploratory laparotomy performed | 36
urinary rupture site surgically corrected | 36
full-thickness urinary bladder biopsy samples obtained | 36
point-of-care ultrasound of the abdomen and chest performed | 36
mild-to-moderate volume of bilateral pleural effusion | 36
complete echocardiogram performed | 36
no evidence of cardiac disease or fluid overload | 36
total fluid balance negative 240 ml | 36
cat appeared clinically euhydrated and euvolemic | 36
thoracocentesis performed | 36
fluid analysis revealed a pure transudate | 36
paired blood sample obtained | 36
creatinine ratio consistent with diagnosis of urothorax | 36
cat recovered uneventfully from surgery | 48
no signs of respiratory distress noted | 48
pleural effusion slowly resolved | 48
culture and sensitivity results from urinary bladder wall showed Klebsiella pneumoniae and Mannheimia haemolytica | 48
enrofloxacin added to treatment protocol | 48
cat discharged 4 days later | 96
no further medical intervention required | 96
point-of-care ultrasound evaluation showed no abdominal or pleural fluid | 168