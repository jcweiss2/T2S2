17 years old | 0
African American | 0
male | 0
admitted to the hospital | 0
past medical history of depression | -672
nonbilious vomiting | -72
new-onset erythematous blanching macular rash | -72
tachycardic | 0
hypertensive | 0
febrile | 0
temperature of 38.5°C | 0
hypotensive | 4
tachycardic | 4
septic shock | 4
blood cultures drawn | 4
empiric antibiotic treatment | 4
hyponatremia | 0
direct hyperbilirubinemia | 0
low lactate dehydrogenase | 0
polymorphic neutrophil dominant leukocytosis | 0
elevated C-reactive protein | 0
sterile pyuria | 0
direct hyperbilirubinemia continued to rise | 192
γ-glutamyl transferase remained within normal limits | 192
lipase remained within normal limits | 192
amylase remained within normal limits | 192
transaminases remained within normal limits | 192
alanine aminotransferase at the high end of the normal range | 192
ultrasound showed an over distended gallbladder | 192
computed tomography was negative | 192
magnetic resonance cholangiopancreatography was negative | 192
infectious disease workup was negative | 192
hypotensive | 0
tachycardic | 0
S3 gallop | 0
orthopnea | 0
elevated brain natriuretic peptide | 0
respiratory distress | 0
bilateral lower lobe pleural effusions | 0
mild decrease in left ventricular function | 0
mild mitral and tricuspid valve regurgitation | 0
small posterior pericardial effusion | 0
transferred to the pediatric intensive care unit | 0
heart failure stabilized | 24
respiratory distress stabilized | 24
new-onset microcytic anemia | 24
thrombocytosis | 24
elevated ferritin | 24
low albumin | 24
diagnosed with incomplete Kawasaki disease | 24
incomplete Kawasaki disease | 24
Kawasaki disease shock syndrome | 24
treated with ursodiol | 24
treated with intravenous immunoglobulin | 24
treated with aspirin | 24
improved | 96
discharged from the hospital | 96
scleral icterus | 96
direct bilirubin remained elevated | 96
discharged on low-dose aspirin | 96
discharged on ursodiol | 96
follow-up | 240
minimal residual peeling of his palms and soles | 240
bilirubin normalized | 240
echocardiogram demonstrated grossly normal coronary arteries | 240
previous abnormalities were no longer appreciated | 240