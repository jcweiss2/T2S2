40 years old | 0
female | 0
admitted to the emergency room | 0
diffuse abdominal pain | 0
tested positive for pregnancy | -192
vaginal spotting | -96
incomplete abortion | -96
D&C | -96
discharged | -96
symptoms persisted | -72
nausea | -72
non-bilious vomiting | -72
abdominal distention | -72
sought medical attention | -72
abdominal distention | -72
rigidity | -72
diffuse tenderness | -72
guarding | -72
severe and stabbing pain | -72
paraumbilical region | -72
uterine perforation suspected | -72
computed tomography scan | -72
rim-enhancing collection | -72
multiple collections | -72
pneumoperitoneum | -72
small bowel perforation suspected | -72
conservative treatment | -72
nothing by mouth | -72
broad-spectrum antibiotics | -72
prophylactic proton-pump inhibitor | -72
mild tachycardia | -72
pigtail catheter inserted | -48
purulent fluid drained | -48
follow-up CT scan | -24
mural defect in duodenum | -24
extravasation of oral contrast | -24
perforated stress ulcer | -24
surgical exploration | 0
repair with omental patch | 0
mild shortness of breath | -72
COVID-19 antigen test negative | -72
RT-PCR test positive | -24
respiratory team consulted | -24
COVID-19 management plan | -24
respiratory condition deteriorated | 72
vigorous treatment plan | 72
improved | 120
residual mild tachycardia | 120
residual tachypnea | 120
deteriorated again | 144
cardiac arrest | 144
died | 144