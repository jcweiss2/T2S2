29 years old | 0
male | 0
admitted to emergency department | 0
severe headaches | 0
confusion | 0
visual disorders | 0
history of deafness | -100000
deafness from childhood | -100000
temporospatial disorientation | 0
ophthalmologic examination | 0
fundoscopic examination | 24
retinal fluorescein angiography | 24
diagnosis of hearing loss | -100000
otolaryngologist opinion | 24
bilateral sensorineural deafness | -100000
cerebrospinal fluid analysis | 24
elevated protein level | 24
lymphocytic pleocytosis | 24
normal glucose level | 24
negative screening of oligoclonal bands | 24
normal laboratory tests | 24
blood screening for infections | 24
blood screening for common vasculitis | 24
angio-computed tomography | 24
normal angio-computed tomography | 24
brain MRI | 24
multiple small lesions | 24
central lesions in corpus callosum | 24
periventricular lesions in hemispheres | 24
lesions in deep gray nuclei | 24
lesions in midbrain | 24
high-signal abnormalities on T2 | 24
high-signal abnormalities on FLAIR | 24
no restriction on diffusion-weighted imaging | 24
no enhancement on T1 post-contrast sequences | 24
Susac syndrome diagnosis | 24
neurological status worsened | 48
second MRI | 72
extensive lesions | 72
corticosteroid therapy | 72
intravenous methylprednisolone | 72
pulse of intravenous immunoglobulin | 72
unconscious | 96
respiratory distress | 96
transfer to intensive care | 96
intubated | 96
sepsis | 120
death | 672
encephalopathy | 0
sensorineural hearing loss | -100000
branch retinal artery occlusions | 0
magnetic resonance imaging features | 24
involvement of corpus callosum | 24
characteristic imaging keys | 24
accurate diagnosis | 24
differential diagnosis | 24
therapy in severe cases | 72
fatal course | 672
inflammatory disorder of CNS | 0
characteristic clinical triad | 0
radiological findings | 24
brain MRI | 24
callosal lesions | 24
differential diagnoses | 24
evolution | 672
aggressive therapy | 672