56 years old | 0
male | 0
diagnosed as pancreatic cancer | -672
multiple liver metastases | -672
received chemotherapy | -672
chemotherapy was not effective | -672
stent insertion | -336
biliary tract obstruction | -336
febrile sense | -336
chills | -336
antipyretics | -336
analgesics | -336
admitted to nursing care hospital | -168
visited emergency room | -168
complaining of unresolved fever | -168
complaining of chill | -168
complaining of abdominal pain | -168
diabetes mellitus | 0
vidagliptin/metformin | 0
blood pressure 100/60 mmHg | 0
decreased to 90/60 mmHg | 1
respiratory rate 20 breaths per minute | 0
pulse rate 90 beats per minute | 0
body temperature 38.8°C | 0
white blood cell count 1,250/mm3 | 0
neutrophils 92.5% | 0
lymphocytes 4.0% | 0
hemoglobin 5.9 g/dL | 0
platelet count 14,000/mm3 | 0
C-reactive protein 19.75 mg/dL | 0
aspartate aminotransferase 274 UI/L | 0
alanine aminotransferase 143 IU/L | 0
total/direct bilirubin 4.11/2.71 mg/dL | 0
total protein 4.4 g/dL | 0
albumin 2.0 g/dL | 0
prothrombin time 25.3 second | 0
active partial thromboplastin time 60.7 second | 0
blood urea nitrogen 34.5 mg/dL | 0
creatinine 1.9 mg/dL | 0
arterial blood gas analysis | 0
pH 7.515 | 0
pCO2 31.6 mmHg | 0
pO2 78.8.0 mmHg | 0
HCO3 25.5 mmol/L | 0
O2 saturation 96.9% | 0
abdomen computed tomography | 0
pancreatic cancer | 0
multiple liver metastases | 0
metallic stent | 0
acute cholangitis | 0
septic shock | 0
intravenous piperacillin/tazobactam | 0
teicoplanin | 0
norepinephrine | 0
packed red cells | 0
platelets | 0
admitted to intensive care unit | 8
APACHE II score 19 | 8
predicted death rate 32.2% | 8
WBC count deteriorated | 48
platelet count deteriorated | 48
died of refractory septic shock | 120
carbapenem-resistant K. pneumoniae | 120
antimicrobial susceptibility testing | 120
resistance to all beta-lactams | 120
resistance to carbapenems | 120
resistance to tigecycline | 120
MCR1 possessing ST307/Tn4401a[blaKPC2] K. pneumonia | 120
multilocus sequence typing | 120
isotyping the Tn4401 | 120
PCR | 120
agarose gel electrophoresis | 120
antimicrobial susceptibility testing for carbapenems | 120
antimicrobial susceptibility testing for tigecycline | 120
antimicrobial susceptibility testing for colistin | 120
amikacin | 120
gentamicin | 120
amoxicillin/Clavulanic acid | 120
ampicillin | 120
aztreonam | 120
cefazolin | 120
cefepime | 120
cefoxitin | 120
ceftazidime | 120
ciprofloxacin | 120
cotrimoxazole | 120
piperacillin/tazobactam | 120
ertapenem | 120
imipenem | 120
meropenem | 120
doripenem | 120
tigecycline | 120
colistin | 120
minimum inhibitory concentrations | 120
broth microdilution method | 120
Korea-Centers for Disease Control and Prevention | 120
MCR1 gene | 120
E. coli | 120
K. pneumoniae | 120
plasmid-mediated colistin resistance | 120
community-onset infections | 120
inter-regional spread | 120
inter-facility spread | 120
contact precaution | 120
ICU | 120
APACHE II score | 8
predicted death rate | 8
inappropriate antimicrobial treatment | 120
mortality | 120
KPC-KP bacteremia | 120
screening | 120
detection | 120
preemptive isolation | 120
outbreak | 120
inter-facility communications | 120
nationwide epidemiologic data | 120
prompt identification | 120
species | 120
antimicrobial susceptibilities | 120
successful treatment | 120