61 years old | 0
male | 0
hypertension | 0
obesity | 0
hyperlipidemia | 0
emergency department presentation | 0
COVID-19 pandemic onset | 0
progressive shortness of breath | -336
cough | -336
generalized fatigue | -336
muscle aches | -336
denied chest pain | 0
denied arm pain | 0
denied jaw pain | 0
denied pressure | 0
denied diabetes mellitus | 0
denied cardiovascular disease | 0
denied chronic lung disease | 0
denied liver disease | 0
denied kidney disease | 0
denied tobacco use | 0
visibly distressed | 0
tachypneic | 0
hypoxic | 0
hypotension | 0
tachycardia | 0
alert | 0
diaphoretic | 0
respiratory distress | 0
weak peripheral pulses | 0
cool extremities | 0
SARS-CoV-2 infection suspected | 0
negative pressure isolation room | 0
sedation | 0
intubation | 0
circulatory support | 0
norepinephrine | 0
vasopressin | 0
dobutamine | 0
sepsis workup | 0
septic shock workup | 0
positive SARS-CoV-2 | 0
negative other respiratory pathogens | 0
elevated D-dimer | 0
elevated cardiac troponin I | 0
elevated WBC | 0
normal platelet | 0
normal hemoglobin | 0
normal creatinine | 0
elevated INR | 0
elevated CRP | 0
elevated LDH | 0
elevated IL-6 | 0
elevated ferritin | 0
normal CK | 0
new diffuse bilateral airspace opacities | 0
pulmonary infection | 0
PE suspected | 0
heparin infusion | 0
transthoracic echocardiography | 0
normal right ventricle size | 0
normal systolic pressure | 0
mildly elevated pulmonary arterial pressure | 0
moderate global hypokinesis | 0
reduced LV systolic function | 0
EF 30-35% | 0
previous echocardiography EF 62% | -2928
ECG ST elevation | 0
anterolateral leads | 0
leads I | 0
leads II | 0
leads V2-V6 | 0
ischemic changes | 0
STEMI suspected | 0
acute coronary syndrome treatment | 0
dual antiplatelet therapy | 0
aspirin | 0
ticagrelor | 0
coronary angiography deferred | 0
myocarditis suspected | 0
thrombolytics not advised | 0
new ST elevation in lead aVF | 24
worsening ST elevation in lead II | 24
worsening ST elevation in anterolateral leads | 24
ventricular tachycardia episodes | 24
emergent LHC | 48
coronary angiography | 48
patent coronaries | 48
no epicardial stenosis | 48
no thrombosis | 48
no delayed coronary filling | 48
left ventriculography | 48
diffuse hypokinesis | 48
EF 409-45% | 48
LV end-diastolic pressure 22 mm Hg | 48
Takotsubo cardiomyopathy excluded | 48
epicardial coronary thrombosis excluded | 48
STEMI excluded | 48
SARS-CoV-2-induced fulminant myocarditis suspected | 48
steroid therapy | 72
cardiac arrest | 96
failed resuscitation | 96
expired | 96
autopsy patent coronaries | 96
no acute myocardial infarct | 96
scattered focal ischemic changes | 96
hypereosinophilic myocytes | 96
nuclear degeneration | 96
no neutrophil infiltrates | 96
no myocarditis | 96
no pericarditis | 96
interstitial edema | 96
increased macrophages | 96
left atrial thrombus | 96
left pulmonary artery thromboembolism | 96
pulmonary vascular microthrombi | 96
pulmonary consolidation | 96
hemorrhage | 96
early hyaline membrane formation | 96
