44 years old | 0
    female | 0
    admitted to the hospital | 0
    hoarseness | -4320
    occasional loss of voice | -4320
    progressively worsening reduction in effort tolerance | -4320
    shortness of breath | -4320
    unintentional weight loss | -1440
    loss of appetite | -1440
    frequent laryngeal irritation | -1440
    globus sensation in the throat | -1440
    recurrent non-productive cough | -1440
    occasional choking | -1440
    coughing on swallowing liquids | -1440
    denied dysphagia | 0
    denied odynophagia | 0
    breathing difficulties | -2880
    noisy breathing | -2880
    treated for bronchial asthma | -2880
    repeat symptoms two weeks later | -2160
    readmitted | -2160
    intensive care unit admission | -2160
    acute exacerbation of bronchial asthma | -2160
    otolaryngology consult obtained | -2160
    referred to UKM Medical Centre | -2160
    apyrexial | 0
    hemodynamically stable | 0
    biphasic stridor at rest | 0
    able to count up to 10 in a single breath | 0
    no respiratory distress | 0
    cardiopulmonary assessment unremarkable | 0
    bulky right false cord | 0
    limited mobility of right vocal cord | 0
    severe bilateral subcordal edema | 0
    nasal and oral cavities normal | 0
    VHI-10 score 24/40 | 0
    EAT-10 score 20/40 | 0
    microcytic hypochromic anemia | 0
    hemoglobin 9.0 g/dl | 0
    immunological screening negative | 0
    chest x-ray unremarkable | 0
    MRI neck thickening | 0
    endolaryngeal microsurgery | 0
    firm mass right ventricle | 0
    carbon dioxide laser ablation | 0
    dilation to 30 French Bougie | 0
    worsening inspiratory stridor | 6
    tachypnea | 6
    emergency tracheostomy | 6
    neoplastic cells infiltrating muscle fibers | 0
    immunohistochemical reactivity | 0
    bone marrow biopsy confirmed AML | 0
    chemotherapy with HiDAC protocol | 0
    mass not visualized after chemotherapy | 0
    neutropenic sepsis | 0
    invasive pulmonary aspergillosis | 0
    refractory AML | 0
    passed away | +24
    