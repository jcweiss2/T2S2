34 years old | 0
male | 0
admitted to the emergency department | 0
cough with expectoration | -720
breathlessness | -240
right-sided chest pain | -720
loss of weight | -720
loss of appetite | -720
pulse rate of 110/min | 0
blood pressure of 120/80mmhg | 0
respiratory rate of 28/min | 0
oxygen saturation of 90% in room air | 0
absent right-sided air entry | 0
crepitation in the left lung mammary area | 0
point-of-care ultrasound (POCUS) of the Right lung | 0
hydro point | 0
defective barcode sign | 0
oxygen support | 0
symptomatically better | 0
chest X-ray | 1
hydropneumothorax confirmed | 1
low-flow oxygen | 1
empirical antibiotics | 1
right intercostal drainage tube | 1
transferred to the intensive care unit | 1
antitubercular drugs | 1
targeted antibiotics | 1
sputum acid-fast bacilli smear | 1
pleural fluid culture | 1
severe sepsis | 24
died | 24
written informed consent from the patient's wife | 0 
tuberculosis | -720 
necrotizing pneumonia | -720 
malignancy | -720 
pleural fistula | -720 
iatrogenic causes | -720 
connective tissue disorders | -720 
cystic lung disease | -720 
diaphragmatic eventration | -720 
diaphragmatic hernia | -720 
giant bronchogenic cyst | -720 
pneumothorax | 0 
pleural effusion | 0 
hydrothorax | 0 
pyopneumothorax | 0 
hemopneumothorax | 0 
dynamic air–fluid interface sign | 0 
sonographic hydro point | 0 
radiographic hydro point | 0 
barcode sign | 0 
hydro point - effusion sign | 0 
defective barcode sign | 0 
M-mode | 0 
respirophasic motion of hydro point | 0 
sequential assessment of pneumothorax | 0 
pleural effusion assessment | 0 
interface assessment | 0 
bedside POCUS | 0 
chest X-rays | 1 
mobilizing the patient | 1 
validation research studies | 24 
conceptualization | -720 
resources | -720 
visualization | -720 
writing-original draft | -720 
writing - reviewing and editing | -720 
conflicts of interest | 0 
declaration of patient consent | 0 
funding | 0 
images | 0 
clinical information | 0 
patient's name | 0 
patient's initials | 0 
anonymity | 0 
guarantee | 0 
patient's wife | 0 
consent form | 0 
journal | 0 
publication | 0 
identity | 0 
efforts | 0 
conceal | 0