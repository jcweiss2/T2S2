63 years old | 0
    male | 0
    peripheral vascular disease (PVD) | 0
    claudication | 0
    hypertension | 0
    diabetes mellitus type-2 | 0
    chronic low back pain | 0
    presented to the emergency room | 0
    dyspepsia | 0
    three days of melanic stools | -72
    taking 800 mg ibuprofen three times daily | -17520
    sinus tachycardia (115 bpm) | 0
    hypotension (90/60 mm Hg) | 0
    left lower extremity weakness | 0
    pallor | 0
    pulselessness | 0
    diffuse skin pallor | 0
    severe anemia (hemoglobin/hematocrit 8.1 gL/dL/22.5 L%) | 0
    leukocytosis (white blood cell = 21,000 Hk/cmm) | 0
    lactic acidosis (lactic acid = 6.2 mmol/L) | 0
    acute renal failure (urea nitrogen/creatinine = 53 mg/dl/1.6 mg/dl) | 0
    hyponatremia (sodium = 124 mmol/L) | 0
    hypokalemia (potassium = 3.1 mmol/L) | 0
    positive occult blood | 0
    positive blood cultures (methicillin sensitive Staphylococcus aureus) | 0
    no coagulopathy | 0
    no thrombocytopenia | 0
    chest radiograph unremarkable | 0
    electrocardiogram (ECG) sinus tachycardia | 0
    computed tomography (CT) abdomen and pelvis with intravenous contrast | 0
    no retroperitoneal hematoma | 0
    no bowel perforation | 0
    admitted to MICU | 0
    standard management for upper GI bleeding | 0
    resuscitation for acute renal failure | 0
    pantoprazole continuous infusion | 0
    packed red blood cells | 0
    crystalloid | 0
    gastroenterology consultation | 0
    bacteremia | 0
    vancomycin | 0
    piperacillin/tazobactam | 0
    ischemic left lower extremity | 0
    vascular surgery consultation | 0
    CT angiogram left lower extremity | 0
    good distal runoff | 0
    opacification to ankle | 0
    downward trending hemoglobin/hematocrit | 0
    worsening lactic acidosis | 0
    emergent EGD | 0
    bleeding duodenal ulcers | 0
    largest ulcer 30 mm x 30 mm | 0
    ulcers cauterized | 0
    epinephrine injection for hemostasis | 0
    tolerated procedure well | 0
    no new complaints post-procedure | 0
    eight hours post-procedure worsening abdominal pain | 8
    abdominal distension | 8
    diaphoresis | 8
    tachypnea | 8
    temperature 95.0 F | 8
    blood pressure 143/83 | 8
    heart rate 142 | 8
    respiratory rate 48 | 8
    oxygen saturation 92% on non-rebreather mask | 8
    diffuse abdominal guarding | 8
    rebound tenderness | 8
    abdominal distension | 8
    mixed respiratory and metabolic acidosis (ABG 7.05/60.4/72.6/16.5) | 8
    STAT abdominal radiograph | 8
    pneumo-peritoneum | 8
    chest radiograph | 8
    free air under diaphragm | 8
    emergently intubated | 8
    general surgery consultation | 8
    CT abdomen and pelvis with oral contrast | 8
    confirmed pneumo-peritoneum | 8
    duodenal perforation | 8
    unclear cause of perforation | 8
    smaller size of perforation | 8
    hypotensive | 8
    norepinephrine infusion | 8
    vasopressin infusion | 8
    hemodynamic instability | 8
    multiple comorbidities | 8
    general surgery recommended non-operative management | 8
    strict bowel rest | 8
    intravenous antibiotics | 8
    intravenous fluconazole | 8
    intubated | 8
    six days intubated | 8
    renal function worsened | 8
    urine output worsened | 8
    acute tubular necrosis | 8
    septic shock | 8
    compartment syndrome | 8
    bladder pressure >15 mm Hg | 8
    oxygen requirements improved | 8
    vasopressor requirements improved | 8
    extubation hospital day 7 | 168
    metabolic derangements | 168
    worsening renal function | 168
    severe tachypnea | 168
    reintubated | 180
    acute renal failure | 180
    oliguria | 180
    hemodialysis initiated hospital day 8 | 192
    intubated | 192
    intermittent hemodialysis | 192
    broad spectrum antibiotics | 192
    micafungin | 192
    stable condition | 192
    off vasopressors | 192
    left lower extremity cold | 192
    pulselessness | 192
    concern for necrosis | 192
    vascular surgery recommended against intervention | 192
    self-extubated hospital day 15 | 360
    requested no re-intubation | 360
    no aggressive measures | 360
    compartment syndrome | 360
    bladder pressure 15-19 mm Hg | 360
    pain management priority | 360
    palliative care approach | 360
    expired hospital day 19 | 456
