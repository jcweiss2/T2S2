49 years old | 0
female | 0
admitted to the hospital | 0
low back pain | -504
intractable cough | -504
productive of green sputum | -504
no chest pain | -504
no shortness of breath | -504
no fevers | -504
no paraesthesia | -504
no weakness of the lower limbs | -504
no urinary symptoms | -504
no bowel symptoms | -504
completed a course of oral cephalexin | -504
hypertension | -504
chronic low-back pain | -504
smoked 20 cigarettes per day | -504
15 pack year smoking history | -504
no respiratory distress | 0
normal vital signs | 0
bronchial breath sounds in the right lung mid to lower zones | 0
coarse crepitations | 0
soft and non-tender abdomen | 0
antalgic gait | 0
normal sensation, power and reflexes in the lower limbs | 0
white cells 19.2 × 10^9/L | 0
neutrophilia | 0
chest radiograph demonstrated an obscured right heart border | 0
community acquired pneumonia of the right middle lobe | 0
cough precipitated the low back pain | 0
commenced on benzyl penicillin | 0
commenced on doxycycline | 0
commenced on analgesics | 0
admitted under the medical team | 0
medical emergency team review | 24
hypotension | 24
presyncope | 24
new onset epigastric/chest pain | 24
back pain | 24
pale | 24
heart rate 78 bpm | 24
blood pressure 66/38 mmHg | 24
unchanged chest examination | 24
soft abdomen | 24
haemoglobin dropped from 115 g/L to 77 g/L | 24
in shock | 24
likely haemorrhagic | 24
aortic dissection suspected | 24
rupture of an aortic aneurysm suspected | 24
haemorrhage from a peptic ulcer suspected | 24
sepsis secondary to pneumonia suspected | 24
obstructive shock secondary to pulmonary embolism suspected | 24
bilateral large bore intravenous access obtained | 24
fluid resuscitation commenced | 24
transfusion of red blood cells | 24
given intravenous ceftriaxone | 24
moved to the high dependency unit | 24
surgical review obtained | 24
haemodynamically responsive to resuscitation | 24
urgent computed tomography scan with contrast of her chest and abdomen | 24
ruptured spleen | 24
large perisplenic haematoma | 24
large haemoperitoneum | 24
active bleeding in portal venous sequences | 24
bilateral pulmonary consolidation | 24
no pulmonary embolism | 24
taken to the operating theatre for an emergency laparotomy | 24
vertical midline upper abdominal laparotomy | 24
large haematoma removed | 24
ongoing bleeding | 24
spleen nearly avulsed | 24
splenophrenic ligament incomplete | 24
partial rupture of the spleen under the ligament | 24
splenonephric ligament absent or avulsed | 24
mobile spleen with medial lie | 24
Ligasure division of the short gastric and splenic arteries and veins | 24
spleen removed | 24
satisfactory haemostasis | 24
splenic artery oversewn | 24
Blake’s drain placed in the left subdiaphragmatic space | 24
abdomen closed | 24
transfusion of six units of red blood cells | 24
transfusion of two units of fresh frozen plasma | 24
transfer to the nearest intensive care unit | 48
successfully extubated | 48
discharged home | 96
investigations for pneumonia did not reveal a causative organism | 96
negative findings for influenza A and B | 96
negative findings for RSV direct antigen tests | 96
negative findings for respiratory virus PCR | 96
negative findings for sputum microscopy and culture | 96
negative findings for urinary antigen testing for legionella and pneumococcus | 96
negative findings for serologic testing for chlamydia, EBV and legionella | 96
histopathology revealed a 95 g spleen | 96
spleen measuring 65 × 60 × 30 mm | 96
25 mm defect consistent with possible site of rupture | 96
pulp architecture preserved | 96
no evidence of malignancy | 96
uncomplicated recovery | 168
pneumonia resolved | 168
surgical wounds healing well | 168
resumed nearly all activities | 168
persisting back pain | 168
immunised against Pneumococcus | 168
immunised against Meningococcus | 168
immunised against Haemophilus influenza type b | 168
declined the trivalent influenza vaccine | 168
commenced on prophylactic amoxicillin | 168
added to the splenectomy register | 168