26 years old | 0
female | 0
twin pregnancy | 0
36 weeks and one day gestation | 0
gravida 1 | 0
0 abortions | 0
admitted to the hospital | 0
malaise | -144
fever | -144
non-productive cough | -144
febrile | 0
tachycardic | 0
hypoxic | 0
O2 saturation of 92% | 0
diffuse rhonchi on auscultation | 0
increased erythrocyte sedimentation rate | 0
non-stress-test reactive for both fetuses | 0
biophysical profiles were 6/8 | 0
decreased fetal movement | 0
multifocal sub-pleural patchy consolidative opacities on both lung fields | 0
COVID-19 pneumonia | 0
cesarean section | 0
both infants in good condition | 0
first minute APGAR score of 9/10 | 0
isolated from their mother | 0
transferred to the Neonatal Intensive Care Unit | 0
COVID-19 infection confirmed in the mother | 0
RT-PCR positive | 0
nasopharynx specimens negative in both infants | 0
asymptomatic at the two-week follow-up | 336
Meropenem started | 0
azithromycin started | 0
hydroxychloroquine started | 0
supplemental oxygen started | 0
lack of favorable response to treatment | 144
plasma transfusion | 144
Favipiravir added | 144
clinical course improved | 168
second CT scan performed | 288
very faint residual ground-glass opacities | 288
dramatic response to therapy | 288
discharged | 336
COVID-19 with pulmonary involvement | 0 
Favipiravir treatment | 144
convalescent plasma therapy | 144 
no COVID-19 symptoms in newborns | 336
negative PCR results in newborns | 336