64 years old | 0
woman | 0
brought to the emergency room | 0
unresponsive | 0
found slumped on the couch | 0
eyes open but speechless | 0
unable to follow commands | 0
no injury | 0
no incontinence | 0
no other signs of seizure | 0
stroke code activated | 0
lethargic | 0
lack of interest in environment | 0
slow responses to stimulation | 0
tendency to fall asleep | 0
blood pressure 131/91 mm Hg | 0
pulse rate 78 beats/min | 0
respiratory rate 15 breaths/min | 0
oxygen saturation 99.8% | 0
afebrile (37.1 °C) | 0
no signs of meningeal irritation | 0
pupils 4 mm and equally reactive to light | 0
no evidence of ophthalmoplegia | 0
no facial asymmetry | 0
no other cranial nerve deficits | 0
moved all extremities spontaneously | 0
reflexes 1+ | 0
no ankle clonus | 0
Babinski sign absent | 0
past history of atrial fibrillation | -35040
past history of right frontal ischemic stroke | -35040
no history of seizures/epilepsy | -35040
survived cardiac arrest 4 years prior | -35040
pacemaker/defibrillator implanted | -35040
computed tomography (CT) head showed encephalomalacia in right frontal lobe | 0
electrocardiogram showed regular atrial-sensed ventricular-paced rhythm | 0
nonconvulsive seizures/status epilepticus ruled out by stat EEG | 0
blood counts normal | 0
blood chemistry normal | 0
chest X-ray normal | 0
no clear evidence of new stroke | 0
tissue plasminogen activator not administered | 0
became stuporous (GCS = 10) | 12
intubated for airway protection | 12
admitted to intensive care unit | 12
magnetic resonance imaging not performed due to pacemaker | 12
repeat head CT 12 hours later revealed bilateral paramedian thalamic infarcts | 12
CT angiography showed filling defects at top of basilar artery and P1 segments | 12
possibility of occluded artery of Percheron could not be ruled out | 12
telemetry showed regular ventricular-paced rhythm | 12
pulse oximetry oxygen saturations ≥99.0% | 12
transthoracic echocardiography with bubble study unrevealing | 12
transesophageal echocardiography attempted but aborted | 12
clopidogrel added to aspirin | 12
intravenous levetiracetam administered | 12
cEEG over 48 hours showed diffuse slowing | 12
no signs of abnormal cortical hyperexcitability | 12
methylphenidate started on day 3 | 72
became more alert | 72
started following simple commands | 72
extubation attempted on day 6 | 144
extubation failed due to upper airway edema | 144
tracheostomy performed | 216
percutaneous endoscopic gastrostomy performed | 216
patient lapsed into stupor again (GCS = 9) on day 12 | 288
blood pressure 144/95 mm Hg | 288
pulse rate 72 beats/min | 288
respiratory rate 18 breaths/min | 288
oxygen saturation 99.1% | 288
telemetry showed normal rate and rhythm | 288
blood test results normal | 288
change in mental status not due to toxic, metabolic, or septic encephalopathy | 288
husband noticed 30-second episode of bilateral leg jerking | 288.5
EEG recording showed sustained generalized epileptiform discharges | 289.33
Salzburg criteria for NCSE satisfied | 289.33
initially awake and motionless | 289.33
extremities started jerking (rhythmic pronation-supination of forearms) | 289.33
rhythmic hip and knee flexion-extension | 289.33
clonic/convulsive seizure lasting 28 seconds | 289.33
EEG obscured by muscle artifact | 289.33
lorazepam 2 mg injected | 289.33
attenuation and dissipation of epileptiform discharges | 289.33
stupor attributed to NCSE | 289.33
midbrain infarction concern | 289.33
family decided against further invasive interventions | 289.33
signs of right third nerve palsy (ptosis and dilated nonreactive pupil) | 291
stat CT head showed same infarct in paramedian thalami | 291
repeat CT head 22 hours after onset of stupor showed midbrain infarct | 312
cEEG showed waxing-waning generalized epileptiform discharges | 312
relapsing and remitting cortical hyperexcitability or NCSE | 312
cEEG periods of generalized slowing without epileptiform discharges | 312
build-up of rhythmic delta activity | 312
increasing density of sharp waves | 312
evolution toward organized 1.5 to 2.5 Hz high-voltage sharp and slow wave complexes | 312
epileptiform discharges persist for hours | 312
patient more somnolent during high-voltage rhythmic discharges | 312
husband witnessed 2 more episodes of bilateral leg jerking | 312
last episode recorded with no EEG change | 312
increasing dose of levetiracetam | 312
phenytoin added | 312
intermittent boluses of lorazepam | 312
temporary suppression of NCSE | 312
NCSE reemerged | 312
generalized rhythmic delta activity | 312
gain in "ictal" features | 312
cEEG omitted for 5 days | 312
patient in and out of NCSE over 3 weeks | 504
family refused induction of coma with anesthesia | 504
sodium valproate added | 504
suppression of epileptiform activity | 504
became more alert and responsive | 504
remained nonverbal | 504
followed simple commands | 504
discharged on hospital day 33 | 792
