55 years old | 0
    female | 0
    admitted to the hospital | 0
    abdominal distension | -336
    ovarian cancer | -9600
    hysterectomy | -9600
    bilateral salpingo-oophorectomy | -9600
    five cycles of chemotherapy | -9600
    normochromic normocytic anemia | 0
    healthy liver function | 0
    healthy kidney function | 0
    normal clotting limits | 0
    significant ascites | 0
    moderate right pleural effusion | 0
    pelvic mass at the distal ileum | 0
    normal liver parenchyma | 0
    DLBCL (diffuse large B-cell lymphoma) | 0
    pleural effusion drained | 0
    ascites drained | 0
    persistent tachycardia | 168
    respiratory failure | 168
    intubation | 168
    ventilation | 168
    metabolic acidosis | 168
    respiratory compensation | 168
    pH 7.29 | 168
    CO2 29mmHg | 168
    pO2 77mmHg | 168
    BE -11.7 | 168
    HCO3-13mmol/L | 168
    lactate 5.7mmol/L | 168
    anion gap 18 | 168
    pneumoperitoneum | 168
    left lower zone lung consolidation | 168
    exploratory laparotomy | 168
    septic shock | 168
    perforated gut | 168
    drowsy | 168
    tachycardic (170 bpm) | 168
    hypotensive (82/50 mmHg) | 168
    fluid boluses | 168
    blood pressure increased to 90/60 mmHg | 168
    noradrenaline infusion | 168
    mean arterial pressure 65mmHg | 168
    pelvic lymphoma | 168
    perforated distal ileum | 168
    feculent peritonitis | 168
    bowel resection | 168
    temporary abdominal closure | 168
    broad-spectrum antibiotics (vancomycin, caspofungin, meropenem) | 168
    hospital-acquired pneumonia | 168
    fentanyl infusion | 168
    noradrenaline weaned off | 192
    mean arterial pressure >65mmHg | 192
    urine output 0.5-1ml/kg/hr | 192
    PlasmaLyte infusion | 192
    20% human albumin solution | 192
    positive fluid balance | 192
    tachycardia persisted | 192
    lactic acidosis persisted | 192
    left shift neutrophilia | 192
    normal liver function | 192
    normal renal function | 192
    respiratory failure resolved | 240
    hyperlactatemia plateaued | 240
    Type A LA contributory | 240
    Type B LA from intra-abdominal sepsis | 240
    Klebsiella pneumoniae isolated | 240
    Candida tropicalis isolated | 240
    meropenem changed to ceftazidime-avibactam | 240
    respiratory wean attempted | 240
    tachypnea (351-45 bpm) | 240
    pain excluded | 240
    pulmonary embolism excluded | 240
    hypoxia excluded | 240
    medications reviewed | 240
    vancomycin continued | 240
    caspofungin continued | 240
    ceftazidime-avibactam continued | 240
    fentanyl continued | 240
    second laparotomy | 264
    bowel ischemia ruled out | 264
    loculated collections ruled out | 264
    intra-abdominal pressure normal (12mmHg) | 264
    double barrel stoma created | 264
    permanent abdominal closure | 264
    daily blood investigations | 264
    biomarkers downward trend | 264
    serum LDH elevated (1002 units/L) | 264
    DLBCL activity high | 264
    CRRT (continuous renal replacement therapy) | 264
    cyclophosphamide started | 264
    rituximab started | 264
    etoposide started | 264
    Type B LA resolved | 336
    extubated | 336
    transferred out of ICU | 336
    succumbed to DLBCL | 3024
    <|eot_id|>
    