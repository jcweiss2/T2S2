60 years old | 0
male | 0
gastroesophageal reflux disease | 0
5-month history of gradually worsening symptoms | -3600
diffuse joint pain | -3600
joint swelling | -3600
diffuse rash | -3600
headaches | -3600
generalized weakness | -3600
subjective fevers | -3600
chills | -3600
profuse night sweats | -3600
unintentional 30-pound weight loss | -3600
pruritic rash | -3600
rash started on face | -3600
rash spread throughout body | -3600
headaches with bilateral eye pain | -3600
eye swelling | -3600
double vision | -3600
mild vision blurriness | -3600
muscle weakness | -3600
lower extremity weakness | -3600
bilateral weakness | -3600
hip flexion and extension weakness (3/5) | -3600
knee flexion and extension weakness (4-/5) | -3600
ankle dorsiflexion and plantarflexion weakness (4-/5) | -3600
dysphagia for solids and liquids | -3600
febrile | 0
mildly toxic appearance | 0
diffuse alopecia | 0
adjacent scarring | 0
polymorphous rash on face, back, and extremities | 0
hypopigmentation | 0
hyperpigmentation | 0
eczematous-like macules and patches on extremities and hips | 0
edematous and tender joints (hands, elbows, shoulders) | 0
symmetrical facial weakness | 0
decreased facial sensation in cranial nerve V2 and V3 distribution | 0
proximal and distal muscle weakness | 0
decreased muscle bulk | 0
increased muscle tone | 0
bilateral positive Babinski reflex | 0
hyperreflexive joint reflexes | 0
normocytic anemia | 0
thrombocytopenia | 0
elevated liver enzymes | 0
normochromic anemia | 0
mild leukopenia | 0
erythrocyte sedimentation rate elevated (55 mm/hr) | 0
C-reactive protein elevated (1.4 mg/dL) | 0
lactate dehydrogenase elevated (373 U/L) | 0
aspartate transaminase elevated (278 U/L) | 0
alanine transaminase elevated (105 U/L) | 0
mild muscle pain in proximal lower extremities | 24
subcutaneous edema | 24
myositis in anterior compartment muscles of left thigh | 24
focal myopathy | 24
denervation atrophy (severe, type II) | 24
seronegative dermatomyositis | 24
high-dose parenteral steroids | 24
immunosuppressive therapy with hydroxychloroquine | 24
transferred to medical intensive care unit | 840
worsening respiratory distress | 840
severe sepsis | 840
intubated | 864
questionable intraperitoneal air on imaging | 864
ejection fraction of 65% | 888
oliguria | 912
acute kidney injury | 912
patient expired | 1008
final muscle biopsy showed gelsolin amyloidosis | 1056
gingival mucosal biopsy showed amyloid deposition | 1056
homozygous missense mutation C>G1375 in exon 10 | 1056
proline 459 to arginine in gelsolin domain 4 | 1056
wild-type exon 4 sequence | 1056
