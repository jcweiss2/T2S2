50 years old | 0
female | 0
admitted to the hospital | 0
altered mental status | 0
acute alcohol intoxication | 0
binge drinking | -12
wine consumption | -12
normal vital signs except for low blood pressure | 0
drowsy | 0
arousable | 0
partially oriented | 0
blood alcohol level of 353 mg/dl | 0
anion gap of 17 | 0
lactate of 4.5 mmol/L | 0
beta hydroxybutyrate of 0.7 mmol/L | 0
positive urine ketones | 0
serum glucose of 80 mg/dl | 0
serum osmolality of 383 mOsm/kg | 0
normal serum osmolal gap | 0
undetectable levels of methanol | 0
undetectable levels of isopropanol | 0
undetectable levels of acetone | 0
received 7 L of normal saline | 0
hypotension | 0
normalized serum alcohol | 12
normalized anion gap | 12
normalized lactate | 12
normalized serum ketones | 12
normalized mental status | 12
unresponsive | 24
found on the floor of her hospital room | 24
blood pressure of 93/60 mm of Hg | 24
Glasgow Coma Score of 3 | 24
required fluid resuscitation | 24
required intubation | 24
unremarkable CT of the head | 24
increased lactate | 24
increased anion gap | 24
extubated | 48
normalized serum lactate | 48
normalized anion gap | 48
alert and fully oriented | 48
unresponsive again | 72
found next to an open and empty bottle of ethanol based hospital hand sanitizer | 72
normal vital signs | 72
Glasgow Coma Score of 3 | 72
lactate of 3.9 mmol/L | 72
anion gap of 15 | 72
serum ethanol of 362 mg/dl | 72
methanol of 0 mg/dl | 72
acetone of 11 mg/dl | 72
isopropanol of 14 mg/dl | 72
arterial blood gas showed a pH of 7.32 | 72
PaCO2 of 43 mm Hg | 72
PaO2 of 73 mm Hg | 72
bicarbonate of 22 mmol/L | 72
admitted to the intensive care unit | 72
required nasopharyngeal airway | 72
supportive care | 72
normalized mental status | 78
normalized lactate levels | 78
normalized metabolic acidosis | 78
admitted to drinking ethanol based hospital hand sanitizer | 78
denied suicidality | 78
hand sanitizers removed from her room | 78
one-to-one monitoring | 78
discharged to an in-patient alcohol treatment program | 96