62 years old | 0
female | 0
primary progressive multiple sclerosis | -672
altered level of consciousness | -168
hypoxemia | -168
shock | -168
tested positive for severe acute respiratory syndrome coronavirus-2 | -168
admitted to the hospital | 0
initial blood pressure 55/32 mm Hg | 0
heart rate 120 beats/min | 0
respiratory rate 32 breaths/min | 0
oxygen saturation 95% on 100% oxygen | 0
dense airspace opacities in the right lung | 0
ground-glass opacity in the left lung | 0
sinus tachycardia with diffuse anterolateral ST-elevation | 0
high-sensitivity cardiac Troponin T 4986 ng/L | 0
N-terminal pro-B-type natriuretic peptide 51,439 ng/L | 0
ferritin 3067 U/L | 0
C-reactive protein 68.2 mg/L | 0
D-dimer 6920 ng/mL | 0
lactate dehydrogenase 1094 U/L | 0
lactate 2.4 mmol/L | 0
creatinine 252 umol/L | 0
resuscitated with intravenous fluids | 0
received dexamethasone | 0
received ceftriaxone | 0
received azithromycin | 0
no intubation | 0
no inotropes | 0
point-of-care ultrasound demonstrated severe left ventricular dysfunction | 0
lung ultrasound findings consistent with pneumonia | 0
urgent cardiac magnetic resonance imaging | 24
CMR findings consistent with acute myocarditis | 24
global hypokinesia | 24
relative sparing of the basal segments | 24
extensive sub-epicardial LGE in the anterolateral and inferolateral left ventricular walls | 24
elevation in tissue mapping-based markers of inflammatory injury | 24
native T1 and T2 values elevated | 24
expansion of the extracellular volume | 24
left ventricular ejection fraction 24% | 24
anakinra administered | 24
rapid clinical improvement | 48
reduced oxygen requirements | 48
improved blood pressure | 48
reduction in heart rate | 48
renal function improved | 48
progressive reduction in inflammatory markers | 48
anakinra treatment continued for 5 days | 120
repeat CMR imaging | 336
marked improvement in left ventricular ejection fraction | 336
reduction in LGE signal intensity | 336
global reductions in myocardial T1 and T2 values | 336
global reductions in extracellular volume | 336
small pericardial effusion | 336
enhancement of the parietal pericardium | 336
resolution of pulmonary consolidation | 336
resolution of pleural effusions | 336
discharged from the hospital | 360