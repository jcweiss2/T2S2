12 years old | 0
male | 0
Maori | 0
admitted to hospital | 0
acute otitis media | -24
perforation | -24
neck swelling | -24
neck pain | -24
septic shock | 0
endotracheal intubation | 0
computed tomography scan | 0
retropharyngeal phlegmon | 0
obstructive thrombi | 0
internal jugular vein | 0
pulmonary septic emboli | 0
pulmonary lesions | 0
Lemierre’s syndrome | 0
antibiotics started | 0
cefotaxime | 0
metronidazole | 0
flucloxacillin | 0
lincomycin | 0
MSSA | 0
blood cultures positive | 0
high-frequency ventilation | 24
hypoxia | 24
mean airway pressure increased | 24
inspired oxygen fraction | 24
oxygenation index | 24
repeat CT scan | 72
jugular clots | 72
pulmonary emboli | 72
pulmonary cavitating lesions | 72
noradrenaline | 72
adrenaline | 72
vasopressin | 72
ECLS | 72
femoral veno-arterial cannulation | 72
rest ventilation | 72
pressure control ventilation | 72
positive end-expiratory pressure | 72
right-sided pneumothorax | 120
pneumothorax drained | 120
left-sided pneumothorax | 144
hemoserous drain losses | 168
inflammatory markers high | 192
inotropic support | 192
CT imaging | 192
abscess formation | 192
osteomyelitis | 192
opacified left mastoid | 192
abscess drained | 192
open incision | 192
cortical mastoidectomy | 192
heparin stopped | 192
tranexamic acid | 192
bleeding controlled | 192
peri-procedure bleeding | 192
red blood cells transfused | 192
platelet transfused | 192
fibrinogen high | 192
cryoprecipitate not required | 192
concentrated fibrinogen not required | 192
tranexamic acid | 192
thrombelastogram | 192
hyperfibrinolysis | 192
cultures from abscess | 192
MSSA growth | 192
cortical mastoidectomy results | 192
middle ear process | 192
negative pressure vacuum dressing | 192
delayed primary closure | 240
CT imaging | 240
lung abscesses | 240
bronchopleural fistula | 240
abscess drainage deferred | 240
pulmonary gas exchange improved | 240
ECLS weaned | 384
decannulation | 384
magnetic resonance imaging | 384
no further abscesses | 384
invasive mechanical ventilation | 552
non-invasive ventilation | 552
high-flow nasal cannula oxygen | 552
secondary pseudomonal sepsis | 552
critical illness myopathy | 552
CT imaging | 552
pathological fractures | 552
lateral masses of C1 | 552
ICU discharge | 1032
follow-up imaging | 1032
lung fields improved | 1032
cavitations improved | 1032
fluid collections resolved | 1032
thrombi persisted | 1032
jugular veins | 1032
venous sinuses | 1032
intravenous flucloxacillin | 1032
intravenous Bactrim | 1032
oral Bactrim | 1032
oral flucloxacillin | 1032
CNS imaging | 1032
mastoid | 1032
C1 collections | 1032
intracranial abscesses | 1032
inflammatory response | 1032
MRI | 1032
resolution of abnormal findings | 1032
gliosis | 1032
cerebellum | 1032
halo-thoracic jacket | 1032
osteomyelitis | 1032
C1 | 1032
C2 | 1032
fractures | 1032
lateral masses of C1 | 1032
neurocognitive assessment | 1032
motor | 1032
cognitive | 1032
behavioural performance | 1032
normal outcomes | 1032
Pediatric Overall Performance Category Assessment | 1032
good overall performance | 1032
audiological assessment | 1032
mild conductive loss | 1032
left ear | 1032
bilateral sensorineural mid to high frequency loss | 1032
hospital discharge | 1248
halo-thoracic jacket removal | 1248