9 years old | 0
    Afghan girl | 0
    severely injured in a car accident | -4320
    admitted to a teaching hospital in southeast Germany | 0
    surgery at an Indian hospital | -4320
    left leg stabilized with external fixation | -4320
    external fixation substituted by femur nail | -4320
    general condition dramatically deteriorated | 0
    dehydrated | 0
    undernourished | 0
    130 cm height | 0
    25 kg body weight | 0
    decreased serum concentration of total protein | 0
    decreased creatinine | 0
    anemia | 0
    several decubitus dorsal ulcers | 0
    stage 2 ulcers | 0
    stage 3 ulcers | 0
    both legs showed multiple wounds | 0
    extended areas of scab | 0
    secretion of large amounts of yellow pus | 0
    pus secreted from a fistula of left hip joint | 0
    MRSA isolated | 0
    carbapenem resistant Pseudomonas aeruginosa isolated | 0
    Gram negative bacteria with ESBL isolated | 0
    Citrobacter sedlakii isolated | 0
    Escherichia coli isolated | 0
    Proteus mirabilis isolated | 0
    Klebsiella pneumoniae isolated | 0
    methicillin susceptible S. aureus isolated | 0
    non ESBL Proteus mirabilis isolated | 0
    Enterococcus faecalis isolated | 0
    Enterococcus hirae isolated | 0
    Bacteroides fragilis isolated | 0
    peptostreptococci isolated | 0
    bacterial identification performed | 0
    antibiotic susceptibility testing performed | 0
    admitted to pediatric surgery ward | 336
    16 surgeries | 336
    approximately 60 dressing changes | 336
    each requiring general anesthetics | 336
    received cefazoline | 0
    received imipenem | 0
    received meropenem | 0
    received ampicillin | 0
    received clindamycin | 0
    received amoxicillin | 0
    received ceftazidime | 0
    received ceftaroline | 0
    received cefuroxime | 0
    MRSA frequently isolated within first 3 weeks | 168
    two decolonization cycles | 168
    MRSA not found in swabs from nose | 168
    MRSA not found in swabs from throat | 168
    MRSA not found in biopsy specimen | 168
    no further proof of MRSA | 168
    MRSA found in nose swab on March 20, 2014 | 4560
    decolonization measures for seven days | 4560
    MRSA found in biopsy sample on May 16, 2014 | 6000
    MRSA found in swabs from nose | 6000
    MRSA found in swabs from throat | 6000
    amputation of lower legs on June 3, 2014 | 6384
    MRSA detected in biopsy of infected limb | 6384
    treated in intensive care unit for 9 days | 6384
    deterioration in general condition | 6384
    systemic inflammatory response syndrome | 6384
    increased heart rate | 6384
    white blood cell count increased | 6384
    decreased blood pressure | 6384
    body temperature rose to 40.3°C | 6384
    C-reactive protein increased to 265.5 mg/L | 6384
    MRSA found in blood culture | 6384
    septic infection | 6384
    antibiotic treatment with ceftaroline | 6384
    continuous improvement of general condition | 6384
    final revision surgery on June 18, 2014 | 6528
    removal of condylar cartilage | 6528
    debridement of necrotic tissue | 6528
    MRSA detected in biopsy specimen | 6528
    no increase of inflammation parameters | 6528
    circulation not impaired | 6528
    ceftaroline application stopped | 6528
    no further MRSA found | 6528
    discharged from hospital | 8760
    MRSA typing performed | 8760
    informed consent given | 8760
    ethics approval not deemed necessary | 8760
    severe infection of both legs | 0
    presence of MRSA | 0
    sepsis caused by MRSA | 6384
    endogenous MRSA infection | 8760
    screening suggested successful MRSA decolonization | 168
    risk of MRSA recolonization | 8760
    infection treated with ceftaroline | 6384
    increased MIC for MRSA | 8760
    reduced antibiotic susceptibility to ceftaroline | 8760
    increased ceftaroline MICs reported | 8760
    ceftaroline resistance in MRSA | 8760
    diagnostic challenges in susceptibility testing | 8760
    preserved ceftaroline as potent antibiotic | 8760
    speaker’s honorarium from AstraZeneca | 8760
    no other conflicts of interest | 8760