78 years old | 0
male | 0
laparoscopic-assisted total gastrectomy | 0
type II diabetes mellitus | 0
ischemic heart disease | 0
previous myocardial infarction | -105216
occasional ongoing angina | 0
benign prostatic hypertrophy | 0
open cholecystectomy | - (unknown)
general anesthesia | 0
epidural analgesia | 0
adhesions around cholecystectomy site | 0
dense perisplenic capsular adhesions | 0
fatty liver | 0
bulky left lobe of liver | 0
Nathanson retractor insertion | 0
retraction of left liver lobe | 0
reverse Trendelenburg position | 0
laparoscopic mobilization of stomach and omentum | 0
duodenum division | 0
stapling device use | 0
oversewing duodenum | 0
splenic capsular bleeding | 0
conservative techniques attempted | 0
laparoscopic division of splenic vessels | 0
splenectomy | 0
epigastric transverse incision | 0
removal of stomach and spleen | 0
Roux-en-Y esophagojejunostomy | 0
feeding jejunostomy tube | 0
total laparoscopic time 3.5 hours | 210
intensive care unit admission | 0
hypotension | 0
increasing inotropic support | 0
blood pressure stabilization | 24
serum AST elevation at 5 hours postoperation | 5
AST peak >20 times normal | 5
AST gradual decrease over 2 days | (5 to 53)
alkaline phosphatase rise | (unknown)
gamma-glutamyltransferase rise | (unknown)
total bilirubin rise | (unknown)
C-reactive protein rise | (unknown)
jejunostomy feed started | 24
tachycardia | 48
fever 38°C | 48
rapid deterioration over next 6 hours | 48 to 54
large inotrope doses | 54
ventilatory assistance | 54
suspicion of anastomotic dehiscence | 54
urgent noncontrast abdominal CT | 54
CT showing liver destruction | 54
intraparenchymal gas loculations | 54
portal radical gas | 54
exploratory laparotomy | 54
left lateral sectionectomy | 54
inotropic support continued | 54
myocardial infarction | 68
death | 68
