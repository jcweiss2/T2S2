73 years old | 0
female | 0
hypertension | -8760
diabetes mellitus type 2 | -8760
diabetic nephropathy | -8760
chronic renal impairment | -8760
dual pacemaker | -8760
sick sinus syndrome | -8760
ST elevation myocardial infarction | -720
three drug-eluting stents | -720
left main coronary artery | -720
proximal right coronary artery | -720
proximal circumflex artery | -720
PEG | -4320
refusal to eat | -4320
true bulbar palsy | -4320
early signs of Alzheimer's disease | -4320
furosemide | -8760
carvedilol | -8760
spironolactone | -8760
clopidogrel | -8760
admitted to the hospital | 0
hypotension | 0
pulmonary edema | 0
ventilator support | 0
tracheal intubation | 0
inotropes | 0
renal replacement therapy | 0
improvement | 72
extubated | 72
acute on chronic renal failure | 72
restart of renal replacement therapy | 72
severe global hypokinesia of the left ventricle | 0
low ejection fraction | 0
bilateral lung ultrasonic B lines | 0
bilateral mild pleural effusions | 0
low cardiac output | 0
generalized edema | 0
noradrenaline | 0
dobutamine | 0
discontinued | 120
hemodialysis | 165
hypotension | 168
noradrenaline infusion | 168
tachypnea | 168
vague abdominal pain | 168
blood pressure 105/45 mm Hg | 168
heart rate 93 beats/min | 168
abdomen slightly distended | 168
hypoactive bowel sounds | 168
elevations of alanine aminotransferase | 168
elevations of aspartate aminotransferase | 168
elevations of lactate dehydrogenase | 168
elevations of white blood cell count | 168
elevations of C-reactive protein | 168
anion gap metabolic acidosis | 168
lactic acidosis | 168
restart of noradrenaline and dobutamine infusions | 168
reintubated | 168
POCUS | 168
sluggish movement of the intestines | 168
bedside echocardiography | 168
severely impaired systolic function | 168
hyperechoic dot artifacts | 168
air extending to the periphery of the liver and hilum | 168
portal venous gas | 168
pneumatosis intestinalis | 168
CT of the abdomen | 168
intravenous and oral contrast | 168
portal venous gas in its tributaries | 168
superior mesenteric vein | 168
bowel ischemia | 168
foci of gas in the walls of the stomach | 168
right side of the colon | 168
small bowel loops | 168
marked atherosclerotic changes | 168
attenuated hepatic artery | 168
superior mesenteric artery | 168
celiac trunk | 168
nonvisualized inferior mesenteric artery | 168
minimal fluid in the pelvis | 168
extensive calcification of the superior mesenteric artery | 168
no occlusive thrombosis | 168
no significant luminal narrowing | 168
nonocclusive diffuse intestinal ischemia | 168
surgeon evaluated | 168
no further interventions | 168
passed away | 192