73 years old | 0
male | 0
myocardial infarction | -720
percutaneous coronary intervention | -720
stent inserted into left circumflex artery | -720
fever | -72
chills | -72
anorexia | -72
nauria | -72
diarrhea | -72
admitted to the hospital | 0
oxygen saturation 85% | 0
high-resolution computed tomography of the chest | 0
ground-glass opacity | 0
Tamiflu | 0
hydroxychloroquine | 0
KALETRA | 0
levofloxacin | 0
linezolid | 0
throat swab sample analyzed | 0
RT-PCR positive for COVID-19 | 0
breathing harder | 24
O2 saturation reduced to 94% | 24
nasal cannula | 24
facial mask | 48
non-rebreather mask | 48
respiratory distress | 72
oxygen saturation below 90% | 72
impairments of consciousness | 72
transferred to ICU | 72
meropenem | 72
impairments of consciousness more pronounced | 96
systolic blood pressure fluctuated | 96
difficult to maintain oxygen saturation over 89% | 96
severe sepsis | 96
septic shock | 96
endotracheal intubation | 144
ventilator with high positive end-expiratory pressure | 144
fraction of inspired oxygen 100% | 144
O2 saturation did not exceed 90% | 144
creatinine level increased | 144
acute kidney damage | 144
jugular vein access | 144
symptoms getting worse in an episodic manner | 144
temperature increased to 39°C | 144
chills | 144
tachycardia | 144
respiratory distress | 144
O2 saturation drop | 144
diarrhea | 144
blood pressure became more unstable | 144
hemoperfusion | 144
Heparin 50 mg/kg | 144
Heparin 15-20 mg/kg/h | 144
symptoms improved significantly | 144
need for oxygen therapy reduced | 144
fever disappeared | 144
heart rate decreased | 144
respiratory rate decreased | 144
second hemoperfusion | 168
mechanical ventilation support reduced | 168
extubated | 192
breathing independently | 192
discharged | 312
fever | 624
decreased oxygen saturation | 624
CT scan | 624
segmental pulmonary thromboembolism | 624
anticoagulant therapy | 624
Enoxaparin | 624
Rivaroxaban | 624
condition became stable | 630