60 years old | 0
male | 0
allergic to bee venom | 0
prostate cancer | 0
hypertension | 0
hypothyroidism | 0
eye surgery | 0
ankle surgery | 0
stung by bees | -24
injected epinephrine | -24
right-sided leg pain | 0
extreme tenderness | 0
diaphoretic | 0
morbidly obese | 0
blood pressure 155/83 mmHg | 0
heart rate 112 beats/min | 0
respiratory rate 16 breaths/min | 0
oxygen saturation 97% | 0
temperature 36.6°C | 0
temperature 38.5°C | 1
ALT 60 U/L | 0
AST 42 U/L | 0
bilirubin 1.5 mg/dL | 0
WBC 9.8 E9/L | 0
neutrophils 93.4% | 0
platelets 120 E9/L | 0
CT scan | 0
gas within the anterior compartment | 0
necrotizing fasciitis | 0
clindamycin 900 mg IV | 0
piperacillin-tazobactam 4.5 g IV | 0
vancomycin 2.5 g IV | 0
surgery for right leg debridement | 1.17
Bovie-cut | 1.17
fasciotomy | 1.17
compartment syndrome | 1.17
debridement | 1.17
wound cultures | 24
Clostridium perfringens | 24
vancomycin discontinued | 24
ertapenem 500 mg IV | 96
excisional debridement | 96
wound vac | 96
topical negative-pressure therapy | 96
hyperbaric oxygen therapy | 96
intermittent hemodialysis | 48
tunneled dialysis catheter | 96
discharged | 264
hyperbaric oxygen therapy continued | 264
dialysis catheter removed | 720
HBO therapy completed | 864
wound healing | 864
able to walk | 864