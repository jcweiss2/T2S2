57 years old | 0
male | 0
obese | 0
body mass index = 39 | 0
admitted to the hospital | 0
breathing constrained disturbances | 0
dyspnea | 0
severe back pain | 0
left knee pain | 0
left knee swelling | 0
asymptomatic consumption of domestic poultry | -720
domestic animals | 0
transferred from another hospital | 0
treated with bed rest for 2 weeks | -336
spine fracture | -336
misdiagnosis | -336
physical examination | 0
no pathologic neurological findings | 0
left osteoarthritic knee | 0
swollen left knee | 0
pleural effusion | 0
chest roentgenogram | 0
lateral plain roentgenogram | 0
computed tomography (CT)-scan | 0
destruction of the T12-vertebral body | 0
intervertebral discs T11-T12 and T12-L1 | 0
paravertebral abscess formation | 0
white blood cells (WBC’s) = 17.5 k/Μl | 0
C-reactive protein (CRP) = 23.1 mg/dL | 0
ESR = 86 mm/1st h | 0
tuberculosis antibody test | 0
virological laboratory tests | 0
rheumatologic laboratory tests | 0
Widal-Wright | 0
urine and stool cultures | 0
blood cultures revealed SE | 0
thoracic drainage tube inserted | 0
3000 cc of seropurulent fluid evacuated | 0
knee puncture | 0
120 cc of purulent fluid evacuated | 0
percutaneous transpedicular biopsy | 0
specimen culture | 0
all cultures isolated SE | 0
quinolone and 3rd generation cephalosporin given | 0
T12 biopsy disclosed chronic osteomyelitis | 0
thoracotomy | 24
left lung stuck to the parietal pleura | 24
residual empyema | 24
7 ml of purulent material evacuated | 24
T12-vertebrectomy | 24
disc resection | 24
bone debridement | 24
expandable titanium mesh cage (TMC) inserted | 24
spine stabilized | 24
knee fused | 720
superficial wound infection | 720
Acinetobacter | 720
local debridement | 720
secondary closure | 720
left knee fused completely | 2160
IV antibiotic treatment | 0
3 months IV antibiotic treatment | 0
discharged | 2160
monthly check of inflammatory markers | 2160
CRP and ESR within normal limits | 4320
radiograms and CT scan showed good result of fusion | 4320
patient free of pain | 4320
patient returned to daily routine | 4320
no sign of recurrence | 4320
anxious | 5040
altered state of consciousness | 5040
cognition | 5040
intubated | 5040
transferred to intensive care unit | 5040
brain CT scan revealed edema | 5040
hydrocephalus | 5040
drainage tube installation | 5040
lumbar puncture | 5040
cerebrospinal fluid indicative of viral infection | 5040
EEG showed slow waves | 5040
blood cultures revealed SE | 5040
patient did not recover | 5280
disconnected from ventilator | 5280
clinically dead | 5280