67 years old| 0
man| 0
admitted to the hospital| 0
sudden onset confusion| -336
dysarthria| -336
tested positive for SARS-CoV-2| -336
sore throat| -336
headache| -336
fever| -336
body aches| -336
diarrhea| -336
hypoxic| 0
oxygen saturation of 75%| 0
supplemental oxygen application| 0
oxygen saturation improved to 95%| 0
lymphocytopenia| 0
thrombocytopenia| 0
borderline lactic acidosis| 0
mixed respiratory acidosis| 0
metabolic acidosis| 0
prothrombin time-international normalized ratio| 0
platelet count| 0
sequential organ failure assessment score| 0
SIC score of 5| 0
bilateral airspace opacities| 0
generalized seizure| 24
cardiac arrest| 24
resuscitation| 24
admitted to the intensive care unit| 24
heparin anticoagulation| 24
vasopressors| 24
mechanical ventilation| 24
ventilator set to airway-pressure-release-ventilation mode| 24
poor ventilator synchrony| 48
switched to pressure-control mode| 48
positive end-expiratory pressure of 5 cm H2O| 48
FiO2 at 50%| 48
respiratory rate of 8 breaths/min| 48
inspiratory pressure of 10 cm H2O| 48
focal region wedge-shaped low attenuation in the left temporal region| 24
acute infarct| 24
diffuse subpleural pneumonitis| 24
ground-glass opacities| 24
consolidation| 24
paraseptal emphysema| 24
acute bilateral pulmonary emboli| 24
right ventricular dysfunction| 24
increasing vasopressor requirements| 120
increasing oxygen demands| 120
unchanged chest radiograph| 120
terminally extubated| 120
hypertension | 0
dyslipidemia | 0
sudden onset confusion | 0
dysarthria | 0
tested positive for SARS-CoV-2 | -336
sore throat | -336
headache | -336
fever | -336
body aches | -336
diarrhea | -336
sudden onset confusion| 0
dysarthria| 0
ventilator set to airway-pressure-release5 mode| 24
