49 years old | 0
    woman | 0
    fell while bathing | -72
    struck face on bath tap faucet | -72
    5 cm partial thickness laceration below left eye | -72
    laceration adjacent to medial canthus | -72
    laceration extending to left malar prominence | -72
    attended local A&E department | -72
    laceration debrided | -72
    laceration irrigated | -72
    laceration sutured | -72
    medical history: Elhers-Danlos syndrome | 0
    medical history: ischemic heart disease | 0
    medical history: previous anaphylaxis to penicillin | 0
    returned to A&E | -48
    complaining of pain below left eye | -48
    complaining of swelling below left eye | -48
    left eye partially closed | -48
    lower lid swelling | -48
    eye examination normal | -48
    no deficit in visual acuity | -48
    systemically well | -48
    discharged | -48
    oral clarithromycin | -48
    possible wound infection | -48
    re-attended A&E | -24
    pyrexial (38.7°C) | -24
    tachycardic (102/min) | -24
    rigors | -24
    confusion | -24
    extensive left-sided facial swelling | -24
    complete closure of left eye | -24
    involvement of soft tissues of left neck | -24
    reduction in left visual acuity | -24
    urgent blood results | -24
    marked neutrophilia | -24
    raised C-reactive protein | -24
    acute bacterial infection | -24
    laceration opened | -24
    necrotic skin edges | -24
    absence of bleeding | -24
    severe facial necrotizing fasciitis | -24
    admitted | 0
    underwent immediate widespread local excision | 0
    excision of necrotic tissue from left lower eyelid | 0
    excision of necrotic tissue from left cheek | 0
    excision of necrotic tissue from soft tissues overlying left angle of mandible | 0
    excision of necrotic tissue from lateral aspect of upper neck | 0
    peri-operative IV clindamycin | 0
    peri-operative IV gentamicin | 0
    post-operative IV clindamycin | 0
    post-operative IV gentamicin | 0
    transferred to ICU | 0
    post-operative support | 0
    remained clinically septic | 24
    extension of necrotic tissue beyond surgical margins | 24
    left eye involvement suspected | 24
    urgent CT scan | 24
    left retro=orbital necrosis | 24
    further surgical excision | 24
    excision of necrotic tissue from left forehead | 24
    excision of necrotic tissue from left temporal region | 24
    excision of necrotic tissue from left upper eyelid | 24
    excision of necrotic tissue from left commissure | 24
    exenteration of left orbital contents | 24
    blood samples sent to microbiology | 24
    tissue samples sent to microbiology | 24
    florid growth of Group A beta-hemolytic Streptococci | 24
    facial necrotizing fasciitis confirmed | 24
    transferred to ICU | 24
    2-week period in ICU | 336
    transferred to surgical high dependency | 336
    3 weeks of ward-based care | 504
    oral clindamycin continued | 504
    initial split thickness skin graft from right thigh | 504
    unsuccessful graft | 504
    second graft required | 504
    wound healing concerns | 504
    graft failure concerns | 504
    abnormal collagen synthesis in Ehlers-Danlos syndrome | 504
    patient reluctance for further surgery | 504
    limited reconstructive attempts | 504

    