84 years old | 0
male | 0
dementia | 0
fever | -48
upper respiratory infection | -48
treatment for upper respiratory infection | -48
decline in blood pressure | -48
decrease in SpO2 | -48
loss of consciousness | -48
admitted to the hospital | 0
respiratory failure | 0
shock | 0
blood pressure 77/48 mmHg | 0
pulse rate 107 beats per minute | 0
SpO2 84% | 0
oxygen administration 10 L/min | 0
respiratory rate 32 breaths per minute | 0
body temperature 38.3℃ | 0
coarse crackles on bilateral lung fields | 0
altered level of consciousness | 0
Japan Coma Scale III-200 | 0
Glasgow Coma Scale 3 | 0
chest radiograph | 0
CT scan | 0
diffuse consolidation in both lungs | 0
leukocytosis | 0
neutrophilia | 0
high C-reactive protein level | 0
elevation of liver and biliary enzyme levels | 0
hypoproteinemia | 0
renal dysfunction | 0
high creatine kinase levels | 0
thrombocytopenia | 0
prolonged prothrombin time | 0
elevated fibrin degradation products | 0
disseminated intravascular coagulopathy | 0
septic shock | 0
aspiration pneumonia | 0
APACHEII score 30 | 0
Sequential Organ Failure Assessment score 15 | 0
meropenem hydrate | 0
dopamine hydrochloride | 0
nafamostat mesylate | 0
nasogastric feeding tube insertion | 48
enteral nutrition | 72
polymeric formula | 72
fever 39.5℃ | 216
decrease in SpO2 | 216
white blood cell count increased | 216
chest radiograph | 216
fresh infiltrations in the right lower field | 216
aspiration from gastric feed reflux | 216
gastric feeding intolerance | 216
nasojejunal tube insertion | 240
gastric decompression function | 240
fluoroscopic guidance | 240
contrast medium | 240
enteral feeding | 240
gastric drainage | 240
dopamine hydrochloride discontinued | 72
nafamostat mesylate discontinued | 120
meropenem hydrate discontinued | 336
sulfamethoxazole | 336
percutaneous endoscopic gastrostomy | 528
swallowing therapy | 1008
discharged | 1032