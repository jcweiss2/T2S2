25 years old | 0
mother | 0
hypothyroidism | 0
meconium-stained amniotic fluid | 0
membranes ruptured | -1
vaginal birth | 0
term baby boy | 0
39w + 4d | 0
birth weight normal | 0
head circumference normal | 0
length normal | 0
good muscle tone | 0
cried vigorously | 0
1st minute Apgar score 9 | 0
respiratory distress | 2
cyanosis | 2
5th minute Apgar score 6 | 2
oxygen saturation level 60% | 2
NCPAP administered | 2
SpO2 level rose | 2
transferred to NICU | 2
SpO2 level dropped | 2
tachypnea | 2
mild intercostal retraction | 2
moderate subcostal retraction | 2
nasal flaring | 2
grunting | 2
full and symmetrical pulses | 2
temperature 37.1°C | 2
respiratory rate 70 breaths/min | 2
heart rate 152 bpm | 2
blood pressure 69/42 mmHg | 2
SpO2 60-65% | 2
decreased sucking | 2
normal grasp | 2
normal Moro reflexes | 2
NCPAP failure | 2
NIPPV administered | 2
SpO2 did not increase | 2
endotracheal suctioning | 2
intubated | 2
sepsis workup | 2
CXR performed | 2
diffuse patchy granular infiltrates | 2
MAS suspected | 2
surfactant administered | 2
respiratory acidosis | 2
VBG revealed | 2
peak inspiratory pressure increased | 4
positive end-expiratory pressure reduced | 4
second dose of surfactant administered | 10
SpO2 increased | 24
VBG improved | 24
COVID-19 RT-PCR performed | 4
COVID-19 RT-PCR result positive | 24
remdesivir administered | 24
IVIG administered | 24
methylprednisolone administered | 24
liver and kidney function tests performed | 24
ferritin level requested | 24
inotropes tapered | 96
fentanyl dosage reduced | 96
extubation prepared | 96
ventilatory support decreased | 120
extubated | 120
NIPPV initiated | 120
SpO2 90-95% | 120
inotropes ceased | 120
CXR repeated | 120
significant improvement | 120
COVID-19 PCR repeated | 120
COVID-19 PCR negative | 120
methylprednisolone tapered | 168
methylprednisolone discontinued | 336
nebulized magnesium sulfate initiated | 168
SpO2 drops stopped | 192
tachypnea improved | 192
magnesium sulfate stopped | 312
discharged | 312
no need for oxygen therapy | 312
follow-up visits planned | 312
last follow-up visit | 744
no respiratory problem | 744
mother tested for COVID-19 | 24
mother COVID-19 positive | 24
mother asymptomatic | 24
mother silent carrier | 480