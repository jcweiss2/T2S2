54 years old | 0
female | 0
admitted to hospital | 0
allergic reaction | -6
amoxicillin | -6
upper respiratory tract infection | -6
transient episodes of turning pale | -648
feeling lightheaded | -648
diffuse non-blanching rash | -6
intravenous adrenaline | -6
hydrocortisone | -6
chest tightness | 0
diffuse mottled vasculitic rash | 0
livedo reticularis | 0
pyrexial | 0
hypertensive | 0
persistently tachycardic | 0
elevated white cell count | 0
C reactive protein | 0
deranged liver function | 0
coagulation profile | 0
biochemical evidence of acute kidney injury | 0
broad spectrum antibiotics | 0
intravenous fluids | 0
supportive therapy | 0
restless | 72
agitated | 72
altered level of consciousness | 72
global encephalopathy | 72
CT head | 72
lumbar puncture | 72
septic screen | 72
CT abdomen | 72
10 cm heterogeneous right adrenal mass | 72
atrial fibrillation | 72
fast ventricular rate | 72
drop in blood pressure | 72
noradrenaline | 72
labile blood pressure | 144
discontinued noradrenaline | 144
intravenous phentolamine | 144
pheochromocytoma crisis | 144
24-h urinary metanephrine measurement | 144
blood pressure stabilized | 180
oral phenoxybenzamine | 192
cardiac arrest | 240
cardiopulmonary resuscitation | 240
ejection fraction of 40% | 240
endocrine surgical opinion | 240
emergency adrenalectomy | 240
multi-organ failure | 240
low Glasgow Coma Scale | 240
deterioration | 384
death | 384