44 years old | 0
female | 0
ECOG performance status 0 | 0
admitted to the hospital | 0
ulcerated MM | -672
Breslow thickness of 1.2 mm | -672
mitosis between 1 and 6 per mm2 | -672
absence of intense intra-tumor lymphocyte infiltrate | -672
Stage III C | -672
BRAF-V600E specific mutation | -672
Pembrolizumab 200 mg flat dose | 0
treatment cycles | 0
severe grade 3 diarrhea | 120
abdominal pain | 120
weight loss | 120
fever | 120
neutropenia | 120
hospitalization | 120
Loperamide and hydration | 120
intravenous antibiotic therapy | 120
Piperacillin/Tazobactam | 120
Vancomycin | 120
antimycotic treatment | 120
bone marrow biopsy | 120
severe hypocellularity | 120
marked reduction of maturing granulopoiesis | 120
normal erythroid component | 120
autoimmune neutropenia | 120
high dose of corticosteroids | 120
methylprednisolone 2 mg/kg | 120
granulocyte colony-stimulating factor (GCSF) | 120
oxygen therapy | 120
Venturi mask | 120
high flow oxygenation ventilation device | 120
hypoxemic respiratory failure | 120
alkalosis | 120
intensive care unit (ICU) | 120
corticosteroid-resistant colitis | 168
Vedolizumab | 168
300 mg flat dose | 168
induction scheme | 168
reduction of symptoms | 168
steroids tapering | 168
disappearance of symptoms | 192
reduction of CRP | 192
reduction of calprotectin | 192
sigmoidoscopy | 336
biopsies | 336
mucosal healing | 336
HLA class I and II | 336
HLA A*02 *02 | 336
HLA B*14 *35 | 336
HLA C *04*08 | 336
HLA DRB *01 *07 | 336
Pembrolizumab therapy discontinued | 336
clinical and instrumental follow-up | 336
Vedolizumab treatment ongoing | 336
maintenance scheme | 336
good general conditions | 744
no signs of disease progression | 744
endoscopic appearance of remission | 744