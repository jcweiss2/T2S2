33 years old | 0
female | 0
admitted to the hospital | 0
cardiac arrest | -1
attempted suicide by hanging | -1
advanced cardiovascular life support | -1
left leg IO needle placement | -1
intubated | 0
admitted to the neurologic intensive care unit | 0
left leg pain | 48
severe tenderness at the left shin IO site | 48
decreased strength on ankle dorsal and plantar flexion | 48
mild dorsal foot swelling | 48
conventional radiograph of the left leg | 48
small, shallow, and linear cortical defect in the proximal diaphysis of the lateral tibial cortex | 48
moderate localized soft tissue swelling | 48
increased swelling and erythema of the left leg | 96
differential considerations: deep venous thrombosis, infection, or sequela of possible blunt soft tissue trauma | 96
elevated D-dimer | 96
pulmonary CT angiography | 96
negative for pulmonary embolism | 96
ultrasound for DVT | 96
negative for DVT | 96
CT of the lower extremities | 96
small, shallow, and linear cortical defect in the anterolateral tibia | 96
asymmetric soft tissue swelling of the left tibialis anterior muscle | 96
left lower extremity magnetic resonance imaging | 96
small, partial-thickness cortical defect along the anterior lateral aspect of the proximal tibia | 96
marked distention of the anterior muscle compartment | 96
abnormally increased T1 and T2 signal consistent with early subacute intramuscular hemorrhage | 96
surgical consultation for a potential fasciotomy | 96
watchful waiting approach | 96
pain and swelling gradually decreased | 120
discharged from the hospital | 120