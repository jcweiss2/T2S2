urinary tract infection | -120
fever | -120
dysuria | -120
clean catch urine specimen collected | -120
started on cephalexin | -120
urine analysis positive for large leukocyte esterase and bacteria | -120
urine culture grew Escherichia coli | -120
cephalexin 500 mg three times daily | -120
extensive erythematous rash | -48
rash developed into sloughing of the skin | -48
discontinued cephalexin | -24
transferred to local burn intensive care unit | -24
admitted to hospital | 0
difficulty swallowing | 0
endotracheal tube placed | 0
diagnosed with toxic epidermal necrolysis syndrome | 0
pulmonary infiltrates | 0
respiratory failure | 0
intubated | 0
two peripheral blood cultures obtained | 0
skin surveillance cultures of nares, axilla, and groin | 0
urine culture from newly placed indwelling Foley catheter | 0
chest radiograph revealed right pleural effusion | 0
right lower and left basilar opacities | 0
norepinephrine and vasopressin drips | 0
continuous infusion of albumin 25% | 0
lactated Ringer’s | 0
tetanus–diphtheria toxoids vaccine | 0
gentamicin 120 mg | 0
fluconazole 100 mg | 0
WBC 5.4 × 103/mm3 | 24
SCr 1.98 mg/dL | 24
venous serum lactate 1.8 mmol/L | 24
random serum gentamicin level 2.4 mg/dL | 24
redosed with 120 mg of gentamicin | 27
supportive continuous renal replacement therapy | 24
fluconazole continued at 200 mg IV every 24 h | 24
Gram’s stain of the tracheal aspirate showed heavy growth of pleomorphic Gram-negative rods and diphtheroid-like Gram-positive rods | 24
wide complex tachycardia | 96
amiodarone restarted | 96
gentamicin held | 96
physical examination revealed sloughing of skin | 120
culture and sensitivity results of the tracheal aspirate grew Pseudomonas aeruginosa | 120
gentamicin administered | 120
patient expired | 144
autopsy performed | 144
necrotizing bronchopneumonia | 144
Severity of Illness Score for TEN calculated | 144
predicted mortality of 62% | 144