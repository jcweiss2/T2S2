50 years old | 0
male | 0
admitted to the hospital | 0
alcoholism | 0
complaining of worsening pain | -48
complaining of redness of the right elbow | -48
history of trivial trauma | -48
X-ray of the elbow was negative | -48
discharged with non-steroidal anti-inflammatory drugs (NSAIDs) | -48
returned to the emergency department | -24
persistent erythema | -24
persistent tenderness around his elbow | -24
no systemic inflammatory symptoms | -24
skin erythema | -24
edema | -24
warmness | -24
tenderness | -24
no axillar lymphadenopathy | -24
white blood cell count of 7770/μL | -24
CRP 533.6 mg/L | -24
hemoglobin 14.8 g/dL | -24
glucose 0.83 g/L | -24
creatinine 1.4 mg/dL | -24
sodium 133 mmol/L | -24
LRINEC score of 6 | -24
kidney function tests were normal | -24
liver function tests were normal | -24
blood culture was negative | -24
diagnose of cellulitis | -24
treated with intravenous antibiotics | -24
Cefazoline 4 g daily | -24
Metronidazole 1500 mg daily | -24
condition continued to deteriorate | -120
intense pain | -120
significant edema | -120
tenderness of his right elbow | -120
wound culture revealed a Streptococcus pyogenes infection | -120
brought to our hospital for a surgical advice | -120
febrile | 0
blood pressure was 148/83 mmHg | 0
white blood cell count of 16000/μL | 0
CRP 95 mg/L | 0
LRINEC score of 3 | 0
blood endotoxin was negative | 0
margins of tenderness and erythema spread | 0
phlyctens | 0
areas of necrosis | 0
emergency aggressive debridement of necrotic tissues | 0
skin swabs taken during the operation were negative | 0
underlying muscles were intact | 0
transferred to the intensive care unit | 0
respiratory support | 0
renal support | 0
circulatory support | 0
treated with intravenous penicillin | 0
underwent multiple sets of vacuum-assisted closure (VAC) technique | 24
underwent hyperbaric oxygen therapy (HBOT) | 24
wound was closed by split-thickness skin graft | 168
postoperatively no complications | 168
discharged | 192
stiff elbow | 192
regained an acceptable range of motion of his right arm | 384
no sign of infection recurrence | 720