70 years old | 0
    male | 0
    admitted to the hospital | 0
    hypoesthesia in the fingers of each hand | -24
    proximal paresis of both legs (motor strength 2/5) | -24
    pronounced dysfunction of gait and standing | -24
    recent-onset bladder incontinence | -24
    rheumatoid arthritis | -24
    asthma | -24
    osteoporosis | -24
    ventral fusion and osteosynthetic stabilization | 0
    induction of anaesthesia with propofol and sufentanil | 0
    total intravenous anaesthesia with propofol infusion | 0
    sufentanil intermittent injections | 0
    mask ventilation | 0
    rocuronium administration | 0
    direct laryngoscopy oral intubation | 0
    Cormack–Lehane grade 1 | 0
    unremarkable oropharyngeal anatomy | 0
    continuous tracheal tube cuff pressure monitoring | 0
    cuff pressure approached 40 mmHg | 0
    splitting of sternocleidomastoid muscle compartment | 0
    lateral displacement of carotid sheath | 0
    microdiscectomy | 0
    polyetheretherketone (PEEK) cage fusion | 0
    osteosynthetic stabilisation | 0
    unremarkable intra-operative course | 0
    unusually large hyoid bone | 0
    no other significant surgical observations | 0
    total operating time 195 minutes | 0
    post-operative swelling of left side of throat | 24
    initial suspicion of surgery-induced hematoma | 24
    palpable laryngeal structures | 24
    probable intra-operative laryngeal dislocation | 24
    postponed extubation | 24
    computed tomography (CT) scan performed | 24
    fixation of overly elongated hyoid bone | 24
    leftward dislocation of entire larynx | 24
    ruled out large hematoma | 24
    transferred to neurosurgical intensive care unit | 24
    referred for Otolaryngology opinion | 24
    failed endolaryngeal repositioning attempt | 24
    indication for open repositioning next day | 24
    reopened wound full depth | 72
    hyoid bone released from entrapment | 72
    subsequent CT scan showed normal laryngeal position | 72
    substantial oedema formation | 72
    mucous membranes tightly surrounded endotracheal tube | 72
    continued intubation | 72
    anti-oedema therapy with dexamethasone | 72
    extubated on sixth post-operative day | 144
    respiratory insufficiency | 144
    reintubation necessary | 144
    bilateral pleural effusions | 144
    decreasing level of consciousness | 144
    conventional open tracheotomy performed | 288
    septic due to ventilator-associated pneumonia | 288
    responded to antibiotic therapy | 288
    decreased level of consciousness | 288
    neurological improvement slow | 288
    discharged into neurological early rehabilitation | 696
    awake and oriented | 696
    followed simple commands | 696
    could breathe using T-piece | 696