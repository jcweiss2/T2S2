56 years old | 0
female | 0
admitted to the hospital | 0
left-sided liver mass | -24
abdominal ultrasound scan | -24
denies previous history of chronic hepatitis | -24
denies alcohol abuse | -24
denies blood transfusion | -24
transabdominal subtotal hysterectomy | -24
concomitant unilateral ophorectomy | -24
utERine leiomyoma | -24
benign ovarian cyst | -24
physical examination unremarkable | -24
routine laboratory tests normal | -24
serum alpha-fetoprotein level 3.2 ng/mL | -24
CA19-9 level 488.43 U/mL | -24
contrast-enhanced upper abdominal ultrasonography | -24
multiple liver tumors | -24
left liver lobe and left-right lobe junction | -24
maximum dimensions 12.1 cm ×7.1 cm | -24
magnetic resonance cholangiopancreatography | -24
diagnosis of left-sided liver cancer | -24
Child-Pugh class A | -24
elective laparotomy | -24
left-sided hepatectomy | -24
hilar lymphadenectomy | -24
concomitant cholecystectomy | -24
histology moderately differentiated ICC | -24
chronic cholecystitis | -24
uneventful postoperative course | -24
follow-up upper abdominal ultrasonography | -56
recurrent diseases in right lobe | -56
Couinaud segments V, VII, and VIII | -56
sizes 1.5 cm ×1.3 cm, 1.2 cm ×1.0 cm, and 0.9 cm ×1.0 cm | -56
liver function reserve class A | -56
serum alpha-fetoprotein level 2.9 ng/mL | -56
Doppler ultrasound-guided RFA | 0
LDRF-120S | 0
conscious sedation anesthesia | 0
puncture through right subcostal margin | 0
three sessions of RFA | 0
initial power 78 W | 0
total duration 16 minutes | 0
follow-up ultrasound scan | 72
filling defect in ablated area | 72
hypoechogenic residual mass | 72
repeated liver and coagulation function tests | 72
no clinically significant abnormality | 72
second RFA | 120
initial power 50 W | 120
total duration 7 minutes | 120
febrile | 144
hemoglobin 80 g/L | 144
white cell count 10.4×10^9/L | 144
liver biochemistry abnormal | 144
alanine transferase 5,304 IU/L | 144
aspartate transferase 7,906 IU/L | 144
albumin 30.7 g/L | 144
total bilirubin 38.9 μmol/L | 144
prothrombin time 22.4 seconds | 144
international normalized ratio 1.91 | 144
emergency contrast-enhanced magnetic resonance imaging | 144
extensive liver necrosis | 144
diagnosis of RFA-associated ALF | 144
symptomatic treatment | 144
prophylactic antimicrobial therapy | 144
blood transfusion | 144
nutritional liver support | 144
lactose enemas | 144
intravenous infusion of aspartic acid, ornithine, and arginine | 144
hyperammonemia | 144
respiratory distress | 144
agitated | 144
confused | 144
heart rate increased | 144
pulse oxygen saturation deteriorating | 144
arterial blood gas analysis | 144
PO2 71 mmHg | 144
PCO2 50 mmHg | 144
pH 7.32 | 144
chest X-ray | 144
bilateral pulmonary extensive inflammatory changes | 144
pleural effusion | 144
contrast echocardiogram | 144
diagnosis of HPS | 144
transnasal intubation | 144
respiratory care unit | 144
mechanical ventilation | 144
tracheostomy | 144
repeated chest X-ray | 240
ultrasound scan | 240
progressively improving pulmonary sepsis | 240
pleural effusion | 240
weaned from ventilator | 336
liver function test improvement | 360
discharged | 792
follow-up at outpatient clinic | 8760
survived free of recurrence | 8760