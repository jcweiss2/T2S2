21 years old | 0
African American | 0
male | 0
admitted to the hospital | 0
GSW to the right posterior thorax | -1
no medical history | 0
tachycardia | 0
hypotension | 0
pain in the right posterior thorax | 0
shortness of breath | 0
decreased breath sounds in the right thorax | 0
right-sided pleural effusion | 0
right pneumothorax | 0
shrapnel material overlying the right inferior thorax | 0
right-sided chest tube placement | 0
1,000 mL of blood drained | 0
heart rate normalized | 1
blood pressure normalized | 1
CT of the chest and abdomen | 2
metallic fragment within the right atrium | 2
right atrial exploration | 4
thoracic IVC repair | 4
general endotracheal anesthesia | 4
left radial and right femoral arterial catheters insertion | 4
right internal jugular central venous catheter insertion | 4
sternotomy | 4
cardiopulmonary bypass initiation | 4
volatile agents administration | 4
opiates administration | 4
benzodiazepines administration | 4
crystalloid administration | 4
blood products administration | 4
vasopressor agents administration | 4
TEE before sternotomy | 4
normal left ventricle | 4
suspicious for IVC or right atrial hematoma | 4
no intracardiac bullet fragments identified | 4
IVC repair | 6
good right ventricular and left ventricular function | 6
radiolucent particle within the intrahepatic IVC | 6
portable intraoperative CXR | 6
shrapnel material lying within the hepatic IVC | 6
weaned from cardiopulmonary bypass | 8
chest closure | 8
transferred to a hybrid operating suite | 8
inferior venacavagraphy | 10
successful removal of a 2-cm bullet fragment | 10
fluoroscopic images | 10
hemodynamically stable | 10
estimated blood loss of approximately 300 mL | 10
transferred to the cardiothoracic intensive care unit | 12
sudden output of roughly 2.5 L of bloody discharge | 12
transfused 6 U of packed red blood cells | 12
transfused 4 U of fresh frozen plasma | 12
transfused 1 U of cryoprecipitate | 12
transfused one pack of pooled platelets | 12
coagulopathy corrected | 12
chest tube output decreased | 12
chest packed and remained open overnight | 12
chest closed | 24
sedation weaned | 48
extubated | 48