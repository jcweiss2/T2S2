24 years old | 0
male | 0
obese | 0
admitted to the hospital | 0
nausea | 0
nonbilious vomiting | 0
hematemesis | 0
fever | -72
fatigue | -72
dry cough | -72
chills | -72
diabetes mellitus type 1 | -8760
hyperlipidemia | -8760
noncompliant with medications | -72
temperature 36.4°C | 0
pulse rate 122 beats/min | 0
blood pressure 141/84 mmHg | 0
respiratory rate 16 breaths/min | 0
oxygen saturation 95% | 0
hypothermic | 2
temperature 32.9°C | 2
Foley probe temperature 36.8°C | 2
mild distress | 0
lethargic | 0
delayed responses | 0
dry mucous membranes | 0
blood glucose 507 mg/dL | 0
hemoglobin A1c 15.8% | -720
ketonuria 160 mg/dL | 0
elevated creatinine 1.4 mg/dL | 0
anion gap 30.6 mEq/L | 0
DKA with metabolic encephalopathy | 0
sepsis | 0
vancomycin | 0
cefepime | 0
sodium bicarbonate infusion | 0
potassium repletion | 0
insulin intravenously | 0
lethargic | 24
fell asleep | 24
DKA with anion gap metabolic acidosis | 24
acute kidney injury | 24
oxygen saturation 99% | 24
increased leukocyte count | 24
cardiac troponins negative | 24
respiratory distress | 48
febrile | 48
tachypneic | 48
SARS-CoV-2 nasopharyngeal swab positive | 48
intubated | 48
mechanically ventilated | 48
chest X-ray showed mild perihilar patchy areas of opacity | 48
azithromycin | 72
hydroxychloroquine | 72
febrile | 96
tachycardic | 96
attempt to titrate FiO2 to 60% | 96
oxygen saturation dropped to 86% | 96
arterial blood gas testing showed improvements | 96
desaturated to 75% | 168
leukocyte count increased | 168
sputum sample collected | 168
vancomycin and cefepime discontinued | 168
meropenem | 168
voriconazole | 168
sputum results showed yeast isolates | 192
chest X-ray showed interval worsening of infiltrates | 192
intermittently febrile | 216
attempts to titrate FiO2 unsuccessful | 216
desaturations | 216
arterial blood gasses revealed worsening hypercapnia | 216
chest X-ray showed diffuse fluffy infiltrates | 216
ARDS | 216
severely hypotensive | 216
bradycardia | 216
pulseless | 216
advanced cardiovascular life support protocol initiated | 216
death | 216