71 years old | 0
male | 0
hypertension | 0
type 2 diabetes mellitus | 0
admitted to the hospital | 0
COVID-19 pneumonia | 0
transferred to our hospital | -48
tocilizumab | -48
corticosteroid | -48
initial COVID-19 RT-PCR test | 0
SARS-CoV-2 positive | 0
no COVID-19 vaccine | 0
hypoxemic respiratory insufficiency | 0
pulmonary involvement by COVID-19 | 0
CT findings (CO-RADS 5-6) | 0
intubated | 0
PaO2/FIO2 ratio of 120 | 0
mechanical ventilation initiated | 0
leukocytosis (29,000 k/uL) | 0
lymphopenia (0.40 K/uL) | 0
C-reactive protein (44 mg/L) | 0
IL-6 (4365 pg/mL) | 0
ferritin (>2000 ng/mL) | 0
D-dimer (6520 ng/mL) | 0
LDH (785 U/L) | 0
creatinine (2.1 mg/dL) | 0
culture samples taken | 0
empiric antibiotic therapy (imipenem, levofloxacin) | 0
renal function deteriorated | 168
four hemofiltration sessions | 168
chest radiography (CXR) revealed cavitary image | 168
hemoculture (no bacterial growth) | 168
urine culture (no bacterial growth) | 168
broad-spectrum antibiotics (meropenem, vancomycin) | 168
antifungal fluconazole | 168
bronchoscopy procedure performed | 168
erythematous lesions in the bronchial tree | 168
abundant purulent secretions | 168
cavitary lesion in the right bronchial tree | 168
BAL isolated Klebsiella pneumoniae | 312
BAL isolated Pseudomonas aeruginosa | 312
BAL fungal culture isolated Trichosporon asahii | 312
BAL negative for ZN stain | 312
BAL negative for GeneXpert MTB/RIF | 312
Löwenstein-Jensen culture negative | 312
ceftazidime/avibactam | 312
colistin | 312
voriconazole | 312
disease progression | 360
septic shock | 360
multi-organ failure | 360
died | 384
fever | -48
cough | -48
dyspnea | -48
oxygen therapy with noninvasive mechanical ventilation | 0
ceftazidime | 0
corticosteroids | 0
invasive mechanical ventilation | 24
septic shock | 24
renal failure (eGFR 27.5 mL/min/1.73 m2) | 24
imipenem/cilastatin | 24
levofloxacin | 24
antithrombotic | 24
eGFR (16.6 mL/min/1.73 m2) | 72
oligoanuria | 72
metabolic acidosis | 72
hemodiafiltration started | 96
second hemodiafiltration session | 120
urea (16) | 120
creatinine (1.9) | 120
improved metabolic acidosis | 120
diuresis | 120
third hemodiafiltration session | 144
leukocytosis | 144
neutrophilia | 144
elevated inflammatory markers | 144
CXR cavitary image in right upper lobe | 144
respiratory weaning failure | 288
sedation | 288
relaxation | 288
paralysis | 288
ventilator strategy protection | 288
FiO2 100% | 312
tidal volume 7-8 mL/kg | 312
respiratory rate 20 per minute | 312
PEEP 5 cm H2O | 312
pressure limit 60 cm H2O | 312
maximum inspiratory flow rate 50 | 312
ramp wave | 312
leak compensation | 312
BAL sample isolation | 336
treatments with ceftazidime/avibactam | 336
colistin | 336
voriconazole | 336
patient deceased | 384
