28 years old | 0 | 0 
male | 0 | 0 
admitted to the hospital | 0 | 0 
fatigue | -48 | 0 
anosmia | -48 | 0 
dyspnea | -48 | 0 
SpO2 levels 55% | -48 | -48 
nasal cannula oxygen therapy | -48 | 0 
chest radiography | 0 | 0 
bilateral lung infiltrates | 0 | 0 
RT-PCR swab tested positive for SARS-CoV-2 infection | 0 | 0 
admitted in a COVID-19 infirmary unit | 0 | 0 
non-invasive ventilation support | 0 | 24 
intubation | 24 | 24 
invasive mechanical ventilation | 24 | 168 
ventral decubitus positioning | 24 | 168 
Escherichia coli detected on sputum culture | 48 | 48 
methicillin-sensitive Staphylococcus aureus detected on sputum culture | 48 | 48 
superinfection | 48 | 48 
amoxicillin prescribed | 48 | 168 
blood culture revealed methicillin-resistant Staphylococcus aureus | 48 | 48 
steady clinical improvement | 168 | 168 
extubated | 168 | 168 
discharged | 168 | 168 
retrosternal thoracalgia | 168 | 168 
thoracalgia irradiating to the left upper limb | 168 | 168 
abduction and external rotation limited due to pain | 168 | 168 
soft tissue swelling of the shoulder and arm | 168 | 168 
fever | 168 | 168 
increased levels of C-reactive protein | 168 | 168 
admitted for further investigation and treatment planning | 168 | 168 
gentamicin prescribed | 168 | 240 
thoracic CT with intravenous contrast administration | 216 | 216 
scapulohumeral synovitis | 216 | 216 
intra-muscular collections | 216 | 216 
glenohumeral joint fluid | 216 | 216 
bilateral shoulder magnetic resonance imaging (MRI) with intravenous contrast administration | 240 | 240 
infraspinatus fossa and subscapular fossa collections | 240 | 240 
capsular thickening and increased signal intensity post-gadolinium administration | 240 | 240 
septic arthritis and rotator cuff collections | 240 | 240 
myonecrosis | 240 | 240 
aspiration of the infraspinatus fossa collection | 252 | 252 
seropurulent fluid sent for analysis | 252 | 252 
drainage catheter left on the left infraspinatus collection | 252 | 252 
drainage catheter removed | 264 | 264 
physical rehabilitation exercises | 264 | 312 
improvement of left shoulder range of motion | 312 | 312 
transferred to another hospital | 312 | 312 
indication to continue physical therapy and rehabilitation exercises | 312 | 312