40 years old | 0
female | 0
admitted to the hospital | 0
swelling in the right side of the face | -264
extraction of an upper right back tooth | -264
feeling normal | -264
pain | -264
unhealed socket | -264
decreased mouth opening | -264
referred to the medical school | -264
toxic | 0
Glasgow coma scale score of 11 | 0
temperature of 40 | 0
tender swelling | 0
fluctuant swelling | 0
necrosis over the right infraorbital region | 0
diplopia | 0
dilated pupil | 0
proptosis | 0
periorbital ecchymosis | 0
loss of vision | 0
abducens nerve palsy | 0
chemosis of the right eye | 0
maxillary tuberosity fractured | 0
necrosis of the palatal mucosa | 0
necrosis of the upper right vestibule | 0
random blood sugar value of 311 mg/dL | 0
total leucocyte count of 18,200 cubic millimeter of blood | 0
polymorph value of 92% | 0
mucosal thickening involving the bilateral maxillary and right ethmoidal sinuses | 0
venous dilatation of the right superior ophthalmic vein | 0
abscess in the right side of the buccal and temporal spaces | 0
intravenous antibiotics | 0
imipenem | 0
clindamycin | 0
ceftriaxone | 0
chloramphenicol | 0
metronidazole | 0
furosemide | 0
mannitol | 0
dexamethasone | 0
nonsteroidal anti-inflammatory drugs | 0
paracetamol | 0
human mixtard insulin | 0
low molecular weight heparin | 0
provisional diagnosis of CST | 0
emergency incision and drainage of the right buccal and temporal spaces | 24
admitted to the intensive care unit | 24
chemosis in the left eye | 48
paralysis of the contralateral side of the body | 48
Glasgow coma scale score of 7 | 48
ventilator | 48
meningitis | 72
septic emboli | 72
blindness | 72
cranial nerve palsies | 72
sepsis | 72
shock | 72
died | 72