48 years old | 0
    male | 0
    admitted to the emergency room | 0
    asthenia | -720
    daily fever | -720
    night sweats | -720
    weight loss of 6 kg | -720
    cough | -120
    dyspnea on exertion | -120
    pancytopenia | -168
    severe neutropenia | -168
    hemoglobin 6.0 g/dL | -168
    leukocyte count 0.8 × 10^9/L | -168
    neutrophil count 0.14 × 10^9/L | -168
    lymphocyte count 0.48 × 10^9/L | -168
    monocyte count 0.17 × 10^9/L | -168
    platelet count 70.0 × 10^9/L | -168
    no adenopathy | 0
    no hepatosplenomegaly | 0
    negative family history for hematological disorders | 0
    negative family history for neoplasms | 0
    bacterial pneumonia | 0
    hospitalized in semi-intensive care unit | 0
    negative blood cultures | 0
    negative serum galactomannan test | 0
    bone marrow aspirate | 0
    lymphoid cells with hairy cell morphology | 0
    immunophenotyping confirmation of HCL | 0
    negative BRAF V600E mutation | 0
    septic shock | 24
    ARDS | 24
    acute renal injury | 24
    hemodialysis | 24
    orotracheal intubation | 24
    negative tracheal aspirate cultures | 24
    broadened antibiotic regimen | 24
    meropenem | 24
    liposomal amphotericin B | 24
    vancomycin | 24
    filgrastim | 24
    IFN-α started | 24
    weaning of vasoactive drugs | 168
    extubated | 168
    increasing neutrophil count | 168
    filgrastim administered for seven days | 168
    two packed red blood cell units provided | 0
    hemoglobin 8.2 g/dL | 168
    leukocyte count 2.68 × 10^9/L | 168
    neutrophil count 1.1 × 10^9/L | 168
    lymphocyte count 1.4 × 10^9/L | 168
    monocyte count 0.1 × 10^9/L | 168
    platelet count 0.63 × 10^9/L | 168
    recovery of renal function | 168
    cladribine prescribed | 216
    discharged | 240
    complete blood count recovery | 240
    satisfactory general condition | 240
    bone marrow biopsy confirming complete response | 4320
    