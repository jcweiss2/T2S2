47 years old | 0
male | 0
admitted to the hospital | 0
pain | -336
massive cervical swelling | -336
oral antibiotic therapy | -336
difficulty in breathing | 0
difficulty in swallowing | 0
necrotic soft tissue areas | 0
pus presence | 0
computed tomography of neck and chest | 0
extensive soft tissue emphysema | 0
left third molar infection | 0
no mediastinal inflammatory involvement | 0
extraction of third molar | 0
drainage | 0
surgical debridement of necrotic tissue | 0
gauze dressing | 0
necrotizing fasciitis diagnosis | 0
fever | 12
necrotic tissue on wound margins | 12
second-look surgery | 12
aggressive surgical debridement | 12
handcrafted vacuum device | 12
NPWT | 12
intensive care unit | 12
drainage tube connected to central negative pressure system | 12
changing dressing twice a day | 12
irrigation with saline solution | 12
calcium alginate within the wound | 24
NPWT device installed | 48
free movement | 48
easily reinserted in society | 48
bacteriological examination | 48
antibiogram | 48
released from hospital | 48
ambulatory treatment | 48
methicillin-sensitive Staphylococcus aureus (MSSA) | 48
Clindamycin | 48
NPWT unit changed every four days | 48
NPWT unit changed every seven or ten days | 96
wound completely healed | 840
no skin graft or reconstruction surgery | 840
silicone scar sheet recommended | 840
follow-up outpatient | 1296