42 years old | 0
male | 0
transferred to intensive care unit | 0
acute necrotizing pancreatitis | 0
catheter-guided implantation of self-expanding nitinol stent | -336
portal vein thrombosis | -336
superior mesenteric artery thrombosis | -336
splenic artery thrombosis | -336
sigmoid colon perforation | -288
resection of sigmoid colon | -288
transversostoma application | -288
postoperative course uneventful | -264
extubated | -264
initial laboratory parameters improved | -216
increased white blood cell count | -72
increased C-reactive protein | -72
fever | -72
computed tomography on day 24 | 0
peripancreatic abscess | 0
left psoas muscle abscess | 0
computed tomography on day 37 | 312
CT-guided percutaneous catheter drainage | 408
drained brownish pus | 408
culture on Columbia blood agar | 408
culture on chocolate agar | 408
culture on MacConkey agar | 408
culture on Kimmig agar | 408
culture on ChromID Candida | 408
Candida albicans identified | 432
Bordetella hinzii identified | 432
deep skin swab sample positive for Bordetella hinzii | 432
intra-abdominal abscess no significant change | 456
Staphylococcus epidermidis detected | 456
Bordetella hinzii detected | 456
16S ribosomal RNA gene sequencing confirmed Bordetella hinzii | 456
antimicrobial susceptibility testing | 432
cefotaxime resistant | 432
levofloxacin resistant | 432
trimethoprim/sulfamethoxazole resistant | 432
piperacillin/tazobactam susceptible | 432
ceftazidime susceptible | 432
meropenem susceptible | 432
tigecycline susceptible | 432
empirical therapy with piperacillin/tazobactam initiated | 408
allergic skin reactions | 408
pruritus | 408
exanthema | 408
switched to meropenem | 408
allergic skin reactions to meropenem | 408
levofloxacin administered | 408
anaphylactic reaction | 408
hypotension | 408
tachycardia | 408
tigecycline initiated | 408
aspartate aminotransferase results available | 408
defervescence | 408
reduction of drained secretion | 408
intravenous tigecycline stopped | 408
whole genome sequencing performed | 432
no acquired antimicrobial resistance genes | 432
extensive alcohol abuse | 0
fatty liver disease | 0
