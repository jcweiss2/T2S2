 The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole or in part. The authors confirm that the images are original with no duplication and have not been previously published in whole