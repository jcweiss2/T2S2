54 years old | 0
    male | 0
    alcoholic cirrhosis (Child A) | 0
    diabetes mellitus | 0
    admitted | 0
    altered sensorium | -48
    fever | -48
    no headache | 0
    no vomiting | 0
    no seizures | 0
    no decreasing urine output | 0
    febrile | 0
    disoriented | 0
    pulse rate 100/min | 0
    blood pressure 150/70 mmHg | 0
    mild icterus | 0
    pedal edema | 0
    no focal neurological deficit | 0
    no signs of meningism | 0
    no papilledema | 0
    no retinitis | 0
    bilateral pupils equal | 0
    bilateral pupils reacting to light | 0
    free fluid | 0
    no organomegaly | 0
    Hb 9.6 gm/dL | 0
    total leukocyte count (TLC) 16 800/mm3 | 0
    normal eosinophil counts | 0
    platelet count 1.1 lac/mm3 | 0
    normal coagulation profile | 0
    INR 1.3 | 0
    serum bilirubin 3.0 mg/dL | 0
    AST 87 IU/L | 0
    ALT 96 IU/L | 0
    arterial ammonia 239 μg/dL | 0
    IgM anti-HEV positive | 0
    HBsAg negative | 0
    anti-HCV negative | 0
    IgM anti-HAV negative | 0
    HIV negative | 0
    high ascites | 0
    high serum, ascites albumin gradient | 0
    normal ascitic cell counts | 0
    ultrasonography abdomen suggestive of chronic liver disease | 0
    coarse echotexture | 0
    normal bilateral kidneys | 0
    normal renal functions | 0
    1+ proteinuria | 0
    full field leucocytes | 0
    8-10 RBC/high-power field on urine analysis | 0
    urine culture positive for enterococcus faecalis | 0
    sensitivity to linezolid only | 0
    altered sensorium persisted | 0
    hepatic encephalopathy | 0
    uro-sepsis | 0
    lactulose | 0
    supportive care for liver failure | 0
    linezolid 600 mg twice a day started | 0
    pruritus developed | 72
    erythematous macular rash developed | 72
    rash involving all extremities | 72
    rash involving trunk | 72
    peripheral blood smear showed eosinophilia | 72
    absolute eosinophil count 2125 cells/mm3 | 72
    serum IgE levels elevated (430 IU/mL) | 72
    2+ proteinuria | 72
    15-20 leukocytes | 72
    WBC casts | 72
    RBC casts | 72
    no eosinophils in urine | 72
    serum creatinine rose to 5.2 mg/dL | 72
    decreasing urine output | 72
    dialytic support required | 72
    DRESS syndrome diagnosed | 72
    linezolid stopped | 72
    rash subsided | 96
    fever subsided | 96
    renal functions remained deranged | 96
    hepatic encephalopathy recovered | 96
    liver functions improved | 96
    ANA negative | 96
    ANCA negative | 96
    normal complement levels | 96
    renal biopsy performed | 168
    normal glomeruli on light microscopy | 168
    interstitium edema | 168
    moderate inflammatory infiltrate | 168
    predominantly mononuclear cells | 168
    few eosinophils | 168
    proximal tubular dilatation | 168
    patchy tubular necrosis | 168
    birefringent oxalate crystals present in tubules | 168
    oxalate crystals present in interstitium | 168
    foreign body giant cell reaction | 168
    no granuloma formation | 168
    arterioles unremarkable | 168
    no vasculitis | 168
    no thrombosis | 168
    no immune complex deposition | 168
    acute tubulointerstitial nephritis diagnosed | 168
    prednisolone course for 2 weeks | 168
    serum creatinine decreased to 1.4 mg/dL | 336
    estimated creatinine clearance 56 mL/min | 336
    no deterioration in renal functions | 336