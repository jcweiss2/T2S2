52 years old | 0
female | 0
admitted for D10 neurofibroma excision | 0
pre-operative fasting (solid food) | -7
pre-operative fasting (clear water) | -2
uneventful laminectomy and tumor excision | 0
general anesthesia | 0
prone position | 0
surgery duration | 4
intraoperative fentanyl | 0
paracetamol administration | -0.5
reversal of neuromuscular blockade | 0
extubation | 0
shifted to PACU | 0
nausea | 0.5
abdominal pain | 0.5
agitation | 0.5
tachypnea | 0.5
dry mouth, tongue, lips | 0.5
hypotension | 0.5
tachycardia | 0.5
afebrile | 0.5
blood glucose 464 mg/dl | 0.5
ABG analysis (pH 7.12) | 0.5
high anion gap metabolic acidosis | 0.5
bicarbonate 8 mmol/L | 0.5
base deficit 18 | 0.5
AG 22 | 0.5
potassium 4.2 mmol/L | 0.5
sodium 132 mmol/L | 0.5
urinary glucose | 0.5
urinary ketones | 0.5
serum β-hydroxybutyrate 5.8 mmol/L | 0.5
DKA diagnosis | 0.5
fluid resuscitation (0.9% NS) | 0.5
insulin bolus 6 U | 0.5
continuous insulin infusion | 0.5
electrolyte correction | 0.5
serum amylase 210 U/L | 0.5
lipase 155 U/L | 0.5
resolution of ketoacidosis | 0.5
subcutaneous insulin initiation | 0.5
shifted to ward | 72
HbA1c 7.2% | 72
sterile blood cultures | 72
sterile urine cultures | 72
blood glucose normalization | 72
discharged | 168
pre-operative fasting (solid food) | -168
pre-operative fasting (clear water) | -120
