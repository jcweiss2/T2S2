62 years old | 0
female | 0
total abdominal hysterectomy | -18360
bilateral salpingo-oophorectomy | -18360
uterine fibroid | -18360
endometrial polyp | -18360
ovarian cyst | -18360
incisional hernia | -504
laparoscopic dual mesh repair | -504
abdominal pain | 0
abdominal wall tenderness | 0
erythema | 0
urinary bladder perforation | 0
subcutaneous collection | 0
calcification anterior bladder wall | 0
calcification collection | 0
surgical emphysema | 0
necrotizing fasciitis | 0
emergency debridement | 0
mesh erosion into urinary bladder | 0
vesico-cutaneous fistula | 0
urethral catheter insertion | 0
septic shock | 24
intensive care | 24
inotropic support | 24
mechanical ventilation | 24
sepsis improvement | 168
repeated debridement | 168
mesh removal | 168
urinary bladder defect repair | 168
abdominoplasty | 672
cystogram confirmed no leakage | 672
wound healing well | 672
- Total abdominal hysterectomy | -26280
Bilateral salpingo-oophorectomy | -26280
Uterine fibroid | -26280
Endometrial polyp | -26280
Ovarian cyst | -26280
Incisional hernia | -15120 (time of repair? Or earlier?)
Laparoscopic dual mesh repair | -15120
total abdominal hysterectomy | -26280
bilateral salpingo-oophorectomy | -26280
uterine fibroid | -26280
endometrial polyp | -26280
ovarian cyst | -26280
incisional hernia | -15120
laparoscopic dual mesh repair | -15120
