59 years old | 0
African American | 0
female | 0
admitted to the hospital | 0
altered mental status | -8
bizarre behavior | -8
slow irrational speech | -8
delusions | -8
abnormal movements | -8
somnolent | -8
headaches | -8
worsening dyspnea | -8
hypertension | -672
hyperlipidemia | -672
type 2 diabetes mellitus | -672
end-stage renal disease | -672
diabetes mellitus nephropathy | -672
amlodipine | -672
carvedilol | -672
lisinopril | -672
hydralazine | -672
isosorbide dinitrite | -672
insulin | -672
methadone | -672
restless | 0
stereotypical movement | 0
episodes of staring | 0
nonsensical involuntary movements | 0
disoriented | 0
incomprehensible sounds | 0
Glasgow Coma Scale 8/15 | 0
bibasilar rales | 0
nasogastric tube | 24
hydralazine | 24
labetalol | 24
hemodialysis | 24
severe agitation | 24
elevated BUN | 24
elevated creatinine | 24
cardiology consultation | 24
clonidine | 48
repeat CT scan | 120
cerebral spinal fluid studies | 120
electroencephalography | 216
levetiracetam | 216
more alert | 240
oriented | 240
followed verbal commands | 240
GCS improved | 240
lethargic | 288
febrile | 288
elevated white counts | 288
neutrophilia | 288
atelectatic changes | 288
intravenous meropenem | 288
acyclovir | 288
magnetic resonance imaging | 336
PRES diagnosis | 336
labetalol infusion | 336
blood pressure control | 336
repeat CSF viral panel PCR | 336
autoimmune encephalopathy markers | 336
acyclovir discontinued | 336
meropenem continued | 336
cultures negative | 336
leukocytosis resolved | 360
alert | 432
oriented | 432
obeying commands | 432
GCS 15/15 | 432
steady blood pressure | 432
hemodialysis sessions | 432
outpatient antihypertensive regimen | 432
counseled on adherence | 432
repeat MRI | 432
increased late subacute hemorrhage | 432
encephalomalacia | 432
discharged | 432
subacute rehabilitation facility | 432
modified Rankin scale 4 | 432
follow-up | 744
repeat MRI | 744
residual brain abnormalities | 744
long-term oral levetiracetam | 744