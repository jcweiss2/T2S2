72 years old | 0
male | 0
Caucasian | 0
current smoker | 0
admitted to the emergency department | 0
dysuria | 0
subjective fever | 0
mild confusion | 0
dizziness | 0
denied shortness of breath | 0
denied loss of consciousness | 0
foley catheter removal | -48
obstructive uropathy | -48
benign prostatic hyperplasia | -48
stage II chronic kidney disease | 0
multiple kidney stones | 0
status post lithotripsy | 0
road traffic accident | -131040
surgery | -131040
right hip osteoarthritis | 0
avascular necrosis | 0
status post replacement | 0
nonalcoholic | 0
denied illicit substance use | 0
mild fever | 0
tachycardia | 0
hypotension | 0
tachypnea | 0
bilateral edematous swelling | 0
normal arterial blood gases | 0
inspired oxygen fraction of 28% | 0
leukocyte count 15.9 × 103/μL | 0
neutrophils 85% | 0
hemoglobin 10.9 mg/dl | 0
normal hematologic and coagulation parameters | 0
serum bicarbonate 22 mEq/L | 0
creatinine 3.4 mg/dl | 0
blood urea nitrogen 39 mg/dl | 0
lactic acid 3.2 mg/dl | 0
normal serum chemistries | 0
normal liver function tests | 0
urinalysis positive for leukocyte esterase | 0
high white cell count | 0
normal electrocardiogram | 0
normal serum troponin levels | 0
septic shock suspected | 0
blood cultures ordered | 0
broad spectrum intravenous antibiotics started | 0
proper fluid replacement | 0
persistent hypotension | 0
central venous catheter placed | 0
high doses of intravenous norepinephrine | 0
bedside ultrasonography performed | 0
good cardiac contractility | 0
no intra-abdominal bleeding | 0
bilateral noncompressible femoral veins | 0
deep vein thrombosis suspected | 0
echocardiogram performed | 0
ejection fraction 60% | 0
normal right ventricular ejection fraction | 0
normal right ventricular dimensions | 0
computed tomography pulmonary embolism protocol negative | 0
bilateral nonobstructive renal stones | 0
stranding suspicious for small retroperitoneal hematoma | 0
re-evaluation of patient presentation | 0
IVC filter placement 15 years ago | -131040
obstructive shock secondary to IVC obstruction suspected | 0
venography performed | 0
almost complete occlusion of the IVC | 0
filling defects within the distal IVC | 0
bilateral common and external iliac veins | 0
common femoral veins compatible with thrombus | 0
hypertrophy of the collateral arising from the left common iliac vein | 0
mechanical thrombectomy performed | 24
350 mL thrombus removed | 24
unfractionated heparin started | 24
closely monitored | 24
stranding in the retroperitoneum considered edema | 24
hemoglobin did not drop | 24
discharged on Rivaroxaban | 72
no recurrence of thrombosis for 3 months | 216
IVC filter removal not recommended | 72
anticoagulation for life | 72