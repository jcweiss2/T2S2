100 years old | 0
male | 0
admitted to the hospital | 0
anterior neck swelling | 0
dysphagia | 0
muffled voice | 0
oral steroid for presumed lymphadenitis | -336
symptoms did not abate with the steroids | -336
unable to wear dentures | -336
only could swallow liquids | 0
hyperlipidemia | 0
benign prostatic hyperplasia | 0
hypertension | 0
no history of alcohol | 0
no history of tobacco | 0
no history of illicit drug use | 0
physical exam | 0
respiratory distress | 0
discomfort secondary to pain | 0
heart rate 89 beats/min | 0
blood pressure 131/81 mmHg | 0
oxygen saturation 94% on room air | 0
respiratory rate 18 breaths/min | 0
severely limited mouth-opening | 0
inter-incisor gap of 1 cm | 0
could not extend neck | 0
white blood count 28,000/ μL | 0
hemoglobin 12.1 g/dL | 0
platelet count 225,000/μL | 0
computerized tomography neck scan | 0
peripherally enhanced loculated fluid collection | 0
surrounding soft tissue edema | 0
resilient mass effect | 0
narrowing of oropharynx | 0
no significant lymphadenopathy | 0
dental caries | 0
lucency suggested dental abscess | 0
oral and maxillofacial surgeon notified | 0
surgical drainage of abscess | 0
airway secured with awake fiberoptic intubation | 0
denitrogenated with 100% oxygen | 0
glycopyrrolate administered | 0
nasal decongestant oxymetazoline administered | 0
topical lidocaine administered | 0
ketamine administered | 0
fiberoptic scope advanced through nares | 0
tracheal intubation successful | 0
7.5 mm cuffed endotracheal tube placed | 0
fentanyl administered | 0
propofol administered | 0
sevoflurane as anesthetic gas | 0
dexamethasone administered | 0
surgical procedure completed | 0
incision and drainage of abscess | 0
collection of cultures | 0
shifted to intensive care unit | 0
elective postoperative ventilation | 0
extubated successfully | 24
surgical cultures revealed Streptococcus viridans | 24
surgical cultures revealed Streptococcus intermedius | 24
discharged | 48