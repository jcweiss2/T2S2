60 years old | 0
female | 0
bipolar disorder | -672
hyperlipidemia | -672
osteoporosis | -672
renal stone | -672
water pipe smoker | -672
history of suicidal behavior | -672
admitted to the hospital | 0
dizziness | 0
drowsiness | 0
drug poisoning | 0
amphetamine in urine | 0
benzodiazepine in urine | 0
Glasgow Coma Scale score 11 | 0
Glasgow Coma Scale score decreased to 9 | 24
Glasgow Coma Scale score fell to 3 | 48
cardiac analysis | 24
right bundle branch block | 24
complete bundle branch block | 24
amphetamine overdose | 24
therapeutic hemodialysis | 48
severe abdominal distension | 72
lack of defecation | 72
absence of bowel sound | 72
abdominal-pelvic sonography | 72
multiloculated fluid collection | 72
GI perforation | 72
severe peritonitis | 72
laparotomy | 72
perforation of the stomach | 72
acute peritonitis | 72
bowel adhesion | 72
stomach perforation repair | 72
retro-gastric fluid collection | 72
sub-diaphragmatic fluid collection | 72
generalized peritonitis | 72
drainage | 72
gall bladder specimen | 72
severe acute or chronic acalculous cholecystitis | 72
focal mucosal necrosis | 72
severe constipation | 336
abdominal distention | 336
ascites | 336
edema | 336
second abdominal-pelvic sonography | 336
multicoated fluid collection | 336
septation | 336
second laparotomy | 336
sepsis | 336
disseminated intravascular coagulation | 336
increase in serum BUN | 336
increase in serum creatinine | 336
renal failure | 336
cardiorespiratory arrest | 336
patient death | 336
CMV infection | -672
CMV gastritis | 72
gastric ulceration | 72
foreign body-type giant cell reaction | 72
CMV immunoreactivity | 72
CMV DNA in gall bladder specimens | 72
CMV DNA in gastric wall biopsy | 72
amphetamine use | -672
amphetamine-induced toxicity | 0
immunosuppression | 0 
low immunity | 0