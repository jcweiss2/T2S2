36 years old | 0
male | 0
admitted to the hospital | 0
severe lower abdominal pain | 0
fever | 0
ulcerative colitis | -8760
mesalazine | -8760
abdominal tenderness | 0
mild abdominal muscle tension | 0
no percussion pain | 0
leukocytes:13.62×10^9/L | 0
neutrophils:90.10% | 0
c-reactive protein:176.50 mg/L | 0
glucose:10.6 mmol/L | 0
lactate:3.0 mmol/L | 0
prothrombin time 16.1S | 0
international normalized ratio 1.43 | 0
activated partial thromboplastin time 32.0S | 0
plasma fibrinogen 2.5 g/L | 0
calcitoninogen 8.967 ng/mL | 0
enlarged and abnormally thick spleen | 0
gastrointestinal perforation | 0
rehydration | 0
anti-infective treatment with imipenem cistatin | 0
emergency surgery | 12
pelvic abscess cavity | 12
dense adhesions | 12
omental necrosis | 12
intestinal wall edema | 12
thickened intestinal wall | 12
gray-white attachments | 12
appendix occluded and swollen with pus | 12
partial sigmoid resection | 12
pelvic-abdominal adhesion release | 12
incidental appendectomy | 12
pelvic abscess incision and drainage | 12
partial resection of the greater omentum | 12
temporary colostomy | 12
rupture of the sigmoid colon | 12
hemorrhage | 12
necrosis | 12
inflammatory cell infiltration | 12
inflammatory exudate | 12
granulation tissue | 12
glandular hyperplasia | 12
thrombosis | 12
negative cut margins | 12
enlarged spleen | 24
heterogeneous density | 24
large air shadow | 24
splenic abscess | 24
fever | 24
blood cultures | 24
imipenemcitabine | 24
ultrasound-guided puncture and drainage | 48
infection index | 48
platelet count | 48
prothrombin time | 48
coagulation routine | 48
hypoproteinemia | 72
coagulation | 72
splenectomy | 96
abdominal drainage | 96
splenic gangrene | 96
red-brown purulent effusion | 96
peripheral yellow-brown effusion | 96
yellow-brown pelvic effusion | 96
partial necrotic hemorrhage | 96
symptomatic treatment | 120
imaging and test indexes | 120
discharged | 168