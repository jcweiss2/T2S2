86 years old | 0
female | 0
nausea | -2
vomiting | -2
right upper quadrant abdominal pain | -2
coronary artery disease | 0
pulmonary hypertension | 0
mitral regurgitation | 0
atrial fibrillation | 0
chronic kidney disease | 0
tachycardic | 0
hypotensive | 0
right upper quadrant tenderness | 0
positive Murphy’s sign | 0
elevated liver enzymes | 0
alkaline phosphatase 387 U/L | 0
alanine aminotransferase 89 U/L | 0
aspartate aminotransferase 78 U/L | 0
total bilirubin 5.9 mg/dL | 0
direct fraction of 5.2 mg/dL | 0
elevated creatinine | 0
elevated white blood cell count | 0
normal lipase | 0
distended gallbladder | 0
cholelithiasis | 0
wall thickness of 3 mm | 0
14-mm dilated common bile duct | 0
sepsis | 0
acute cholecystitis | 0
choledocholithiasis | 0
acute kidney injury | 0
intravenous hydration | 2
empiric antibiotics | 2
endoscopic retrograde cholangiopancreatography | 4
obstructed cystic duct | 4
multiple CBD stones | 4
sphincterotomy | 4
10F x 9 cm plastic stent placement | 4
ultrasound-guided PC tube placement | 96
clinical condition improved | 96
discharged home | 96
multiple evaluations | 192
exchanges of the PC tube | 192
percutaneous cholangiograms | 192
patent cystic duct | 192
occluded biliary stent | 192
contrast reaching the duodenum | 192
another ERCP | 216
biliary stent removal | 216
CBD stones removal | 216
cholangioscope | 216
electrohydraulic lithotripsy | 216
10F X 7 cm plastic stent placement | 216
hybrid percutaneous-endoscopic technique | 432
cholecystostomy drain opening dilation | 432
28F sheath placement | 432
pediatric gastroscope advancement | 432
gallbladder visualization | 432
multiple stones identification | 432
lithotripsy | 432
gallstones removal | 432
Roth net | 432
retrieval basket | 432
sheath removal | 432
20F drainage catheter placement | 432
another ERCP | 672
biliary stent removal | 672
stone removal | 672
12-mm balloon | 672
percutaneous cholangiogram | 680
contrast flow into the duodenum | 680
no significant obstruction | 680
PC tube removal | 680
dilated PC site healed | 680
asymptomatic | 1152
asymptomatic | 2080