51 years old | 0
male | 0
admitted to the hospital | 0
chest tightness | -720
atrial fibrillation diagnosis | -720
moderate to severe mitral stenosis | -720
mild to moderate regurgitation | -720
mild aortic valve insufficiency | -720
mild tricuspid valve insufficiency | -720
decreased left ventricular function | -720
small amount of pericardial effusion | -720
diarrhoea | -720
anti-diarrhoea medication use | -720
temperature 36.5°C | 0
heart rate 91 bpm | 0
respiratory rate 15 cpm | 0
blood pressure 131/79 mmHg | 0
severe diastolic murmur in mitral region | 0
systolic murmur in tricuspid valve | 0
enlarged cardiac border | 0
slurred speech | 24
shallow left nasolabial fold | 24
grade 4 muscle strength in left limb | 24
acute cerebral infarction in right frontotemporal occipital lobe | 24
small amount of post-infarct blood leakage | 24
high fever 38.6°C | 216
heart rate 170 bpm | 216
blood pressure 90/60 mmHg | 216
respiratory rate 25 cpm | 216
white blood cell count 7010/mm3 | 216
85.6% neutrophils | 216
lactate level 2.8 mmol/L | 216
calcitonin level 0.98 Pg/L | 216
vegetation on anterior leaflet of mitral valve | 216
acute cerebral haemorrhage | 216
septic shock | 216
fluid replacement | 216
volume expansion | 216
norepinephrine 18 μg/min | 216
vancomycin 1 g q12h | 216
mitral bioprosthetic valve replacement | 216
tricuspid valvuloplasty | 216
radiofrequency ablation of atrial fibrillation | 216
left atrial auricular resection | 216
levosimendan 1 mg/h | 216
norepinephrine 24 μg/min | 216
warfarin 2.5 mg qd | 216
fever persisted | 240
levosimendan discontinued | 240
norepinephrine discontinued | 240
piperacillin tazobactam 4.5 g q8h | 240
vancomycin 1 g q12h | 240
fever resolved | 288
neutrophil percentage normalized | 288
blood cultures positive | 240
blood cultures negative | 408
discharged | 408
asymptomatic at follow-up | 1464
normal biologic valve function | 1464
no abnormal echogenicity | 1464
