59 years old | 0
male | 0
admitted to the hospital | 0
chronic hepatitis B viral infection | 0
cirrhosis | 0
hypertension | 0
liver mass | 0
hepatocellular carcinoma | 0
non-tumorous portal vein thrombosis | 0
MELD score 18 | 0
living related liver transplant | 0
extended right lobe graft | 0
compatible blood group | 0
no anatomical variation | 0
right hepatic vein reconstruction | 0
middle hepatic vein reconstruction | 0
portal vein thromboendovenectomy | 0
right lobe graft anastomosed to inferior vena cava | 0
right lobe graft anastomosed to portal vein | 0
intra-operative portal vein anastomosis balloon dilatation | 0
stent placement | 0
right hepatic artery anastomosed to common hepatic artery | 0
hepaticojejunostomy | 0
extubated | 48
transferred from intensive care unit | 72
AST level decreased | 72
ALT level decreased | 72
general clinical condition improved | 72
hypertension | 216
sudden chest pain | 216
collapsed | 216
cardio-pulmonary resuscitation | 216
spontaneous circulation returned | 216
aortic dissection Stanford A | 216
ascending aortic replacement | 216
circulatory arrest | 216
clinical condition improved | 240
liver function improved | 240
intra-abdominal collection | 240
biliary leakage | 240
sepsis | 240
massive upper gastrointestinal hemorrhage | 984
hemodynamic unstable | 984
gastro-duodeno scope | 984
massive bleeding from duodenum | 984
angiogram | 984
bleeding from pseudoaneurysm of gastroduodenal artery | 984
thromboses of hepatic artery proper | 984
coil embolization | 984
bleeding stopped | 984
vital signs returned to normal | 984
liver function worsened | 984
re-operate | 1008
re-anastomose hepatic artery inflow | 1008
extensively thrombosed | 1008
portal vein arterialization | 1008
common hepatic artery connected to splenic vein | 1008
liver function improved | 1032
no deceased donor | 1032
another massive upper gastrointestinal hemorrhage | 1232
bleeding from portal hypertensive gastropathy | 1232
embolization | 1232
unnamed vein embolization | 1232
splenic artery embolization | 1232
died | 1368
recurrent upper gastrointestinal hemorrhage | 1368
uncontrolled intra-abdominal sepsis | 1368
liver abscess | 1368