55 years old | 0
male | 0
admitted to the hospital | 0
malaise | -336
fever | -336
weakness | -336
weight loss | -336
sore throat | -336
dry cough | -336
distant history of stab wounds | -10080
splenectomy | -10080
denies tick bites | -336
febrile | 0
tachypneic | 0
tachycardic | 0
jaundice | 0
acute renal injury | 0
elevated creatinine | 0
mild liver injury | 0
elevated INR | 0
mixed hyperbilirubinemia | 0
elevated lactate dehydrogenase | 0
undetectable haptoglobin | 0
intracellular parasites | 0
parasitemia | 0
B. microti detected by PCR | 0
fulminant babesiosis infection | 0
multi-organ systemic failure | 0
Atovaquone treatment | 0
azithromycin treatment | 0
transferred to medical intensive care unit | 0
positive c-ANCA | 24
positive ANA | 24
low complement levels | 24
exchange transfusions | 24
parasitemia level dropped | 48
clinical status improved | 48
laboratory parameters improved | 48
discharged | 168
follow up | 1440
resolution of parasitemia | 1440
creatinine level improved | 1440
c-ANCA level negative | 1440