84 years old | 0
    female | 0
    Caucasian | 0
    generalized abdominal pain | -48
    vomiting | -48
    diarrhea | -48
    no prior symptoms | -48
    afebrile prior to presentation | -48
    altered general status | 0
    respiratory distress | 0
    tachypneic | 0
    use of accessory muscles | 0
    febrile | 0
    tachycardic | 0
    tachypneic | 0
    desaturation | 0
    hypotensive | 0
    primary metabolic acidosis | 0
    anion gap | 0
    oxygen saturation increased | 0
    hydration | 0
    systolic blood pressure increased | 0
    right upper quadrant tenderness | 0
    positive Murphy’s sign | 0
    blood cultures taken | 0
    urine cultures taken | 0
    Amikacin | 0
    Vancomycin | 0
    Tazocin | 0
    COVID-19 PCR negative | 0
    elevated C-reactive protein | 0
    elevated lactate dehydrogenase | 0
    elevated ferritin | 0
    elevated fibrinogen | 0
    elevated erythrocyte sedimentation rate | 0
    lymphopenic | 0
    elevated amylase | 0
    elevated bilirubin | 0
    normal aspartate aminotransferase | 0
    normal alanine aminotransferase | 0
    CT chest-abdomen-pelvis | 0
    patchy consolidations | 0
    air bronchograms | 0
    ground glass opacities | 0
    COVID-19 pneumonia | 0
    gallbladder distended | 0
    enhancing wall | 0
    focal defects | 0
    fat stranding | 0
    peri-vesicular fluid | 0
    pericholecystic abscesses | 0
    acute ischemic gangrenous cholecystitis | 0
    scheduled for percutaneous drainage | 0
    repeat COVID-19 PCR | 0
    hypotensive again | 0
    refractory to IV fluids | 0
    Dopamine | 0
    systolic blood pressure elevated | 0
    deteriorated | 24
    hypotensive | 24
    desaturated | 24
    double oxygen source | 24
    non-rebreather face mask | 24
    nasal cannula high flow oxygen | 24
    saturation did not improve | 24
    remained hypotensive | 24
    intubated | 24
    cardio-pulmonary arrest | 24
    resuscitation failed | 24
    pronounced dead | 24
    repeat PCR positive | 24
    blood cultures negative | 24
    urine culture negative | 24
    