46 years old | 0 | 0 
female | 0 | 0 
obesity | 0 | 0 
psoriatic arthritis | 0 | 0 
hypoparathyroidism | -7200 | 0 
hypothyroidism | -7200 | 0 
total thyroidectomy | -7200 | -7200 
multinodular goitre | -7200 | -7200 
elective sleeve gastrectomy | 0 | 0 
gastric perforations | 0 | 0 
friable mucosa | 0 | 0 
abdominal sepsis | 4 | 4 
transfer to intensive care | 4 | 4 
critically low calcium level | 4 | 4 
intravenous calcium gluconate infusion | 4 | 192 
normocalcaemia | 4 | 192 
prolonged ICU admission | 4 | 192 
abdominal operations | 4 | 192 
weight loss | 4 | 192 
Endocrinology advice | 14 | 192 
hypothyroidism management | 14 | 192 
intravenous triiodothyronine | 14 | 192 
euthyroidism | 14 | 192 
high dose intravenous calcium | 14 | 192 
ionised calcium measurement | 14 | 192 
serum phosphate level | 14 | 192 
intravenous calcitriol | 42 | 47 
limited stock | 47 | 47 
high cost | 47 | 47 
intramuscular cholecalciferol | 56 | 56 
low 1,25(OH)vitamin D3 level | 56 | 79 
normal renal function | 56 | 192 
eGFR > 90 mL/min/1.73 m2 | 56 | 192 
reduced calcium gluconate requirements | 84 | 192 
intravenous thyroxine | 88 | 192 
maintenance schedule | 88 | 192 
discharge | 192 | 192 
oral intake | 192 | 192 
normocalcaemia | 192 | 288 
follow-up | 288 | 288 
weight | 288 | 288 
BMI | 288 | 288 
calcium replacement | 0 | 192 
parenteral treatment | 0 | 192 
hypoparathyroidism management | 0 | 192 
elective bariatric surgery | 0 | 0 
complications | 0 | 192 
difficulties in managing hypocalcaemia | 0 | 192 
impaired gastrointestinal absorption | 0 | 192 
subcutaneous recombinant PTH | 0 | 0 
approval | 0 | 0 
future management | 0 | 0 
research | 0 | 0 
funding | 0 | 0 
author contribution | 0 | 0 
declaration of interest | 0 | 0 
conflict of interest | 0 | 0 
impartiality | 0 | 0 
clinical care | 0 | 192 
writing of manuscript | 0 | 192 
surgical hypoparathyroidism | -7200 | 0 
parathyroidectomy | -7200 | -7200 
bariatric surgery | 0 | 192 
gastrointestinal disorders | 0 | 192 
malabsorption | 0 | 192 
international guidelines | 0 | 0 
recommendation | 0 | 0 
use of PTH 1–84 | 0 | 0 
government subsidised | 0 | 0 
Australian Register of Therapeutic Goods | 0 | 0 
enteral absorption | 0 | 192 
calcium and calcitriol | 0 | 192 
gastrostomy tube insertion | 0 | 0 
pancreatic enzyme supplementation | 0 | 0 
abdominal sepsis | 4 | 4 
friable mucosa | 0 | 0 
gastric bypass surgery | 0 | 0 
pre-existing hypoparathyroidism | 0 | 0 
hypocalcaemia management | 0 | 192 
potential difficulties | 0 | 0 
approval of subcutaneous recombinant PTH | 0 | 0 
hypoparathyroidism in Australia | 0 | 0 
future management | 0 | 0 
elective bariatric surgery | 0 | 0 
patients with pre-existing hypoparathyroidism | 0 | 0 
careful consideration | 0 | 0 
hypocalcaemia | 4 | 192 
impaired gastrointestinal absorption | 0 | 192 
complications | 0 | 192 
subcutaneous recombinant PTH | 0 | 0 
hypoparathyroidism management | 0 | 192 
parenteral treatment | 0 | 192 
calcium replacement | 0 | 192 
intravenous calcium gluconate | 4 | 192 
intravenous calcitriol | 42 | 192 
intramuscular cholecalciferol | 56 | 56 
intravenous thyroxine | 88 | 192 
maintenance schedule | 88 | 192 
discharge | 192 | 192 
follow-up | 288 | 288 
weight | 288 | 288 
BMI | 288 | 288 
normocalcaemia | 192 | 288 
oral intake | 192 | 192 
hypoparathyroidism | -7200 | 0 
hypothyroidism | -7200 | 0 
total thyroidectomy | -7200 | -7200 
multinodular goitre | -7200 | -7200 
elective sleeve gastrectomy | 0 | 0 
gastric perforations | 0 | 0 
friable mucosa | 0 | 0 
abdominal sepsis | 4 | 4 
transfer to intensive care | 4 | 4 
critically low calcium level | 4 | 4 
intravenous calcium gluconate infusion | 4 | 192 
normocalcaemia | 4 | 192 
prolonged ICU admission | 4 | 192 
abdominal operations | 4 | 192 
weight loss | 4 | 192 
Endocrinology advice | 14 | 192 
hypothyroidism management | 14 | 192 
intravenous triiodothyronine | 14 | 192 
euthyroidism | 14 | 192 
high dose intravenous calcium | 14 | 192 
ionised calcium measurement | 14 | 192 
serum phosphate level | 14 | 192 
intravenous calcitriol | 42 | 47 
limited stock | 47 | 47 
high cost | 47 | 47 
intramuscular cholecalciferol | 56 | 56 
low 1,25(OH)vitamin D3 level | 56 | 79 
normal renal function | 56 | 192 
eGFR > 90 mL/min/1.73 m2 | 56 | 192 
reduced calcium gluconate requirements | 84 | 192 
intravenous thyroxine | 88 | 192 
maintenance schedule | 88 | 192 
discharge | 192 | 192 
oral intake | 192 | 192 
normocalcaemia | 192 | 288 
follow-up | 288 | 288 
weight | 288 | 288 
BMI | 288 | 288 
calcium replacement | 0 | 192 
parenteral treatment | 0 | 192 
hypoparathyroidism management | 0 | 192 
elective bariatric surgery | 0 | 0 
complications | 0 | 192 
difficulties in managing hypocalcaemia | 0 | 192 
impaired gastrointestinal absorption | 0 | 192 
subcutaneous recombinant PTH | 0 | 0 
approval | 0 | 0 
future management | 0 | 0 
research | 0 | 0 
funding | 0 | 0 
author contribution | 0 | 192 
declaration of interest | 0 | 0 
conflict of interest | 0 | 0 
impartiality | 0 | 0 
clinical care | 0 | 192 
writing of manuscript | 0 | 192 
surgical hypoparathyroidism | -7200 | 0 
parathyroidectomy | -7200 | -7200 
bariatric surgery | 0 | 192 
gastrointestinal disorders | 0 | 192 
malabsorption | 0 | 192 
international guidelines | 0 | 0 
recommendation | 0 | 0 
use of PTH 1–84 | 0 | 0 
government subsidised | 0 | 0 
Australian Register of Therapeutic Goods | 0 | 0 
enteral absorption | 0 | 192 
calcium and calcitriol | 0 | 192 
gastrostomy tube insertion | 0 | 0 
pancreatic enzyme supplementation | 0 | 0 
abdominal sepsis | 4 | 4 
friable mucosa | 0 | 0 
gastric bypass surgery | 0 | 0 
pre-existing hypoparathyroidism | 0 | 0 
hypocalcaemia management | 0 | 192 
potential difficulties | 0 | 0 
approval of subcutaneous recombinant PTH | 0 | 0 
hypoparathyroidism in Australia | 0 | 0 
future management | 0 | 0 
elective bariatric surgery | 0 | 0 
patients with pre-existing hypoparathyroidism | 0 | 0 
careful consideration | 0 | 0 
hypocalcaemia | 4 | 192 
impaired gastrointestinal absorption | 0 | 192 
complications | 0 | 192 
subcutaneous recombinant PTH | 0 | 0 
hypoparathyroidism management | 0 | 192 
parenteral treatment | 0 | 192 
calcium replacement | 0 | 192 
intravenous calcium gluconate | 4 | 192 
intravenous calcitriol | 42 | 192 
intramuscular cholecalciferol | 56 | 56 
intravenous thyroxine | 88 | 192 
maintenance schedule | 88 | 192 
discharge | 192 | 192 
follow-up | 288 | 288 
weight | 288 | 288 
BMI | 288 | 288 
normocalcaemia | 192 | 288 
oral intake | 192 | 192 
hypoparathyroidism | -7200 | 0 
hypothyroidism | -7200 | 0 
total thyroidectomy | -7200 | -7200 
multinodular goitre | -7200 | -7200 
elective sleeve gastrectomy | 0 | 0 
gastric perforations | 0 | 0 
friable mucosa | 0 | 0 
abdominal sepsis | 4 | 4 
transfer to intensive care | 4 | 4 
critically low calcium level | 4 | 4 
intravenous calcium gluconate infusion | 4 | 192 
normocalcaemia | 4 | 192 
prolonged ICU admission | 4 | 192 
abdominal operations | 4 | 192 
weight loss | 4 | 192 
Endocrinology advice | 14 | 192 
hypothyroidism management | 14 | 192 
intravenous triiodothyronine | 14 | 192 
euthyroidism | 14 | 192 
high dose intravenous calcium | 14 | 192 
ionised calcium measurement | 14 | 192 
serum phosphate level | 14 | 192 
intravenous calcitriol | 42 | 47 
limited stock | 47 | 47 
high cost | 47 | 47 
intramuscular cholecalciferol | 56 | 56 
low 1,25(OH)vitamin D3 level | 56 | 79 
normal renal function | 56 | 192 
eGFR > 90 mL/min/1.73 m2 | 56 | 192 
reduced calcium gluconate requirements | 84 | 192 
intravenous thyroxine | 88 | 192 
maintenance schedule | 88 | 192 
discharge | 192 | 192 
oral intake | 192 | 192 
normocalcaemia | 192 | 288 
follow-up | 288 | 288 
weight | 288 | 288 
BMI | 288 | 288 
calcium replacement | 0 | 192 
parenteral treatment | 0 | 192 
hypoparathyroidism management | 0 | 192 
elective bariatric surgery | 0 | 0 
complications | 0 | 192 
difficulties in managing hypocalcaemia | 0 | 192 
impaired gastrointestinal absorption | 0 | 192 
subcutaneous recombinant PTH | 0 | 0 
approval | 0 | 0 
future management | 0 | 0 
research | 0 | 0 
funding | 0 | 0 
author contribution | 0 | 192 
declaration of interest | 0 | 0 
conflict of interest | 0 | 0 
impartiality | 0 | 0 
clinical care | 0 | 192 
writing of manuscript | 0 | 192 
surgical hypoparathyroidism | -7200 | 0 
parathyroidectomy | -7200 | -7200 
bariatric surgery | 0 | 192 
gastrointestinal disorders | 0 | 192 
malabsorption | 0 | 192 
international guidelines | 0 | 0 
recommendation | 0 | 0 
use of PTH 1–84 | 0 | 0 
government subsidised | 0 | 0 
Australian Register of Therapeutic Goods | 0 | 0 
enteral absorption | 0 | 192 
calcium and calcitriol | 0 | 192 
gastrostomy tube insertion | 0 | 0 
pancreatic enzyme supplementation | 0 | 0 
abdominal sepsis | 4 | 4 
friable mucosa | 0 | 0 
gastric bypass surgery | 0 | 0 
pre-existing hypoparathyroidism | 0 | 0 
hypocalcaemia management | 0 | 192 
potential difficulties | 0 | 0 
approval of subcutaneous recombinant PTH | 0 | 0 
hypoparathyroidism in Australia | 0 | 0 
future management | 0 | 0 
elective bariatric surgery | 0 | 0 
patients with pre-existing hypoparathyroidism | 0 | 0 
careful consideration | 0 | 0 
hypocalcaemia | 4 | 192 
impaired gastrointestinal absorption | 0 | 192 
complications | 0 | 192 
subcutaneous recombinant PTH | 0 | 0 
hypoparathyroidism management | 0 | 192 
parenteral treatment | 0 | 192 
calcium replacement | 0 | 192 
intravenous calcium gluconate | 4 | 192 
intravenous calcitriol | 42 | 192 
intramuscular cholecalciferol | 56 | 56 
intravenous thyroxine | 88 | 192 
maintenance schedule | 88 | 192 
discharge | 192 | 192 
follow-up | 288 | 288 
weight | 288 | 288 
BMI | 288 | 288 
normocalcaemia | 192 | 288 
oral intake | 192 | 192 
hypoparathyroidism | -7200 | 0 
hypothyroidism | -7200 | 0 
total thyroidectomy | -7200 | -7200 
multinodular goitre | -7200 | -7200 
elective sleeve gastrectomy | 0 | 0 
gastric perforations | 0 | 0 
friable mucosa | 0 | 0 
abdominal sepsis | 4 | 4 
transfer to intensive care | 4 | 4 
critically low calcium level | 4 | 4 
intravenous calcium gluconate infusion | 4 | 192 
normocalcaemia | 4 | 192 
prolonged ICU admission | 4 | 192 
abdominal operations | 4 | 192 
weight loss | 4 | 192 
Endocrinology advice | 14 | 192 
hypothyroidism management | 14 | 192 
intravenous triiodothyronine | 14 | 192 
euthyroidism | 14 | 192 
high dose intravenous calcium | 14 | 192 
ionised calcium measurement | 14 | 192 
serum phosphate level | 14 | 192 
intravenous calcitriol | 42 | 47 
limited stock | 47 | 47 
high cost | 47 | 47 
intramuscular cholecalciferol | 56 | 56 
low 1,25(OH)vitamin D3 level | 56 | 79 
normal renal function | 56 | 192 
eGFR > 90 mL/min/1.73 m2 | 56 | 192 
reduced calcium gluconate requirements | 84 | 192 
intravenous thyroxine | 88 | 192 
maintenance schedule | 88 | 192 
discharge | 192 | 192 
oral intake | 192 | 192 
normocalcaemia | 192 | 288 
follow-up | 288 | 288 
weight | 288 | 288 
BMI | 288 | 288 
calcium replacement | 0 | 192 
parenteral treatment | 0 | 192 
hypoparathyroidism management | 0 | 192 
elective bariatric surgery | 0 | 0 
complications | 0 | 192 
difficulties in managing hypocalcaemia | 0 | 192 
impaired gastrointestinal absorption | 0 | 192 
subcutaneous recombinant PTH | 0 | 0 
approval | 0 | 0 
future management | 0 | 0 
research | 0 | 0 
funding | 0 | 0 
author contribution | 0 | 192 
declaration of interest | 0 | 0 
conflict of interest | 0 | 0 
impartiality | 0 | 0 
clinical care | 0 | 192 
writing of manuscript | 0 | 192 
surgical hypoparathyroidism | -7200 | 0 
parathyroidectomy | -7200 | -7200 
bariatric surgery | 0 | 192 
gastrointestinal disorders | 0 | 192 
malabsorption | 0 | 192 
international guidelines | 0 | 0 
recommendation | 0 | 0 
use of PTH 1–84 | 0 | 0 
government subsidised | 0 | 0 
Australian Register of Therapeutic Goods | 0 | 0 
enteral absorption | 0 | 192 
calcium and calcitriol | 0 | 192 
gastrostomy tube insertion | 0 | 0 
pancreatic enzyme supplementation | 0 | 0 
abdominal sepsis | 4 | 4 
friable mucosa | 0 | 0 
gastric bypass surgery | 0 | 0 
pre-existing hypoparathyroidism | 0 | 0 
hypocalcaemia management | 0 | 192 
potential difficulties | 0 | 0 
approval of subcutaneous recombinant PTH | 0 | 0 
hypoparathyroidism in Australia | 0 | 0 
future management | 0 | 0 
elective bariatric surgery | 0 | 0 
patients with pre-existing hypoparathyroidism | 0 | 0 
careful consideration | 0 | 0 
hypocalcaemia | 4 | 192 
impaired gastrointestinal absorption | 0 | 192 
complications | 0 | 192 
subcutaneous recombinant PTH | 0 | 0 
hypoparathyroidism management | 0 | 192 
parenteral treatment | 0 | 192 
calcium replacement | 0 | 192 
intravenous calcium gluconate | 4 | 192 
intravenous calcitriol | 42 | 192 
intramuscular cholecalciferol | 56 | 56 
intravenous thyroxine | 88 | 192 
maintenance schedule | 88 | 192 
discharge | 192 | 192 
follow-up | 288 | 288 
weight | 288 | 288 
BMI | 288 | 288 
normocalcaemia | 192 | 288 
oral intake | 192 | 192 
hypoparathyroidism | -7200 | 0 
hypothyroidism | -7200 | 0 
total thyroidectomy | -7200 | -7200 
multinodular goitre | -7200 | -7200 
elective sleeve gastrectomy | 0 | 0 
gastric perforations | 0 | 0 
friable mucosa | 0 | 0 
abdominal sepsis | 4 | 4 
transfer to intensive care | 4 | 4 
critically low calcium level | 4 | 4 
intravenous calcium gluconate infusion | 4 | 192 
normocalcaemia | 4 | 192 
prolonged ICU admission | 4 | 192 
abdominal operations | 4 | 192 
weight loss | 4 | 192 
Endocrinology advice | 14 | 192 
hypothyroidism management | 14 | 192 
intravenous triiodothyronine | 14 | 192 
euthyroidism | 14 | 192 
high dose intravenous calcium | 14 | 192 
ionised calcium measurement | 14 | 192 
serum phosphate level | 14 | 192 
intravenous calcitriol | 42 | 47 
limited stock | 47 | 47 
high cost | 47 | 47 
intramuscular cholecalciferol | 56 | 56 
low 1,25(OH)vitamin D3 level | 56 | 79 
normal renal function | 56 | 192 
eGFR > 90 mL/min/1.73 m2 | 56 | 192 
reduced calcium gluconate requirements | 84 | 192 
intravenous thyroxine | 88 | 192 
maintenance schedule | 88 | 192 
discharge | 192 | 192 
oral intake | 192 | 192 
normocalcaemia | 192 | 288 
follow-up | 288 | 288 
weight | 288 | 288 
BMI | 288 | 288 
calcium replacement | 0 | 192 
parenteral treatment | 0 | 192 
hypoparathyroidism management | 0 | 192 
elective bariatric surgery | 0 | 0 
complications | 0 | 192 
difficulties in managing hypocalcaemia | 0 | 192 
impaired gastrointestinal absorption | 0 | 192 
subcutaneous recombinant PTH | 0 | 0 
approval | 0 | 0 
future management | 0 | 0 
research | 0 | 0 
funding | 0 | 0 
author contribution | 0 | 192 
declaration of interest | 0 | 0 
conflict of interest | 0 | 0 
impartiality | 0 | 0 
clinical care | 0 | 192 
writing of manuscript | 0 | 192 
surgical hypoparathyroidism | -7200 | 0 
parathyroidectomy | -7200 | -7200 
bariatric surgery | 0 | 192 
gastrointestinal disorders | 0 | 192 
malabsorption | 0 | 192 
international guidelines | 0 | 0 
recommendation | 0 | 0 
use of PTH 1–84 | 0 | 0 
government subsidised | 0 | 0 
Australian Register of Therapeutic Goods | 0 | 0 
enteral absorption | 0 | 192 
calcium and calcitriol | 0 | 192 
gastrostomy tube insertion | 0 | 0 
pancreatic enzyme supplementation | 0 | 0 
abdominal sepsis | 4 | 4 
friable mucosa | 0 | 0 
gastric bypass surgery | 0 | 0 
pre-existing hypoparathyroidism | 0 | 0 
hypocalcaemia management | 0 | 192 
potential difficulties | 0 | 0 
approval of subcutaneous recombinant PTH | 0 | 0 
hypoparathyroidism in Australia | 0 | 0 
future management | 0 | 0 
elective bariatric surgery | 0 | 0 
patients with pre-existing hypoparathyroidism | 0 | 0 
careful consideration | 0 | 0 
hypocalcaemia | 4 | 192 
impaired gastrointestinal absorption | 0 | 192 
complications | 0 | 192 
subcutaneous recombinant PTH | 0 | 0 
hypoparathyroidism management | 0 | 192 
parenteral treatment | 0 | 192 
calcium replacement | 0 | 192 
intravenous calcium gluconate | 4 | 192 
intravenous calcitriol | 42 | 192 
intramuscular cholecalciferol | 56 | 56 
intravenous thyroxine | 88 | 192 
maintenance schedule | 88 | 192 
discharge | 192 | 192 
follow-up | 288 | 288 
weight | 288 | 288 
BMI | 288 | 288 
normocalcaemia | 192 | 288 
oral intake | 192 | 192 
hypoparathyroidism | -7200 | 0 
hypothyroidism | -7200 | 0 
total thyroidectomy | -7200 | -7200 
multinodular goitre | -7200 | -7200 
elective sleeve gastrectomy | 0 | 0 
gastric perforations | 0 | 0 
friable mucosa | 0 | 0 
abdominal sepsis | 4 | 4 
transfer to intensive care | 4 | 4 
critically low calcium level | 4 | 4 
intravenous calcium gluconate infusion | 4 | 192 
normocalcaemia | 4 | 192 
prolonged ICU admission | 4 | 192 
abdominal operations | 4 | 192 
weight loss | 4 | 192 
Endocrinology advice | 14 | 192 
hypothyroidism management | 14 | 192 
intravenous triiodothyronine | 14 | 192 
euthyroidism | 14 | 192 
high dose intravenous calcium | 14 | 192 
ionised calcium measurement | 14 | 192 
serum phosphate level | 14 | 192 
intravenous calcitriol | 42 | 47 
limited stock | 47 | 47 
high cost | 47 | 47 
intramuscular cholecalciferol | 56 | 56 
low 1,25(OH)vitamin D3 level | 56 | 79 
normal renal function | 56 | 192 
eGFR > 90 mL/min/1.73 m2 | 56 | 192 
reduced calcium gluconate requirements | 84 | 192 
intravenous thyroxine | 88 | 192 
maintenance schedule | 88 | 192 
discharge | 192 | 192 
oral intake | 192 | 192 
normocalcaemia | 192 | 288 
follow-up | 288 | 288 
weight | 288 | 288 
BMI | 288 | 288 
calcium replacement | 0 | 192 
parenteral treatment | 0 | 192 
hypoparathyroidism management | 0 | 192 
elective bariatric surgery | 0 | 0 
complications | 0 | 192 
difficulties in managing hypocalcaemia | 0 | 192 
impaired gastrointestinal absorption | 0 | 192 
subcutaneous recombinant PTH | 0 | 0 
approval | 0 | 0 
future management | 0 | 0 
research | 0 | 0 
funding | 0 | 0 
author contribution | 0 | 192 
declaration of interest | 0 | 0 
conflict of interest | 0 | 0 
impartiality | 0 | 0 
clinical care | 0 | 192 
writing of manuscript | 0 | 192 
surgical hypoparathyroidism | -7200 | 0 
parathyroidectomy | -7200 | -7200 
bariatric surgery | 0 | 192 
gastrointestinal disorders | 0 | 192 
malabsorption | 0 | 192 
international guidelines | 0 | 0 
recommendation | 0 | 0 
use of PTH 1–84 | 0 | 0 
government subsidised | 0 | 0 
Australian Register of Therapeutic Goods | 0 | 0 
enteral absorption | 0 | 192 
calcium and calcitriol | 0 | 192 
gastrostomy tube insertion | 0 | 0 
pancreatic enzyme supplementation | 0 | 0 
abdominal sepsis | 4 | 4 
friable mucosa | 0 | 0 
gastric bypass surgery | 0 | 0 
pre-existing hypoparathyroidism | 0 | 0 
hypocalcaemia management | 0 | 192 
potential difficulties | 0 | 0 
approval of subcutaneous recombinant PTH | 0 | 0 
hypoparathyroidism in Australia | 0 | 0 
future management | 0 | 0 
elective bariatric surgery | 0 | 0 
patients with pre-existing hypoparathyroidism | 0 | 0 
careful consideration | 0 | 0 
hypocalcaemia | 4 | 192 
impaired gastrointestinal absorption | 0 | 192 
complications | 0 | 192 
subcutaneous recombinant PTH | 0 | 0 
hypoparathyroidism management | 0 | 192 
parenteral treatment | 0 | 192 
calcium replacement | 0 | 192 
intravenous calcium gluconate | 4 | 192 
intravenous calcitriol | 42 | 192 
intramuscular cholecalciferol | 56 | 56 
intravenous thyroxine | 88 | 192 
maintenance schedule | 88 | 192 
discharge | 192 | 192 
follow-up | 288 | 288 
weight | 288 | 288 
BMI | 288 | 288 
normocalcaemia | 192 | 288 
oral intake | 192 | 192 
hypoparathyroidism | -7200 | 0 
hypothyroidism | -7200 | 0 
total thyroidectomy | -7200 | -7200 
multinodular goitre | -7200 | -7200 
elective sleeve gastrectomy | 0 | 0 
gastric perforations | 0 | 0 
friable mucosa | 0 | 0 
abdominal sepsis | 4 | 4 
transfer to intensive care | 4 | 4 
critically low calcium level | 4 | 4 
intravenous calcium gluconate infusion | 4 | 192 
normocalcaemia | 4 | 192 
prolonged ICU admission | 4 | 192 
abdominal operations | 4 | 192 
weight loss | 4 | 192 
Endocrinology advice | 14 | 192 
hypothyroidism management | 14 | 192 
intravenous triiodothyronine | 14 | 192 
euthyroidism | 14 | 192 
high dose intravenous calcium | 14 | 192 
ionised calcium measurement | 14 | 192 
serum phosphate level | 14 | 192 
intravenous calcitriol | 42 | 47 
limited stock | 47 | 47 
high cost | 47 | 47 
intramuscular cholecalciferol | 56 | 56 
low 1,25(OH)vitamin D3 level | 56 | 79 
normal renal function | 56 | 192 
eGFR > 90 mL/min/1.73 m2 | 56 | 192 
reduced calcium gluconate requirements | 84 | 192 
intravenous thyroxine | 88 | 192 
maintenance schedule | 88 | 192 
discharge | 192 | 192 
oral intake | 192 | 192 
normocalcaemia | 192 | 288 
follow-up | 288 | 288 
weight | 288 | 288 
BMI | 288 | 288 
calcium replacement | 0 | 192 
parenteral treatment | 0 | 192 
hypoparathyroidism management | 0 | 192 
elective bariatric surgery | 0 | 0 
complications | 0 | 192 
difficulties in managing hypocalcaemia | 0 | 192 
impaired gastrointestinal absorption | 0 | 192 
subcutaneous recombinant PTH | 0 | 0 
approval | 0 | 0 
future management | 0 | 0 
research | 0 | 0 
funding | 0 | 0 
author contribution | 0 | 192 
declaration of interest | 0 | 0 
conflict of interest | 0 | 0 
impartiality | 0 | 0 
clinical care | 0 | 192 
writing of manuscript | 0 | 192 
surgical hypoparathyroidism | -7200 | 0 
parathyroidectomy | -7200 | -7200 
bariatric surgery | 0 | 192 
gastrointestinal disorders | 0 | 192 
malabsorption | 0 | 192 
international guidelines | 0 | 0 
recommendation | 0 | 0 
use of PTH 1–84 | 0 | 0 
government subsidised | 0 | 0 
Australian Register of Therapeutic Goods | 0 | 0 
enteral absorption | 0 | 192 
calcium and calcitriol | 0 | 192 
gastrostomy tube insertion | 0 | 0 
pancreatic enzyme supplementation | 0 | 0 
abdominal sepsis | 4 | 4 
friable mucosa | 0 | 0 
gastric bypass surgery | 0 | 0 
pre-existing hypoparathyroidism | 0 | 0 
hypocalcaemia management | 0 | 192 
potential difficulties | 0 | 0 
approval of subcutaneous recombinant PTH | 0 | 0 
hypoparathyroidism in Australia | 0 | 0 
future management | 0 | 0 
elective bariatric surgery | 0 | 0 
patients with pre-existing hypoparathyroidism | 0 | 0 
careful consideration | 0 | 0 
hypocalcaemia | 4 | 192 
impaired gastrointestinal absorption | 0 | 192 
complications | 0 | 192 
subcutaneous recombinant PTH | 0 | 0 
hypoparathyroidism management | 0 | 192 
parenteral treatment | 0 | 192 
calcium replacement | 0 | 192 
intravenous calcium gluconate | 4 | 192 
intravenous calcitriol | 42 | 192 
intramuscular cholecalciferol | 56 | 56 
intravenous thyroxine | 88 | 192 
maintenance schedule | 88 | 192 
discharge | 192 | 192 
