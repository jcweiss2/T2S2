27 years old | 0
female | 0
emergency cesarean section due to arrest of labor | 0
bradycardia | -0.5
hypotension | -0.5
postpartum hemorrhage | 0
hypoxemia | 24
refractory hypotension | 24
hemoglobin 115 g/L | 24
platelet count 81 × 10E9/L | 24
fibrinogen 0.4 g/L | 24
international normalized ratio 1.8 | 24
creatinine 130 μmol/L | 24
pH 7.38 | 24
pCO2 26 mm Hg | 24
pO2 91 mm Hg | 24
HCO3 15 mmol/L | 24
lactate 1.7 mmol/L | 24
sinus tachycardia | 24
nonspecific T-wave changes | 24
troponin level elevated 492 ng/L | 24
RV dilation | 24
reduced RV systolic function | 24
McConnell’s sign | 24
moderate tricuspid regurgitation | 24
IVC thrombus | 24
pulmonary embolism | 24
gonadal vein thrombosis | 24
bilateral renal cortical necrosis | 24
norepinephrine initiation | 48
epinephrine administration | 24
dobutamine administration | 24
unfractionated heparin initiation | 48
hemodynamic improvement | 72
pressor support weaning | 72
continuous renal replacement therapy initiation | 48
intermittent hemodialysis transition | 144
discharge | 288
3-month follow-up | 2160
repeat echocardiogram normal biventricular function | 2160
no dialysis dependence | 2160
