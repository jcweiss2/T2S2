57 years old | 0
female | 0
menopausal | 0
admitted to the gynecological emergency unit | 0
left lower quadrant abdominal pain | -504
pelvic heaviness | -504
urinary frequency | -504
past history of 5 miscarriages | -10000
tubal ligation | -10000
active smoker | 0
no medication | 0
large and painful mass | 0
pelvic MRI | 0
mass measuring 18 × 17 × 12 cm | 0
well-delimited, polylobed, poorly vascularized | 0
central fluid component | 0
seemingly located on the left ovary | 0
extending up to the umbilicus | 0
no lymphadenopathy | 0
no ascites | 0
no peritoneal implants | 0
uterus and adnexa were normal | 0
serum tumor markers were negative | 0
surgical pelvic exploration | 672
30-centimeter mass of the left broad ligament | 672
no ascites | 672
no peritoneal carcinomatosis | 672
uterus and right adnexa were normal | 672
total hysterectomy with adnexectomy | 672
removal of the mass | 672
definitive histological diagnosis was leiomyosarcoma | 672
isolated fever | 48
fever of 39 °C | 48
major inflammatory syndrome | 48
leukocytes 15,000/μL | 48
C-reactive protein 317 mg/dL | 48
contrast-enhanced computed tomography scan | 48
bilobed air and fluid collection | 48
abscess | 48
retroperitoneum | 48
left psoas muscle | 48
Douglas pouch | 48
blood pressure dropped | 48
74/46 mmHg | 48
intravenous volume replacement | 48
2 L of Ringer Lactate | 48
vasopressor therapy | 48
continuous infusion of noradrenaline | 48
blood pressure stabilization | 48
100/60 mmHg | 48
emergency revision surgery | 72
peritoneal cavity exploration | 72
moderately abundant non-purulent serosanginous peritoneal fluid | 72
adhesions to the Douglas pouch | 72
peritonitis | 72
antibacterial treatment | 72
piperacillin/tazobactam | 72
gentamicin | 72
microbiological samples | 72
extubated | 72
hemodynamic support | 72
noradrenaline | 72
transferred to the intensive care unit | 72
clinically improved | 96
noradrenaline requirement decreased | 96
discontinuation of noradrenaline | 96
decrease in inflammatory markers | 96
microbiological analysis of the peritoneal fluid | 96
Gardnerella vaginalis | 96
gentamicin discontinued | 96
metronidazole added | 96
Atopobium vaginae | 120
antibacterial susceptibility testing | 120
Garderella vaginalis resistant to metronidazole | 120
Garderella vaginalis resistant to ciprofloxacin | 120
Garderella vaginalis susceptible to penicillin G | 120
Garderella vaginalis susceptible to amoxicillin/clavulanate | 120
Garderella vaginalis susceptible to cefotaxim | 120
Garderella vaginalis susceptible to clindamicin | 120
Garderella vaginalis susceptible to vancomycin | 120
Atopobium vaginae susceptible to all tested antibacterials | 120
Atopobium vaginae susceptible to metronidazole | 120
piperacillin/tazobactam active against both bacteria | 120
discharged from the intensive care unit | 120
antibacterial therapy stopped | 168