14 years old | 0
    male | 0
    presented to the pediatric OPD | 0
    fever | -96
    abdominal pain | -72
    cough | -24
    chills | -96
    sweating | -96
    no rigors | -96
    periumbilical region pain | -72
    movement-aggravated pain | -72
    rest-relieved pain | -72
    coughing multiple episodes | -24
    dry cough | -24
    fast breathing | -24
    no noisy breathing | -24
    no chest indrawing | -24
    no bluish discoloration of skin | -24
    no recent travel | 0
    no known sick contacts | 0
    no chronic medications | 0
    no drug allergies | 0
    no dust allergies | 0
    no food allergies | 0
    thinly built | 0
    weight <3rd centile | 0
    febrile | 0
    tachypneic | 0
    respiratory rate 42 breaths/min | 0
    hypotension | 0
    blood pressure 90/48 (61) mm Hg | 0
    oxygen saturation maintained | 0
    right inguinal lymph nodes enlarged | 0
    non-tender lymph nodes | 0
    soft abdomen | 0
    distended abdomen | 0
    liver palpable 3 cm | 0
    liver span 12 cm | 0
    fluid thrill present | 0
    no splenomegaly | 0
    decreased air entry right mammary area | 0
    neutrophilia | 0
    lymphopenia | 0
    thrombocytopenia | 0
    elevated liver enzymes | 0
    low serum albumin | 0
    deranged liver function test | 0
    normal renal function test | 0
    arterial blood gas pH 7.43 | 0
    arterial blood gas Pco2 27 | 0
    arterial blood gas Po2 135 | 0
    arterial blood gas HCO3 20 | 0
    urine pus cells | 0
    urine culture no growth | 0
    negative scrub typhus test | 0
    chest X-ray diffuse coalescent opacities | 0
    chest X-ray volume loss left | 0
    ultrasound gross ascites | 0
    ultrasound minimal pleural effusion | 0
    echocardiography minimal pericardial effusion | 0
    echocardiography mild tricuspid regurgitation | 0
    echocardiography mild mitral regurgitation | 0
    ascitic fluid elevated WBC count | 0
    ascitic fluid lymphocytosis | 0
    ascitic fluid high ADA | 0
    ascitic fluid TC-300/mm3 | 0
    ascitic fluid N-2% | 0
    ascitic fluid L-98% | 0
    ascitic fluid glucose 92mg/dL | 0
    ascitic fluid protein 4g/dL | 0
    ascitic fluid ADA-54U/L | 0
    ascitic fluid LDH-1080IU/L | 0
    ascitic fluid gram stain no organisms | 0
    ascitic fluid culture no growth | 0
    normal peripheral blood smear | 0
    negative troponin marker | 0
    CK-MB 18IU/L | 0
    admitted to pediatric ICU | 0
    intravenous antibiotics | 0
    ceftriaxone | 0
    metronidazole | 0
    intravenous fluids | 0
    vasopressors | 0
    dobutamine | 0
    dopamine | 0
    albumin administration | 0
    CT scan subpleural reticular opacities | 0
    CT scan ground glass opacity | 0
    CT scan mild hepatomegaly | 0
    positive Covid-antibody | 0
    intravenous immunoglobulin | 0
    high dose methylprednisolone | 0
    suspected MIS-C | 0
    diuretics | 24
    low molecular weight heparin | 24
    BIPAP respiratory support | 24
    upgraded antibiotics | 96
    clindamycin | 96
    piperacillin-tazobactam | 96
    positive troponin marker | 120
    CK-MB 26 IU/L | 120
    improved condition | 120
    tapered inotropes | 120
    weaned oxygen | 120
    afebrile | 192
    oxygen saturation maintained | 192
    stopped low molecular heparin | 192
    stopped intravenous diuretics | 192
    oral rivaroxaban | 192
    oral diuretics | 192
    feeding initiated | 192
    shifted to pediatric ward | 312
    oxygen saturation room air | 312
    dilated IVC | 312
    dilated left ventricle | 312
    no diastolic dysfunction | 312
    minimum pericardial effusion | 312
    coronary artery diameter 3mm | 312
    ejection fraction 65% | 312
    improved platelet count | 312
    discharged | 336
    afebrile at discharge | 336
    feeding well | 336
    clinically stable | 336
    oral antibiotics | 336
    oral steroids | 336
    oral anticoagulants | 336
    oral diuretics | 336
    oral multivitamins | 336
    follow-up after 2 weeks | 336
    normal chest x-ray | 1344

<|eot_id|>