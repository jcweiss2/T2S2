11 years old | 0
female | 0
systemic methicillin-resistant staph aureus infection | -1008
right knee pain | -1008
back pain | -1008
fevers | -1008
purulent spider bite | -1008
COVID-19 infection | -1008
dehydration | -1008
altered mental status | -1008
incontinence | -1008
febrile | -1008
tachypneic | -1008
tachycardic | -1008
hypoxic | -1008
admitted to the pediatric intensive care unit | -1008
blood culture positive for MRSA | -1008
intravenous antibiotic therapy | -1008
magnetic resonance imaging of the spine | -1008
computed tomography of her chest, abdomen and pelvis | -1008
multifocal fluid collections | -1008
inflammation involving the right psoas muscle | -1008
right thoracolumbar paraspinal soft tissues | -1008
cervical and thoracic prevertebral soft tissues | -1008
multifocal septic arthritis | -1008
bilateral pleural effusions | -1008
multifocal opacities | -1008
multiple pulmonary nodules | -1008
septic emboli | -1008
MRI of the brain | -1008
signs of meningitis | -1008
ventriculitis | -1008
cerebrospinal fluid positive for MRSA | -1008
multiarticular surgical washouts | -1008
washout of her paraspinal abscesses | -1008
bilateral chest tubes | -1008
empyema | -1008
clearing of her blood cultures | -792
transferred to our facility for rehabilitation | -792
clinically well appearing | 0
afebrile | 0
normal vital signs | 0
CT imaging of her chest, abdomen, and pelvis | 192
increased size of the right psoas collection | 192
MRI showing increased T1 signal intensity | 192
CT angiography | 192
enhancing lesions in the left medial lower lobe | 192
right posterior mediastinum | 192
right psoas | 192
pseudoaneurysms | 192
retrospective review of the prior imaging | 192
hematocrit level remained stable | 192
interventional radiology service consulted | 192
embolization | 192
access obtained to the right common femoral vein | 192
left pulmonary artery selectively catheterized | 192
diagnostic angiogram | 192
pseudoaneurysm arising from a medial branch | 192
embolization coils | 192
postembolization angiography | 192
access obtained to the left common femoral artery | 192
diagnostic angiography of the right L2-L3 lumbar artery | 192
pseudoaneurysm arising from a superior intramuscular branch | 192
coil embolized | 192
pseudoaneurysm in the posterior mediastinum | 192
active hemorrhage | 192
embolized | 192
postembolization angiography | 192
completion fluoroscopic images | 192
embolization coils at the sites of all 3 treated pseudoaneurysms | 192
returned to the PICU | 192
clinically stable | 192
transferred back to the rehabilitation medicine service | 216
CT angiogram | 432
stable position of embolization coils | 432
no evidence of recurrent pulmonary, lumbar, or intercostal PSA | 432
marked decrease in the size of her right psoas collection | 432
discharged | 504
follow-up CT angiogram | 1224
further decrease in the size of her multifocal fluid collections | 1224
no evidence of new or recurrent PSAs | 1224