34 years old| 0
female | 0
COVID-19 infection | 0
cough | -72
fever | -72
COVID-19 positive | 0
admitted to another hospital | 0
chest CT showing bilateral and peripheral ground-glass opacity | 0
moderate COVID-19 pneumonia | 0
intravenous remdesivir | 0
oral dexamethasone | 0
discharged | 240
chest pain | 24
ECG ST elevation in leads II, III, and aVF | 24
inferior-wall acute myocardial infarction | 24
emergency coronary angiography showing embolic occlusion in left circumflex branch | 24
anticoagulation with heparin sodium | 24
contrast-enhanced CT showing right renal infarction | 24
brain MRI showing acute multi-territory ischemic stroke | 24
fever of 38.9℃ | 24
blood culture positive for Gram-positive coccus | 24
transthoracic echocardiography showing 11-mm vegetation on posterior mitral valve leaflet | 24
left ventricular ejection fraction 60% | 24
native mitral valve IE causing multiple embolisms | 24
intravenous vancomycin | 24
cefazolin | 24
transferred to university hospital | 24
clear consciousness | 0
no neurological deficit | 0
blood pressure 74/48 mmHg | 0
pulse 69 beats/minute | 0
body temperature 39.1℃ | 0
conjunctiva petechiae | 0
hemorrhagic spots on soft palate | 0
grade II/VI pansystolic murmur | 0
white blood cell count 20.9 K/μL | 0
C-reactive protein 10.12 mg/dL | 0
Troponin T 0.627 ng/mL | 0
NT-proBNP 4,041 pg/mL | 0
lactate 2.9 mmol/L | 0
chest X-ray no cardiac enlargement | 0
ECG sinus rhythm | 0
transthoracic echocardiography showing 13.8×6.8 mm vegetations on mitral posterior leaflet | 0
severe mitral regurgitation | 0
MSSA infection | 0
antimicrobial therapy continued | 0
antimicrobial refractory IE | 0
septic shock | 0
surgical mitral valve replacement | 168
discharged | 600
