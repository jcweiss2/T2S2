18 years old | 0
male | 0
admitted to the hospital | 0
COVID-19 pneumonia | 0
acute respiratory failure | 0
oxygen therapy | 0
nonrebreather mask oxygen | 0
SpO2 89% | 0
pH 7.45 | 0
PaCO2 36 | 0
PaO2 65 | 0
PaO2/FiO2 175.7 | 0
awake prone position | 0
noninvasive mechanical ventilation | -672
nasal high-flow therapy | -672
intubation | 24
ventilator-free days | 72
ICU stay | 120
short-term mortality | 672
discharged | 720
SpO2 95% | 24
pH 7.46 | 24
PaCO2 37 | 24
PaO2 82 | 24
PaO2/FiO2 190.2 | 24
intubation requirement | 24
mortality rate | 672
diabetes | -672
hypertension | -672
coronary artery disease | -672
chronic obstructive pulmonary disease | -672
congestive heart failure | -672
chronic renal failure | -672
cancer | -672
other comorbidities | -672