33 years old | 0
male | 0
renal transplant recipient | 0
admitted to the hospital | 0
severe upper abdominal pain | -72
nausea | -72
upper abdominal pain radiating towards his back | -72
immunosuppressive therapy with methylprednisolone, tacrolimus, and mycophenolate mofetil (MMF) | -4320
end-stage renal disease | -4320
parent-to-child kidney transplantation | -4320
analgesic treatment | -72
abdominal computed tomography (CT) | -72
ultrasonography | -72
aspartate aminotransferase (AST) increased | -72
alanine aminotransferase (ALT) increased | -72
referred to the hospital | -72
complained of nausea | 0
complained of upper abdominal pain | 0
diagnosis of acute abdominal pain | 0
diagnosis of liver damage | 0
flurbiprofen tapes for pain relief | 0
intravenous magnesium isoglycyrrhizinate against liver damage | 0
empirical antimicrobial therapy with intravenous cefoperazone sodium and sulbactam sodium | 0
septic shock | 24
multiple organ dysfunction syndrome (MODS) | 24
liver dysfunction | 24
acute kidney injury | 24
transferred to the intensive care unit (ICU) | 24
lethargic | 0
heart rate of 136 beats/min | 0
respiratory rate of 23 breaths/min | 0
blood pressure of 83/42 mmHg | 0
body temperature of 36.8 °C | 0
abdominal tenderness in the upper quadrants | 0
no muscle guarding or rebound tenderness | 0
high levels of ALT | 0
high levels of AST | 0
high levels of alkaline phosphatase | 0
high levels of gamma-glutamyltransferase | 0
high concentrations of C-reactive protein | 0
high concentrations of procalcitonin | 0
high concentrations of creatinine | 0
prolonged activated partial thromboplastin time | 0
prolonged thrombin time | 0
low fibrinogen | 0
serological tests for hepatitis A, B, and C viruses | 0
serological tests for human immunodeficiency virus | 0
serological tests for treponema pallidum | 0
hepatitis B surface and core antibodies | 0
immunoglobulin (Ig) M antibodies against toxoplasma | 0
immunoglobulin (Ig) M antibodies against rubella virus | 0
immunoglobulin (Ig) M antibodies against cytomegalovirus | 0
immunoglobulin (Ig) M antibodies against herpes simplex virus 2 | 0
blood culture | 0
polymerase chain reaction (PCR) of Epstein-Barr virus DNA | 0
abdominal ultrasonography | 0
abdominal and pelvic CT | 0
chest X-ray | 0
electrocardiogram | 0
next-generation sequencing (NGS) | 24
real-time PCR for VZV | 24
VZV IgG-negative | 24
visceral disseminated VZV infection | 24
septic shock | 24
MODS with liver dysfunction and acute kidney injury | 24
antiviral therapy with intravenous acyclovir | 24
intravenous meropenem | 24
intravenous linezolid | 24
intravenous caspofungin | 24
noradrenaline | 24
terlipressin | 24
intravenous sodium bicarbonate | 24
acute liver failure | 40
disseminated intravascular coagulation | 40
acute respiratory failure | 40
acute renal injury | 40
died | 40