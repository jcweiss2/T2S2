76 years old | 0
male | 0
diabetic | 0
hypertensive | 0
post-coronary artery bypass graft surgery | 0
admitted to the hospital | 0
fever | -120
myalgia | -120
tested positive for SARS-CoV-2 infection | -120
ICD implantation | -2628
CT coronary angiography | -432
patent grafts | -432
asymptomatic | -432
metoprolol XL | -432
telmisartan | -432
spironolactone | -432
multiple ICD shocks | -6
stable vital signs | 0
oxygen saturation of 97% | 0
normal sinus rhythm | 0
no ST-T changes | 0
QTc interval of 464 milliseconds | 0
global hypokinesia | 0
left ventricular ejection fraction of 30% | 0
elevated C-reactive protein | 0
elevated ferritin | 0
elevated creatine kinase | 0
elevated troponin T | 0
elevated N-terminal pro-brain natriuretic peptide | 0
monomorphic VTs | 0
ventricular ectopic | 0
anti-tachycardia pacing | 0
ICD-delivered shocks | 0
amiodarone infusion | 0
metoprolol doses increased | 0
VT storm controlled | 24
symptomatic treatment for COVID-19 infection | 0
recovered | 240
discharged | 240
amiodarone | 240
metoprolol XL | 240
telmisartan | 240
torsemide-spironolactone | 240
aspirin | 240
statins | 240
oral hypoglycemics | 240
no episodes of VT | 2160
asymptomatic | 2160