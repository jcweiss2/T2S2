22 years old | 0
male | 0
admitted to the hospital | 0
fever | -96
myalgia | -96
arthralgia | -96
sore throat | -96
vomiting | -48
diarrhoea | -48
intensive care admission | 24
high-dose intravenous steroids | 24
severe global left ventricular impairment | 24
elevated troponin | 24
myocarditis | 24
cardiac MRI | 96
severe global left ventricular systolic impairment | 96
elevated ferritin | 288
maculopapular rash | 384
rheumatology review | 384
Adult-onset Still’s disease | 384
pulsed i.v. methylprednisolone | 408
tocilizumab | 408
clinical and biochemical improvement | 408
transitioned to oral prednisone | 576
discharged home | 600
clinical and biochemical relapse | 888
tocilizumab dose escalation | 1008
biochemical remission | 1512
ceased prednisone | 4320
transitioned to fortnightly subcutaneous adalimumab | 7200
repeat cardiac MRI | 12960
no evidence of on-going inflammation | 12960
non-smoker | 0
no regular medications | 0
no past medical history | 0
no recreational drug history | 0
no family history | 0
fever of 38.4°C | 0
pulse 89 beats per minute | 0
blood pressure 77/34 mmHg | 0
respiratory rate 18 breaths per minute | 0
oxygen saturations 98% | 0
normal haemoglobin | 0
mild thrombocytopaenia | 0
leukocytosis | 0
neutrophilia | 0
monocytosis | 0
lymphopaenia | 0
normal eosinophils | 0
normal basophils | 0
acute kidney injury | 0
mildly deranged liver function tests | 0
high-sensitivity troponin T elevated | 0
elevated NT-proBNP | 0
C-reactive protein elevated | 0
lactate raised | 0
mild hyponatraemia | 0
normal potassium | 0
sinus rhythm | 0
right-axis deviation | 0
diffuse ST-segment elevation | 0
unremarkable chest radiograph | 0
septic shock | 24
vasopressor support | 24
empiric broad-spectrum antibiotics | 24
high-dose intravenous dexamethasone | 24
clinical and biochemical improvement | 24
transthoracic echocardiography | 24
severe global left ventricular systolic impairment | 24
moderate systolic impairment | 24
no significant valvular pathology | 24
no pericardial effusion | 24
endomyocardial biopsy | 24
subtle interstitial lymphocytes | 24
oedema | 24
no myonecrosis | 24
no giant cells | 24
no eosinophils | 24
no granulomas | 24
no fibrosis | 24
negative stains for amyloid and iron | 24
cardiac MRI | 96
high myocardial T2 signal | 96
myocardial oedema | 96
extensive circumferential late gadolinium enhancement | 96
subepicardial distribution | 96
consistent with acute myocarditis | 96
attempt to de-escalate intravenous to oral steroid therapy | 240
unsuccessful | 240
clinical and biochemical deterioration | 240
re-attempt to de-escalate intravenous to oral steroid therapy | 336
unsuccessful | 336
clinical and biochemical deterioration | 336
rheumatology review | 384
strong suspicion for diagnosis of Adult-onset Still’s disease | 384
new maculopapular rash | 408
consistent with AOSD diagnosis | 408
commencement of pulsed i.v. methylprednisolone | 408
initial infusion of tocilizumab | 408
first signs of sustained clinical and biochemical improvement | 408
transitioned to oral prednisone | 576
discharged home | 600
signs of clinical and biochemical relapse | 888
second infusion of tocilizumab | 1008
tocilizumab dose escalation | 1008
third infusion of tocilizumab | 1008
biochemical remission | 1512
ceased prednisone | 4320
transitioned to fortnightly subcutaneous adalimumab | 7200
repeat cardiac MRI | 12960
no evidence of on-going inflammation | 12960