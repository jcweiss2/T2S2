spleen removal due to idiopathic thrombocytopenic purpura and menometrorhagia | -15552
vaccination with PPV23 | -15552
vaccination response test | -4
general body malaise | -48
diarrhea | -48
vomiting | -48
influenza-like symptoms | -48
confusion | -24
hospital admission | 0
fever | 0
hypotension | 0
bradycardia | 0
tachypnea | 0
decreased oxygen saturation | 0
cyanosis | 0
no sign of neck stiffness | 0
no meningeal reactions | 0
normal cardiac and pulmonic auscultations | 0
soft and not tender abdomen | 0
diagnosis of severe sepsis | 0
volume therapy | 0
broad-spectrum antimicrobial therapy | 0
hydrocortisone | 0
laboratory studies | 0
white blood cell count | 0
neutrophils | 0
hemoglobin | 0
thrombocytes | 0
C-reactive protein | 0
P-lactate | 0
aB-P-O2 | 0
aB-P-CO2 | 0
aB-pH | 0
Streptococcus pneumococcal urinary antigen test | 0
chest x-ray | 0
discrete pulmonic stasis | 0
transfer to ICU | 0
disseminated intravascular coagulation | 24
microthrombi in hands and feet | 24
blood cultures showed growth of S. pneumoniae | 48
antimicrobial treatment changed to penicillin G | 48
suspicion of endocarditis | 72
trans-thoracic echocardiography | 72
modest hypokinesia of left ventricle | 72
ejection fraction of 45% | 72
no endocarditis | 72
necrosis of fingertips and toes | 72
renal insufficiency | 72
hemodialysis | 72
antibiotic therapy altered to ceftriaxone | 72
leucocytes and CRP decreased | 96
fever dissolved | 96
tracheal secret culture negative | 96
transfer from ICU to medical department | 216
antibiotics stopped | 216
serological analysis of pneumococcal isolate | 216
serotype 12F | 216
afebrile with fluctuating CRP | 270
clinical condition improved | 270
discharge with oral dicloxacillin | 528
necrotic fingers and toes amputated | 2160
readmission with severe sepsis | 2160
sepsis regimen and ceftriaxone therapy | 2160
transesophageal echocardiography | 2160
endocarditis with moving elements on aortic valve | 2160
blood cultures showed growth of S. pneumoniae | 2160
antimicrobial treatment altered to penicillin G | 2160
conservative treatment with penicillin G | 2160
recovery | 2268
serological tests of pneumococcal capsule polysaccharides | 0
antibody response test | -15552
antibody response test | -4
antibody response test | 2160
antibody response test | 3720