73 years old | 0
male | 0
admitted to the hospital | 0
huge mass in left scrotum | 0
intolerable lower abdominal pain | 0
groin pain | 0
duration of 2 weeks | -336
left inguinoscrotal hernia diagnosis | -14400
refusal of early surgical intervention | -14400
general weakness | -144
decreased urine output | -144
pitting edema of bilateral lower limbs | 0
tenderness in left lower abdomen | 0
tenderness in inguinal region |8
large irreducible inguinoscrotal hernia | 0
bilateral inguinal ecchymosis | 0
white blood cell count 21.57 × 10³/μL | 0
92.3% neutrophils | 0
thrombocytopenia | 0
platelet count 90 × 10³/μL | 0
C-reactive protein 35.32 mg/dL | 0
procalcitonin 24.96 ng/mL | 0
serum creatinine 2.3 mg/dL | 0
abdominal CT scan without contrast | 0
herniation of small intestine | 0
herniation of colon | 0
small number of ascites | 0
incarcerated inguinal hernia | 0
sepsis | 0
intravenous administration of Flomoxef | 0
emergency surgery | 0
supine position under general anesthesia | 0
inguinal incision on left side | 0
hernial sac filled with ileum | 0
hernial sac filled with sigmoid colon | 0
failure to reduce contents into abdominal cavity | 0
mini-midline incision | 0
incarcerated organs pulled out | 0
adhesion separation | 0
hernial contents grossly inflamed | 0
mild swelling | 0
erythematous appearance | 0
incarcerated organs reduced into abdomen | 0
hernial repair with tension-free techniques | 0
unabsorbable polypropylene mesh sutured | 0
Jackson-Pratt drain placement | 0
transfer to intensive care unit | 0
no complications during early postoperative period | 24
adequate infection control | 336
recovered and discharged | 336
no evidence of relapse at 3-month follow-up | 2160
