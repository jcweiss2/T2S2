51 years old | 0
male | 0
non-smoker | 0
admitted to the emergency room | 0
abdominal pain | -72
no medical history | 0
no drug history | 0
denies significant family history of the disease | 0
diaphoretic | 0
uncomfortable | 0
severe distress | 0
blood pressure 156/87 mm Hg | 0
respiratory rate 19 breaths/minute | 0
heart rate 132 beats/minute | 0
temperature within normal limits | 0
oxygen saturation 93% on room air | 0
distended abdomen | 0
severely tender to palpation | 0
IV fluids started | 0
IV ondansetron for nausea | 0
morphine sulfate for pain | 0
leukocytosis | 0
WBC count 14.5 thou/cm | 0
laparotomy | 0
small and large intestine normal | 0
vasculature normal | 0
discharged | 48
nausea | 72
abdominal pain | 72
dyspnea | 72
tachypnea | 72
tachycardia | 72
low-grade fever | 72
lung CT | 72
abdominopelvic CT | 72
intubated | 72
Covid-19 RT-PCR | 72
CBC | 72
WBC 17000 per microliter | 72
Hb 12.8.7 g/dL | 72
Plt 350,000 per microliter | 72
urea 170 mg/dL | 72
Cr 4.2 mg/dL | 72
LDH 504 U/L | 72
CRP 47mg/L | 72
negative viral disease | 72
hydroxychloroquine sulfate | 72
lopinavir/ritonavir | 72
ribavirin | 72
β interferon | 72
fecaloid discharged from abdominal suture | 120
sepsis | 120
CBC | 120
WBC 24000 per microliter | 120
Hb 12 g/dL | 120
Plt 347000 per microliter | 120
urea 206 mg/dL | 120
Cr 3.2 mg/dL | 120
amylase 67 U/L | 120
re-laparotomy | 120
serosanguinous secretions | 120
necrotic changes in the small intestine | 120
small intestine resected | 120
ileostomy | 120
pathological study | 120
intravascular thrombosis | 120
mesenteric tissue necrotic margin | 120
RT-PCR of covid-19 positive | 120
heparin infusion | 120
broad-spectrum antibiotics | 120
extubated | 192
hemodynamic stable | 192
platelet count decreased | 192
gastrointestinal bleeding | 216
CBC | 216
WBC 7100 per microliter | 216
Hb 8.7 g/dL | 216
plt 162000 per microliter | 216
Cr 1.3 mg/dL | 216
amylase 65 U/L | 216
Plt decreased | 216
Cr decreased | 216
PT normal | 216
PTT normal | 216
D-dimer 2500 ng/mL | 216
fibrinogen 150 mg/dL | 216
PT 44 sec | 216
PTT 44 sec | 216
INR 1.7 | 216
no schistocyte | 216
treatment-resistant sepsis | 216
DIC | 216
death | 216