24 years old | 0 | 0 | Factual
primigravida | 0 | 0 | Factual
37 weeks of gestation | 0 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
high grade fever | -72 | 0 | Factual
decreased urine output | -72 | 0 | Factual
yellowish discolouration | -72 | 0 | Factual
altered sensorium | -72 | 0 | Factual
disoriented | 0 | 0 | Factual
febrile | 0 | 0 | Factual
icteric | 0 | 0 | Factual
sub-conjunctival haemorrhages | 0 | 0 | Factual
fine basal crepitations | 0 | 0 | Factual
receiving intravenous artesunate | -72 | 0 | Factual
receiving ceftriaxone | -72 | 0 | Factual
receiving doxycycline | -72 | 0 | Factual
anaemia | 0 | 0 | Factual
jaundice | 0 | 0 | Factual
deranged liver function | 0 | 0 | Factual
coagulopathy | 0 | 0 | Factual
thrombocytopenia | 0 | 0 | Factual
increased total leucocyte count | 0 | 0 | Factual
elevated blood urea nitrogen | 0 | 0 | Factual
elevated serum creatinine | 0 | 0 | Factual
singleton pregnancy | 0 | 0 | Factual
adequate liquor | 0 | 0 | Factual
umbilical artery systolic-diastolic ratio of 2:1 | 0 | 0 | Factual
mild hepato-splenomegaly | 0 | 0 | Factual
non-reassuring fetal heart rate | 0 | 0 | Factual
aspiration prophylaxis | 0 | 0 | Factual
high-risk consent | 0 | 0 | Factual
rapid sequence intubation | 0 | 0 | Factual
cricoid pressure | 0 | 0 | Factual
thiopental | 0 | 0 | Factual
succinylcholine | 0 | 0 | Factual
right internal jugular vein cannulation | 0 | 0 | Factual
left radial artery cannulation | 0 | 0 | Factual
anaesthesia maintained with isoflurane | 0 | 2 | Factual
N2O-O2 mixture | 0 | 2 | Factual
atracurium | 0 | 2 | Factual
delivery of a 2.25 kg baby | 2 | 2 | Factual
fentanyl | 2 | 2 | Factual
oxytocin infusion | 2 | 24 | Factual
Apgar score of 6 | 2 | 2 | Factual
Apgar score of 8 | 7 | 7 | Factual
cord blood pH of 7.28 | 2 | 2 | Factual
base deficit of 5.4 | 2 | 2 | Factual
blood sugar level of 50 mg/dl | 2 | 2 | Factual
hypotension | 2 | 24 | Factual
blood loss | 2 | 24 | Factual
packed red blood cells transfusion | 2 | 24 | Factual
fresh frozen plasma transfusion | 2 | 24 | Factual
platelets transfusion | 2 | 24 | Factual
noradrenaline infusion | 2 | 24 | Factual
mild acidosis | 24 | 24 | Factual
normal electrolytes | 24 | 24 | Factual
normal serum glucose | 24 | 24 | Factual
intensive care unit | 24 | 144 | Factual
post-operative analgesia | 24 | 144 | Factual
ultrasound guided bilateral transverse abdominis plane block | 24 | 144 | Factual
pulmonary haemorrhage | 48 | 48 | Factual
blood products transfusion | 48 | 48 | Factual
fibre-optic bronchoscopy | 48 | 48 | Factual
erythematous mucosa | 48 | 48 | Factual
blood clots | 48 | 48 | Factual
active oozing | 48 | 48 | Factual
diffuse bleeding | 48 | 48 | Factual
broncho alveolar lavage | 48 | 48 | Factual
Factor VIIa administration | 48 | 48 | Factual
bleeding cessation | 60 | 60 | Factual
reduction of inspired oxygen fraction | 60 | 60 | Factual
bilateral non-homogeneous opacities | 48 | 48 | Factual
clear chest radiograph | 60 | 60 | Factual
acute kidney injury | 0 | 144 | Factual
severe hyperbilirubinemia | 0 | 144 | Factual
haemolytic uremic syndrome | 0 | 144 | Factual
high serum lactate dehydrogenase | 0 | 144 | Factual
schistocytes in peripheral blood | 0 | 144 | Factual
nephrology opinion | 72 | 72 | Factual
plasmapheresis | 72 | 72 | Factual
dialysis | 72 | 72 | Factual
computed tomography of the brain | 72 | 72 | Factual
diffuse cerebral oedema | 72 | 72 | Factual
cerebroprotective measures | 72 | 144 | Factual
head elevation | 72 | 144 | Factual
not rotating neck | 72 | 144 | Factual
maintain serum sodium 145-155 Meq/L | 72 | 144 | Factual
keeping blood partial pressure of carbondioxide 32-40 mmHg | 72 | 144 | Factual
stress ulcer prevention | 24 | 144 | Factual
deep vein thrombosis prophylaxis | 24 | 144 | Factual
glycemic control | 24 | 144 | Factual
reducing fever | 96 | 96 | Factual
improving consciousness | 96 | 96 | Factual
inotropic support tapered | 96 | 96 | Factual
improving urine output | 96 | 96 | Factual
improving liver function test | 96 | 96 | Factual
improving coagulation parameters | 96 | 96 | Factual
improving Pao2/Fio2 ratio | 96 | 144 | Factual
extubation | 144 | 144 | Factual
discharged from the hospital | 168 | 168 | Factual