68 years old| 0
    male| 0
    no previous medical history| 0
    no known history of allergy| 0
    no known history of asthma| 0
    brought to the emergency department| 0
    near cardiac arrest| 0
    persistent severe hypotension| 0
    made spicy pork kidneys| -24
    dinner| -24
    found gasping on the armchair| -24
    telephone-assisted CPR| -24
    CPR performed for 15 minutes| -24
    spontaneous circulation restored| -24
    severely hypotensive| -24
    norepinephrine administration| -24
    afebrile| 0
    tachycardic| 0
    tachypneic| 0
    oxygen saturation of 85%| 0
    drowsy| 0
    awake| 0
    Glasgow coma scale of 4-5-6| 0
    heart auscultation no murmurs| 0
    lung sounds clear| 0
    abdomen soft| 0
    no tenderness| 0
    no guarding| 0
    skin examination no efflorescence| 0
    tick embedded in the skin extracted| 0
    mechanical ventilation initiated| 0
    sinus tachycardia| 0
    no signs of acute ischaemia| 0
    white cell count 14,700 per cubic millimeter| 0
    predominantly neutrophils| 0
    C-reactive protein elevated to 64 mg/l| 0
    procalcitonin 0.1 ng/ml| 0
    renal functions normal| 0
    hepatic enzymes normal| 0
    lactate elevated 6.3 mmol/l| 0
    echocardiography no hypovolemia| 0
    no regional dyskinesis| 0
    no akinesis| 0
    no signs of right ventricular strain| 0
    no LVOTO| 0
    high left ventricle ejection fraction| 0
    hyperkinetic circulation| 0
    whole-body CT consolidation lower lobe left lung| 0
    pneumonia suspicion| 0
    treating for pneumonia| 0
    treating for septic shock| 0
    started to feel itches all over after lunch| -24
    precipitous speed of deterioration| 0
    postprandial timing| 0
    itchy skin| 0
    protracted anaphylaxis diagnosis| 0
    serum tryptase elevated 52.9 mcg/l| 0
    total IgE levels elevated| 0
    investigation of potential trigger| 0
    spices| -24
    pork kidneys| -24
    delayed allergic reaction| 0
    alpha-gal syndrome considered| 0
    specific IgE against alpha-gal positive 85 kIU/l| 0
    allergologist consultation requested| 0
    alpha-gal syndrome diagnosed| 0
    vasoplegic shock| 0
    rapid progression to cardiac arrest| 0
    tick-borne anaphylaxis| 0
    severe protracted anaphylaxis| 0
    alpha-gal syndrome| 0
    life-threatening protracted delayed vasoplegic shock| 0
    idiopathic anaphylaxis| 0
    vasoplegia| 0
    diagnostic errors| 0
    tick-borne diseases| 0
    written informed consent obtained| 0