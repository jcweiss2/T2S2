57 years old | 0
female | 0
admitted to the hospital | 0
medical history of diabetes | 0
medical history of hypertension | 0
high-grade fever | -72
history of fall | -336
initial treatment at a primary health center | -336
ambulating well at home | -336
conscious and oriented | 0
febrile | 0
hypotensive | 0
minimal respiratory distress | 0
diagnosis of sepsis | 0
fluid resuscitation | 0
cultures | 0
imaging | 0
broad-spectrum antibiotics | 0
leukocytosis | 0
toxic neutrophil granulation | 0
normal renal panel | 0
normal liver panel | 0
normal coagulation panel | 0
right axis deviation | 0
S1Q3T3 pattern | 0
no right heart strain | 0
no lower limb deep venous thrombosis (DVT) | 0
CT pulmonary angiogram | 0
no pulmonary embolism (PE) | 0
unfractionated heparin for DVT prophylaxis | 0
blood cultures grew methicillin-sensitive Staphylococcus aureus (MSSA) | 24
antibiotic de-escalation | 24
gradually improving | 24
CT abdomen | 24
fracture of body of D8 vertebra | 24
transesophageal echocardiography | 24
no infective endocarditis | 24
acute left lower limb swelling | 48
pain | 48
redness | 48
acute DVT | 48
therapeutic anticoagulation with intravenous heparin infusion | 48
magnetic resonance imaging of the spine | 72
moderate wedging of T8 and T11 vertebral body | 72
no cord edema or mass | 72
compression of the left common iliac vein by the right common iliac artery | 72
acute thrombus in the left common iliac vein | 72
May-Thurner syndrome (MTS) | 72
catheter-based thrombolysis suggested | 96
venous stenting suggested | 96
placement of filter in the inferior vena cava (IVC) | 120
long-term anticoagulation with factor Xa inhibitor (Rivaroxaban) | 120
afebrile and stable at discharge | 168
asymptomatic during subsequent follow-up | 720