80 years old | 0\
female | 0\
non-smoker | 0\
hypertension | 0\
acute dyspnea | -24\
fecal incontinence | -7.4\
left hemiplegia | -7.4\
dextroversion | -7.4\
dysarthria | -7.4\
vomiting | -7.4\
impaired consciousness | -7.4\
transported to the emergency department | -7.4\
right thalamus and putamen bleeding | -7.4\
conservative treatment | -7.4\
poor oral hygiene | -7.4\
diminished breath sounds on the left side | -7.4\
coarse crackles in the right lung | -7.4\
decrease in breath sounds in the front of the chest | -7.4\
respiratory condition deteriorated | -7.4\
endotracheal intubation | -7.4\
mechanical ventilation | -7.4\
bilateral infiltration | -7.4\
admitted to the intensive care unit | -7.4\
decreased leukocyte count | -7.4\
mildly elevated C-reactive protein level | -7.4\
respiratory failure | -7.4\
partial pressure of oxygen in arterial blood | -7.4\
normal hepatorenal function | -7.4\
extensive infiltration shadows | -7.4\
hematoma extending from the right basal ganglia and putamen to the thalamus | -7.4\
cerebral edema | -7.4\
consolidations admixture with ground-glass opacities | -7.4\
Mendelson's syndrome | -7.4\
aspiration of gastric contents | -7.4\
bacterial aspiration pneumonia | -7.4\
Streptococcus agalactiae | -7.4\
Klebsiella oxytoca | -7.4\
leukocytopenia | -7.4\
low serum CRP level | -7.4\
respiratory viral pneumonia | -7.4\
management in the ventilator mode | 0\
meropenem | 0\
levofloxacin | 0\
prednisolone | 0\
synchronous intermitted mandatory ventilation with pressure control ventilation | 0\
intravenous Sivelestat sodium hydrate | 0\
lung-protection strategies | 0\
low tidal volume strategy with permissive hypercapnia | 0\
partial pressure of oxygen in arterial blood/fraction of inspired oxygen | 0\
P/F ratio | 0\
moderate severity | 0\
no fever | 0\
temperature never exceeded 37 °C | 0\
infiltration shadows improved | 288\
P/F ratio improved | 288\
extubated | 288\
transferred to the Department of Neurosurgery | 528\
transferred to a rehabilitation hospital | 528