73 years old | 0
male | 0
admitted to the hospital | 0
huge mass in left scrotum | 0
intolerable lower abdominal and groin pain | 0
duration of approximately 2 weeks | -336
diagnosed with huge left inguinoscrotal hernia | -1440
refused early surgical intervention | -1440
general weakness | -168
decreased urine output | -168
history of left inguinal hernia | -1440
no history of chronic diseases | 0
no history of surgeries | 0
working as a security guard | 0
lifting and carrying packages | 0
no relevant family history | 0
body temperature 36°C | 0
blood pressure 106/73 mmHg | 0
heart rate 95 beats/min | 0
respiratory rate 22 breaths/min | 0
pitting edema of bilateral lower limbs | 0
tenderness in left lower abdomen and inguinal region | 0
large irreducible inguinoscrotal hernia | 0
bilateral inguinal ecchymosis | 0
white blood cell count 21.57 × 10^3/μL | 0
neutrophils 92.3% | 0
thrombocytopenia | 0
platelet count 90 × 10^3/μL | 0
C-reactive protein 35.32 mg/dL | 0
procalcitonin 24.96 ng/mL | 0
serum creatinine 2.3 mg/dL | 0
abdominal computed tomography scan | 0
huge left inguinal hernia | 0
herniation of small intestine and colon | 0
small number of ascites | 0
intravenously administered antibiotics | 0
Flomoxef 1g every 12 h | 0
emergency surgery | 0
ingual incision on left side | 0
hernial sac filled with ileum and sigmoid colon | 0
mini-midline incision | 0
incarcerated organs pulled out | 0
adhesion between hernial contents separated | 0
hernial contents grossly inflamed | 0
hernial repair using tension-free techniques | 0
unabsorbable polypropylene mesh | 0
Jackson-Pratt drain placed | 0
transferred to intensive care unit | 0
no complications during early postoperative period | 336
discharged | 336
outpatient follow-up examination | 720
no evidence of relapse of hernia | 720