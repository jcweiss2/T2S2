59 years old | 0
male | 0
admitted to the medical intermediate unit | 0
acute progressive dyspnea | 0
new-onset ascites | 0
low albumin gradient (SAAG < 1.1 g/dL) | 0
high protein ascites | 0
type 2 diabetes | 0
hypertension | 0
old pulmonary tuberculosis | 0
end-stage renal disease | 0
no residual urine output | 0
hemodialysis three times a week | 0
triple vessel disease | 0
left ventricular ejection fraction 27% | 0
peripheral artery disease | 0
chronic limb ischemia | 0
dry gangrene | 0
left percutaneous transluminal angioplasty stent | 0
femoral artery endarterectomy | 0
dyspnea on day 3 | -72
emergency MDCT angiography | -72
right atrial thrombus (1.9 × 0.7 cm2) | -72
enoxaparin 40 mg SC OD started | -72
SC injection at abdominal wall | -72
anti-Xa level measured after 6th dose | 96
anti-Xa level 0.72 IU/mL | 96
peripheral edema | 0
ascites | 0
weight gain (6 kg) | 0
abdominal paracentesis | 0
TCC removal surgery on day 11 | 192
enoxaparin held for 4 days (day 10 to 13) | -24 to 96
bleeding in endotracheal tube | 192
enoxaparin withheld for 2 more days | 192 to 240
persistent right atrial thrombus | 192
repeated echocardiogram | 192
enoxaparin restarted 40 mg SC OD | 240
anti-Xa level after 5th dose (0.3 IU/mL) | 408
enoxaparin dose increased to 60 mg SC OD | 408
anti-Xa level 0.25 IU/mL after increased dose | 456
SC injection site switched to deltoid | 456
peak anti-Xa levels 0.45 and 0.51 IU/mL at deltoid | 504 and 672
hemodialysis | varies (see table)
vasopressor (norepinephrine) use | 0
hemodynamic instability | 0
fungemia | 0
right-side heart failure | 0
suspected DIC | 0
hypoalbuminemia | 0
enoxaparin maintained at 60 mg SC OD | 504
