70 years old | 0
male | 0
hypertension | 0
diabetes | 0
auricular fibrillation | 0
oral anticoagulation | 0
adenocarcinoma of the sigmoid colon | 0
T4aN1M0 | 0
laparoscopic exploration | 0
perforated neoplasm of the sigma | 0
infiltrating terminal ileum and right colon | 0
open surgery | 0
total oncologic colectomy | 0
ileo-rectal stapled anastomosis | 0
abdominal bleeding | -48
self-limited | -48
high dose of low molecular weight heparin (LMWH) | -48
hiccups | -48
haloperidol | -48
chlorpromazine | -48
CT scan | -24
absence of intraabdominal complication | -24
admitted to the intensive unit care | -24
fever peaks | -12
bacteraemia related to CVC | -12
inflammatory signs on the right jugular venous access | -12
cervicothoracic CT | -12
thrombus and air bubbles into the right jugular vein | -12
dilatation of an area of the vein intimately related to the phrenic nerve | -12
septic thrombosis of the jugular vein | -12
treatment with LMWH and antibiotics | 0
catheter removal | 168
discharged from the intensive care unit | 168
isolated fever peaks | 168
catheter removal | 192
3 weeks’ intravenous antibiotic cycle | 192
discharged from the hospital | 360