60 years old | 0
male | 0
admitted to the hospital | 0
severe epigastric dilation | 0
stomachache | 0
fever | 0
epigastric pain | -48
vomiting | -24
abdominal pain | -24
high fever | -24
pancreatic cancer | -336
obstructive jaundice | -336
endoscopic biliary stenting | -336
abdominal distention | 0
hepatomegaly | 0
liver span of 2 cm below the right costal margin | 0
epigastric tenderness | 0
mild rebounding pain | 0
almost no gurgling sound | 0
increased WBC count | 0
low hemoglobin | 0
low platelet count | 0
irregular gas-containing lesions in the liver | 0
liver parenchymal moth-eaten destruction | 0
pneumatized bile duct | 0
no obvious inflammation around | 0
stent in the common bile duct | 0
no obstruction | 0
severe intrahepatic infection | 0
enterogenous aerogenes | 0
multiorgan deficiency | 0
hepatic injury | 0
renal injury | 0
cardiac injury | 0
coagulopathy | 0
biapenem treatment | 0
ornidazole treatment | 0
vigorous fluid resuscitation | 0
inotropic support | 10
norepinephrine infusion | 10
blood pressure falling | 10
multiorgan failure | 20
sudden cardiac arrest | 20
death | 20
blood specimen culture | 0
gram-positive bacilli | 24
Clostridium perfringens infection | 24
phospholipase C lecithinase production | 24
hemolysis | 24
gas gangrene | 24
capillary leakage | 24
Clostridium perfringens liver abscess | 24
pneumocholangiosis | -336
ERCP | -336
bile duct stenting | -336
Vater’s ampulla damage | -336
local infection in the liver parenchyma | -336
high-dose penicillin treatment | 20
surgical debridement | 20
hyperbaric oxygen therapy | 20
deteriorated condition | 20
multiorgan insufficiency | 20
dreadful prognosis | 20