77 years old | 0
woman | 0
admitted to undergo posterior lumbar interbody fusion | 0
hypertension | 0
amlodipine | 0
carvedilol | 0
preoperative leukocyte count 7,770/ml | 0
hemoglobin level 14.1 mg/dl | 0
hematocrit 40.1% | 0
platelet count 268,000/ml | 0
chest radiography normal | 0
electrocardiogram normal | 0
physical examination normal | 0
central venous catheter inserted | -24
surgery | 0
patient arrived in operating room | 0
BP 130/90 mmHg | 0
heart rate 75 beats/min | 0
peripheral oxygen saturation 100% | 0
anesthesia induced | 0
propofol | 0
remifentanil | 0
rocuronium 50 mg administered | 0
endotracheal intubation | 0
BP 130/70 mmHg | 0
heart rate 80 beats/min | 0
right radial artery cannula inserted | 0
central venous pressure monitored | 0
FloTrac/EV1000 device used | 0
cardiac index 2.8 L/min/m2 | 0
SVR index 2,394 dynes·sec/cm5/m2 | 0
mean arterial BP 95 mmHg | 0
heart rate 77 beats/min | 0
SVV 12% | 0
central venous pressure 13 mmHg | 0
arterial blood gas analysis pH 7.455 | 0
pCO2 32.9 mmHg | 0
pO2 203.7 mmHg | 0
hematocrit 34% | 0
mean arterial BP decreased to 56 mmHg | 45
SVRI decreased to 1,932 dynes·sec/cm5/m2 | 45
phenylephrine 50 µg administered | 45
mean arterial BP increased to 123 mmHg | 47
SVRI increased to 4,254 dynes·sec/cm5/m2 | 47
nicardipine HCl 500 µg administered | 47
mean arterial BP decreased to 47–59 mmHg | 47
SVV 15% | 47
cardiac index 2.7–3.3 L/min/m2 | 47
SVRI 1,079–1,242 dynes·sec/cm5/m2 | 47
phenylephrine bolus repeated | 47
mean arterial BP not above 60 mmHg | 47
packed red blood cells transfused | 47
hemoglobin level 11.0 mg/dl | 47
hematocrit 31.5% | 47
platelet count 144,000/ml | 47
mean arterial BP 47–58 mmHg | 47
SVRI 1,097–1,550 dynes·sec/cm5/m2 | 47
cardiac index 2.2–2.8 L/min/m2 | 47
norepinephrine 0.1 µg/kg/min | 47
norepinephrine increased to 0.3 µg/kg/min | 47
mean arterial BP 60 mmHg | 47
SVRI 1,239 dynes·sec/cm5/m2 | 47
no skin rash | 47
no urticaria | 47
no change in peak airway pressure | 47
sugammadex 140 mg administered | 47
spontaneous breathing resumed | 47
patient recovered consciousness | 47
endotracheal tube removed | 47
transferred to PACU | 47
BP 82/64 mmHg | 47
HR 78 beats/min | 47
peripheral oxygen saturation 100% | 47
vasopressin initiated at 2 U/h | 47
BP increased to 104/64 mmHg | 47
BP decreased to 82/57 mmHg | 47
12-lead ECG normal | 47
transthoracic echocardiography normal | 47
left ventricular ejection fraction 65% | 47
no regional wall motion abnormality | 47
no pericardial effusion | 47
no hematoma | 47
cardiogenic shock ruled out | 47
anaphylactic shock ruled out | 47
hypovolemic shock ruled out | 47
vasoplegic syndrome diagnosed | 47
methylene blue 0.5 mg/kg administered | 47
BP increased to 112/66 mmHg | 47
vomiting occurred | 47
methylene blue discontinued | 47
total methylene blue dose 26 mg | 47
systolic BP above 110 mmHg | 47
transferred to ICU | 47
norepinephrine 0.2 µg/kg/min | 47
vasopressin 2 U/h | 47
systolic BP maintained above 110 mmHg | 24
heart rate 80 beats/min | 24
norepinephrine tapered | 24
vasopressin tapered | 24
norepinephrine stopped | 24
vasopressin stopped | 24
transferred to general ward | 48
discharged | 384
no complications | 384
