48 years old|0
male|0
Caucasian|0
chest pain (CCS III)|0
dyspnoea (NYHA III)|0
bilateral sensorineural hypacusis|0
hearing aids since age 40|0
regular heart rhythm|0
no extra heart sounds|0
blood pressure ∼115/80 mmHg|0
similar blood pressure in both arms|0
excluded uncontrolled arterial hypertension|0
electrocardiogram (ECG)|0
short PR interval (PQ 94 ms)|0
narrow QRS complex|0
inversion of T-waves in V4–V6, I, aVL|0
non-significant depression of ST segments (−0.12 mV) in I, II, aVL|0
elevated high sensitive troponin T (0.046 ng/L)|0
elevated N-terminal proBNP (252 pg/mL)|0
normal creatinine kinase (121 ng/L)|0
HbA1c 7.3 mmol/L (prediabetic)|0
slightly elevated ferritin (674 ng/mL)|0
excluded relevant iron overload|0
excluded coronary artery disease|0
symmetric non-obstructive HCM|0
diffuse reduced LVEF (48%)|0
symmetric increased myocardial wall thickness (IVS 15 mm, LVPW 14 mm)|0
LV wall thickness unexplained by physical training or valve disease|0
excluded arterial hypertension|0
LV intracavitary gradient below 30 mmHg at rest|0
LV intracavitary gradient below 30 mmHg during Valsalva manoeuver|0
increase of E/e` (17.5)|0
elevated left ventricular mass index (178 g/m²)|0
inconspicuous strain analysis|0
no typical 'apical sparing' pattern|0
global longitudinal strain −18.3%|0
normal right ventricle diameter and function|0
TAPSE 27 mm|0
cardiac MRI confirmed mildly reduced LV function (LVEF 48%)|0
LV end-diastolic volume 170 mL|0
LV end-systolic volume 88 mL|0
cardiac index 2.94 L/min/m2|0
RV wall thickness 3 mm|0
RV end-diastolic volume 130 mL|0
RV end-systolic volume 51 mL|0
RV cardiac index 2.85 L/min/m2|0
myocardial fibrosis detected by late gadolinium enhancement (LGE)|0
LGE predominantly mid-myocardial and epicardial|0
progressive myocardial fibrosis|0
ruled out cardiac amyloidosis|0
negative genetic testing for sarcomeric genes (MYBPC3, MYH7, TNNT2, TNNI3)|0
endomyocardial biopsy (EMB)|0
hypertrophy of cardiomyocytes|0
diffuse fibrosis|0
excluded infiltrative or active inflammatory disease|0
excluded storage diseases|0
normal α-D-galactosidase-A activity (0.150 mU/mL)|0
negative next-generation sequencing (NGS) for sarcomeric genes|0
advanced genetic testing|0
m.3243A > G mutation in 25% of mitochondrial DNA|0
no ventricular tachycardia on Holter monitoring|0
estimated 5-year SCD risk 2.43%|0
ICD not recommended|0
family members with m.3243A > G mutation|0
clinical screening of family members|0
father (KS) with ischemic cardiomyopathy (iCM)|0
mother (EM) with dilative cardiomyopathy (DCM)|0
half-brother (JF) with DCM|0
half-brother (KF) with HCM|0
sister (MS) with m.3243A > G mutation|0
half-nephews (Je, Mo) with m.3243A > G mutation|0
mother (EM) died from sepsis-induced multiple organ dysfunction syndrome|0
JF died suddenly at 53|0
KF's HCM diagnosed in 2013|0
KF's LVEF 28% in 2019|0
KF's ICD terminated ventricular tachycardia in 2016|0
KF's QRS broadened into left branch bundle block (161 ms)|0
KF's ICD upgraded to CRT-D|0
index patient's symptoms unchanged at 6-month follow-up|0
LV wall thickness unchanged|0
LVEF unchanged|0
estimated 5-year SCD risk 2.27%|0
ICD not recommended at follow-up|0
heart failure medications intended to improve symptoms|0
next follow-up scheduled at 3 months|0
m.3243A > G mutation associated with mitochondrial disorder|0
maternally inherited diabetes and deafness (MIDD)|0
hearing loss before diabetes|0
progression of myocardial fibrosis and scarring|0
recommendations for repeated cardiac MRIs every 3–5 years|0
intra-familial phenotypic cardiomyopathy variability|0
heterogeneous cardiomyopathies in family members|0
chest pain and dyspnoea in 2012 (42 years old)|0
TTE diagnosis of non-obstructive HCM in 2012|0
chest pain and dyspnoea in 2015 (45 years old)|0
cardiac MRI and genetic testing for sarcomeric genes in 2015|0
chest pain and dyspnoea in 2018 (48 years old)|0
cardiac MRI and coronary angiography in 2018|0
myocardial biopsy in 2018|0
advanced genetic testing in 06/2019|0
clinical and genetic screening of family members in 10/2019|0
hearing loss in 2000 (30 years old)|0
bilateral hearing aids in 2010 (40 years old)|0
mother (EM) heart failure diagnosis in 1988 (52 years old)|0
LV dysfunction and dilatation in 1988|0
LV thrombus in 1988|0
cardioembolic stroke in 1988|0
sepsis-induced multiple organ dysfunction syndrome in 1988|0
KF's HCM diagnosis in 2013|0
KF's initial ECG findings in 2013|0
KF's LVEF 28% in 2013|0
KF's coronary angiography in 2016|0
KF's ICD termination of ventricular tachycardia in 2016|0
KF's QRS broadening over time|0
KF's CRT-D upgrade|0
index patient's follow-up in 06/2019|0
scheduled follow-up in outpatient clinic|0
