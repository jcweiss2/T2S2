29 years old | 0
male | 0
lumberjack | 0
alcohol consumer | 0
fever | -336
cough | -336
septic shock | 0
confused state | 0
Glasgow Coma Scale E4V2M5 | 0
temperature 38.0°C | 0
blood pressure 85/42 mmHg | 0
pulse rate 135 b.p.m | 0
neck stiffness | 0
bilateral upper and lower limbs power 3 | 0
normal heart sounds | 0
bilateral lung crepitations | 0
fluid resuscitation | 0
vasopressor | 0
mechanical ventilator | 0
anaemia | 0
thrombocytopenia | 0
normal total white cells | 0
normal renal function | 0
splenic microabscesses | 0
bilateral lung fields consolidation | 0
normal CT brain | 0
no cerebrospinal fluid inflammation | 0
B. pseudomallei in blood culture | 0
IV ceftazidime | 0
IV C-penicillin | 0
IV noradrenaline | 0
ventilator-associated pneumonia | 72
multidrug-resistant Acinetobacter baumanii | 72
IV imipenem | 96
high-grade temperature | 96
leukopenia | 96
oral trimethoprim-sulfamethoxazole | 168
sepsis-induced supraventricular tachycardia | 168
left-sided hemiparesis | 504
pansystolic murmur | 504
thrills at the apex of the heart | 504
right corona radiata infarct | 504
high parietal petechia haemorrhage | 504
thickened mitral valve | 504
oscillating mass at the posterior mitral valve leaflet | 504
moderate eccentric mitral regurgitation | 504
IV gentamicin | 504
intensive phase therapy for 6 weeks | 504
eradication phase therapy | 1008
discharged | 1008
minimal residual left sided weakness | 1008
Modified Rankin Score of 2 | 1008
follow-up at 9 months | 1944
vegetation on mitral valve resolved | 1944
residual moderate mitral regurgitation | 1944
left ventricular ejection fraction of 66.5% | 1944
Modified Rankin Score of 2 | 1944