17 years old | 0 | 0 
male | 0 | 0 
Caucasian | 0 | 0 
admitted to the hospital | 0 | 0 
throat pain | -168 | 0 
odynophagia | -168 | 0 
blood tests | 0 | 0 
Hemoglobin: 7.0 g/dL | 0 | 0 
Hematocrit: 21% | 0 | 0 
WBC: 33 x 10^9 cells/L | 0 | 0 
platelets: 38 x 10^9 cells/L | 0 | 0 
Acute promyelocytic leukemia (M3) | 0 | 0 
daunorubicin plus vesanoid | 0 | 0 
necrotic lesion in the M. palatoglossus | 0 | 0 
necrotic lesion in the soft palate | 0 | 0 
necrotic lesion in the uvula | 0 | 0 
necrotic lesion in the right tonsil | 0 | 0 
unpleasant odor | 0 | 0 
biopsy | 0 | 0 
culture | 0 | 0 
nonspecific chronic diffuse inflammation | 0 | 0 
necrotic areas | 0 | 0 
numerous bacteria | 0 | 0 
Enterococcus spp | 0 | 0 
Staphylococcus aureus | 0 | 0 
Candida SP | 0 | 0 
noma-like lesion | 0 | 0 
antibiotic therapy | 0 | 0 
ceftazidime | 0 | 0 
amicacin | 0 | 0 
vancomycin | 0 | 0 
fluconazole | 0 | 0 
penicillin G | 0 | 0 
pneumonia | 0 | 45 
sepsis | 0 | 45 
intensive care unit | 0 | 45 
total recovery | 45 | 45 
extensive loss of soft palate tissue | 45 | 45 
mucocutaneous leishmaniasis | 0 | 0 
lupus erythematosus | 0 | 0 
leprosy | 0 | 0 
agranulocytic ulcerations | 0 | 0 
physical trauma | 0 | 0 
syphilis | 0 | 0 
oral cancer | 0 | 0 
yaws | 0 | 0 
infections of the oral cavity | 0 | 0 
early diagnosis | 0 | 0 
accurate diagnosis | 0 | 0 
treatment | 0 | 45 
conflict-of-interest disclosure | 0 | 0 
no competing financial interest | 0 | 0