36 years old | 0
female | 0
pregnant | 0
admitted to the hospital | 0
severe pre-eclampsia | 0
obesity class 3 | 0
oligohydramnios | 0
intrauterine growth restriction | 0
COVID-19 | -672
estimated fetal weight 2200 g | 0
attended 10 regular antenatal visits | -672
blood pressure normal | -672
blood pressure 170/110 mm Hg | -24
urinary protein +2 | -24
MgSO4 treatment | 0
IgG antibody to SARS-CoV-2 reactive | 0
chest radiograph normal | 0
reverse transcription PCR test for SARS-CoV-2 | 0
fetal well-being tests abnormal | 0
non-stress test low variability and late deceleration | 0
caesarean section | 0
sterilisation | 0
meconium-stained amniotic fluid | 0
baby born with birth weight 2190 g | 0
Apgar scores 7 and 8 | 0
maternal COVID-19 molecular test negative | 24
maternal condition deteriorated | 24
fluid resuscitation | 24
severe anaemia | 48
exploratory laparotomy | 72
Couvelaire uterus | 72
haematoma in the left adnexa | 72
supracervical hysterectomy | 72
total blood loss 1200 mL | 72
fluid input 2300 mL | 72
whole blood transfusion | 72
ventilator support | 72
oxygen saturation 97%-100% | 72
GCS E4VxM6 | 72
anaemia | 72
hypoalbuminaemia | 72
thrombocytopenia | 72
hyponatraemia | 72
hypokalaemia | 72
non-steroidal anti-inflammatory drugs | 72
ceftriaxon | 72
albumin | 72
packed red cell transfusion | 72
serum electrolyte correction | 72
rhonchi detected | 96
pulmonary oedema suspected | 96
furosemide | 96
intravenous meropenem | 96
SARS-CoV-2 molecular test positive | 168
COVID-19 pneumonia | 168
bacterial pneumonia | 168
remdesivir | 168
isosorbide dinitrate | 168
nicardipine | 168
ventilator maintained | 168
unstable respiratory function | 168
oxygenation parameter | 168
NRBM | 192
oxygen saturation 97%-98% | 192
heparin | 216
D-dimer levels increased | 216
fever | 216
antipyretics | 216
incisional wound bleeding | 264
wound care | 264
convalescent plasma transfusion | 264
ultrasound | 264
haematoma superficial to fascia | 264
heparin stopped | 312
incisional site bleeding stopped | 312
RT-PCR results negative | 360
blood culture showed Enterococcus gallinarum | 432
antibiotics changed | 432
levofloxacin | 432
ciprofloxacin | 432
patient's condition improved | 576
stable vital signs | 576
incisional wound healed | 576
discharged | 600