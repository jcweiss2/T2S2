32 years old | 0
male | 0
presented to the emergency department | 0
fracture of the right sacroiliac joint | 0
open wound of right tibial fracture |8
elective surgery |0
sacroiliac disruption |0
pubic diastasis |0
high-grade fever (102°F) |72
tachycardia |72
hypotension |72
increasing pain |72
progressive swelling |72
erythema |72
crepitus over the right calf leg |72
unable to move his right lower extremity |72
no sensation below the knee joint level |72
severely swollen |72
brownish skin of the right lower extremity |72
necrotic wound along the fracture site |72
foul smelling wound |72
X-ray gas in the interfacial planes |72
extensive gas formation throughout all the muscle compartments |72
increased total leukocyte counts (TLCs) (24, 270/cubic mm3) |72
erythrocyte sedimentation rate (122 mm/h) |72
C-reactive-protein (17.13 mg/dl) |72
presumptive diagnosis of gas gangrene |72
emergency surgical debridement |72
wound debrided extensively |72
pus pockets removed |72
necrosed medial gastrocnemius muscle debrided |72
tissue and pus sample sent for gram-stain and culture |72
Gram-positive rods in the smear |72
anaerobic blood agar plate growth |72
identified as C. sordelli |72
started clindamycin 300 mg |72
started linezolid 600 mg |72
antibiotics deescalated |72
started metronidazole 750 mg |72
started clindamycin 300 mg intravenously |72
improved after 48 h |120
six sittings of hyperbaric oxygen therapy (HOBT) |120
wound healed well |480
repeated pus culture sterile |240
discharged |480
