79 years old | 0 | 0 
male | 0 | 0 
hypertension | 0 | 0 
ischemic heart disease | 0 | 0 
admitted to the hospital | 0 | 0 
severe symptomatic aortic stenosis | 0 | 0 
coronary artery bypass graft surgery | -7920 | -7920 
mitral valve repair | -7920 | -7920 
preprocedural transthoracic echocardiography | -1 | 0 
severe aortic stenosis | -1 | 0 
left ventricular ejection fraction of 45% | -1 | 0 
induction of general anesthesia | 0 | 0 
TEE probe insertion | 0 | 0 
SAPIEN 3 valve deployment | 0 | 1 
postprocedural TEE | 1 | 1 
prosthesis in good position | 1 | 1 
no visible paravalvular leak | 1 | 1 
gastric aspiration | 1 | 1 
blood-tinged secretions | 1 | 1 
extubation | 1 | 1 
transferred to the intensive care unit | 1 | 1 
progressive chest pain | 2 | 2 
shivering | 2 | 2 
computed tomography | 2 | 2 
pneumomediastinum | 2 | 2 
right hydropneumothorax | 2 | 2 
esophageal perforation suspected | 2 | 2 
right thoracic drain insertion | 2 | 2 
serosanguinous liquid drained | 2 | 2 
esophagogastroscopy | 2 | 2 
4-cm vertical perforation of the middle third of the esophagus | 2 | 2 
right thoracotomy | 7 | 7 
repair of esophageal perforation | 7 | 7 
primary closure of the esophageal wall | 7 | 7 
intercostal muscular flap mobilized | 7 | 7 
thoracic drains left in place | 7 | 7 
transferred to the intensive care unit | 7 | 7 
pneumonia | 7 | 720 
severe delirium | 7 | 720 
congestive heart failure | 7 | 720 
pulmonary edema | 7 | 720 
withdrawal of care | 720 | 720 
died | 720 | 720 
prominent anterior thoracic osteophytes | -1 | 0 
vertebral osteophytes compressing the esophagus | -1 | 0 
anatomic proximity of thoracic osteophytes to the esophagus | -1 | 0 
esophageal laceration | 0 | 1 
transesophageal probe manipulation | 0 | 1 
esophageal perforation | 1 | 2 
esophageal injury | 1 | 2 
repeated insertion and withdrawal of the probe | 0 | 1 
extensive transesophageal probe manipulation | 0 | 1 
preoperative imaging | -1 | 0 
chest CT | -1 | 0 
vertebral osteophytes | -1 | 0 
anatomic relation to the esophagus | -1 | 0 
safe performance of TEE | 0 | 0 
relative contraindication to TEE | 0 | 0 
elderly patients | 0 | 0 
interventional cardiologic procedures | 0 | 0 
general anesthesia | 0 | 0 
MitralClip implantation | 0 | 0 
left atrial appendage occlusion | 0 | 0 
guide catheter–based procedures | 0 | 0 
probe manipulations | 0 | 1 
repeated motion | 0 | 1 
esophageal injury | 0 | 1 
procedural duration | 0 | 1 
contributing factor | 0 | 1 
preoperative pulmonary radiography | -1 | 0 
CT | -1 | 0 
anatomic proximity of thoracic osteophytes to the esophagus | -1 | 0 
safe performance of TEE | 0 | 0 
routine investigation | -1 | 0 
chest CT | -1 | 0 
vertebral osteophytes | -1 | 0 
anatomic relation to the esophagus | -1 | 0 
esophageal perforation | 1 | 2 
iatrogenic esophageal perforation | 1 | 2 
transesophageal echocardiography | 0 | 1 
rare event | 0 | 0 
high mortality rate | 0 | 0 
incidence | 0 | 0 
complication | 1 | 2 
adverse effect | 1 | 2 
adverse event | 1 | 2 
laceration | 1 | 2 
rupture | 1 | 2 
tear | 1 | 2 
injury | 1 | 2 
perforation | 1 | 2 
osteophyte | -1 | 0 
hyperostosis | -1 | 0 
exostoses | -1 | 0 
diffuse idiopathic skeletal hyperostosis | -1 | 0 
spine | -1 | 0 
vertebral column | -1 | 0 
preexisting esophageal pathologies | 0 | 0 
esophageal stricture | 0 | 0 
Zenker's diverticulum | 0 | 0 
fibrosis | 0 | 0 
prior chest radiation | 0 | 0 
ulceration | 0 | 0 
medication | 0 | 0 
severe cardiomegaly | 0 | 0 
large calcified lymph nodes | 0 | 0 
mechanical compression | 0 | 1 
mucosal and muscular fibers | 0 | 1 
esophagus | 0 | 1 
vertebral osteophytes | -1 | 0 
common radiologic findings | -1 | 0 
elderly population | -1 | 0 
diffuse idiopathic skeletal hyperostosis | -1 | 0 
dysphagia | -1 | 0 
aspiration | -1 | 0 
anterior cervical osteophytes | -1 | 0 
thoracic region | -1 | 0 
tracheal bifurcation | -1 | 0 
diaphragmatic hiatus | -1 | 0 
anatomic space | -1 | 0 
vertebral column | -1 | 0 
esophagus | -1 | 0 
symptoms | -1 | 0 
extrinsic esophageal compression | -1 | 0 
lower thoracic region | -1 | 0 
supine position | -1 | 0 
weight of thoracic organs | -1 | 0 
esophagus | -1 | 0 
osteophytes | -1 | 0 
preoperative imaging | -1 | 0 
chest CT | -1 | 0 
anatomic proximity of thoracic osteophytes to the esophagus | -1 | 0 
safe performance of TEE | 0 | 0 
relative contraindication to TEE | 0 | 0 
elderly patients | 0 | 0 
interventional cardiologic procedures | 0 | 0 
general anesthesia | 0 | 0 
MitralClip implantation | 0 | 0 
left atrial appendage occlusion | 0 | 0 
guide catheter–based procedures | 0 | 0 
probe manipulations | 0 | 1 
repeated motion | 0 | 1 
esophageal injury | 0 | 1 
procedural duration | 0 | 1 
contributing factor | 0 | 1 
preoperative pulmonary radiography | -1 | 0 
CT | -1 | 0 
anatomic proximity of thoracic osteophytes to the esophagus | -1 | 0 
safe performance of TEE | 0 | 0 
routine investigation | -1 | 0 
chest CT | -1 | 0 
vertebral osteophytes | -1 | 0 
anatomic relation to the esophagus | -1 | 0 
esophageal perforation | 1 | 2 
iatrogenic esophageal perforation | 1 | 2 
transesophageal echocardiography | 0 | 1 
rare event | 0 | 0 
high mortality rate | 0 | 0 
incidence | 0 | 0 
complication | 1 | 2 
adverse effect | 1 | 2 
adverse event | 1 | 2 
laceration | 1 | 2 
rupture | 1 | 2 
tear | 1 | 2 
injury | 1 | 2 
perforation | 1 | 2 
osteophyte | -1 | 0 
hyperostosis | -1 | 0 
exostoses | -1 | 0 
diffuse idiopathic skeletal hyperostosis | -1 | 0 
spine | -1 | 0 
vertebral column | -1 | 0 
preexisting esophageal pathologies | 0 | 0 
esophageal stricture | 0 | 0 
Zenker's diverticulum | 0 | 0 
fibrosis | 0 | 0 
prior chest radiation | 0 | 0 
ulceration | 0 | 0 
medication | 0 | 0 
severe cardiomegaly | 0 | 0 
large calcified lymph nodes | 0 | 0 
mechanical compression | 0 | 1 
mucosal and muscular fibers | 0 | 1 
esophagus | 0 | 1 
vertebral osteophytes | -1 | 0 
common radiologic findings | -1 | 0 
elderly population | -1 | 0 
diffuse idiopathic skeletal hyperostosis | -1 | 0 
dysphagia | -1 | 0 
aspiration | -1 | 0 
anterior cervical osteophytes | -1 | 0 
thoracic region | -1 | 0 
tracheal bifurcation | -1 | 0 
diaphragmatic hiatus | -1 | 0 
anatomic space | -1 | 0 
vertebral column | -1 | 0 
esophagus | -1 | 0 
symptoms | -1 | 0 
extrinsic esophageal compression | -1 | 0 
lower thoracic region | -1 | 0 
supine position | -1 | 0 
weight of thoracic organs | -1 | 0 
esophagus | -1 | 0 
osteophytes | -1 | 0 
preoperative imaging | -1 | 0 
chest CT | -1 | 0 
anatomic proximity of thoracic osteophytes to the esophagus | -1 | 0 
safe performance of TEE | 0 | 0 
relative contraindication to TEE | 0 | 0 
elderly patients | 0 | 0 
interventional cardiologic procedures | 0 | 0 
general anesthesia | 0 | 0 
MitralClip implantation | 0 | 0 
left atrial appendage occlusion | 0 | 0 
guide catheter–based procedures | 0 | 0 
probe manipulations | 0 | 1 
repeated motion | 0 | 1 
esophageal injury | 0 | 1 
procedural duration | 0 | 1 
contributing factor | 0 | 1 
preoperative pulmonary radiography | -1 | 0 
CT | -1 | 0 
anatomic proximity of thoracic osteophytes to the esophagus | -1 | 0 
safe performance of TEE | 0 | 0 
routine investigation | -1 | 0 
chest CT | -1 | 0 
vertebral osteophytes | -1 | 0 
anatomic relation to the esophagus | -1 | 0 
esophageal perforation | 1 | 2 
iatrogenic esophageal perforation | 1 | 2 
transesophageal echocardiography | 0 | 1 
rare event | 0 | 0 
high mortality rate | 0 | 0 
incidence | 0 | 0 
complication | 1 | 2 
adverse effect | 1 | 2 
adverse event | 1 | 2 
laceration | 1 | 2 
rupture | 1 | 2 
tear | 1 | 2 
injury | 1 | 2 
perforation | 1 | 2 
osteophyte | -1 | 0 
hyperostosis | -1 | 0 
exostoses | -1 | 0 
diffuse idiopathic skeletal hyperostosis | -1 | 0 
spine | -1 | 0 
vertebral column | -1 | 0 
preexisting esophageal pathologies | 0 | 0 
esophageal stricture | 0 | 0 
Zenker's diverticulum | 0 | 0 
fibrosis | 0 | 0 
prior chest radiation | 0 | 0 
ulceration | 0 | 0 
medication | 0 | 0 
severe cardiomegaly | 0 | 0 
large calcified lymph nodes | 0 | 0 
mechanical compression | 0 | 1 
mucosal and muscular fibers | 0 | 1 
esophagus | 0 | 1 
vertebral osteophytes | -1 | 0 
common radiologic findings | -1 | 0 
elderly population | -1 | 0 
diffuse idiopathic skeletal hyperostosis | -1 | 0 
dysphagia | -1 | 0 
aspiration | -1 | 0 
anterior cervical osteophytes | -1 | 0 
thoracic region | -1 | 0 
tracheal bifurcation | -1 | 0 
diaphragmatic hiatus | -1 | 0 
anatomic space | -1 | 0 
vertebral column | -1 | 0 
esophagus | -1 | 0 
symptoms | -1 | 0 
extrinsic esophageal compression | -1 | 0 
lower thoracic region | -1 | 0 
supine position | -1 | 0 
weight of thoracic organs | -1 | 0 
esophagus | -1 | 0 
osteophytes | -1 | 0 
preoperative imaging | -1 | 0 
chest CT | -1 | 0 
anatomic proximity of thoracic osteophytes to the esophagus | -1 | 0 
safe performance of TEE | 0 | 0 
relative contraindication to TEE | 0 | 0 
elderly patients | 0 | 0 
interventional cardiologic procedures | 0 | 0 
general anesthesia | 0 | 0 
MitralClip implantation | 0 | 0 
left atrial appendage occlusion | 0 | 0 
guide catheter–based procedures | 0 | 0 
probe manipulations | 0 | 1 
repeated motion | 0 | 1 
esophageal injury | 0 | 1 
procedural duration | 0 | 1 
contributing factor | 0 | 1 
preoperative pulmonary radiography | -1 | 0 
CT | -1 | 0 
anatomic proximity of thoracic osteophytes to the esophagus | -1 | 0 
safe performance of TEE | 0 | 0 
routine investigation | -1 | 0 
chest CT | -1 | 0 
vertebral osteophytes | -1 | 0 
anatomic relation to the esophagus | -1 | 0 
esophageal perforation | 1 | 2 
iatrogenic esophageal perforation | 1 | 2 
transesophageal echocardiography | 0 | 1 
rare event | 0 | 0 
high mortality rate | 0 | 0 
incidence | 0 | 0 
complication | 1 | 2 
adverse effect | 1 | 2 
adverse event | 1 | 2 
laceration | 1 | 2 
rupture | 1 | 2 
tear | 1 | 2 
injury | 1 | 2 
perforation | 1 | 2 
osteophyte | -1 | 0 
hyperostosis | -1 | 0 
exostoses | -1 | 0 
diffuse idiopathic skeletal hyperostosis | -1 | 0 
spine | -1 | 0 
vertebral column | -1 | 0 
preexisting esophageal pathologies | 0 | 0 
esophageal stricture | 0 | 0 
Zenker's diverticulum | 0 | 0 
fibrosis | 0 | 0 
prior chest radiation | 0 | 0 
ulceration | 0 | 0 
medication | 0 | 0 
severe cardiomegaly | 0 | 0 
large calcified lymph nodes | 0 | 0 
mechanical compression | 0 | 1 
mucosal and muscular fibers | 0 | 1 
esophagus | 0 | 1 
vertebral osteophytes | -1 | 0 
common radiologic findings | -1 | 0 
elderly population | -1 | 0 
diffuse idiopathic skeletal hyperostosis | -1 | 0 
dysphagia | -1 | 0 
aspiration | -1 | 0 
anterior cervical osteophytes | -1 | 0 
thoracic region | -1 | 0 
tracheal bifurcation | -1 | 0 
diaphragmatic hiatus | -1 | 0 
anatomic space | -1 | 0 
vertebral column | -1 | 0 
esophagus | -1 | 0 
symptoms | -1 | 0 
extrinsic esophageal compression | -1 | 0 
lower thoracic region | -1 | 0 
supine position | -1 | 0 
weight of thoracic organs | -1 | 0 
esophagus | -1 | 0 
osteophytes | -1 | 0 
preoperative imaging | -1 | 0 
chest CT | -1 | 0 
anatomic proximity of thoracic osteophytes to the esophagus | -1 | 0 
safe performance of TEE | 0 | 0 
relative contraindication to TEE | 0 | 0 
elderly patients | 0 | 0 
interventional cardiologic procedures | 0 | 0 
general anesthesia | 0 | 0 
MitralClip implantation | 0 | 0 
left atrial appendage occlusion | 0 | 0 
guide catheter–based procedures | 0 | 0 
probe manipulations | 0 | 1 
repeated motion | 0 | 1 
esophageal injury | 0 | 1 
procedural duration | 0 | 1 
contributing factor | 0 | 1 
preoperative pulmonary radiography | -1 | 0 
CT | -1 | 0 
anatomic proximity of thoracic osteophytes to the esophagus | -1 | 0 
safe performance of TEE | 0 | 0 
routine investigation | -1 | 0 
chest CT | -1 | 0 
vertebral osteophytes | -1 | 0 
anatomic relation to the esophagus | -1 | 0 
esophageal perforation | 1 | 2 
iatrogenic esophageal perforation | 1 | 2 
transesophageal echocardiography | 0 | 1 
rare event | 0 | 0 
high mortality rate | 0 | 0 
incidence | 0 | 0 
complication | 1 | 2 
adverse effect | 1 | 2 
adverse event | 1 | 2 
laceration | 1 | 2 
rupture | 1 | 2 
tear | 1 | 2 
injury | 1 | 2 
perforation | 1 | 2 
osteophyte | -1 | 0 
hyperostosis | -1 | 0 
exostoses | -1 | 0 
diffuse idiopathic skeletal hyperostosis | -1 | 0 
spine | -1 | 0 
vertebral column | -1 | 0 
preexisting esophageal pathologies | 0 | 0 
esophageal stricture | 0 | 0 
Zenker's diverticulum | 0 | 0 
fibrosis | 0 | 0 
prior chest radiation | 0 | 0 
ulceration | 0 | 0 
medication | 0 | 0 
severe cardiomegaly | 0 | 0 
large calcified lymph nodes | 0 | 0 
mechanical compression | 0 | 1 
mucosal and muscular fibers | 0 | 1 
esophagus | 0 | 1 
vertebral osteophytes | -1 | 0 
common radiologic findings | -1 | 0 
elderly population | -1 | 0 
diffuse idiopathic skeletal hyperostosis | -1 | 0 
dysphagia | -1 | 0 
aspiration | -1 | 0 
anterior cervical osteophytes | -1 | 0 
thoracic region | -1 | 0 
tracheal bifurcation | -1 | 0 
diaphragmatic hiatus | -1 | 0 
anatomic space | -1 | 0 
vertebral column | -1 | 0 
esophagus | -1 | 0 
symptoms | -1 | 0 
extrinsic esophageal compression | -1 | 0 
lower thoracic region | -1 | 0 
supine position | -1 | 0 
weight of thoracic organs | -1 | 0 
esophagus | -1 | 0 
osteophytes | -1 | 0 
preoperative imaging | -1 | 0 
chest CT | -1 | 0 
anatomic proximity of thoracic osteophytes to the esophagus | -1 | 0 
safe performance of TEE | 0 | 0 
relative contraindication to TEE | 0 | 0 
elderly patients | 0 | 0 
interventional cardiologic procedures | 0 | 0 
general anesthesia | 0 | 0 
MitralClip implantation | 0 | 0 
left atrial appendage occlusion | 0 | 0 
guide catheter–based procedures | 0 | 0 
probe manipulations | 0 | 1 
repeated motion | 0 | 1 
esophageal injury | 0 | 1 
procedural duration | 0 | 1 
contributing factor | 0 | 1 
preoperative pulmonary radiography | -1 | 0 
CT | -1 | 0 
anatomic proximity of thoracic osteophytes to the esophagus | -1 | 0 
safe performance of TEE | 0 | 0 
routine investigation | -1 | 0 
chest CT | -1 | 0 
vertebral osteophytes | -1 | 0 
anatomic relation to the esophagus | -1 | 0 
esophageal perforation | 1 | 2 
iatrogenic esophageal perforation | 1 | 2 
transesophageal echocardiography | 0 | 1 
rare event | 0 | 0 
high mortality rate | 0 | 0 
incidence | 0 | 0 
complication | 1 | 2 
adverse effect | 1 | 2 
adverse event | 1 | 2 
laceration | 1 | 2 
rupture | 1 | 2 
tear | 1 | 2 
injury | 1 | 2 
perforation | 1 | 2 
osteophyte | -1 | 0 
hyperostosis | -1 | 0 
exostoses | -1 | 0 
diffuse idiopathic skeletal hyperostosis | -1 | 0 
spine | -1 | 0 
vertebral column | -1 | 0 
preexisting esophageal pathologies | 0 | 0 
esophageal stricture | 0 | 0 
Zenker's diverticulum | 0 | 0 
fibrosis | 0 | 0 
prior chest radiation | 0 | 0 
ulceration | 0 | 0 
medication | 0 | 0 
severe cardiomegaly | 0 | 0 
large calcified lymph nodes | 0 | 0 
mechanical compression | 0 | 1 
mucosal and muscular fibers | 0 | 1 
esophagus | 0 | 1 
vertebral osteophytes | -1 | 0 
common radiologic findings | -1 | 0 
elderly population | -1 | 0 
diffuse idiopathic skeletal hyperostosis | -1 | 0 
dysphagia | -1 | 0 
aspiration | -1 | 0 
anterior cervical osteophytes | -1 | 0 
thoracic region | -1 | 0 
tracheal bifurcation | -1 | 0 
diaphragmatic hiatus | -1 | 0 
anatomic space | -1 | 0 
vertebral column | -1 | 0 
esophagus | -1 | 0 
symptoms | -1 | 0 
extrinsic esophageal compression | -1 | 0 
lower thoracic region | -1 | 0 
supine position | -1 | 0 
weight of thoracic organs | -1 | 0 
esophagus | -1 | 0 
osteophytes | -1 | 0 
preoperative imaging | -1 | 0 
chest CT | -1 | 0 
anatomic proximity of thoracic osteophytes to the esophagus | -1 | 0 
safe performance of TEE | 0 | 0 
relative contraindication to TEE | 0 | 0 
elderly patients | 0 | 0 
interventional cardiologic procedures | 0 | 0 
general anesthesia | 0 | 0 
MitralClip implantation | 0 | 0 
left atrial appendage occlusion | 0 | 0 
guide catheter–based procedures | 0 | 0 
probe manipulations | 0 | 1 
repeated motion | 0 | 1 
esophageal injury | 0 | 1 
procedural duration | 0 | 1 
contributing factor | 0 | 1 
preoperative pulmonary radiography | -1 | 0 
CT | -1 | 0 
anatomic proximity of thoracic osteophytes to the esophagus | -1 | 0 
safe performance of TEE | 0 | 0 
routine investigation | -1 | 0 
chest CT | -1 | 0 
vertebral osteophytes | -1 | 0 
anatomic relation to the esophagus | -1 | 0 
esophageal perforation | 1 | 2 
iatrogenic esophageal perforation | 1 | 2 
transesophageal echocardiography | 0 | 1 
rare event | 0 | 0 
high mortality rate | 0 | 0 
incidence | 0 | 0 
complication | 1 | 2 
adverse effect | 1 | 2 
adverse event | 1 | 2 
laceration | 1 | 2 
rupture | 1 | 2 
tear | 1 | 2 
injury | 1 | 2 
perforation | 1 | 2 
osteophyte | -1 | 0 
hyperostosis | -1 | 0 
exostoses | -1 | 0 
diffuse idiopathic skeletal hyperostosis | -1 | 0 
spine | -1 | 0 
vertebral column | -1 | 0 
preexisting esophageal pathologies | 0 | 0 
esophageal stricture | 0 | 0 
Zenker's diverticulum | 0 | 0 
fibrosis | 0 | 0 
prior chest radiation | 0 | 0 
ulceration | 0 | 0 
medication | 0 | 0 
severe cardiomegaly | 0 | 0 
large calcified lymph nodes | 0 | 0 
mechanical compression | 0 | 1 
mucosal and muscular fibers | 0 | 1 
esophagus | 0 | 1 
vertebral osteophytes | -1 | 0 
common radiologic findings | -1 | 0 
elderly population | -1 | 0 
diffuse idiopathic skeletal hyperostosis | -1 | 0 
dysphagia | -1 | 0 
aspiration | -1 | 0 
anterior cervical osteophytes | -1 | 0 
thoracic region | -1 | 0 
tracheal bifurcation | -1 | 0 
diaphragmatic hiatus | -1 | 0 
anatomic space | -1 | 0 
vertebral column | -1 | 0 
esophagus | -1 | 0 
symptoms | -1 | 0 
extrinsic esophageal compression | -1 | 0 
lower thoracic region | -1 | 0 
supine position | -1 | 0 
weight of thoracic organs | -1 | 0 
esophagus | -1 | 0 
osteophytes | -1 | 0 
preoperative imaging | -1 | 0 
chest CT | -1 | 0 
anatomic proximity of thoracic osteophytes to the esophagus | -1 | 0 
safe performance of TEE | 0 | 0 
relative contraindication to TEE | 0 | 0 
elderly patients | 0 | 0 
interventional cardiologic procedures | 0 | 0 
general anesthesia | 0 | 0 
MitralClip implantation | 0 | 0 
left atrial appendage occlusion | 0 | 0 
guide catheter–based procedures | 0 | 0 
probe manipulations | 0 | 1 
repeated motion | 0 | 1 
esophageal injury | 0 | 1 
procedural duration | 0 | 1 
contributing factor | 0 | 1 
preoperative pulmonary radiography | -1 | 0 
CT | -1 | 0 
anatomic proximity of thoracic osteophytes to the esophagus | -1 | 0 
safe performance of TEE | 0 | 0 
routine investigation | -1 | 0 
chest CT | -1 | 0 
vertebral osteophytes | -1 | 0 
anatomic relation to the esophagus | -1 | 0 
esophageal perforation | 1 | 2 
iatrogenic esophageal perforation | 1 | 2 
transesophageal echocardiography | 0 | 1 
rare event | 0 | 0 
high mortality rate | 0 | 0 
incidence | 0 | 0 
complication | 1 | 2 
adverse effect | 1 | 2 
adverse event | 1 | 2 
laceration | 1 | 2 
rupture | 1 | 2 
tear | 1 | 2 
injury | 1 | 2 
perforation | 1 | 2 
osteophyte | -1 | 0 
hyperostosis | -1 | 0 
exostoses | -1 | 0 
diffuse idiopathic skeletal hyperostosis | -1 | 0 
spine | -1 | 0 
vertebral column | -1 | 0 
preexisting esophageal pathologies | 0 | 0 
esophageal stricture | 0 | 0 
Zenker's diverticulum | 0 | 0 
fibrosis | 0 | 0 
prior chest radiation | 0 | 0 
ulceration | 0 | 0 
medication | 0 | 0 
severe cardiomegaly | 0 | 0 
large calcified lymph nodes | 0 | 0 
mechanical compression | 0 | 1 
mucosal and muscular fibers | 0 | 1 
esophagus | 0 | 1 
vertebral osteophytes | -1 | 0 
common radiologic findings | -1 | 0 
elderly population | -1 | 0 
diffuse idiopathic skeletal hyperostosis | -1 | 0 
dysphagia | -1 | 0 
aspiration | -1 | 0 
anterior cervical osteophytes | -1 | 0 
thoracic region | -1 | 0 
tracheal bifurcation | -1 | 0 
diaphragmatic hiatus | -1 | 0 
anatomic space | -1 | 0 
vertebral column | -1 | 0 
esophagus | -1 | 0 
symptoms | -1 | 0 
extrinsic esophageal compression | -1 | 0 
lower thoracic region | -1 | 0 
supine position | -1 | 0 
weight of thoracic organs | -1 | 0 
esophagus | -1 | 0 
osteophytes | -1 | 0 
preoperative imaging | -1 | 0 
chest CT | -1 | 0 
anatomic proximity of thoracic osteophytes to the esophagus | -1 | 0 
safe performance of TEE | 0 | 0 
relative contraindication to TEE | 0 | 0 
elderly patients | 0 | 0 
interventional cardiologic procedures | 0 | 0 
general anesthesia | 0 | 0 
MitralClip implantation | 0 | 0 
left atrial appendage occlusion | 0 | 0 
guide catheter–based procedures | 0 | 0 
probe manipulations | 0 | 1 
repeated motion | 0 | 1 
esophageal injury | 0 | 1 
procedural duration | 0 | 1 
contributing factor | 0 | 1 
preoperative pulmonary radiography | -1 | 0 
CT | -1 | 0 
anatomic proximity of thoracic osteophytes to the esophagus | -1 | 0 
safe performance of TEE | 0 | 0 
routine investigation | -1 | 0 
chest CT | -1 | 0 
vertebral osteophytes | -1 | 0 
anatomic relation to the esophagus | -1 | 0 
esophageal perforation | 1 | 2 
iatrogenic esophageal perforation | 1 | 2 
transesophageal echocardiography | 0 | 1 
rare event | 0 | 0 
high mortality rate | 0 | 0 
incidence | 0 | 0 
complication | 1 | 2 
adverse effect | 1 | 2 
adverse event | 1 | 2 
laceration | 1 | 2 
rupture | 1 | 2 
tear | 1 | 2 
injury | 1 | 2 
perforation | 1 | 2 
osteophyte | -1 | 0 
hyperostosis | -1 | 0 
exostoses | -1 | 0 
diffuse idiopathic skeletal hyperostosis | -1 | 0 
spine | -1 | 0 
vertebral column | -1 | 0 
preexisting esophageal pathologies | 0 | 0 
esophageal stricture | 0 | 0 
Zenker's diverticulum | 0 | 0 
fibrosis | 0 | 0 
prior