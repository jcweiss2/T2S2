77 years old | 0
male | 0
admitted to hospital | 0
anorexia | 0
deranged liver enzymes | 0
no significant past medical history | 0
no significant risk factors for liver disease | 0
does not take regular medications | 0
denied abdominal pain | 0
denied altered bowel habits | 0
afebrile | 0
hemodynamically stable | 0
unremarkable abdominal examination | 0
elevated alkaline phosphatase | 0
elevated gamma-glutamyl transferase | 0
elevated total bilirubin | 0
raised white blood cell count | 0
raised neutrophil count | 0
abdominal ultrasound showed no visible gallstones | 0
became febrile | 336
worsening ALP | 336
worsening GGT | 336
Escherichia Coli bacteraemia | 336
Klebsiella pneumoniae bacteraemia | 336
hypodense focal liver lesions | 336
multiple thrombosed portal vein branches | 336
pneumobilia | 336
infra-renal abdominal aortic aneurysm | 336
commenced on Piperacillin-Tazobactam | 336
commenced on Rivaroxaban | 336
portal vein thrombosis | 336
responded well to medical therapy | 336
hematemesis | 672
clinically unstable | 672
interval increase in infra-renal AAA | 672
impending rupture | 672
aortoenteric fistula | 672
Rivaroxaban ceased | 672
large blood clots in gastric fundus | 672
large blood clots in gastric body | 672
pulsatile lesion at D2 | 672
emergency endovascular aneurysm repair | 672
admitted to ICU | 672
acute right lower limb pain | 840
acute right lower limb swelling | 840
extensive deep vein thrombosis | 840
intravenous heparin infusion | 840
second episode of hematemesis | 912
bleeding duodenal fistula | 912
cholecystoduodenal fistula | 912
second laparotomy | 912
fistula between gallbladder and duodenum | 912
stones in gallbladder | 912
sludge in gallbladder | 912
6 mm stone in ampulla | 912
fistula repaired | 912
adjacent duodenal wall repaired | 912
cholecystectomy | 912
further hematemesis | 936
third laparotomy | 936
deep ulcer in D3 | 936
aortoenteric fistula with D3 | 936
aneurysm sac bleeding into duodenum | 936
iliolumbar arteries closed | 936
inferior mesenteric artery closed | 936
discharged from hospital | 0
re-admitted | 504
passed away | 504
