66 years old | 0
woman | 0
visited hospital's Department of Urology | 0
haematuria | 0
nausea | 0
hypercalcaemia | -72
calcium 22.6 mg/dL | 0
alkaline phosphatase 152 U/L | 0
amylase 1046 U/L | 0
lipase 499 U/L | 0
creatinine 2.42 mg/dL | 0
troponin T 1415.8 U/L | 0
C-reactive protein 17.79 mg/dL | 0
white blood cell count 30 000/μL | 0
ECG negative for ischemic heart disease | 0
ultrasound negative for ischemic heart disease | 0
CT scan demonstrated severe pancreatitis | 0
thyroid or parathyroid tumour | 0
blood pressure gradually dropped | 0
diagnosed with septic shock due to pancreatitis | 0
admitted to the intensive care unit | 0
noradrenaline | 0
adrenaline | 0
calcitonin 80 U/day | 0
isotonic fluids | 0
calcium levels did not decrease | 0
intact parathyroid hormone level 2204 pg/mL | 24
ultrasound imaging showed 40-mm hypoechoic heterogeneous tumour with ill-defined borders | 24
suspected parathyroid carcinoma | 24
hypercalcaemia | 24
severe pancreatitis | 24
enhanced CT scan not performed due to renal dysfunction | 24
plain CT scan showed pancreatitis (CT grade 2) | 24
over 3 points of negative prognostic factors | 24
shock | 24
Cr > 2 mg/dL | 24
CRP 15 mg/dL | 24
diagnosed with severe pancreatitis | 24
hypercalcaemia persisted (15 mg/dL) | 48
continuous hemodiafiltration (CHDF) | 48
zoledronic acid | 48
evocalcet | 48
altered mentation | 48
circulatory function decline | 48
respiratory function decline | 48
ventilator support initiated | 48
ECMO-assisted surgery scheduled | 48
administration of elcatonin 60 U/day | 48
isotonic fluids | 48
CHDF initiated | 48
hypercalcaemia persisted | 48
operation assisted by ECMO | 72
initiated V-A ECMO | 72
parathyroidectomy | 72
left thyroidectomy | 72
left recurrent laryngeal nerve resection | 72
intact parathyroid hormone (PTH) dropped remarkably | 96
circulatory function improved | 96
terminated ECMO use | 96
calcium levels decreased gradually | 96
treated pancreatitis using i.v. fluids | 96
antibiotics | 96
dialysis due to renal dysfunction | 96
noradrenaline | 96
de-escalated | 120
stopped 1 month after surgery | 744
ventilatory support weakened respiratory muscles | 744
transferred to another hospital for rehabilitation | 744
