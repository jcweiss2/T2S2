69 years old | 0
male | 0
admitted to the hospital | 0
primary arterial hypertension | 0
dyslipidemia | 0
ischemic heart disease | 0
severe heart ejection fraction 15–20% | 0
mechanical aortic valve | 0
stage 4 chronic kidney disease | 0
early-stage Alzheimer’s dementia | 0
non-bloody diarrhea | -96
diffuse abdominal pain | -96
dyspnoea | -96
unquantified fever | -96
prostrated | 0
hypotensive | 0
homogeneous opacity involving the middle and lower lobes of the right hemithorax | 0
pleural effusion | 0
protein C-reactive protein was 27 mg/dL | 0
serum creatinine was 6 mg/dl | 0
hypoxemic respiratory failure | 0
lactate level at admission was 1,37 mmol/L | 0
septic shock | 0
multiorgan dysfunction | 0
empirical antibiotic therapy with ceftriaxone | 0
vasopressor support | 0
invasive mechanical ventilation | 0
continuous renal function replacement technique | 0
transferred to the ICU | 0
antibiotic therapy escalated to meropenem and linezolid | 0
L. monocytogenesis identified in blood cultures | 24
L. monocytogenesis identified in pleural fluid | 24
HIV negative | 24
extensive multiloculated right pleural effusion | 48
pleural decortication | 48
hemothorax | 48
linezolid changed to ampicillin | 48
meropenem continued | 48
decrease in inflammatory parameters | 72
ampicillin treatment | 48
piperacillin-tazobactam added | 312
inflammatory parameters increased | 312
pleural imaging worsened | 312
suspension of invasive measures | 600
died | 720