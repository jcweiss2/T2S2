22 years old | 0
female | 0
multiparous | 0
pregnant | 0
24 week gestation | 0
altered consciousness | 0
vomiting | 0
bleeding per vaginum | 0
PV manipulation by a local health worker | -24
pale | 0
dehydrated | 0
tender abdomen | 0
distended abdomen | 0
BP 80/46 mm Hg | 0
HR 130/min | 0
respiratory rate 35/min | 0
Glasgow coma score 8 | 0
no neck rigidity | 0
normal reflexes | 0
gangrenous bowel loops protruding from vagina | 0
abdominal skiagram showed gas under diaphragm | 0
electrocardiogram showed prolonged PR interval | 0
wide QRS complex | 0
peaked T wave | 0
rehydrated with normal saline | 0
hypoxia | 0
invasive positive pressure ventilation (SIMV) | 0
Ryle's tube | 0
Foley's catheterization | 0
central venous cannulation | 0
Midazolam infusion | 0
Fentanyl infusion | 0
severe anaemia | 0
deranged renal functions | 0
metabolic acidosis |"0
hyperkalaemia | 0
hyponatraemia | 0
nebulised with Salbutamol | 0
dextrose-insulin infusion | 0
unsafe abortion | -24
uterine perforation | -24
bowel perforation | -24
continued fluid replacement | 0
BP returned to 116/62 mm Hg | 2
emergency laparotomy | 2
general anaesthesia | 2
sudden hypotension | 2
cardiac arrest | 2
fluid mixed blood clots expulsion | 2
feculent matter expulsion | 2
external cardiac massage | 2
colloid bolus | 2
Inj. adrenaline | 2
revived after 2 minutes | 2
Dopamine infusion | 2
vitals remained stable | 2
no further episodes of arrhythmia | 2
Anaesthesia maintained with Ketamine | 2
nitrous oxide-oxygen combination | 2
neuromuscular blockade by Atracurium | 2
6-month-old dead foetus extracted | 2
uterine perforation (3 cm × 4 cm) | 2
gangrenous bowel loops (ileum, transverse and sigmoid colon) | 2
resection anastomosis | 2
subtotal hysterectomy | 2
end-colostomy | 2
blood transfusion | 2
fluid transfusion | 2
surgery lasted approximately four hours | 6
shifted to ICU | 6
maintained in SIMV mode | 6
dopamine infusion tapered over twenty-four hours | 30
extubated after two days | 54
survived with no major organ failure | 240
no neurological deficit | 240
discharged on tenth post-operative day | 240
