52 years old | 0
female | 0
admitted to the hospital | 0
colicky left flank pain | 0
no medical history of chronic or immunodeficiency diseases | 0
no previous history of urolithiasis or urinary tract infections | 0
stable vital signs | 0
blood pressure 110/70 mmHg | 0
respiratory rate 20/min | 0
pulse rate 69/min | 0
temperature 37.0℃ | 0
left flank pain | 0
left costovertebral angle tenderness | 0
white blood cells 9970/mm3 | 0
neutrophils 84.4% | 0
lymphocytes 6.4% | 0
hemoglobin 10.6 g/dL | 0
platelet count 142,000/mm3 | 0
C-reactive protein 57.5 mg/dL | 0
blood urea nitrogen 19 mg/dL | 0
creatinine 0.8 mg/dL | 0
total protein 6.5 g/dL | 0
albumin 3.2 g/dL | 0
total bilirubin 2.2 mg/dL | 0
aspartate aminotransferase 34 IU/L | 0
alanine aminotransferase 47 IU/L | 0
no WBCs in urinalysis | 0
red blood cells over 100 per high-power field | 0
urinary stone in the left ureter | 0
ESWL | 72
ESWL aggravated flank pain | 72
ESWL aggravated costovertebral angle tenderness | 72
body temperature rose to 39.9℃ | 120
blood pressure fell to 70/50 mmHg | 168
heart rate 125/min | 168
respiratory rate 26/min | 168
body temperature 39.0℃ | 168
oxygen saturation 80% | 168
mechanical ventilation | 168
shock management | 168
WBCs 18,400/mm3 | 168
neutrophils 90.4% | 168
lymphocytes 5.5% | 168
hemoglobin 11 g/dL | 168
platelet count 92,000/mm3 | 168
CRP 240 mg/dL | 168
BUN 56 mg/dL | 168
creatinine 2.4 mg/dL | 168
cefepime administration | 168
vancomycin administration | 168
computed tomography | 168
4 mm left proximal ureter stone | 168
hydroureteronephrosis | 168
no WBCs or RBCs in urine | 168
blood cultures positive for gram-negative bacilli | 168
Achromobacter xylosoxidans identified | 168
antibiotics changed to imipenem | 216
blood cultures no longer revealed A. xylosoxidans | 336
renal function worsened | 336
continuous renal replacement therapy | 336
Burkholderia cepacia isolated from blood cultures | 384
central venous catheter removed | 384
tip culture negative | 408
repeated blood cultures negative | 408
respiratory failure | 504
bilateral opacities on chest imaging | 504
passed away from septic shock and multiple organ failure | 696
16S rRNA sequencing identified A. xylosoxidans | 696