58 years old | 0
female | 0
hypertension | 0
stage 3 chronic kidney disease | 0
undisclosed muscle spasticity | 0
admitted to the emergency department | 0
complaint of worsening upper extremities tremors | 0
paresthesia | 0
limb weakness | 0
pins and needle sensation | 0
temperature of 103 F | 0
tachycardia to 103 beats per minute | 0
hypertensive to 150/90 mmHg | 0
tachypneic to 21 breaths per minute | 0
saturating 97% in room air | 0
coarse tremors | 0
neurology examination revealed ⅗ strength in bilateral upper extremities | 0
neurology examination revealed ⅘ strength in bilateral lower extremities | 0
decreased sensation in all 4 extremities | 0
lungs were clear to auscultation | 0
initial impression was sepsis | 0
initial impression was fever of unknown origin | 0
started on broad spectrum antibiotics | 0
started on cefepime | 0
started on vancomycin | 0
started on metronidazole | 0
laboratory work including white blood cell (WBC) count | 0
laboratory work including lactic acid | 0
laboratory work including inflammatory markers | 0
blood cultures were negative | 0
urine cultures were negative | 0
respiratory cultures were negative | 0
lumbar puncture | 0
cerebrospinal fluid analysis ruled out meningitis | 0
chest x-ray | 0
abdominal ultrasound | 0
magnetic resonance imaging of head | 0
magnetic resonance imaging of spine | 0
neurology consultation | 0
electroencephalography (EEG) | 0
EEG ruled out seizure disorder | 0
ruling out Guillain Barre Syndrome | 0
ruling out Alcohol withdrawal syndrome | 0
toxicology consultation | 0
concern of anticholinergic toxicity | 0
anticholinergic toxicity was ruled out | 0
persistent fever | 72
worsening mental status | 72
visual hallucinations | 72
hyperpyrexia | 72
ocular clonus | 72
profound muscle rigidity | 72
somnolent | 72
unable to follow command | 72
continuous tremors | 72
given lorazepam | 72
given phenobarbital | 72
given intravenous haloperidol | 72
rapid response was called | 72
evaluated by the intensive care unit (ICU) team | 72
minimally responsive | 72
tachypnea to 40 breaths/minute | 72
ABG showed pH of 7.3 | 72
ABG showed PCO2 of 28.6 | 72
ABG showed PaO2 of 70 on room air | 72
intubated | 72
transferred to the ICU | 72
possible diagnosis of neuroleptic malignant syndrome | 72
possible diagnosis of baclofen withdrawal | 72
laboratory work for serum creatinine kinase | 72
laboratory work for lactic acid | 72
started bromocriptine | 72
history and home medications were reviewed | 72
patient was on oral baclofen 10 mg 3 times a day | 0
patient was not taking baclofen for the last 3 days | -72
baclofen was restarted | 96
resolution of fever | 120
improvement in mental status | 120
complete cessation of tremors | 120
extubated | 120
transferred to the medical floor | 120
discharged to an acute rehabilitation facility | 144
on oral baclofen for the last 2 years | -2880