38 years old | 0
male | 0
obese | 0
BMI 35.93 kg/m2 | 0
admitted to the hospital | 0
fever | -48
dry cough | -48
shortness of breath | -48
positive COVID-19 PCR test | 0
no known medical or surgical history | 0
no immunization against COVID-19 | 0
vital stability | 0
normal chest examination | 0
normal cardiovascular examination | 0
no abdominal tenderness | 0
patch of pneumonic consolidation | 0
left lower lobe of the lung | 0
respiratory distress | 96
tachycardia | 96
tachypnea | 96
hypotension | 96
hypoxia | 96
bilateral crepitations | 96
soft and lax abdomen | 96
increasing bilateral patchy infiltrates | 96
severe COVID-19 pneumonia | 96
enoxaparin | 96
severe persistent abdominal pain | 120
diaphoresis | 120
vomiting | 120
GCS 15/15 | 120
lax abdomen | 120
mild tenderness in the epigastrium | 120
elevated D-dimer | 120
hypodense filling defect of the superior mesenteric artery | 120
venous thrombosis | 120
ischemic changes of the small bowel loops | 120
exploratory laparotomy | 120
ischemic nonviable bowel | 120
duodenojejunal flexure | 120
mid transverse colon | 120
ischemic bowel resection | 120
postoperative sepsis | 168
multiorgan failure | 168
pulseless ventricular tachycardia | 168
resuscitation | 168
death | 216
passing away | 216