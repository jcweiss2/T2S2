61 years old | 0
female | 0
admitted to emergency | 0
soft tissue infection of left buttock | 0
soft tissue infection of posterior thigh | 0
chronic left perineum sinus | -8760
excision of chronic left perineum sinus | -8760
CT scan | -8760
colonoscopy | -8760
asymptomatic sigmoid diverticulosis | -8760
left maxillary sinus mass | -7200
granulomatosis with polyangiitis | -7200
osteomyelitis | -7200
left-sided hydronephrosis | -7200
inflammatory changes in sigmoid diverticulitis | -7200
ureteric stenting | -7200
conservative management of diverticulitis | -7200
colorectal carcinoma ruled out | -5760
repeat colonoscopy | -5760
blistering rash over left buttock | -672
blistering rash over gluteal fold | -672
treated with acyclovir | -672
new painful induration over left buttock | -72
diagnosed as early abscess | -72
prescribed amoxicillin–clavulanate | -72
enlarged induration | -24
serous discharge | -24
chills | -24
leukocytosis | 0
acute kidney injury | 0
creatinine of 191 μmol/L | 0
non-contrast CT scan | 0
performed sigmoid diverticulitis | 0
free air tracking inferiorly into left pelvis | 0
abscess | 0
subcutaneous emphysema | 0
wide debridement of left buttock | 12
wide debridement of perineum | 12
wide debridement of leg | 12
laparotomy | 12
washout | 12
left hemicolectomy | 12
antibiotic treatment with piperacillin/tazobactam | 12
antibiotic treatment with clindamycin | 12
antibiotic treatment with vancomycin | 12
further debridement | 36
drainage of retroperitoneal abscesses | 36
drainage of pre-rectal abscesses | 36
end colostomy creation | 36
polymicrobial gut flora | 36
negative pressure wound therapy | 48
transfer to rehabilitation hospital | 432
delayed wound closure | 144
rotational flap on left buttock | 144
left ureteric stent removed | 156
resolution of hydronephrosis | 156
ulcerating lesions over left hip | 4320
biopsied | 4320
pyoderma gangrenosum | 4320
consulted to dermatology | 4320
treated with prednisone | 4320
treated with colchicine | 4320
treated with azathioprine | 4320
chronically maintained with mycophenolic acid | 9000
intralesional triamcinolone injections | 9000
investigations for immunodeficiency syndromes | 9000