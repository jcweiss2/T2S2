48 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
admitted to the Emergency Service | 0 | 0 | Factual
toothache | -96 | 0 | Factual
dyspnea | -96 | 0 | Factual
chest pain | -96 | 0 | Factual
sweating | -96 | 0 | Factual
tachyarrhythmia | -96 | 0 | Factual
sore throat | -96 | 0 | Factual
fever | -96 | 0 | Factual
gross swelling of the lower right cheek | 0 | 0 | Factual
submandibular and mental regions were erythematous and warm on palpation | 0 | 0 | Factual
difficulties in opening the jaw | 0 | 0 | Factual
inflammatory changes of the mucous membrane of his oral cavity | 0 | 0 | Factual
treated at home with ceftriaxone-steroids-based | -96 | 0 | Factual
ineffective treatment | -48 | 0 | Factual
condition of the patient worsened | -48 | 0 | Factual
dyspnea | -48 | 0 | Factual
chest pain | -48 | 0 | Factual
increase in the amount of white blood cells | 0 | 0 | Factual
neutrophils | 0 | 0 | Factual
C-reactive protein | 0 | 0 | Factual
urgent orotracheal intubation | 0 | 0 | Factual
left pleural effusion | 0 | 0 | Factual
mediastinitis | 0 | 0 | Factual
right parapharyngeal abscess | 0 | 0 | Factual
possible complication of an odontogenic infection | 0 | 0 | Possible
drainage of the right neck | 0 | 0 | Factual
left chest drain | 0 | 0 | Factual
intravenous antibiotic therapy | 0 | 0 | Factual
piperacillin sodium plus tazobactam sodium | 0 | 48 | Factual
clinical condition of the patient worsened | 48 | 48 | Factual
transferred to an Intensive Care Unit | 48 | 48 | Factual
air collection in the right submandibular | 48 | 48 | Factual
air collection in the left carotid | 48 | 48 | Factual
air collection in the retroesophageal and pretracheal spaces | 48 | 48 | Factual
cervical necrotizing fasciitis with DNM | 48 | 48 | Factual
bilateral pleural effusions | 48 | 48 | Factual
additive pleural drain | 72 | 72 | Factual
abscesses in the cervical spaces | 72 | 72 | Factual
extensive mediastinal empyema | 72 | 72 | Factual
left pleural effusion | 72 | 72 | Factual
right hydropneumothorax | 72 | 72 | Factual
aggressive mediastinal debridement | 72 | 72 | Factual
VATS | 72 | 72 | Factual
incision and drainage of the neck abscesses | 72 | 72 | Factual
oral tooth extraction | 72 | 72 | Factual
purulent fluid in the cavity below was drained and packed | 72 | 72 | Factual
Streptococcus anginosus | 72 | 72 | Factual
Gemella morbillorum | 72 | 72 | Factual
Staphylococcus lugdunensis | 72 | 72 | Factual
antibiotic therapy | 72 | 168 | Factual
Amoxicillin | 72 | 168 | Factual
Metronidazole | 72 | 168 | Factual
dismissed in better health conditions | 168 | 168 | Factual