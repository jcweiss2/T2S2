50 years old | 0
male | 0
idiopathic pulmonary fibrosis | -672
hypoxia | -192
acute exacerbation of idiopathic pulmonary fibrosis | -192
broad-spectrum antibiotics | -192
prednisolone | -192
intubated | -192
mechanically ventilated | -192
partial pressure of arterial carbon dioxide (PaCO2) was 88 mmHg | -192
partial pressure of arterial oxygen (PaO2) was 48 mmHg | -192
fraction of inspired oxygen (FIO2) of 1.0 | -192
V-V ECMO | -192
21-Fr drainage cannula was inserted in the left femoral vein | -192
19-Fr return cannula was inserted in the right femoral vein | -192
tracheostomy | -168
sedated | 0
mechanically ventilated | 0
ECMO blood flow around 4 L/min | 0
peripheral capillary oxygen saturation (SpO2) over 85% | 0
sweep gas flow with 100% of oxygen | 0
membrane oxygenator | 0
PaCO2 between 30 mmHg and 35 mmHg | 0
mechanical ventilation settings altered to a “lung rest” setting | 0
driving pressure of 5 cmH2O | 0
positive end-expiratory pressure of 10 cmH2O | 0
FIO2 of 0.4 | 0
heart rate was 50 beats/min | 0
blood pressure was 156/104 mmHg | 0
echocardiography revealed an ejection fraction of 60.7% | 0
tricuspid regurgitation pressure gradient (TR-PG) of 10 mmHg | 0
renal function was normal | 0
anticoagulant with heparin | 0
activated partial thromboplastin time between 50 and 80 seconds | 0
vancomycin prophylaxis | 0
mechanical ventilation was discontinued | 38
tracheostomy tube removed | 42
speech cannula | 42
low-flow or high-flow oxygen therapy | 42
oral intake began | 47
severe respiratory failure persisted | 47
target SpO2 and PaCO2 values achieved | 47
analgesia was induced by the administration of morphine | 47
fully awake, oriented, and communicative | 47
seen daily by a physiotherapist for exercise and respiratory training | 47
clinical decision that the patient's respiratory failure was irreversible | 59
listed on the LTx registry | 284
membrane oxygenator changed 23 times | 0
cannula changed 10 times | 0
oxygenator changed because of gas exchange failure | 0
oxygenator changed because of apparent thrombus on the membrane | 0
oxygenator changed because of acute platelet reduction | 0
average lifespan of the oxygenators was 16 days | 0
cannula changed when the patient was clinically diagnosed with sepsis | 0
double lumen cannula was not available | 0
two-site cannulation mode was necessary for V-V ECMO | 0
right internal jugular vein for drainage | 0
right femoral vein for drainage | 0
left femoral vein for drainage | 0
left internal jugular vein for return | 0
right femoral vein for return | 0
left femoral vein for return | 0
25 or 23-Fr cannula for drainage | 0
23 or 21-Fr cannula for return | 0
no technical complications | 0
complained of dyspnea | 223
SpO2 was around 90% on ECMO with a flow of 5 L/min | 223
echocardiography showed a D shape | 223
TR-PG was 56 mmHg | 223
endothelin-receptor antagonist bosentan | 223
phosphodiesterase type 5 inhibitor sildenafil | 223
right failure became worse | 226
TR-PG increased to 78 mmHg | 226
decision to convert the configuration of ECMO from V-V to venovenous-arterial (VV-A) | 226
condition improved | 226
TR-PG decreased to 43 mmHg | 226
ECMO configuration was converted from VV-A back to V-V | 282
finally listed on the LTx registry | 284
attempted to change the cannula | 305
cannula-related blood stream infection | 305
remaining veins were occluded by thrombosis | 305
could not access them to modify the site of cannulation | 305
used the same cannula that was inserted on day 276 | 305
septic shock | 371
attempted to change the cannula again | 371
no flow in any of the veins | 371
decided not to continue ECMO support | 371
disconnected from ECMO | 403
died soon thereafter | 403