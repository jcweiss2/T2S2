61 years old | 0
man | 0
admitted to hospital | 0
fever | -168
muscle weakness | -168
fatigue | -168
family contacts tested positive for COVID-19 | -168
end-stage renal failure | -168
renal transplant in 2009 | -168
immunosuppressed | -168
type 2 diabetes mellitus | -168
cerebrovascular disease | -168
sleep apnea | -168
orthostatic hypotension | -168
benign prostatic hyperplasia | -168
transurethral resection of the prostate in 2009 | -168
recurrent urinary tract infections | -168
temperature mildly elevated at 37.6°C | 0
pulse 112 beats per minute | 0
blood pressure 111/74 | 0
urinalysis positive for leucocytes | 0
urinalysis positive for nitrites | 0
urinalysis positive for trace amounts of blood | 0
admitted and treated in hospital for urosepsis | 0
developed low oxygen saturations | 0
tested positive for COVID-19 | 0
received treatment with dexamethasone | 0
received treatment with tocilizumab | 0
persistently poor oxygen saturations | 168
limited urine output | 168
transfer to intensive care unit | 168
intubated | 168
hemodialysed | 168
persistent fluctuating low oxygen saturations | 120
computed tomography pulmonary angiogram performed | 120
saddle pulmonary embolus | 120
extension into segmental and subsegmental pulmonary artery branches | 120
bilateral ground-glass attenuation | 120
patchy consolidation | 120
severe COVID-19 pneumonitis | 120
treatment with low molecular weight heparin initiated | 120
diagnosis of saddle pulmonary embolus | 120
bilateral edematous eyelids | 168
ophthalmology opinion sought | 168
ocular examination revealed bilaterally fixed pupils | 168
ocular examination revealed bilaterally constricted pupils | 168
left eye 2 mm | 168
right eye 3 mm | 168
no exophthalmos noted | 168
asymmetrical right-sided conjunctival injection | 168
asymmetrical right-sided chemosis | 168
visual acuity difficult to ascertain | 168
unconscious | 168
receiving invasive ventilation | 168
CT head with orbital imaging performed | 168
expanded and hyperdense right SOV | 168
asymmetrical hyperdensity of right masticator space venous structures | 168
swelling of right pterygoid muscles | 168
effacement of fat planes | 168
acute thrombosis of right SOV | 168
acute thrombosis of right pterygoid venous plexus | 168
left SOV dilated | 168
suspicion of bilateral caroticocavernous fistula | 168
multidisciplinary team decision to treat with low molecular weight heparin | 168
patient made excellent progress | 168
extubated | 408
repeat interval imaging | 408
CT head | 408
computed tomography pulmonary angiogram | 408
complete resolution of right SOV thrombosis | 408
complete resolution of pulmonary embolism | 408
marked improvement in lung parenchymal appearances | 408
completely recovered from illness | 408
no residual abnormalities in SOV thrombosis | 408
preserved range of movement in eyes bilaterally | 408
no diplopia | 408
no deficiency in visual acuity | 408
undergoing speech and language therapy | 408
undergoing physiotherapy | 408
undergoing rehabilitation | 408
prolonged hospital admission with COVID-19 | 408
