75 years old| 0
male| 0
arterial hypertension| 0
chronic atrial fibrillation| 0
type 2 diabetes| -87600
moderate chronic renal failure| 0
myocardial infarction| -96720
coronary artery bypass grafting| -96720
implantable defibrillator| -96720
low left ventricle ejection fraction| -96720
ramipril| 0
cardensiel| 0
aldactone| 0
fluindione| 0
metformin| 0
furosemide| 0
anasarca| -144
worsening exertional dyspnea| -144
increased furosemide| -144
introduction of spironolactone| -144
indwelling urinary catheterization| -144
acute renal failure| -144
dobutamine| -144
arterial hypotension| -144
LVEF of 20%| -144
decreasing aortic velocity integral time| -144
transthoracic echocardiography control| -144
transferred to intensive care unit| 0
confused| 0
hypothermic| 0
atrial tachycardia| 0
capillary blood glucose level of 2.55 g/L| 0
mottling| 0
deep hypotension| 0
dobutamine at 10 µg/kg/min| 0
no functional digestive signs| 0
no hematuria| 0
cloudy urinary residues| 0
foul-smelling urinary residues| 0
