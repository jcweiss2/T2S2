80 years old | 0
female | 0
Alzheimer’s dementia | 0
diabetes mellitus | 0
hypertension | 0
chronic kidney disease | 0
admitted to the intensive care unit | 0
hypotension | -336
lactic acidosis | -336
progressive altered mental status | -336
physical decline | -336
blood pressure 89/56 | 0
normal heart rate | 0
normal oxygen saturation | 0
no fever | 0
no tachypnea | 0
lactic acid 3.6 mmol/L | 0
leukocytosis 14.7 x 10^3 cells/μL | 0
neutrophilic predominance | 0
troponin peaked at 1104 pg/mL | 0
no other laboratory abnormalities | 0
no other clinical abnormalities | 0
Wells score 0 points | 0
D-dimer not obtained | 0
admitted for presumptive septic shock | 0
treated with fluids | 0
treated with broad-spectrum antibiotics | 0
blood pressure improved | 0
lactic acidosis resolved | 0
troponin elevation due to demand ischemia | 0
blood cultures negative | 0
reached pre-hospital baseline | 0
hemodynamic stability | 0
improvement in the ICU | 0
transferred to gerontology unit | 0
discharge planning | 0
afebrile | 0
heart rate 80 | 0
blood pressure 117/62 | 0
SpO2 99% | 0
jugular venous distension | 0
normal cardiopulmonary auscultatory exam | 0
no peripheral edema | 0
no asymmetric lower extremity swelling | 0
cardiac POCUS using HUD | 0
dilated RV | 0
akinesis of mid-RV free wall | 0
apical sparing | 0
McConnell’s sign | 0
diastolic septal flattening | 0
D-sign | 0
IVC dilated to 3.0 cm | 0
minimal inspiratory variation | 0
formal transthoracic echocardiography | 0
electrocardiogram | 0
S1Q3T3 pattern | 0
D-dimer 51190 ng/mL | 0
CT angiography | 0
saddle PE | 0
RV strain | 0
heparin infusion initiated | 0
transitioned to oral apixaban | 0
no hemodynamic compromise | 0
no further complications | 0
megestrol use | 0
no hypercoagulability workup | 0
