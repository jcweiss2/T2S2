25 years old | 0
male | 0
admitted to the hospital | 0
perineal pain | -96
swelling | -96
discharge | -96
high-grade fever | -96
vomiting | -96
visited health center | -96
given po medication | -96
no improvement | -96
no history of trauma | 0
no recent surgery | 0
no history of diabetes | 0
no history of hypertension | 0
no history of chronic illness | 0
no history of chronic alcohol abuse | 0
seronegative for HIV | 0
no history of drug intake | 0
no known drug allergy | 0
temperature 38.8°C | 0
blood pressure 85/46 mmHg | 0
pulse rate 120 beats per minute | 0
respiratory rate 24 breaths per minute | 0
no shortness of breath | 0
body mass index (BMI) 19 kg/m2 | 0
distended abdomen | 0
guarding | 0
rebound | 0
severe direct tenderness in the hypogastrium | 0
normal bowel sounds | 0
bilateral necrotic scrotum | 0
perineum | 0
foul-smelling pus discharge | 0
palpable crepitus | 0
enlarged, edematous and tender scrotum | 0
ruptured perianal abscess | 0
WBC 19,000 | 0
RBC 2.86 | 0
HGB 8.6 g/dl | 0
HCT 23.7 | 0
PLT 377,000 | 0
NEUT 87% | 0
ESR 38 | 0
NA+ 132 | 0
K+ 3.53 | 0
CL 97 | 0
CREAT 1.57 | 0
UREA 64 | 0
ALP 50 | 0
ALB 2.9 | 0
BIL. T 1.0 | 0
RBS 218 | 0
resuscitated with normal saline | 0
started broad spectrum antibiotics | 0
transferred to operation room | 0
operated on under general anesthesia | 0
debridement | 0
necrotic tissue and abscess | 0
thrombosed vessels | 0
debrided thoroughly | 0
wound washed with hydrogen peroxide and normal saline | 0
transfused with 2 units of crossed-matched blood | 0
drain left in the retroperitoneum | 0
re-debridement planned after 24 h | 0
transferred to surgical intensive care unit (ICU) | 0
vital signs monitored continuously | 0
input and output monitoring | 0
antibiotics continued | 0
wound care BID | 0
wound dressing | 0
stayed in surgical ICU for 5 days | 120
transferred to surgical ward | 120
multiple debridements | 120
infection fully controlled | 120
wound granulated well | 120
primary closure of abdominal skin | 120
bilateral testicles buried in the medial thigh | 120
scrotal reconstruction | 120
discharged home improved | 168
follow-up at surgical referral clinic | 168
doing well | 168