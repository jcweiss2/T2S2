37 years old | 0
    female | 0
    admitted to the hospital | 0
    pulmonary arterial hypertension (PAH) | 0
    dyspnoea | -17520
    dizziness | -17520
    syncope | -17520
    weakness | -17520
    fatigue | -17520
    3rd pregnancy | -17520
    gradually worsening symptoms of dyspnoea on exertion | -17520
    initial presentation in a primary care facility | -168
    clinical deterioration (WHO functional Class IV) | -168
    pulmonary embolism ruled out | -168
    echocardiographic diagnosis of severe pulmonary hypertension | -168
    estimated systolic PA pressure 100 mmHg | -168
    transfer to intensive care unit | -168
    initiation of Sildenafil medication | -168
    symptomatic improvement | -144
    estimated systolic PA-pressure lowered to 55 mmHg | -144
    emergent caesarean section | -120
    stand-by mechanical circulatory support | -120
    healthy child delivered | -120
    transfer to standard cardiology ward | -96
    right heart catheterization | -96
    left heart catheterization | -96
    coronary artery disease ruled out | -96
    arteriovenous shunts ruled out | -96
    elevated mean PA pressure | -96
    elevated pulmonary vascular resistance | -96
    left ventricular end diastolic pressure slightly elevated | -96
    secondary aetiologies ruled out | -48
    diagnosis of idiopathic pulmonary hypertension | -48
    sequential therapy with Macicentan initiated | -48
    discharge from hospital | 24
    combination therapy of Sildenafil and Macicentan | 24
    out-patient follow-up | 264
    symptomatic patient (WHO functional Class III) | 264
    elevated systolic PA pressure values of about 60 mmHg | 264
    right heart catheterization with vasodilator testing | 408
    elevated mean PA pressure | 408
    elevated pulmonary vascular resistance | 408
    vasodilator testing with significant positive result | 408
    intravenous Epoprostenol 15 ng/kg/min | 408
    high-dose calcium channel blocker (CCB) therapy initiated | 408
    Sildenafil discontinued | 408
    therapy well tolerated | 492
    symptoms improved significantly | 492
    normal values for pulmonary vascular resistance | 492
    slightly increased values for mean PA pressure | 492
    stable patient | 528
    regular out-patient visits | 528
    WHO functional class improved to I | 528
    natriuretic peptides in normal range | 528
    estimated systolic PA pressure decreased to 40 mmHg | 528
    improvements in 6 min walk test | 528
    improvements in cardiopulmonary exercise testing results | 528
    classified as low risk (<5%) | 528
    no adverse events occurred | 528
    high-dose CCB therapy well tolerated | 528
    shortness of breath (SoB) | 0
    World Health Organisation functional class (WHO FC) IV | 0
    symptom onset during 1st trimester of pregnancy | -672
    mild SoB | -672
    transthoracic echocardiogram showing no abnormalities | -672
    initial electrocardiogram showing right heart strain or pulmonary embolism | -672
    computed tomography (CT) ruled out pulmonary embolism | -672
    signs of right heart stress on CT | -672
    ventilation/perfusion (V/Q) scan not performed | -672
    one healthy child | -17520
    one abortion due to acute toxoplasmosis | -17520
    medical history unremarkable | -17520
    left ventricle normal size | 0
    signs of chronic right heart pressure overload | 0
    estimated systolic pulmonary artery pressure (sPAP 86 mmHg + central vein pressure) elevated | 0
    chest pain | 0
    oxygen supply needed (2 L/min) | 0
    sinus tachycardia (110/min) | 0
    tachypnoea (28/min) | 0
    BNP values above 300 pg/mL | 0
    therapy with Sildenafil initiated | 0
    estimated sPAP gradually reduced to 60 mmHg | 0
    V/Q scan excluded pulmonary embolic disease | 24
    blood work for vasculitis negative | 24
    blood work for connective tissue disease negative | 24
    blood work for overlap syndromes negative | 24
    no signs of chronic infectious disease | 24
    chronic pulmonary disease ruled out | 24
    interstitial lung disease ruled out | 24
    restrictive ventilatory dysfunction ruled out | 24
    obstructive ventilatory dysfunction ruled out | 24
    abdominal ultrasound ruled out portal hypertension | 24
    diagnosis of Idiopathic PAH aggravated by pregnancy | 24
    elevated mean PA pressure of 66 mmHg | 24
    left ventricular end-diastolic pressure (LVEDP) of 16 mmHg | 24
    elevated pulmonary vascular resistance (PVR) of 608 dyn s/cm5 | 24
    classified in intermediate risk (ESC/ERS score 1.55) | 24
    Macitentan added | 24
    discharged in stable condition | 24
    followed up 6 months later | 408
    risk stratification suggested low risk (ESC/ERS score 1.27) | 408
    still in WHO FC III | 408
    elevated sPAP of 58 mmHg | 408
    right heart catheterization | 408
    PVR and mean PA pressure still elevated | 408
    vasodilator testing showed significant response | 408
    high-dose CCB therapy initiated | 408
    Sildenafil discontinued | 408
    therapy well tolerated | 492
    symptoms improved to WHO FC II | 492
    decrease of mean PA pressure to 25 mmHg | 492
    reduction of PVR | 492
    non-invasive estimation of sPAP < 40 mmHg | 528
    stable clinical condition | 528
    WHO FC I | 528
    BNP values <100 pg/mL | 528
    scheduled for follow-up every 6 months | 528
    no adverse events occurred | 528
    high-dose CCB therapy well tolerated | 528
    
    