83 years old | 0
female | 0
admitted to the hospital | 0
abdominal pain | -120
hematochezia | -48
asthenia | -120
cutaneous squamous cell carcinoma | -720
total excision of cSCC | -720
recurrence of squamous cell carcinoma | -360
radiation therapy | -360
radiation therapy completed | -270
CT scan | -90
hypodense structure in pelvic cavity | -90
follow-up | -90
worsening abdominal pain | 0
hematochezia | 0
asthenia | 0
low blood pressure | 0
guarding | 0
rebound tenderness | 0
plasma creatinine level | 0
white blood cell count | 0
hemoglobin level | 0
C-reactive protein level | 0
hyperlactatemia | 0
abdominal CT scan | 0
extraluminal air bubbles | 0
fat stranding | 0
intra-abdominal free fluid | 0
intestinal perforation | 0
fluid resuscitation | 0
proton pump inhibitor therapy | 0
antibiotic treatment | 0
blood cultures | 0
emergency exploratory laparotomy | 0
purulent peritonitis | 0
ileal perforation | 0
segmental resection of ileum | 0
damage control surgical approach | 0
histological analysis | 0
non-keratinizing squamous cell carcinoma | 0
venous invasion | 0
lymph node | 0
septic shock | 0
norepinephrine support | 0
broad-spectrum antibiotic | 0
corticoid administration | 0
death | 24