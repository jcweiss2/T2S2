54 years old | 0
male | 0
uncontrolled diabetes mellitus | -672
admitted to the hospital | 0
complaint of right frontal headache | 0
vomiting | 0
elevated glucose level | 0
normal complete blood count | 0
normal renal profile | 0
normal hepatic profile | 0
negative blood culture | 0
negative HIV serology | 0
normal CD4 count | 0
circumferential mucosal thickening in the sphenoid sinuses | 0
mild scattered mucosal thickening in the other paranasal sinuses | 0
fluid opacification of the mastoid air cells and middle ear cavities | 0
started on insulin | 0
started on Augmentin | 0
sudden loss of vision in the right eye | 120
jaw pain | 120
repeated brain CT scan | 120
progression of the inflammatory changes in the paranasal sinuses | 120
suspected giant cell arteritis | 120
treatment with pulse intravenous methylprednisolone | 120
temporal artery biopsy | 144
corticosteroids discontinued | 144
worsened symptoms | 144
third CT scan brain | 168
progression of the sinusitis to the retropharyngeal abscess | 168
sinonasal biopsy | 168
histopathological examination showed positive GMS stain for fungus | 168
diagnosed with mucormycosis | 168
treated with amphotericin B | 168
developed sepsis | 240
started on broad-spectrum antibiotics | 240
started on vancomycin | 240
started on meropenem | 240
mild bilateral pleural effusions | 240
mucosal edema involving the ascending colon | 240
melena mixed with streaks of blood | 336
hemoglobin dropped | 336
upper GI endoscopy | 336
severe erythematous gastritis | 336
huge gastric ulcer | 336
non-bleeding visible vessel | 336
clipped | 336
sigmoidoscopy | 336
pale mucosa with ischemic changes | 336
biopsies obtained | 336
microscopic examination showed severe acute chronic inflammation | 336
fibrinous exudate | 336
extensive ulceration | 336
numerous fibrin microthrombi | 336
fungal microorganisms in the form of single and clustered small narrow-based budding yeasts | 336
diagnosed with GI cryptococcosis | 336
deteriorated with refractory septic shock | 408
multiorgan failure | 408
passed away | 408