32 years old | 0
male | 0
worsening epigastric pain | -48
ruptured appendicitis | 0
laparoscopic appendectomy | 0
discharged home | 0
fevers | 0
abdominal pain | 0
severe, worsening right upper quadrant epigastric pain | 168
radiating to the back | 168
no guarding | 168
no rebound tenderness | 168
no abdominal ecchymosis | 168
denied alcohol use | 168
denied recreational drug use | 168
no history of oropharyngeal infection | 168
no history of respiratory tract infection | 168
septic shock | 168
temperature 103 °F | 168
pulse 108 beats/minute | 168
mean arterial pressure 47 mmHg | 168
oral examination unremarkable | 168
neck examination unremarkable | 168
respiratory examination unremarkable | 168
cardiovascular examination unremarkable | 168
neurological examination unremarkable | 168
transferred to medical intensive care unit | 168
aggressive fluid resuscitation | 168
vasopressors | 168
initiation of vancomycin | 168
initiation of piperacillin/tazobactam | 168
elevated white blood cell count | 168
absolute neutrophil count 12,400 cells/mm³ | 168
normal platelet count | 168
normal hemoglobin | 168
normal electrolytes | 168
normal renal function | 168
normal pancreatic enzymes | 168
normal liver function tests | 168
negative urine drug screen | 168
negative blood alcohol test | 168
negative HIV ELISA | 168
negative viral hepatitis profile | 168
splenomegaly | 168
acute thrombosis of the proximal main portal vein | 168
acute thrombosis of superior mesenteric vein | 168
acute thrombosis of splenic vein | 168
no hepatic abnormalities | 168
no cirrhosis | 168
no infarct | 168
no abscess | 168
no cavernous transformation | 168
negative hypercoagulability workup | 168
F. necrophorum identification | 144
discontinued vancomycin | 144
added metronidazole | 144
anticoagulated with intravenous heparin | 144
persistent abdominal pain | 144
thrombus progression | 144
cavernous transformation of the portal vein | 144
transhepatic endovascular thrombolysis | 144
successful recanalization of porto-mesenteric veins | 144
discharged home on warfarin | 144
discharged home on clindamycin | 144
complete symptom relief | 144
