46 years old| 0
    female | 0
    underwent elective sleeve gastrectomy | 0
    obesity | 0
    psoriatic arthritis | 0
    multiple immunosuppressants | 0
    surgical hypoparathyroidism | -175200
    hypothyroidism | -175200
    total thyroidectomy | -175200
    multinodular goitre | -175200
    no history of diabetes | 0
    no history of dyslipidaemia | 0
    no history of hypertension | 0
    no history of obstructive sleep apnoea | 0
    hypoparathyroidism managed on oral calcium carbonate | -175200
    hypoparathyroidism managed on calcitriol | -175200
    emergency Roux-en-Y gastric bypass surgery | 0
    multiple gastric perforations | 0
    friable mucosa | 0
    abdominal sepsis | 96
    transfer to intensive care | 96
    nil orally | 96
    calcium level 0.78 mmol/L | 96
    asymptomatic without seizure | 96
    asymptomatic without arrhythmia | 96
    continuous intravenous calcium gluconate infusion | 96
    maintenance intermittent IV calcium boluses | 96
    prolonged ICU admission 6 months | 96
    required more than 20 abdominal operations | 96
    received all medication intravenously | 96
    received nutrition intravenously | 96
    lost 14 kg | 96
    Endocrinology advice for hypoparathyroidism | 96
    Endocrinology advice for hypothyroidism | 96
    TSH 5.83 mU/L | 408
    intravenous triiodothyronine 10 µg BD | 408
    euthyroidism achieved | 408
    high dose intravenous calcium 4.4 mmol five times daily | 408
    serum phosphate level 1.07 mmol/L | 408
    intravenous calcitriol 1 µg alternate daily | 1008
    intravenous calcitriol ceased | 1008
    intramuscular cholecalciferol 150 000 units | 1344
    1,25(OH)vitamin D3 level 31 pmol/L | 1344
    1,25(OH)vitamin D3 level 29 pmol/L | 2184
    eGFR > 90 mL/min/1.73 m² | 2184
    intravenous calcium gluconate 4.4 mmol five times daily | 2184
    intravenous calcitriol recommenced 1 µg alternate daily | 2184
    calcium gluconate requirements reduced to 4.4 mmol three times per day | 2184
    intramuscular thyroxine 600 µg | 2184
    intravenous thyroxine 200 µg alternate daily | 2184
    maintenance schedule established | 2184
    discharged | 5760
    recommenced oral intake | 5760
    calcitriol 0.75 µg daily | 5760
    calcium 1200 mg orally twice daily | 5760
    normocalcaemia 6 weeks post-discharge | 6384
    normocalcaemia 12 weeks post-discharge | 8736
    normocalcaemia 4 months post-discharge | 11040
    weight 71.8 kg | 11040
    BMI 29 kg/m² | 11040

<|eot_id|>
