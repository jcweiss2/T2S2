16 years old | 0 | 0 
primigravida | 0 | 0 
admitted to the emergency room | 0 | 0 
pregnancy diagnosis of 37.6 weeks of gestation | -672 | 0 
viable intrauterine pregnancy | -672 | 0 
fetal heart rate of 143 beats per minute | -672 | 0 
fetus situated longitudinally with cephalic presentation | -672 | 0 
back to the left | -672 | 0 
cervix 6 cm dilated | -5 | 0 
70% effaced | -5 | 0 
station +1 | -5 | 0 
intact membranes | -5 | 0 
mild edema of the extremities | -5 | 0 
normal osteotendinous reflexes | -5 | 0 
obstetrical ultrasound | -5 | 0 
pregnancy of 37+0 weeks of gestation | -5 | 0 
posterior body placenta maturation grade III | -5 | 0 
amniotic fluid index of 8.7 cm | -5 | 0 
biophysical profile of 8/8 | -5 | 0 
Hadlock of 34.2% | -5 | 0 
weight of 3033 grams | -5 | 0 
labor monitoring | 0 | 5 
spontaneous rupture of the membranes | 0 | 0 
labor progressed | 0 | 5 
effective labor | 0 | 5 
4 contractions every 10 minutes | 0 | 5 
contractions lasted 40 to 45 seconds | 0 | 5 
live newborn delivered | 5 | 5 
Apgar scores of 7 and 9 | 5 | 5 
gestational age of 40 weeks | 5 | 5 
height 48 cm | 5 | 5 
weight of 2650 grams | 5 | 5 
placenta came out with normal characteristics | 5 | 5 
grade III uterine inversion | 5 | 5 
manual reinversion maneuvers | 5 | 5 
total blood loss of 1200 mL | 5 | 24 
uterine atony | 5 | 24 
oxytocin | 5 | 24 
carbetocin | 5 | 24 
misoprostol | 5 | 24 
persistent uterine inversion | 5 | 24 
exploratory laparotomy | 5 | 24 
reinversion of the uterus | 10 | 10 
persistent uterine atony | 10 | 24 
persistent postpartum hemorrhage | 10 | 24 
Hayman hemostatic suture | 15 | 15 
bilateral ligation of the anterior trunk of the hypogastric artery | 20 | 20 
recovery of uterine tone | 20 | 20 
cessation of postpartum hemorrhage | 20 | 20 
postligation bleeding of 50 mL | 20 | 24 
transfusion of 2 bags of packed red blood cells | 15 | 24 
transfer to the recovery room | 24 | 24 
transfer to the medical intensive care unit | 24 | 24 
transfer to a hospital room | 48 | 48 
normal diet | 48 | 48 
ambulation | 48 | 48 
spontaneous uresis | 48 | 48 
normal peristalsis | 48 | 48 
breastfeeding | 48 | 48 
discharge from the hospital | 48 | 48