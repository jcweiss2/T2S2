demyelination | 0
destruction of myelin-supporting cells | 0
oligodendrocytes | 0
schwann cells | 0
central nervous system | 0
peripheral nervous system | 0
dysmyelination | 0
genetic defect | 0
synthesis and turnover of myelin membranes | 0
leukodystrophy | 0
central demyelination | 0
peripheral demyelination | 0
Multiple sclerosis | 0
inflammatory demyelination | 0
geographical variation | 0
women | 0
men | 0
age of presentation | 0
Acute-disseminated encephalomyelitis (ADEM) | 0
post-infectious encephalomyelitis | 0
T-cell hypersensitivity reaction | 0
viral infection | 0
measles | 0
mumps | 0
rubella | 0
varicella-zoster | 0
Epstein-Barr virus (EBV) | 0
cytomegalovirus (CMV) | 0
herpes simplex virus | 0
hepatitis A | 0
hepatitis B | 0
Coxsackie virus | 0
influenza A | 0
influenza B | 0
human immunodeficiency virus (HIV) | 0
human T-cell lymphotropic virus-1 (HTLV-1) | 0
bacterial infection | 0
Mycoplasma pneumoniae | 0
Campylobacter jejuni | 0
Leptospira | 0
group A Streptococci | 0
Borrelia | 0
Chlamydia | 0
Legionella | 0
vaccines | 0
diphtheria–tetanus–polio | 0
rabies | 0
hepatitis B | 0
measles | 0
mumps | 0
smallpox | 0
rubella | 0
Japanese B encephalitis | 0
pertussis | 0
influenza | 0
Etanercept | 0
Botulinum Toxin Type A | 0
Adalimumab | 0
Eculizumab | 0
Lansoprazole | 0
Oxcarbazepine | 0
gonadotropins | 0
Acute hemorrhagic leucoencephalitis (AHL) | 0
hyper acute variant | 0
viral infection | 0
M pneumoniae infection | 0
anti-tubercular drugs | 0
inhalational anesthetic agents | 0
isoflurane | 0
desflurane | 0
ulcerative colitis | 0
Crohn's disease | 0
septicemia | 0
Osmotic demyelination syndromes | 0
osmotic stress | 0
disruption of the blood-brain barrier (BBB) | 0
central pontine myelinolysis (CPM) | 0
extrapontine myelinolysis (EPM) | 0
alcoholism | 0
malnutrition | 0
hypoxic-ischemic states | 0
deep burns | 0
intensive care treatment | 0
metabolic disorders | 0
uremia | 0
prolonged diuretic use | 0
dialysis | 0
diabetes | 0
liver transplantation | 0
psychogenic polydipsia | 0
burns | 0
post-pituitary surgery | 0
post-urological surgery | 0
gynecological surgery | 0
glycine infusions | 0
Viral demyelination | 0
Progressive multifocal leukoencephalopathy (PML) | 0
JC papovavirus (JCV) | 0
childhood | 0
adolescence | 0
immunosuppressed conditions | 0
cell-mediated immunity | 0
immunosuppressive drug therapy | 0
antibody-based regimens | 0
autoimmune-disease patients | 0
multiple sclerosis | 0
Crohn's disease | 0
Subacute sclerosing panencephalitis (SSPE) | 0
measles virus infection | 0
neurons | 0
glial cells | 0
oligodendrocytes | 0
immune response | 0
children | 0
young adults | 0
boys | 0
girls | 0
mandatory immunization | 0
Guillain-Barré syndrome | 0
acute-onset immune-mediated disease | 0
infections | 0
Campylobacter jejuni | 0
cytomegalovirus (CMV) | 0
Mycoplasma pneumonia | 0
Epstein-Barr virus | 0
influenza virus | 0
molecular mimicry | 0
epitopes | 0
peripheral nerves | 0
infectious agents | 0
surgery | 0
vaccination | 0
parturition | 0
Acute Inflammatory Demyelinating Polyradiculoneuropathy (AIDP) | 0
Miller Fisher syndrome (MFS) | 0
anti-GQ1b | 0
anti-GT1a | 0
Chronic inflammatory demyelinating polyradiculoneuropathy | 0
acquired demyelinating syndrome | 0
myelin sheaths | 0
peripheral nervous system | 0
cellular immunity | 0
T-cell activation | 0
humoral immune system | 0
immunoglobulin | 0
complement deposition | 0
myelinated nerve fibers | 0
Lewis-Sumner syndrome | 0
multi-focal acquired demyelinating sensory and motor neuropathy (MADSAM) | 0
sensory-predominant CIDP | 0
distal acquired demyelinating sensory neuropathy (DADS) | 0
IgM paraprotein | 0
CIDP with central nervous system involvement | 0
steroids | 0
plasma exchange | 0
IVIg | 0
Paraproteinemic demyelinating neuropathy | 0
paraprotein | 0
immunoglobulin molecule | 0
monoclonal plasma cell expansion | 0
monoclonal gammopathy | 0
MGUS | 0
IgM PDN | 0
IgG | 0
IgA | 0
myelin-associated glycoprotein | 0
anti-myelin-associated antibodies | 0
Charcot Marie Tooth type 1 | 0
Charcot Marie Tooth type X | 0
peripheral nerve myelin protein 22 (PMP22) | 0
GJB1 gene | 0
connexin 32 | 0
X-chromosome | 0
Copper deficiency | 0
copper containing metalloenzymes | 0
superoxide dismutase (SOD) | 0
CNS demyelination | 0
Combined central and peripheral demyelination | 0
Acute combined central and peripheral inflammatory demyelination | 0
MS with idiopathic inflammatory-demyelinating neuropathy | 0
simultaneous GBS and ADEM | 0
pediatric population | 0
cerebral involvement | 0
acute and relapsing polyneuropathy | 0
chronic autoimmune hepatitis | 0
CIDP | 0
central pontine myelinolysis (CPM) | 0
MRI | 0
brain | 0
spinal roots | 0
brachial plexus | 0
lumbosacral plexus | 0
cauda equina | 0
nerve regions | 0
Electrodiagnostic testing | 0
nerve conduction studies | 0
cerebrospinal fluid analysis | 0
brain biopsy | 0
nerve biopsy | 0
laboratory studies | 0