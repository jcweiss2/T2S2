3.28 kg | 0
    female | 0
    born at 40 weeks gestation | 0
    mother with history of two abortions | 0
    third pregnancy | 0
    delivered by caesarean section | 0
    scoliosis | 0
    right hydronephrosis | 0
    active stagnation | 0
    suspected intrauterine infection | 0
    prenatal screening tests unremarkable | 0
    no evidence of C. albicans in vaginal secretion six months previously | 0
    no antibiotics for UTI or other bacterial infection in previous six months | 0
    mother developed fever 38.0°C two hours before birth | -2
    amniotomy performed | -2
    IV oxytocin 2 mU/min | -2
    IV cefuroxime sodium 1.5 g | -2
    Apgar score 8/9 at 1 minute | 0
    Apgar score 8/9 at 5 minutes | 0
    amniotic fluid clear without meconium staining | 0
    severe acute chorioamnionitis | 0
    moderate umbilical vasculitis | 0
    neutrophilic infiltration in placenta | 0
    cellulose attachment in villi | 0
    admitted to NICU | 0
    groaning | 0
    spitting | 0
    generalized erythematous papular eruption | 0
    pustules observed | 72
    desquamation observed | 72
    palms affected | 72
    soles affected | 72
    skin scrapings negative for Candida spp | 72
    no oral thrush | 72
    no perianal thrush | 72
    transient respiratory distress | 0
    low-flow oxygen for two days | 0
    decreased transmittance chest X-ray | 0
    increase in CRP levels 68.2 mg/l | 18
    leucocytosis with left shift | 18
    lumbar puncture | 18
    CSF culture negative | 18
    CSF WBC count 15 cells/mm3 | 18
    CSF protein 63.4 mg/dl | 18
    CSF glucose 2.5 mmol/l | 18
    treated with cefoperazone/sulbactam | 0
    treated with penicillin | 0
    differential diagnosis of rash | 0
    skin rash desquamated | 168
    excoriated lesions persisted | 168
    WBC count normal | 168
    CRP levels normal | 168
    antibiotics stopped | 168
    blood culture positive for C. albicans | 168
    urine culture positive for C. albicans | 168
    skin culture positive for C. albicans | 168
    serum (1–3)-β-D-glucan assay negative | 168
    started on IV fluconazole | 168
    topical miconazole nitrate | 168
    high-throughput DNA sequencing negative | 312
    urine cultures negative | 312
    increase in acute phase reactants | 480
    sepsis suspected | 480
    urinary tract infection | 480
    started on ceftazidime | 480
    IV fluconazole stopped | 480
    oral fluconazole initiated | 480
    persistence of UTI | 672
    E. coli | 672
    Enterococcus faecium | 672
    serial treatment with piperacillin/tazobactam | 672
    started vancomycin | 840
    cutaneous lesions resolved | 528
    recurrent bacterial UTIs | 0
    immune deficiency suspected | 0
    blood immunity-related genetic analysis | 0
    immune function tests | 0
    normal immune function | 0
    excluded chronic granulomatous disease | 0
    excluded galactosemia | 0
    vesicoureteral reflux suspected | 0
    voiding cystourethrography not performed | 0
    repeat urine cultures sterile | 240
    urine routine examinations normal | 240
    audiometry normal | 240
    ophthalmologic examination | 384
    brain MRI normal | 384
    chest CT normal | 312
    liver ultrasonography normal | 72
    renal ultrasonography normal | 72
    bladder ultrasonography normal | 72
    99mTc-DMSA static renal scan normal | 1176
    echocardiogram showed atrial septal defect | 72
    patent foramen ovale | 72
    discharged | 1440
    good development | 1440
    congenital systemic candidiasis | 0
    CCC | 0
    candidemia due to C. albicans | 168
    invasive C. albicans | 168
    treated with IV fluconazole | 168
    treated with topical fluconazole | 168
    total fluconazole treatment six weeks | 0
    resolved UTIs | 240
    small atrial septal defect | 72
    patent foramen ovale without endocarditis | 72
    normal brain MRI | 384
    normal chest CT | 312
    normal liver | 72
    normal renal | 72
    normal bladder | 72
    normal 99mTc-DMSA scan | 1176
    no endocarditis | 72
    