28 years old | 0
male | 0
presented to casualty | 0
near drowning in a paper factory | -120
ventilated | -120
acute respiratory distress syndrome | -120
received ceftriaxone | -120
received empiric antibiotic | -120
received other therapies | -120
presented with high-grade fever | 0
presented with tachypnea | 0
oxygen saturation of 87% | 0
lab investigations revealed leukocytosis (17,200/cumm) | 0
hemoglobin 11.1 g% | 0
normal electrolytes | 0
creatinine of 1.8 mg/dl | 0
endotracheal secretions sent for gram stain | 0
endotracheal secretions sent for fungal stain | 0
endotracheal secretions sent for acid-fast stain | 0
endotracheal secretions sent for cultures | 0
blood sent for gram stain | 0
blood sent for fungal stain | 0
blood sent for acid-fast stain |0
blood sent for cultures |0
urine samples sent for gram stain |0
urine samples sent for fungal stain |0
urine samples sent for acid-fast stain |0
urine samples sent for cultures |0
antibiotic coverage changed to cefoperazone + sulbactam |0
chest X-ray revealed bilateral alveolar shadows |0
chest X-ray revealed cystic lesion in the lung parenchyma |0
CT brain showed multiple ill-defined round hypodense lesions in bilateral cerebral hemispheres |0
CT brain showed surrounding edema |0
CT chest showed multiple well-defined round nodular lesions scattered in both lungs |0
CT chest showed few lesions with central cavitation |0
CT abdomen revealed patchy hypodensities in both kidneys |0
CT abdomen revealed patchy hypodensities in the gluteal muscles bilaterally |0
echocardiography was normal |0
BAL performed |0
transbronchial biopsy performed |0
antibiotic escalated to meropenem |0
all microbiological laboratory reports negative |48
serum galactomannan (1.5) raised |48
endotracheal aspirate fungal stain showed Aspergillus species |48
voriconazole started |48
caspofungin started |48
suspicion of invasive aspergillosis |48
hemodynamic instability |48
developed hemoptysis |48
developed tachycardia |48
developed desaturation |48
controlled with fresh frozen plasma |48
controlled with tranexamic acid |48
developed septic shock |72
requiring vasopressors |72
worsening respiratory acidosis |72
leukopenia (2200/cumm) |72
transbronchial biopsy revealed neutrophilic exudates |72
transbronchial biopsy revealed foci of fungal broad hyphae |72
transbronchial biopsy revealed broad angle branching |72
BAL culture revealed Aspergillus fumigatus growth |72
expired |120
severe multiorgan dysfunction |120
