61 years old | 0
male | 0
presented to hospital | 0
transient loss of consciousness | 0
acute chest discomfort | 0
upper respiratory tract infection | -336
subjective fever | -24
rigors | -24
apyrexic | 0
initial physical examination normal | 0
serum leukocyte count normal | 0
chest radiograph normal | 0
12-lead electrocardiogram demonstrated inferior ST-segment elevation myocardial infarction | 0
no stigmata of endocarditis | 0
no signs of aortic dissection | 0
intravenous thrombolysis administered | 0
transferred to tertiary care hospital | 0
coronary angiography demonstrated occlusion of distal left-dominant posterior descending artery | 0
angioplasty not possible | 0
transthoracic echocardiography showed left ventricular apical-inferior hypokinesis | 0
no valve lesions | 0
cranial computed tomography identified small cerebellar hemorrhage | 0
transferred to cardiac intensive care unit | 0
onset of polymorphic ventricular tachycardia storm | 24
profound shock | 24
admission blood cultures grew methicillin-sensitive Staphylococcus aureus | 0
intravenous antibiotics administered | 0
maximum supportive therapy | 0
died | 48
autopsy revealed acute bacterial myocarditis | 48
multifocal suppuration of lower interventricular septum and inferior ventricles | 48
cardiac valves unremarkable | 48
intramyocardial abscesses contained gram-positive cocci | 48
posterior descending artery exhibited acute bacterial vasculitis | 48
adjacent abscess | 48
microabscesses in brain and spinal cord | 48