76 years old | 0
female | 0
hypertension | -175200
type II diabetes mellitus | -175200
coronary heart disease | -175200
myocardial infarction | -131400
senile dementia | -175200
open cholecystectomy | -2620800
abdominal wall hernia repairs (five occasions) | -175200
morbid obesity | 0
BMI 37.8 kg/m² | 0
no regular alcohol consumption | 0
no smoking | 0
progressive abdominal pain | -120
admission | 0
weak general condition | 0
status febrilis | 0
septico-toxic shock | 0
acute abdomen | 0
eventrated hernia (size of a handball) | 0
local defense musculaire (right subcostal region) | 0
abdominal ultrasonography | 0
laboratory tests | 0
chest X-ray | 0
native abdominal X-ray | 0
central venous access | 0
epidural cannulation | 0
intravesical catheter insertion | 0
urgent right upper transverse laparotomy | 0
general anesthesia | 0
complete muscle relaxation | 0
local feculent peritonitis | 0
subcutaneous inflammatory oedema | 0
incarcerated and perforated ascending colon | 0
perforated terminal ileum | 0
extended right hemicolectomy | 0
resection of terminal ileum (60 cm) | 0
side-to-side ileo-transversostomy | 0
necrectomy | 0
abdominal gap (223 cm²) | 0
closure defect by direct sutures (not possible) | 0
biological graft unavailable | 0
synthetic mesh implantation (not considered) | 0
dermal-subcutaneous pannicule removal | 0
epidermis removal | 0
subcutaneous adipose tissue removal | 0
dermal flaps preparation | 0
first homogeneous dermal graft insertion | 0
dermal graft fixation (interrupted 2/0 non7absorbable stitches) | 0
external dermal graft fixation | 0
external dermal graft perforation | 0
greater omentum spared | 0
no direct abdominal sutures | 0
surgery duration (250 minutes) | 0
dermal graft preparation duration (50 minutes) | 0
intraoperative blood loss (740 mL) | 0
intensive care (first 4 postoperative days) | 24
imipenem/cilastatin antibiotic therapy | 0
enoxaparin thrombosis prophylaxis | 6
fever cessation (4th postoperative day) | 96
bowel movement restart (Mannitol solution) | 120
red blood cell transfusions (5 units) | 120
nasogastric tube (removed on 3rd day) | 72
respiratory function normal | 0
kidney function normal | 0
O2 saturation 92-95% | 0
urine production >1600 mL/day | 0
oral nourishment (160/80 g carbohydrate/protein diet) | 120
mobilization (5th postoperative day) | 120
elastic abdominal belt application | 120
intra-abdominal drain removal (6th day) | 144
left subcutaneous drain removal (7th day) | 168
right subcutaneous drain removal (10th day) | 240
skin sutures removal (15th day) | 360
no seroma | 0
no diffuse subcutaneous fluid accumulation | 0
discharge (18th postoperative day) | 432
enoxaparin s.c. prescribed for 21 days | 432
wound healing per primam intentionem | 432
elastic bandage instruction | 432
avoid bloating food | 432
physical examinations (1st and 3rd month) | 720
blood tests (1st and 3rd month) | 720
abdominal wall ultrasonographies (1st and 3rd month) | 720
abdominal computed tomography (6th month) | 4320
no hernia recurrence | 4320
no subcutaneous fistula | 4320
no seroma formation | 4320
