45 years old | 0
female | 0
history of hypertension | -336
history of type 2 diabetes | -336
presented to emergency department | 0
acute onset of chest pain | 0
chest pain radiating to left arm | 0
diaphoresis | 0
shortness of breath | 0
last seen by primary care physician | -336
routine check-up | -336
medications included metformin | -336
medications included lisinopril | -336
medications included atorvastatin | -336
elevated blood pressure | 0
heart rate of 110 bpm | 0
oxygen saturation of 92% on room air | 0
ECG showed ST-segment elevation | 0
diagnosed with AMI | 0
started on aspirin | 0
started on clopidogrel | 0
started on intravenous heparin | 0
PCI performed | 3
drug-eluting stent placed in LAD artery | 3
transferred to CCU | 3
developed atrial fibrillation | 15
managed with rate control | 15
managed with anticoagulation | 15
discharged on day 5 | 120
new prescription for beta-blocker | 120
continuation of previous medications | 120
referral to cardiac rehabilitation program | 120