58 years old|0
female|0
alcoholism|0
chronic obstructive pulmonary disease|0
tobacco abuse|0
presented with shortness of breath|0
presented with cough|0
admitted to the hospital|0
respiratory rate of 32 breaths/min|0
temperature of 38.0°C|0
heart rate of 115 bpm|0
blood pressure of 73/40 mmHg|0
oxygen saturation of 72% on room air|0
lethargic|0
arousable to voice|0
tachycardic|0
regular rhythm|0
no murmurs|0
mild respiratory distress|0
coarse rhonchi|0
warm extremities|0
strong pulses|0
white blood cell count 12.4×103 cells/uL|0
arterial blood gas pH 7.07|0
arterial blood gas pCO2 106 mmHg|0
arterial blood gas pO2 80 mmHg|0
arterial blood gas bicarbonate 30 mmol/L|0
chest X-ray no acute pathology|0
CT imaging multifocal pneumonia|0
diagnosed with septic shock|0
community-acquired pneumonia|0
started on ceftriaxone|0
started on azithromycin|0
fluid resuscitation with 3 liters of lactated ringers|0
low blood pressure|0
started on norepinephrine|0
SpO2 83% on 15 L O2 via non-rebreather mask|0
intubated|0
blood cultures negative|0
respiratory cultures negative|0
liberated from norepinephrine on hospital day 2|24
FiO2 40% on hospital day 5|120
PEEP 5 cm H2O on hospital day 5|120
FiO2 30% on hospital day 6|144
PEEP 5 cm H2O on hospital day 6|144
extubated on hospital day 6|144
respiratory distress on hospital day 6|144
respiratory rate of 28 breaths/min|144
temperature of 38.2°C|144
heart rate of 112 bpm|144
blood pressure of 80/55 mmHg|144
oxygen saturation of 85% on 60 L heated high-flow oxygen therapy|144
arterial blood gas pH 7.32|144
arterial blood gas pCO2 56 mmHg|144
arterial blood gas pO2 78 mmHg|144
arterial blood gas bicarbonate 24 mmol/L|144
re-intubated|144
restarted on norepinephrine|144
FiO2 100%|144
PEEP 5 cm H2O|144
repeat CXR new left lower lobe infiltrate|144
diagnosed with ventilator-associated pneumonia|144
started on vancomycin|144
started on cefepime|144
MRSA nasal swab negative|144
vancomycin discontinued on hospital day 7|168
continued on cefepime monotherapy|168
fevers up to 38.2°C|168
up-trending leukocytosis|168
ongoing vasopressor need|168
endotracheal aspirate culture positive for MRSA|216
MRSA resistant to oxacillin|216
MRSA resistant to clindamycin|216
MRSA resistant to erythromycin|216
MRSA sensitive to linezolid|216
MRSA sensitive to tetracycline|216
MRSA sensitive to gentamycin|216
MRSA sensitive to trimethoprim/sulfamethoxazole|216
MRSA sensitive to vancomycin|216
blood cultures negative|216
restarted on vancomycin|216
liberated from norepinephrine|216
liberated from ventilator|216
transferred out of ICU|216
completed 7 days of intravenous vancomycin|216
