45 years old | 0
male | 0
chronic smoker | 0
admitted to hospital | 0
blunt chest trauma | -2160
chest pain | -2160
respiratory distress | -2160
two prior admissions | -2160
high-resolution computed tomography (HRCT) | 0
bilateral hydropneumothorax | 0
multiple rib fractures | 0
shifted to intensive care unit (ICU) | 0
signs of respiratory failure | 0
bilateral chest tubes | 0
intermittent non-invasive ventilation (NIV) | 0
antibiotics | 0
adequate analgesia | 0
supportive management | 0
chest tubes removed | 24
minimal fluid on ultrasound chest | 24
dyspnoea persisted | 24
repeat HRCT chest | 24
infective pathology (atypical pneumonia) | 24
lesions in the apical segment of right upper lobe | 24
lymphangitis carcinomatosa | 24
arterial blood gases reported | 24
persistently high pCO2 | 24
mild hypoxia | 24
acute exacerbation of COPD | 24
type 2 respiratory failure | 24
oral steroid started | 24
20-30% improvement in dyspnoea | 48
NIV 3-4 hours/day | 48
echocardiography done | 48
normal echocardiography | 48
repeat contrast-enhanced computed tomography (CECT) lung | 336
spiculated nodule in upper part of right lower lobe | 336
multiple sclerotic lesions in vertebral body of D1 and sternum | 336
lytic lesion in D11 | 336
ultrasound abdomen | 336
hepatomegaly | 336
multiple space-occupying lesions in both lobes of the liver | 336
fine-needle aspiration cytology | 336
adenocarcinoma metastasis | 336
chemotherapy could not be started | 336
poor general condition of patient | 336
expired | 346
occult primary malignancy | 336
pulmonary lymphangitis carcinomatosa (PLC) | 336
liver metastasis | 336