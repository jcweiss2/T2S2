33 years old | 0
male | 0
alcohol use disorder | -672
seizures | -672
admitted to the emergency room | 0
hypothermic | 0
tachypneic | 0
required Bi-level Positive Airway Pressure ventilation | 0
cirrhotic liver | 0
large volume ascites | 0
bilateral pleural effusions | 0
anion gap metabolic acidosis | 0
sepsis | 0
urinary tract infection | 0
cirrhosis | 0
hypoxemic respiratory failure | 0
admitted to the step down unit | 0
thoracentesis | 24
paracentesis | 24
developed melena | 72
gastroenterology consulted | 72
interventional radiology consulted | 72
TIPS procedure planned | 72
MELD score calculated | 216
MELD score 19 | 216
TIPS procedure performed | 216
1 unit of platelets transfused | 216
ultrasound-guided access through the right internal jugular vein | 216
angiography and hepatic venography | 216
TIPs puncture needle rotated and advanced to the portal vein | 216
guidewire inserted to confirm portal vein access | 216
angiographic catheter advanced into the portal vein | 216
venography repeated to visualize varices | 216
track dilated with a balloon catheter | 216
stent deployed | 216
portal pressure measured for gradient reduction | 216
venography repeated to confirm variceal bleeding had stopped | 216
somnolent | 216
systolic blood pressure in the 80s | 216
rapid response called | 216
hemoglobin levels decreased | 216
white blood cell count elevated | 216
2 units of red blood cells transfused | 216
CT abdomen performed | 216
shunt patent | 216
large area of decreased enhancement of the liver | 216
dense material within the lesser sac and along the lateral border of the liver | 216
hemoperitoneum | 216
upgraded to the intensive care unit | 216
4 units of red blood cells transfused | 216
5% albumin transfused | 216
2 units of cryoprecipitate transfused | 216
3 units of fresh frozen plasma transfused | 216
multiple transfusions due to drop in hemoglobin levels | 240
hematology consulted | 240
coagulopathy | 240
prolonged INR/PT and aPTT levels | 240
10 mg of intravenous vitamin K daily for 3 days | 240
cryoprecipitate to achieve a fibrinogen level of 100-120 | 240
platelet count maintained above 50,000 | 240
1000 micrograms of subcutaneous cyanocobalamin once | 240
ferrous sulfate supplementation 3 times a day | 240
folic acid supplementation continued | 240
angiogram performed | 384
no active extravasation | 384
post-TIPs venogram performed | 384
patent TIPs shunt | 384
hemoglobin and hematocrit stabilized | 408
discharged from the hospital | 408
referred for transfer to a liver transplant center | 408
denied transfer | 408
advised to follow up as an outpatient with an end-stage renal disease center | 408