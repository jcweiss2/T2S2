18 years old | 0
male | 0
hypertension | 0
degenerative joint disease | 0
bilateral knee replacement | 0
substance abuse | 0
trauma to his face and chest wall | 0
lightheadedness | 0
fatigue | 0
leukocytosis | 0
hemoglobin | 0
venous lactic acid | 0
intramuscular and subpectoral hematoma | -48
extrapleural extension into the chest | -48
acute right second through fifth anterior rib fractures | -48
bilateral lower lobe bronchopneumonia | -48
blood cultures | -48
empiric antibiotics | -48
afebrile | -48
hypotensive | -48
suspected septic shock | -48
vasopressors | -48
Day 2 of hospitalization | -48
antibiotics broadened | -48
vancomycin | -48
cefepime | -48
metronidazole | -48
repeat blood, urine and sputum cultures | -48
blood and urine cultures negative | -48
sputum cultures grew methicillin-resistant Staphylococcus aureus | -48
antibiotics narrowed | -48
vancomycin | -48
Day 4 of hospitalization | -48
left knee pain | -96
notable swelling on physical exam | -96
concern for infection of his prosthetic knee joint | -96
sterile left knee aspiration | -96
synovial fluid was cloudy, amber colored | -96
white blood cells of 9.28 × 10^3/mcL | -96
6.0 × 10^3/mcL | -96
calcium pyrophosphate crystals | -96
complete washout and debridement of the joint | -96
retention of the prosthesis | -96
operative note described an infected knee with purulence | -96
five cultures from the infected area | -96
joint specimen | -96
tissue specimen | -96
fluid specimen | -96
anaerobic and aerobic media | -96
antibiotic regimen transitioned | -96
cefazolin | -96
postoperative Day 1 | -96
hospitalization Day 7 | -96
C. bifermentans | -96
ampicillin–sulbactam | -96
oral suppression with amoxicillin–clavulanic acid | -96
contrast computerized tomography scan of the abdomen | -96
negative | -96
human immunodeficiency virus screening | -96
negative | -96
clinically improve | -96
discharged to a rehabilitation facility | -96
referral to gastroenterology for outpatient colonoscopy | -96
follow-up with internal medicine | -96
recovered full range of motion of his left knee | -96
no signs of lingering joint or systemic infection | -96
still taking Augmentin | -96
reported medication adherence | -96
colonoscopy to investigate for source of infection | -96
septic arthritis | -672
empyema | -672
osteomyelitis | -672
soft tissue infection | -672
brain abscess | -672
bacteremia | -672
endocarditis | -672
meniscectomy | -672
arthrotomy and debridement of the joint | -672
intra-articular and intravenous penicillin | -672
oral penicillin | -672
debridement, antibiotics and implant retention (DAIR) procedure | -96
stable, well-fixed implant | -96
mechanical loosening or sinus tracts | -96
uniform susceptibility of C. bifermentans to antibiotics | -96
Infectious Diseases Society of America guidelines | -96
2 weeks of intravenous antibiotics | -96
6 months of oral antibiotics | -96
suppressive antibiotics | -96
spore-forming bacterium | -96
resistant to antibiotics when in spore form | -96
treatment failure | -96
4-fold increased risk of treatment failure | -96
discontinuing oral antibiotics | -96
two-stage arthroplasty | -96
PJI with C. bifermentans | -96
DAIR | -96
prosthesis to be retained without complication | -96
immediate postoperative period | -96
further case reports and long-term outcome follow-up | -96
treatment of the joint with DAIR | -96
prosthesis to be retained without complication | -96
immediate postoperative period | -96
long-term outcome follow-up | -96