35 years old | 0
man | 0
admitted to the hospital | 0
coughing | -168
respiratory distress | -24
no fever | 0
no nasal discharge | 0
no chest pain | 0
no hemoptysis | 0
no hematuria | 0
no passage of worms in stool | 0
denied atopy | 0
denied recent travel | 0
denied exposure to pets | 0
denied exposure to birds | 0
denied exposure to cotton | 0
denied exposure to dust | 0
denied exposure to metal fumes | 0
blood pressure 110/70 mmHg | 0
pulse rate 112 beats/minute | 0
respiratory rate 30 breaths/minute | 0
pallor | 0
use of accessory muscles of respiration | 0
no lymphadenopathy | 0
no cyanosis | 0
no clubbing | 0
no pedal edema | 0
no palpable purpura | 0
jugular venous pressure not elevated | 0
bilateral rhonchi | 0
crackles | 0
liver palpable 4 cm | 0
spleen palpable 5 cm | 0
hemoglobin 8.3 g/dL | 0
white cell count 27.6×10^9/L | 0
differential count 39% polymorphs | 0
differential count 11% lymphocytes | 0
differential count 2% monocytes | 0
differential count 48% eosinophils | 0
absolute eosinophil count 13.2×10^9/L | 0
platelet count 420×10^9/L | 0
erythrocyte sedimentation rate 24 mm/hour | 0
lactate dehydrogenase 1000 U/L | 0
uric acid 565 µmol/L | 0
normal renal function | 0
normal liver function | 0
arterial blood gas pH 7.38 | 0
arterial blood gas partial pressure of oxygen 67 mmHg | 0
arterial blood gas partial pressure of carbon dioxide 35.5 mmHg | 0
oxygen saturation 85% | 0
chest X-ray bilateral fluffy alveolar opacities | 0
cardiac size normal | 0
cardiac contour normal | 0
computed tomography symmetrical confluent airspace opacities | 0
computed tomography suggestive of pulmonary edema | 0
troponin I negative | 0
pulmonary capillary wedge pressure 5 mmHg | 0
serum procalcitonin 0.3 µg/L | 0
blood cultures sterile | 0
leptospira serology negative | 0
mycoplasma serology negative | 0
legionella serology negative | 0
filariasis serology negative | 0
strongyloides stercoralis serology negative | 0
legionella urine antigen negative | 0
anti-nuclear antibody negative | 0
anti-neutrophil cytoplasmic antibody negative | 0
stool examination no cysts/ova | 0
serum immunoglobulin E 708 IU/mL | 0
nerve conduction normal | 0
diethylcarbamazine 300 mg | 0
glucocorticoid oral prednisone 60 mg daily | 0
symptoms did not improve | 0
type-1 respiratory failure worsened | 0
bronchoscopy performed | 0
bronchoalveolar lavage eosinophil-rich infiltrate | 0
transbronchial lung biopsy fibroblastic proliferation | 0
transbronchial lung biopsy Masson bodies | 0
transbronchial lung biopsy eosinophils in interstitial spaces | 0
bone marrow examination granulocytic hyperplasia | 0
bone marrow examination marked increase in eosinophils | 0
bone marrow examination no blasts | 0
FIP1L1-PDGFRA mRNA detected | 0
BCR1-ABL1 mRNA not detected | 0
diagnosed with myeloid neoplasm associated with eosinophilia | 0
diagnosed with PDGFRA gene rearrangement | 0
imatinib 100 mg daily | 0
clinical improvement within 1 week | 168
radiological improvement within 1 week | 168
hematological improvement within 1 week | 168
complete hematological remission at 2 weeks | 336
normalization of peripheral blood counts | 336
no splenomegaly | 336
discharged | 336
regular follow-ups | 336
eosinophilia | 0
hypereosinophilic syndrome | 0
end organ damage | 0
myeloid neoplasm with PDGFRA rearrangement | 0
chronic eosinophilia not otherwise specified | 0
idiopathic hypereosinophilic syndrome | 0
hematological system involvement | 0
cardiovascular system involvement | 0
skin involvement | 0
nervous system involvement | 0
pulmonary system involvement | 0
nocturnal coughing | 0
wheezing | 0
productive sputum | 0
dyspnea | 0
radiographic abnormalities | 0
ground glass opacities | 0
patchy consolidation | 0
ARDS | 0
imatinib resistance | 0
molecular remission after imatinib re-initiation | 0
organomegaly | 0
elevated lactate dehydrogenase | 0
FIP1L1-PDGFRA transcripts identified | 0
no mechanical ventilation | 0
