60 years old | 0
female | 0
hepatitis C-related cirrhosis | -6720
recurrent hepatic encephalopathies | -6720
chronic portal vein thrombosis | -6720
liver transplantation | 0
end-to-side anastomosis of the donor portal vein to the superior mesenteric vein | 0
end-to-end bile duct anastomosis | 0
massive venous bleeding from local varices | 0
iliac conduit construction | 0
normal liver graft function | 0
stenosis of the bile duct anastomosis | -720
biliary leakage | -720
elevated liver enzymes | -720
pigtail treatment | -720
FCSCEMS insertion | -504
persisting leakage | -504
stent extraction | -168
hepatitis C reinfection | -168
recurrent stenosis of the biliary anastomosis | -168
ERCP | -168
balloon dilatations | -168
pigtail placements | -168
stent placements | -168
biopsy-proven significant fibrosis | -624
treatment with pegylated interferon and ribavirin | -624
elective ERCP | 0
biliary pigtail exchange | 0
portobiliary fistula diagnosis | 0
hemobilia | 0
FCSEMS placement | 0
prophylactic antibiotic treatment with ciprofloxacin | 0
septic shock | 48
admission to intensive care unit | 48
hemodynamic support | 48
empiric broad-spectrum antibiotic treatment | 48
computed tomography | 48
angiography | 48
chronic obliteration of the iliac conduit | 48
partial perfusion of the hepatic artery by gastroduodenal collaterals | 48
anuric kidney failure | 48
continuous venovenous hemofiltration | 48
intermittent hemodialysis | 48
recovery | 192
FCSEMS replacement | 3456
extraction of the lying FCSEMS | 3456
no evidence of persisting leakage | 3456
no relevant stenosis | 3456
follow-up | 7200
no evidence of recurrent stenosis or portobiliary fistula | 7200