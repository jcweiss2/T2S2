6-year-old girl | 0
    presented to the emergency department | 0
    severe headache | -48
    nausea | -48
    vomiting | -48
    family history of neurological disorders | 0
    no family history of neurological disorders | 0
    normal psychomotor development | 0
    recent episode of mumps infection | -240
    spontaneous resolution of mumps infection | -240
    altered consciousness level | 0
    mildly confused | 0
    Glasgow Coma Scale = E4 V4 M6 | 0
    trunk ataxia | 0
    gait ataxia | 0
    bilateral dysmetria on finger-nose tests | 0
    body temperature 37.5 °C | 0
    normal heart rate | 0
    normal breath rate | 0
    dysautonomic troubles | +few
    heart rate decreased to 55 beats/min | +few
    arterial pressure dropped to 80/50 mmHg | +few
    transferred to the Pediatric Intensive Care Unit | +few
    brain computed tomography scan | +few
    cerebellar ill-defined hypodense lesion | +few
    mass effect on the fourth ventricle | +few
    dilation of the upper ventricular system | +few
    multimodal magnetic resonance imaging performed | +few
    cerebellar high-intensity areas on T2-weighted images | +few
    cerebellar high-intensity areas on FLAIR images | +few
    diffuse edema | +few
    mass effect on the fourth ventricle | +few
    mass effect on the brainstem | +few
    tonsillar herniation | +few
    supratentorial hydrocephalus | +few
    no bleeding on T2* sequence | +few
    no diffusion restriction | +few
    leptomeningeal enhancement along the cerebellar folia | +few
    Magnetic Resonance Spectroscopy | +few
    reduced level of N acetyl aspartate (NAA)/Creatine | +few
    normal Choline/Creatine ratios | +few
    doublet of lactate-lipid peak (1.3 ppm) | +few
    hemoglobin concentration 12.7 g/dL | 0
    white blood cell count 14280/mm3 | 0
    85% neutrophils | 0
    9% lymphocytes | 0
    4.8% monocytes | 0
    platelet count | 0
    erythrocyte sedimentation rate 20 mm/h | 0
    C-reactive protein level above 2 mg/L | 0
    lumbar puncture not performed | 0
    serological tests for Epstein Barr virus | 0
    serological tests for human herpes virus | 0
    serological tests for human immunodeficiency virus | 0
    serological tests for rubella virus | 0
    serological tests for parvovirus B19 | 0
    serological tests for measles virus | 0
    serological tests for Mycoplasma pneumoniae | 0
    serological test for mumps virus positive with IgM and IgG | 0
    control serology done 10 d later | +240
    IgG positive in control serology | +240
    post-infectious acute hemicerebellitis diagnosis | +few
    treated with mannitol | +few
    treated with corticosteroid | +few
    IV methylprednisolone 30 mg/kg per day for 3 d | +few
    oral prednisone 1 mg/kg per day tapered within 1 mo | +few
    discharge | +432
    brain MRI 18 days after discharge | +432+432
    partial resolution of signal alterations in the cerebellar hemispheres | +432+432
    brain MRI performed 3 mo later | +432+432+2160
    complete resolution | +432+432+2160
    final diagnosis: post-infectious acute hemicerebellitis | +few
    treatment with mannitol | +few
    treatment with corticosteroid | +few
    pseudotumoral cerebellitis diagnosis | +few
    risk of cerebellar herniation | 0
    no shortness of breath | 0
    denies chest pain | 0
    normal vital signs | 0
    negative serological tests except mumps | 0
    no history of neurological disorders | 0
    normal psychomotor development | 0
    stable vital signs initially | 0
    no bleeding | +few
    no diffusion restriction | +few
    benign mumps infection | -240
    mumps virus positive serology | 0
    pseudotumoral cerebellitis secondary to mumps infection | +few
    severe headache resolved | +432
    nausea resolved | +432
    vomiting resolved | +432
    trunk ataxia resolved | +432
    gait ataxia resolved | +432
    bilateral dysmetria resolved | +432
    dysautonomic troubles resolved | +432
    heart rate normalized | +432
    arterial pressure normalized | +432
    corticosteroid therapy completed | +432+720
    mannitol therapy completed | +432+720
    MRI follow-up | +432+432
    MRI follow-up complete resolution | +432+432+2160
    neurological symptoms resolved | +432+432
    hydrocephalus resolved | +432+432
    mass effect resolved | +432+432
    edema resolved | +432+432
    leptomeningeal enhancement resolved | +432+432
    tonsillar herniation resolved | +432+432
    supratentorial hydrocephalus resolved | +432+432
    normal neurological examination at discharge | +432
    improved consciousness level | +432
    Glasgow Coma Scale normalized | +432
    no recurrence of symptoms | +432+432+2160
    full recovery | +432+432+2160
    