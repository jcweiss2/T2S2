32 years old | 0
male | 0
admitted to the Emergency Department | 0
tonic-clonic seizures | 0
hypothyroidism | -168
morbid type 3 obesity | -168
gastritis with a gastric ulcer | -168
penicillin allergies | -168
endoscopic procedure | -168
erosive gastropathy | -168
admitted to the Intensive Care Unit (ICU) | 0
hypoxemia | 0
endotracheal tube placement | 0
invasive mechanical ventilation | 0
sedation with midazolam | 0
analgesia with fentanyl | 0
laboratory test results | 0
chest X-ray showed a right basal atelectatic band | 0
computed tomography (CT) scan of the chest showed bilateral basal condensation areas | 0
brain CT scan showed a normal brain | 0
rational antibiotic therapy with piperacillin plus tazobactam and clindamycin | 0
sputum, blood, and urine samples for cultures | 0
sedated with midazolam | 24
sedated with fentanyl | 24
bronchoscopy | 48
reddened mucosa with a cavity | 48
hemorrhagic stitches | 48
active bleeding | 48
bronchioalveolar lavage analysis | 48
MRSA (1×105 colony-forming unit [CFU]/mL) | 48
mecA and luk-PV gene-resistance mechanisms | 48
piperacillin plus tazobactam suspended | 48
intravenous vancomycin | 48
cerebrospinal fluid obtained by lumbar puncture | 0
no bacterial growth | 0
significant clinical improvement | 72
weaning of sedation | 72
weaning of invasive mechanical ventilation | 72
extubated | 72
good ventilatory mechanics | 72
99% saturation | 72
retained oxygen support with a mask | 72
respiratory rate of 19 breaths/min | 72
oriented to time, space, and person | 72
Glasgow Coma Scale score of 15/15 | 72
reactive isochoric pupils | 72
afebrile | 96
awake | 96
breathing ambient air | 96
discharged from the ICU | 144
hospitalized | 144
followed up through the Outpatient Department | 240
in general good health | 4320