31 years old | 0
female | 0
non-smoking | 0
Caucasian | 0
no past medical history | 0
sudden-onset severe headache | -840
left arm numbness | -840
cranial computed tomography (CT) scan | -840
grade 2 (Hunt and Hess scale) SAH | -840
admitted to the neurosurgical ward | 0
digital subtraction angiography (DSA) | 0
ruptured right middle cerebral artery aneurysm | 0
percutaneous endovascular coil embolization | 0
fever | -672
chills | -672
constant abdominal pain | -672
purulent uterine discharge | -672
admitted to the hospital | -672
suspected postpartum endometritis | -672
piperacillin/tazobactam | -672
vancomycin | -672
azithromycin | -672
sepsis | -640
septic shock | -640
transferred to the intensive care unit | -640
body temperature 38.3 °C | -640
invasive blood pressure 90/65 mmHg | -640
heart rate 135/min | -640
arterial oxygen saturation 82 % | -640
mild disorientation | -640
slower capillary refill | -640
coarse rales | -640
sequential organ failure assessment (SOFA) score 4 | -640
hemoglobin 6.8 g/dL | -640
d-dimers 4.58 μg/mL | -640
C-reactive protein 322 mg/L | -640
fibrinogen concentration 6.4 mL | -640
blood culture showed E. coli | -640
chest radiography | -640
pulmonary nodules | -640
CT of the thorax | -640
transvaginal ultrasound | -640
enlarged uterus | -640
complete loss of zonal anatomy | -640
abdominal magnetic resonance imaging (MRI) | -640
enlarged heterogenous myometrial mass | -640
splenic metastatic lesion | -640
serum β-human chorionic gonadotrophin (β-hCG) 232,085 mUI/mL | -640
suction evacuation and curettage | -640
pathology report confirmed choriocarcinoma diagnosis | -640
International Federation of Gynecology and Obstetrics (FIGO) modified WHO prognostic scoring system | -640
total score of 12 | -640
high risk of developing resistance to single-drug chemotherapy | -640
multiagent chemotherapy regimen | 0
low-dose etoposide | 0
cisplatin | 0
EMA/CO regimen | 0
etoposide | 0
methotrexate | 0
actinomycin D | 0
cyclophosphamide | 0
vincristine | 0
six cycles of EMA/CO | 0
β-hCG levels plateaued above normal | 168
restaging with MRI of the brain | 168
18F-fluorodeoxyglucose (FDG) positron emission tomography (PET)/CT scan | 168
decreased pulmonary nodules | 168
decreased uterine mass | 168
low standardized uptake value (SUV) of <3.8 | 168
revised FIGO score 7 | 168
EP/EMA regimen | 168
normalization of β-hCG | 336
grade 3 neutropenia | 168
granulocyte colony stimulating factor (G-SCF) | 168
dose reduction of both etoposide and actinomycin D | 168
grade 2 alopecia | 168
grade 2 nausea | 168
dexamethasone | 168
ondansetron | 168
grade 2 fatigue | 336
male condoms | 0
follow-up | 0
alive 21 months post diagnosis | 1008