77 years old | 0
    male | 0
    admitted to the hospital | 0
    abrupt onset of impaired consciousness | 0
    hypotension | 0
    intermittent mild lower abdominal discomfort | -120
    small amount of bloody, loose stools | -120
    occurring two to four times per day | -120
    for 5 days prior to admission | -120
    prostate cancer | -17544
    complete remission | -17544
    hypertension | -17544
    hyperlipidemia | -17544
    hyperuricemia | -17544
    lumbar spinal stenosis | -17544
    cold limbs | 0
    moist limbs | 0
    body temperature 35.6°C | 0
    pulse rate 42 bpm | 0
    blood pressure 65/36 mmHg | 0
    respiration rate 28 breaths/min | 0
    oxygen saturation 95% | 0
    mild abdominal distension | 0
    normal bowel sounds | 0
    normal white blood cell count | 0
    neutrophils 49.9% | 0
    normal platelet count | 0
    hemoglobin within normal range | 0
    C-reactive protein within normal range | 0
    procalcitonin within normal range | 0
    liver function tests within normal range | 0
    clotting screen within normal range | 0
    arterial blood gases within normal range | 0
    serum creatinine elevated | 0
    lactic acid elevated | 0
    hemoglobin A1c slightly elevated | 0
    no abnormalities on echocardiography | 0
    no abnormalities on abdominal ultrasound | 0
    mild edematous swelling of the small-intestinal wall | 0
    no marked free air | 0
    no ascites | 0
    septic shock | 0
    suspected complicating intra-abdominal infection | 0
    intravenous crystalloid solution administered | 0
    noradrenaline administered | 0
    meropenem initiated | 0
    state of consciousness improved | 72
    vital signs normalized | 72
    body temperature spike to 38.5°C | 72
    blood culture positive for C. paraputrificum | 0
    gram-positive bacillus with terminal spores | 0
    intravenous ampicillin/sulbactam initiated | 72
    treated for 10 days | 72
    laboratory parameters improved | 96
    clinical conditions improved | 96
    discharged from ICU | 96
    frequent loose, small amounts of bloody stools | 96
    low-grade fever | 96
    mild anemia | 96
    Clostridium difficile toxins A and B negative | 96
    glutamate dehydrogenase antigen negative | 96
    stools negative for ova | 96
    stools negative for parasites | 96
    stools negative for culture | 96
    diffuse mucosal inflammation on sigmoidoscopy | 840
    loss of vascular markings | 840
    engorgement of the mucosa | 840
    exudates | 840
    edema | 840
    touch friability | 840
    spontaneous bleeding in the rectum | 840
    crypt disarray | 840
    no signs of crypt abscesses | 840
    epithelial cell abnormalities | 840
    mucin depletion | 840
    neutrophil invasion | 840
    increased lamina propria cellularity | 840
    basal plasmacytosis | 840
    lamina propria eosinophils | 840
    ulcerative colitis | 840
    oral probiotics administered | 840
    intravenous intestinal prokinetic medications administered | 840
    abdominal manifestations persisted | 840
    dilated colon >12 cm in diameter | 1488
    colonic dilatation with no sign of thromboses | 1488
    no mechanical obstruction | 1488
    acute colonic pseudo-obstruction | 1488
    total parenteral nutrition initiated | 1488
    pharmacologic therapy initiated | 1488
    endoscopic decompression therapy initiated | 1488
    treatments unsuccessful | 1488
    dilated colon resected | 2256
    acute colonic pseudo-obstruction in ulcerative colitis | 2256
