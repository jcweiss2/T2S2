2.5 years old | 0  
    male | 0  
    Pearson syndrome | 0  
    Pearson syndrome | 0  
    marrow failure | 0  
    pancytopenia | 0  
    pancreatic insufficiency | 0  
    daily filgrastim therapy (G-CSF) for 2 years before presentation | -17520  
    bone marrow aspirate 2 months before presentation | -1440  
    modest number of blast cells | -1440  
    testing of 20 cells showed 19 had 45 chromosomes, including X and Y, but lacked chromosome 7 (monosomy 7) | -1440  
    scraped left first toe on tricycle 2 weeks before presentation | -336  
    small, erythematous, scabbed lesion on medial aspect of the toe | -336  
    treated with oral clindamycin | -336  
    progressive swelling | 0  
    progressive erythema | 0  
    hospitalization | 0  
    intravenous vancomycin | 0  
    absolute neutrophil count 6895 | 0  
    did not improve over next 2 days | 48  
    cefepime added | 48  
    MRI demonstrated osteomyelitis of distal half of left first metatarsal | 48  
    concern for sepsis of first metatarso-pharyngeal joint | 48  
    voriconazole added | 48  
    ambisome added | 48  
    Orthopedics consulted | 48  
    aspiration of first metatarsal performed | 48  
    serosanguinous fluid obtained | 48  
    fluid culture grew Fusarium species | 48  
    suppurative arthritis | 48  
    proven invasive fungal disease | 48  
    voriconazole continued | 48  
    ambisome continued | 48  
    toe appeared less erythematous after 2 days of treatment | 96  
    severe hypotension | 96  
    transfer to pediatric intensive care unit | 96  
    restoration of perfusion with intravenous fluids | 96  
    restoration of perfusion with dobutamine | 96  
    blood cultures negative for bacteria | 96  
    blood cultures negative for fungi | 96  
    computed tomography scan of chest, abdomen, and pelvis showed no evidence of fungal dissemination | 96  
    patient stabilized | 96  
    edema of foot did not improve | 96  
    erythema of foot did not improve | 96  
    edema and erythema waxing and waning in intensity | 96  
    biopsy of first metatarsal performed | 96  
    washout of joint performed | 96  
    culture negative for fusarium | 96  
    pathology report confirmed presence of fungal elements with appearance of fusarium in bone tissue fragments | 96  
    initial fusarium isolate MIC 16 to voriconazole | 96  
    initial fusarium isolate MIC >16 for posaconazole | 96  
    initial fusarium isolate MIC >16 for itraconazole | 96  
    initial fusarium isolate MIC 2 mcg/mL to amphotericin B | 96  
    voriconazole discontinued | 96  
    amphotericin B continued | 96  
    caspofungin added | 96  
    regimen continued for 3 weeks | 624  
    minimal clinical improvement | 624  
    repeat MRI demonstrated progression of bone destruction | 624  
    repeat MRI demonstrated joint space widening | 624  
    need for eradication of osteomyelitis before bone marrow transplant | 624  
    concern for imminent transformation of monosomy 7 into frank monocytic leukemia | 624  
    partial foot amputation performed 5 weeks after initial presentation | 840  
    Gomori methenamine silver stain positive for fungal hyphae and yeast-like structures compatible with Fusarium species | 840  
    Periodic acid-Schiff stain positive for fungal hyphae and yeast-like structures compatible with Fusarium species | 840  
    osteomyelitis with abscess formation around base of first toe involving phalangeal-metatarsal bones | 840  
    caspofungin discontinued 2 days after amputation | 888  
    amphotericin B discontinued 7 days after amputation | 1128  
    bone marrow transplantation successfully performed | 1128  
    no evidence of recurrent infection in lower extremity over ensuing 7 months | 1128  
    patient passed away after contracting viral respiratory illness | 1128  
    viral respiratory illness progressed to respiratory failure | 1128  
    viral respiratory illness progressed to renal failure | 1128  
    underlying metabolic disorder | 1128