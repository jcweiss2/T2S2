65 years old | 0
    male | 0
    chronic obstructive pulmonary disease | 0
    presented to the emergency department | 0
    weight loss | -6480
    lack of appetite | -6480
    generalized fatigue | -6480
    dehydrated | 0
    cachexic | 0
    fluid-responsive hemodynamics | 0
    heart rate 109 beats per minute | 0
    blood pressure 78/54 mm Hg | 0
    respiratory rate 17 per min | 0
    oxygen saturation 97% | 0
    received 3 L of crystalloids | 0
    blood pressure rose to 93/69 mm Hg | 0
    numerous ecchymoses | 0
    coarse crepitations | 0
    nontender splenomegaly | 0
    palpable periumbilical mass | 0
    anemia 62 g/L | 0
    thrombocytopenia 48 × 10^9/L | 0
    hypoglycemia 2.9 mmol/L | 0
    metabolic acidosis pH 7.22 | 0
    hyperlactatemia 18.8 mmol/L | 0
    admitted to high-dependency unit | 0
    received crystalloids | 0
    blood transfusion | 0
    broad-spectrum antibiotics | 0
    negative blood cultures | 0
    negative urine cultures | 0
    normal D-lactate level | 0
    cervical=mediastinal lymphadenopathy | 0
    nodular consolidative changes | 0
    mesenteric mass 3.9 cm × 1.8 cm | 0
    persistent hypoglycemia 2.5–3.9 mmol/L | 0
    no neuroglycopenic symptoms | 0
    mild hypothyroidism TSH 7.11 mIU/L | 0
    hypothyroidism fT4 7.3 pmol/L | 0
    required dextrose infusion | 0
    oral food intake | 0
    mesenteric mass inaccessible | 0
    bronchoscopy | 0
    gastrointestinal endoscopy | 0
    no malignant cells | 0
    bronchoalveolar lavage negative | 0
    bone marrow aspiration delayed | 0
    bone marrow biopsy delayed | 0
    CD20-positive non-Hodgkin's lymphoma | 264
    diffuse large B-cell lymphoma | 264
    CD10 overexpression | 264
    cyclin D1 overexpression | 264
    lactate levels climbed steadily | 456
    continued dextrose infusions | 456
    initiated prednisone 100 mg daily | 456
    encephalopathy | 432
    nosocomial pneumonia | 432
    sepsis | 432
    tumor lysis syndrome | 432
    multiorgan failure | 432
    transfer to intensive care unit | 432
    mechanical intubation | 432
    vasopressors | 432
    continuous renal replacement therapy | 432
    withdrawal of care | 456
    passed away | 456
    