33 years old | 0
male | 0
polysubstance abuse | -8760
saddle pulmonary embolus | -8760
abdominal pain | -8760
abdominal pain persisted | 0
nausea | 0
weight loss | -8760
methadone | -8760
Eliquis | -8760
pulmonary embolism | -8760
family history of pulmonary embolism | 0
family history of deep vein thrombosis | 0
tachycardia | 0
hypertension | 0
diaphoresis | 0
diffusely tender abdomen | 0
fullness in the epigastrium and upper quadrants | 0
elevated white blood cell count | 0
neutrophilic shift | 0
elevated lactate | 0
CT scan of abdomen and pelvis | 0
mesenteric distortion | 0
infiltration within the right mid abdomen | 0
partial small bowel obstruction | 0
exploratory laparotomy | 12
large mass with indurated mesentery | 12
areas of necrosis | 12
bowel folded upon itself like an accordion | 12
foreshortened and thickened mesentery | 12
adherent to the retroperitoneum | 12
small bowel resection | 12
ileocecal junction resection | 12
proximal ascending colon resection | 12
distal ileum anastomosed to the right colon | 12
postoperative fever | 24
fever workup | 24
discharged | 168
follow-up office appointment | 192
pathology report | 192
torsion of the ileum | 192
early ischemic changes | 192
mesenteric panniculitis | 192
genetic screening panel | 192
heterozygous for FV Leiden | 192
tumor markers | 192
flow cytometry results | 192
Chromogranin A | 192
anticoagulation treatment with apixaban | 192
medication adherence | 192