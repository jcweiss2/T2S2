72 years old | 0
immunocompetent | 0
male | 0
severe high fever | 0
gastrointestinal symptoms | 0
genitourinary symptoms | 0
acute prostatitis | 0
hospitalized | 0
gentamycin | 0
ampicillin-resistant K. pneumoniae isolated | 0
floaters in the right eye | 72
loss of vision | 72
intraocular inflammation | 72
topical therapy with cycloplegics | 72
corticosteroid eye drops | 72
endogenous endophthalmitis suspected | 120
best corrected visual acuity hand motion | 120
intraocular pressure 12 mmHg | 120
marked exudation in the anterior chamber | 120
poorly dilated, round pupil | 120
fibrin on the anterior lens capsule | 120
opaque fundus view | 120
left eye normal status | 120
right eye ultrasound hyper-reflective signal compatible with abscess or hemorrhage | 120
pars plana vitrectomy | 120
vitreous biopsy | 120
intravitreal injection of vancomycin | 120
intravitreal injection of ceftazidime | 120
retina moderately ischemic | 120
signs of vasculitis | 120
infiltrated retina temporal to the central fovea | 120
vitreous samples Gram staining | 120
microbiological cultures for bacteria and fungi | 120
K. pneumoniae growth | 120
inflammation slowly started to subside | 120
K. pneumoniae resistant to ampicillin | 120
K. pneumoniae sensitive to all other tested antibiotics | 120
targeted injection of ceftazidime intravitreally | 168
fever | 168
sepsis suspected | 168
transferred to infectious disease department | 168
examined daily by ophthalmologist | 168
re-deterioration of vision | 216
opacities in the vitreous | 216
retinal detachment temporal to the central fovea | 216
moderate cataract | 216
phacoemulsification | 216
in-the-bag intraocular lens implantation | 216
posterior capsulotomy | 216
pars plana vitrectomy | 216
vitreous cavity highly infiltrated with dense inflammatory cells and fibrin | 216
large retinal necrotic area of 4×5 optic disk diameters | 216
no laser photocoagulation | 216
no cryotherapy | 216
no holes identified intraoperatively | 216
long-lasting tamponading agent (silicone oil) chosen | 216
scar tissue developed in location of necrotic retina | 216
retina flat | 216
inflammation completely disappeared | 216
BCVA improved to 0.2 | 216
retina remained attached | 7200
silicone oil removed | 7200
laser photocoagulation around edges of retinal defects | 7200
visual function improved | 7200
optical coherence tomography scan showed regular foveal contour | 7200
final BCVA stabilized to 0.3 | 2160
