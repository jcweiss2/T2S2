Nijmegen breakage syndrome | 0
male | 0
29 years old | 0
admitted to the hospital | 0
dysphonia | 0
dyspnea | 0
15 kg weight loss | 0
recurrent fever | 0
coughing | -168
fever | -168
leg pain | -168
elevated lactate dehydrogenase | -168
elevated C-reactive protein | -168
elevated uric acid | -168
elevated d-dimer | -168
discharged | -168
elevated lactate dehydrogenase | 0
elevated uric acid | 0
elevated C-reactive protein | 0
cervical and supraclavicular lymphadenopathy | 0
left vocal cord paresis | 0
FDG uptake in masses | 0
FDG-positive cervical lymph node | 0
diffuse large B-cell lymphoma | 0
stage IVB DLBCL | 0
dexamethasone treatment | 0
Rituximab-CHOP regimen | 0
extended antibiotic and antifungal infection prophylaxis | 0
PEGylated granulocyte colony-stimulating factor | 0
complete remission | 144
follow-up | 216
follow-up | 432
follow-up | 648
follow-up | 864
biopsy | 876
chronic inflammation | 876
no signs of neoplasia | 876
diagnosed with NBS | -10440
diagnosed with stage IV nodular sclerosis cHL | -4320
treated with chemotherapy | -4320
complete remission | -2880
registered in the NBS Registry | -10440
selective IgG4 deficiency | -10440
fungal sepsis | -4320
liver failure | -4320
kidney failure | -4320
severe infectious complications | -4320
discharged | -2880
second complete remission | 0