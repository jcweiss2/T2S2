52 years old | 0
male | 0
body mass index 23.6 kg/m2 | 0
no comorbidities | 0
admitted to the hospital | 0
open modified Scopinaro procedure | -7200
weight 216 kg | -7200
BMI 57.4 kg/m2 | -7200
weight reganance | -1200
incisional hernia | -1200
bariatric revisional surgery | -1200
hernia repair | -1200
weight 170 kg | -1200
BMI 45.1 | -1200
gastric pouch leak | -1200
intra-abdominal collections | -1200
sepsis | -1200
conservative management | -1200
open abdomen | -1200
negative wound pressure therapy | -1200
parenteral nutrition | -1200
intravenous antibiotics | -1200
epithelized gastrocutaneous fistula | -600
controlled but persistent drainage | -600
proximal edge of planned ventral hernia | -600
upper endoscopy | -600
fistulous orifice | -600
vertical staple line | -600
esophagogastric junction | -600
extraluminal extravasation | -600
recurrent left subphrenic abscess | -600
endoscopic treatment | -600
argon plasma coagulation | -600
internal drainage | -600
external drainage | -600
clipping | -600
fibrin sealants | -600
e-vac therapy | -600
stenting | -600
multidisciplinary team discussion | 0
decision to proceed with innovative endoscopic technique | 0
placement of CSDO | 0
Occlutech muscular VSD occluder | 0
catheterization laboratory | 0
intravenous sedation | 0
topic anesthesia | 0
fistula cannulation | 0
biliary stent deployment system | 0
direct endoscopic guidance | 0
extraluminal leakage | 0
contrast injection | 0
Amplatz extra stiff guidewire | 0
fluoroscopy | 0
delivery system | 0
CSDO deployment | 0
endoscopic guidance | 0
fluoroscopic guidance | 0
no immediate adverse events | 0
contrast study | 0
no extravasation of contrast material | 0
restricted oral intake | 24
liquid diet | 24
regular diet | 288
pigtail drain | 0
accidental displacement of pigtail | 432
systemic signs of sepsis | 432
computed tomography | 432
fluoroscopy | 432
recurrence of abscess | 432
partial dislodgment of CSDO | 432
second attempt with oversized disc | 432
Occlutech Figulla Flex II UNI | 432
sealing of fistulous orifice | 432
upper endoscopy | 1296
contrast-enhanced CT scan | 1296
device engrafted | 1296
reduction of chronic abscess | 1296
no signs of fistula recurrence | 1296
pigtail removal | 1296
no drainage | 1296