59 years old | 0
male | 0
chronic hepatitis B viral infection | 0
cirrhosis | 0
well controlled hypertension |B0
liver mass found during transabdominal ultrasound screening program | 0
multiphase computed tomography scan | 0
single early hepatocellular carcinoma diagnosed | 0
non-tumorous portal vein thrombosis | 0
MELD score 18 | 0
living related liver transplant decision made | 0
extended right lobe graft from son | 0
son 26 years old male | 0
no underlying medical conditions in son | 0
compatible blood group | 0
no anatomical variation indicated from CTA and MRCP | 0
no post-operative complications | 0
right hepatic vein reconstructed with triangular shape technique | 0
middle hepatic vein reconstructed with triangular shape technique | 0
total hepatectomy performed | 0
portal vein thromboendovenectomy done | 0
right lobe graft anastomosed to inferior vena cava with polypropylene 5/0 continuous technique | 0
right lobe graft anastomosed to portal vein with polypropylene 6/0 continuous technique | 0
doppler ultrasound of portal vein did not show good inflow | 0
intra-operative portal vein anastomosis balloon dilatation | 0
stent placement through inferior mesenteric vein | 0
right hepatic artery anastomosed to common hepatic artery proper using polypropylene 8/0 interrupted technique | 0
