19 years old | 0
male | 0
admitted to the hospital | 0
fever | -48
malaise | -48
headache | -48
vomiting | -48
near-syncope | -48
confusion | 0
maculopapular rash | 0
tender nodule in the left armpit | -48
elevated white count | 0
elevated neutrophils | 0
elevated procalcitonin | 0
elevated lactic acid | 0
normal breath sounds | 0
no lymphadenopathy | 0
started on ceftriaxone and doxycycline | 0
lumbar puncture | 24
cerebrospinal fluid analysis | 24
transthoracic echocardiogram | 24
persistent hypotension | 48
tachycardia | 48
fever to 40 °C | 48
upper and lower extremities weakness | 48
transferred to ICU | 48
elevated liver enzymes | 48
elevated creatinine kinase | 48
elevated troponin | 48
elevated D-dimer | 48
elevated C-reactive protein | 48
elevated erythrocyte sedimentation rate | 48
elevated interleukin-6 | 48
elevated fibrinogen | 48
repeat SAR-CoV-2 RT-PCR | 48
started on IV vancomycin | 96
white count started trending down | 96
lactic acid started trending down | 96
fever decreased | 96
vitals became stable | 96
discharged from ICU | 96
left armpit pain | 96
nodule evolved into an abscess | 96
flushed | 96
nonspecific erythrasma on the lower limbs | 96
deep palmar erythema | 96
incision and drainage of the abscess | 120
abscess culture | 120
rashes started to have central clearance | 120
flaky skin | 120
discharged from hospital | 168
diffuse erythroderma nearly resolved | 168
flakiness in the palms | 168
pinkish coloration in the palms | 168
cultures from the wound showed methicillin-susceptible Staphylococcus aureus | 168
diagnosis of staphylococcal TSS | 168
started on oral amoxicillin-clavulanate | 168