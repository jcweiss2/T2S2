60 years old | 0
female | 0
height: 157 cm | 0
body weight: 45.9 kg | 0
diagnosed with hepatitis B virus-induced liver cirrhosis | -2190
diagnosed with hepatocellular carcinoma | -2190
treated with trans-arterial chemoembolization | -2190
treated with palliative radiotherapy | -2190
used an albuterol inhaler | -8760
umbilical hernia repair | -8760
total thyroidectomy | -7300
papillary thyroid carcinoma | -7300
taking an antiviral agent | -2190
taking warfarin | -2190
taking diuretics | -2190
hospitalization | -168
medication | -168
ascites was refractory | -168
laboratory values had improved slightly | -168
liver cirrhosis progressed | -168
HCC was unresectable | -168
LT was planned | -168
preoperative hematocrit was 0.283% | -24
preoperative hemoglobin was 9.2 g/dl | -24
preoperative platelet count was 63000 /μl | -24
preoperative prothrombin time with an international normalized ratio was 1.17 | -24
preoperative sodium was 133 mmol/L | -24
preoperative model for end-stage liver disease score was 15 points | -24
vital signs were within the normal range | -24
preoperative chest radiography confirmed no active lung lesion | -24
preoperative diaphragm was elevated toward the left side | -24
pulmonary function test showed a combined severe obstructive and moderate restrictive pattern | -24
transthoracic echocardiography showed diastolic dysfunction grade 1 | -24
esophagogastroduodenoscopy revealed esophageal varices | -24
esophagogastroduodenoscopy revealed portal hypertensive gastropathy | -24
esophagogastroduodenoscopy revealed gastric varices at cardia | -24
son was willing to donate his liver | -168
son's blood type was AB | -168
patient's blood type was A | -168
received a single intravenous dose of rituximab | -336
isoagglutinin immunoglobulin M and G titers against B antigen were measured | -336
plasmapheresis was performed | -336
target isoagglutinin titer was less than 1 : 16 | -336
13 units of AB type fresh frozen plasma were used for each plasmapheresis | -336
LT was scheduled | -48
RBC antibody screen was negative | -24
electrocardiography was conducted | 0
pulse oximetry was conducted | 0
non-invasive blood pressure was conducted | 0
two puffs of albuterol were administered | 0
anesthesia was induced | 0
intubation was performed | 0
radial artery cannulation was performed | 0
bispectral index monitoring was started | 0
hospital blood bank informed that her RBC antibody screen test had been positive | 0
RBC antibody screen test was positive | -48
pack of single-donor platelets had been transfused | -1096
pack of single-donor platelets had been transfused | -730
anti-C and anti-M were identified | -730
induction was postponed | 3
four more units of packed RBCs were received | 3
cross-matched | 3
two 20 G catheters were inserted | 3
7 French central catheter was placed | 3
magnetic induction fluid warmer was connected | 3
FloTrac/Vigileo system monitoring started | 3
IVC reconstruction was performed | 3
re-perfused | 3
methylprednisolone was infused | 3
basiliximab was infused | 3
bleeding around the hepatic artery was controlled | 3
diaphragm was repaired | 3
two chest tubes were inserted | 3
patient was transferred to the surgical intensive care unit | 3
wound was closed | 48
wedge biopsy of the transplanted liver was conducted | 48
centrilobular hemorrhagic necrosis of hepatocytes was found | 48
stricture of the hepatic vein was found | 48
tracheostomy was applied | 168
IgM and IgG antibodies gradually increased | 168
re-transplantation was planned | 744
patient expired due to sepsis | 744