75 years old | 0
woman | 0
admitted to the Emergency Department | 0
mildly itching skin rash | -48
fever | -48
shivering | -48
weakness | -48
rash initially noticed on the torso | -48
rash spread to the extremities | -48
self-medication with cetirizine | -48
no signs of respiratory disorders | 0
no signs of gastrointestinal disorders | 0
SARS-CoV-2 polymerase chain reaction test negative | 0
chest X-ray no signs of pulmonary infiltrates | 0
allopurinol prescribed for hyperuricemia | -504
long-term antihypertensive drugs (amlodipine, valsartan) | -504
maculopapulous exanthema covering the whole body | 0
prominent on the back, abdomen, and between the breasts | 0
no oral lesions | 0
skin lesions caused by viral infection | 0
adverse drug reaction induced by allopurinol considered | 0
allopurinol discontinued | 0
oral prednisolone (0.9 mg/kg/d for 2 days) | 0
cetirizine (10 mg/d) | 0
treatment on outpatient basis | 0
patient declined hospitalization | 0
worsening exanthema | 48
hospital admission | 48
maculopapulous exanthema as widespread blistering and skin peeling | 48
oral involvement | 48
mucosal ulceration | 48
erythema of the conjunctiva | 48
fulminant progression | 48
diagnosis of TEN | 48
prednisolone intravenously (3.7 mg/kg/d for 3 days) | 48
cyclosporine (5 mg/kg/d for 10 days) | 48
skin biopsy showed typical signs of TEN | 48
transferred to ICU | 48
daily multidisciplinary supportive team review | 48
SCORTEN assessed on admission | 48
initial SCORTEN predicted 90% mortality | 48
fluid replacement adjusted daily | 48
large blisters decompressed | 48
warm sterile lotions of polyhexanide and octenidine | 48
nonadhesive gauze, antiseptic gel, and sterile compresses | 48
metalline foil used | 48
oral lesions rinsed with saline and antiseptic lotions | 48
intense pain | 48
patient-controlled analgesia | 48
enteral nutrition by nasogastric feeding | 48
prophylactic anticoagulation | 48
bacteriuria treated by antibiotics | 48
ophthalmologic consultations confirmed recovery | 48
gynecological consultations revealed labia minora and introitus necrolysis | 48
no other organ involvement | 48
regression of renal failure | 48
regression of inflammatory markers | 48
transferred to Dermatology Department | 168
recovered completely | 1008
discharged | 1008
adverse drug reaction documented | 1008
communicated to general practitioner | 1008
