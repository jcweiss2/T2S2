41 years old | 0
Caucasian | 0
woman | 0
presented to a regional tertiary hospital | 0
intermittent headaches | -1344
dizziness | -1344
visual disturbance | -1344
headaches localized around the occipital cortex | -1344
gradual onset | -1344
worsening over two weeks | -1344
associated with dizziness | -1344
visual blurriness | -1344
morning emesis | -1344
unintentional weight loss of 10 kg | -1344
Carbamazepine 400 mg twice a day | -1344
epilepsy | -1344
no recent history of seizure relapse | -1344
no history of HIV | -1344
no history of Tuberculosis | -1344
no exposure to pigeons | -1344
no immunosuppressive treatments | -1344
blood tests | 0
biochemical tests | 0
brain computed tomography scan | 0
unremarkable tests | 0
provisional diagnosis of occipital neuralgia | 0
oral Pregabalin 50 mg twice daily | 0
discharged | 0
referral for outpatient Magnetic Resonance Imaging scan | 0
outpatient neurologist review appointment | 0
re-presented | 504
re-admitted | 504
worsening headache | 504
nausea | 504
vomiting | 504
bilateral double vision on lateral gaze | 504
dry cough | 504
shortness of breath | 504
bilateral abducens nerve palsy | 504
chest radiograph showed right middle lobe consolidation | 504
treated for community acquired pneumonia | 504
intravenous ceftriaxone 1 g | 504
doxycycline 100 mg orally | 504
CRP of 46 mg/L | 504
inpatient MRI scan | 504
neurological opinion requested | 504
MRI brain scan showed small meningioma in right frontal cortex | 504
evidence of meningitis | 504
lumbar puncture | 504
high opening pressure (>34 cm H2O) | 504
high protein (1100 mg/L) | 504
low glucose (14 mmol/L) | 504
high white cell count (220 × 106/L) | 504
83% mononuclear cells | 504
positive cryptococcal titer of 1:1024 | 504
cerebrospinal fluid culture showed growth of C. neoformans | 504
commenced on daily IV amphotericin B (AmBisome liposomal 50 mg) | 504
oral 5-fluorocytosine 1500 mg 6-hourly | 504
induction therapy | 504
fluconazole 600 mg daily | 504
chest CT scan showed possible large cryptoccoma | 504
confirmed with bronchoscopy | 504
bronchial lavage | 504
lumbar percutaneous drainage due to high intracranial pressure | 504
percutaneous drainage site infected by MRSA | 504
negative for MRSA colonization previously | 504
treated as hospital acquired infection | 504
removal of the drain | 504
IV vancomycin 1 g twice a day | 504
rifampicin 300 mg daily | 504
initial presenting symptoms began to improve | 504
CSF cryptococcal clearance by week three | 504
transferred to rehabilitation ward | 504
oral Fluconazole 400 mg daily | 504
external ventricular drain inserted | 504
continued deterioration | 504
persistent headaches | 504
visual impairment | 504
ongoing high output EVD | 504
insertion of ventriculoperitoneal shunt | 504
week seven | 1176
fever (38.2°C) | 1176
worsening vision | 1176
confusion | 1176
non-localized headache | 1176
septic screen unremarkable | 1176
repeated CSF analysis | 1176
normal open pressure | 1176
increased protein (4300 mg/L) | 1176
raised white cell count (191 × 106/L) | 1176
repeated MRI brain revealed gyro hyper-intensity on FLAIR | 1176
intensive treatment with IV cefepime 2 g | 1176
IV vancomycin 1 g every 12 hours | 1176
level of consciousness deteriorated | 1176
admitted to ICU | 1176
endotracheal intubation | 1176
monitoring for 48 hours | 1176
CSF culture negative | 1176
IRIS suspected | 1176
high dose IV steroids | 1176
oral prednisolone | 1176
patient improved within next week | 1176
returned to ward | 1176
vision severely impaired | 1176
two visual evoked potential tests | 1176
no abnormal results | 1176
normal baseline visual examination | 1176
ophthalmology review during week ten | 1680
bilateral optic neuropathy confirmed | 1680
declared legally blind | 1680
tested negative for Hepatitis B | 1680
tested negative for HIV | 1680
positive hepatitis C antibodies | 1680
evidence of past infection (IgG) | 1680
normal immunoglobulin levels (IgG, IgA, IgM) | 1680
normal complement levels | 1680
