48 years old | 0
female | 0
admitted to the hospital | 0
sleeve gastrectomy | -480
wound evisceration | -384
reoperated | -384
intravenous cefazolin | -384
systemic hypertension | 0
type 2 diabetes mellitus | 0
chronic obstructive pulmonary disease | 0
sleep apnea syndrome | 0
recurrent fever | -192
blood cultures negative | -192
urine cultures negative | -192
rectal swab cultures negative | -192
Klebsiella pneumonia in catheter tip cultures | -192
Acinetobacter baumannii in catheter tip cultures | -192
intravenous colistin | -192
no clinical improvement | -96
meropenem | -96
blurred vision in the right eye | -72
visual acuity of light perception in the right eye | 0
visual acuity 0.00 logMAR in the left eye | 0
anterior segment examination normal | 0
light reaction normal | 0
vitreous clear | 0
central hemorrhagic hypopigmented lesion in the right fovea | 0
small hypopigmented lesions in both peripheral retinas | 0
hyperreflective vitreous dots on SD-OCT | 0
elevated subfoveal lesion on SD-OCT | 0
early hypofluorescence and late phase leakage on FA | 0
fungal chorioretinitis suspected | 0
intravenous voriconazole | 0
loading dose of voriconazole | 0
maintenance dose of voriconazole | 48
improvement in ocular findings | 72
visual acuity counting fingers from 1 meter in the right eye | 168
decrease in retinal lesions | 168
no growth in final cultures | 240
IV voriconazole treatment for 10 days | 240
oral voriconazole for 4 weeks | 240
visual acuity 0.20 logMAR in the right eye at first-month control | 720
visual acuity 0.00 logMAR in the left eye at first-month control | 720
pigment changes in the right eye fovea | 720
disruption of retinal pigment epithelium layer on SD-OCT | 720
window defect on FA | 720