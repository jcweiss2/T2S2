23 years old | 0
male | 0
history of methicillin-resistant Staphylococcus aureus (MRSA) impetigo | -8760
right tibia fracture | -8760
intramedullary fixation (IMN) | -8760
interlocking screws removed | -744
skin irritation | -744
pain | -744
redness and swelling at the surgical site | -672
stitch abscess | -672
cultures from the surgical site were positive for MRSA | -672
oral antibiotic treatment | -672
fever | -216
right groin pain | -216
viral infection | -216
systemic fever | -168
myalgia | -168
difficult and painful ambulation | -168
right forearm cellulitis | -168
right sudden onset uveitis | -168
systemic rash | -168
right hip lymphadenopathy | -168
increased CRP | -168
elevated WBC count | -168
hepatic enzymes elevation | -168
lactic dehydrogenase (LDH) elevation | -168
creatine phosphokinase (CPK) elevation | -168
intravenous (IV) antibiotics | -168
deterioration of medical condition | -120
positron emission tomography-computed tomography (PET-CT) scan | -120
OIM abscess with systemic manifestations | -120
blood cultures were positive for MRSA bacteria | -120
hemodynamic deterioration | -120
fulminant MRSA sepsis | -120
admitted to the intensive care unit (ICU) | -120
ultrasound-guided drainage | -96
full-body CT scan | -72
enlargement of the abscesses diameter | -72
persistent fever | -72
elevated CRP level | -72
elevated WBC count | -72
surgical intervention | 0
combined approach of Smith-Peterson and modified Stoppa | 0
surgical planning | 0
CT scan findings | 0
comprehensive multidisciplinary discussion | 0
orthopaedic team consultation | 0
general anaesthesia with muscle relaxant | 0
surgical technique | 0
Stoppa approach | 0
Smith-Peterson approach | 0
improvement of general condition | 24
less frequent fever spikes | 24
decrease in CRP and WBC levels | 24
additional antibiotic treatment | 24
almost complete recovery | 144
normal ambulation without pain or functional limitations | 144
return to daily activities | 144