45 years old | 0
male | 0
hypertension | 0
admitted to the hospital | 0
COVID-19 | 0
ground-glass pattern on thoracic CT | 0
nasopharyngeal swab test positive for SARS-CoV-2 RNA | 0
oseltamivir | 0
hydroxychloroquine | 0
broad-spectrum antibiotics | 0
mechanical ventilation | 24
transferred to ICU | 24
endotracheal intubation | 24
favipiravir | 24
rehabilitation program (planned) | 24
ARDS | 24
complications | 24
bed positioning every 2 hours | 24
prone position 12-16 hours | 24
sepsis | 720
continued broad-spectrum antibiotics | 720
tracheostomy | 720
stayed in ICU for two months | 720
mechanical ventilation for 55 days | 720
transferred to ward | 2880
oxygen support needed | 2880
stayed in ward for eight days | 2880
rehabilitation program planned again | 2880
discharged | 3408
PMR outpatient clinic evaluation | 3408
one week later, visited outpatient clinic | 4368
walking disability | 4368
stiffness in hips, elbows, shoulders | 4368
unable to stand up and move comfortably | 4368
completely dependent on daily living activities | 4368
no red, warm, swollen joints | 4368
pain in elbows and hips | 4368
hard, fixed growth masses palpated in hips | 4368
ankylosis of elbows | 4368
decreased shoulder ROM | 4368
flexion deformity in hips | 4368
difficulty lying prone | 4368
normal ROM in other joints | 4368
muscle strength not evaluable in affected limbs | 4368
X-rays showed HO in hips, shoulders, elbows | 4368
increased ALP (291 IU/L) | 4368
normal serum calcium (9.3 mEq/L) | 4368
chronic sensory-motor polyneuropathy | 4368
cranial MRI showed mild cerebral atrophy | 4368
home-based rehabilitation program | 4368
stretching exercises | 4368
submaximal muscle strengthening exercises | 4368
pulmonary exercises | 4368
physiotherapist supervision | 4368
indomethacin 25 mg t.i.d. | 4368
follow-up ongoing | 4368
rehabilitation ongoing | 4368
