18 years old | 0
male | 0
farmer | 0
ingestion of two fresh tablets of Celphos (AlP) | -4
vomiting | -4
pain in the abdomen | -4
agitated | -4
anxious | -4
irritable | -4
pulse rate (PR) was not palpable | -4
blood pressure (BP) was not recordable | -4
heart rate (HR) was 110/minutes | -4
respiratory rate (RR) was 28/min | -4
oxygen saturation (SPO2) was 95% | -4
sinus tachycardia | -4
T wave inversion in lead 3 | -4
intravenous (IV) crystalloids | 0
IV magnesium sulphate 1 gm stat and 8 hourly | 0
IV calcium gluconate 8 hourly | 0
IV hydrocortisone 100 mg stat and 12 hourly | 0
IV dopamine | 0
noradrenaline | 0
immediate gastric lavage with potassium permanganate (KMnO4) | 0
activated charcoal was kept in the stomach, repeated 8 hourly | 0
arterial blood gas (ABG) analysis showed a metabolic acidosis | 0
metabolic acidosis correction was performed as per the protocol | 0
intubated | 0
shifted to an intensive care unit (ICU) | 0
BP was 60–80 mmHg (systolic) | 6
PR was 120/min | 6
RR was 20/min | 6
input/output was 3L/300 ml over the next 24 hours | 24
monomorphic ventricular tachycardia (VT) | 48
DC cardio-version of synchronised 150 J | 48
IV amiodarone 150 mg bolus and infusion continued till the next 48 hours | 48
cardiac bio-markers also raised | 48
normal sinus rhythm was maintained till discharge | 48
ABG showed a pH of 7.4 | 96
HCO3 of 18 mmol/L | 96
CO2 of 42 mmol/L | 96
BP was ranging from 70/50 mmHg to 90/60 mmHg | 96
blood urea was 100 mg/dl | 96
serum creatinine was 4.5 mg/dl | 96
urine output was 400 ml/24 hours | 96
AST/ALT was 80/90 IU/L | 96
ALP was 200 U/L | 96
S bilirubin was 2.5 mg/dl | 96
haemodialysis was performed | 120
haemodialysis was performed | 168
blood urea after haemodialysis was 70 mg/dl | 168
creatinine was 4.0 mg/dl | 168
urine output improved to around 1200 ml/24 hours | 168
extubated | 120
shifted to a step down unit (SDU) | 168
vitals were normal | 168
liver and kidney functions were improving | 168
normal by the 14th day | 168
cardiac arrhythmia (VT) | 48
septicemia | 120
aspiration pneumonitis | 120
electrolyte imbalance | 120
severe hypoxia | 120
gastro-intestinal bleeding | 120
refractory shock | 120
metabolic acidosis | 120
cardiovascular collapse | 48
ventricular tachycardia | 48
metabolic acidosis | 120
low bicarbonate | 120
low pH | 120