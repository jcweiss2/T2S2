60 years old | 0
female | 0
admitted to the hospital | 0
left flank pain | -48
radiating to the groin | -48
vomiting | -48
dizziness | -48
lightheadedness | -48
absence of urinary symptoms | -48
absence of fever | -48
coronary artery disease | -6720
prior angioplasty | -6720
type 2 diabetes mellitus | -6720
insulin glargine | -6720
insulin lispro | -6720
dulaglutide | -6720
empagliflozin | -336
hypertension | -6720
losartan | -6720
hypertriglyceridemia | -6720
icosapent ethyl | -6720
former smoker | -2520
family history for heart disease | -6720
family history for hypertension | -6720
family history for diabetes | -6720
family history for dyslipidemia | -6720
body mass index | 0
costovertebral tenderness | 0
tachycardia | 0
hypotension | 0
lactic acidosis | 0
leukocytosis | 0
left shift | 0
thrombocytopenia | 0
glycosylated hemoglobin A1C | -6720
kidney function compromised | 0
creatinine | 0
blood urea nitrogen | 0
liver function tests abnormal | 0
aspartate aminotransaminase | 0
alanine transaminase | 0
alkaline phosphatase | 0
total bilirubin | 0
serum glucose | 0
urine analysis | 0
glucose in urine | 0
bacteria in urine | 0
white blood cells in urine | 0
emphysematous pyelonephritis | 0
ischemic colitis | 0
portal venous gas | 0
air within branches of the superior mesenteric vein | 0
cefepime | 0
vancomycin | 0
metronidazole | 0
nephrectomy | 24
bowel viable | 24
postoperative management | 24
intensive care unit | 24
pan-susceptible Escherichia coli | 24
antibiotics de-escalated | 24
discharged home | 168
cefpodoxime | 168
empagliflozin discontinued | 168
near-syncope episode | 720
abdominal pain | 720
small bowel obstruction | 720
decompensated | 720
cardiopulmonary arrest | 720
massive emesis | 720
aspiration of gastric contents | 720
resuscitation | 720
ICU stay | 720
anoxic brain injury | 720
withdraw life support | 720
death | 720