59 years old | 0
male | 0
presented to the emergency department | 0
generalized weakness | -12
chest pain | -12
dyspnea | -12
back pain | -12
chronic obstructive pulmonary disease | 0
requiring 3 L nasal cannula oxygen at baseline | 0
coronary artery disease | 0
history of bypass surgery | -8760 (approximated as 1 year prior)
insulin dependent diabetes mellitus | 0
obstructive sleep apnea | 0
morbid obesity | 0
BMI 46.3 | 0
urinary retention | 0
managed with indwelling urinary catheter | 0
Do Not Resuscitate order | 0
prior hospitalization | -8760 (approximated as 1 year prior)
scrotal cystocele decompressed by indwelling urethral catheter | -8760
mild hydronephrosis | -8760
ureters inserting into the bladder cephalad to the symphysis pubis | -8760
tachycardia | 0
hypertensive | 0
increasing oxygen requirements | 0
significant leukocytosis | 0
acute renal insufficiency | 0
CT obtained | 0
distended bladder within the right hemiscrotum | 0
bladder trigone migrated outside of the pelvis | 0
ureters coursing anterior and distal to the pubic symphysis |;0
catheter removed | 0
sterile urinalysis obtained | 0
catheter could not be replaced | 0
became hypotensive | 12 (approximated 12 hours after admission)
transferred to the intensive care unit | 12
bedside ultrasound performed | 12
placed two holding sutures into the anterior scrotum | 12
tenting the bladder anteriorly | 12
placed a 14fr catheter using a Cook One Step Suprapubic Catheter Introducer | 12
stabilized in the ICU | 24 (approximated 24 hours after ICU transfer)
discharged | 120
follow up cystoscopy performed | 144 (approximated 24 hours after discharge)
catheter exchanges performed monthly | N/A (ongoing, no specific timestamp)
no symptomatic infections | N/A (ongoing, no specific timestamp)
scrotal cystocele managed with trans scrotal neocystotomy tube | 12
urosepsis from scrotal cystocele | 0
trans scrotal drainage via neocystotomy | 12
