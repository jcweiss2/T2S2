69 years old | 0
male | 0
Child–Pugh class C cirrhosis | 0
admitted to the Emergency department | 0
slipping on wet grass and falling on his left side | -1
Glasgow coma score 15/15 | 0
vital signs within normal limits | 0
pulse rate 78/min | 0
RR 13/min | 0
BP 113/54 mm Hg | 0
SpO2-100% in air | 0
left hip tenderness | 0
no ecchymosis to the abdomen, flank or thigh | 0
radiograph of his pelvis revealed an undisplaced fracture of his left acetabulum | 0
liver dysfunction | 0
pH 7.271 | 0
base excess minus 7.3 | 0
PT 18.2 | 0
INR-1.5 | 0
APTT ratio 1.42 | 0
platelets 73 | 0
bilirubin 63 mmol/l | 0
Hb 124 g/l | 0
18 g intravenous cannula inserted | 0
warmed Hartmanns one litre infusion commenced | 0
referred to the Orthopaedic on call team | 1
blood pressure dropped to 75/51 mm Hg | 1
tachycardic | 1
serum lactate 9 mmol/l | 1
FAST examination revealed intraabdominal fluid | 1
treated for sepsis | 1
intensive care, orthopaedic and general registrar attended the patient | 2
pH 7.227 | 2
base excess of −17.9 | 2
serum lactate of 16.3 mmol/l | 2
Hb 75 g/l | 2
arterial blood pressure 90/60 mm Hg | 2
pulse rate 90/min | 2
left lower abdominal quadrant and upper thigh swollen with ecchymosis | 2
diagnosis of haemorrhagic shock | 2
massive transfusion pathway activated | 2
four units of Blood transfused | 2
four units of FFP transfused | 2
two adult therapeutic doses of platelets transfused | 2
10 units of cryoprecipitate transfused | 2
noradrenaline infusion commenced | 2
pelvic binder in place | 2
CT scan | 4
CT abdomen confirmed the fracture of the left acetabulum | 4
significant haematoma on left pelvic sidewall adjacent to the fracture | 4
8 mm enhancing nodule suggestive of an internal iliac artery pseudoaneurysm | 4
ill-defined blush of contrast within the haematoma | 4
extra-peritoneal haematoma inseparable from the bladder | 4
cirrhotic liver | 4
6.7 cm infra-renal aortic aneurysm | 4
transferred to the intensive care unit | 4
invasive cardiovascular monitoring | 4
CT Angiogram | 48
no arterial bleed | 48
prophylactic embolization recommended | 48
gelfoam embolization of anterior and posterior division segmental branches of the left internal iliac artery | 48
10 lb skeletal traction applied | 48
discharged to the orthopaedic ward | 120
uncontrollable bleeding from his pin site | 120
skeletal traction removed | 120
continuous pressure applied to the wound | 120
died on 30 January 2017 | 1224
chronic liver disease | 1224