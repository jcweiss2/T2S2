66 years old | 0
male | 0
admitted to the hospital | 0
history of AF | -672
history of common atrial flutter | -672
radiofrequency pulmonary vein isolation procedure | 0
wide defragmentation of the left atrium | 0
creation of a posterior box | 0
sinus rhythm restored | 0
external electric shock | 0
general anesthesia | 0
3D intracardiac navigation | 0
transseptal approach | 0
transoesophageal echocardiography (TEE) | 0
fluoroscopic guidance | 0
oesophageal temperature monitored | 0
discharged from the hospital | 24
anticoagulant treatment | 0
proton pump inhibitors (PPI) | 0
dyspnoea at rest | 336
thoracic discomfort | 336
pericardial involvement | 336
rapid AF | 336
inflammation | 336
C-reactive protein (CRP) > 200 mg/L | 336
hyperleukocytosis | 336
hemodynamically stable | 336
poor tolerance of the arrhythmia | 336
bradycardia with beta-blockers | 336
digoxin | 336
cardioversion attempt with amiodarone | 336
abundant heterogeneous pericardial effusion | 336
circumferential pericardial effusion | 336
systolic–diastolic notch on the left atrium | 336
respiratory variation of the transvalvular flow | 336
cardiac tamponade | 336
pericardiocentesis | 336
cloudy, orange pericardial fluid | 336
purulent fluid | 336
pericardial drain | 336
hemodynamic failure | 336
hypotension | 336
fever | 336
acute respiratory failure | 336
signs of shock | 336
acute anuric renal failure | 336
hepatic failure | 336
hyperlactatemia | 336
severe acute right ventricular dysfunction | 336
broad-spectrum antibiotic treatment | 336
inotropic support with dobutamine | 336
multiphase thoracic–abdominal–pelvic CT scan | 336
minimal hydroaeric pericardial effusion | 336
discontinuity in the anterior oesophageal wall | 336
extraluminal contrast leakage | 336
oesophageal–pericardial fistula | 336
endoscopic management | 360
fistulous orifice | 360
covered oesophageal prosthesis | 360
fluoroscopic guidance | 360
rapid extubation | 384
weaning from amines | 384
altered neurological state | 432
Glasgow Coma Scale | 432
ischaemic strokes of gaseous origin | 432
diffuse intraparenchymal and subarachnoid air embolism | 432
migration of the oesophageal prosthesis | 432
air bubbles in the left ventricle and left auricle | 432
fistula between the esophagus and the right superior pulmonary vein | 432
brain MRI | 456
poor prognosis | 456
brain damage | 456
multiple ischaemic lesions | 456
gas emboli | 456
mesencephalic involvement | 456
diffuse supra-tentorial cerebral edema | 456
subfalcine herniation | 456
brain death | 480