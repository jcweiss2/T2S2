25 years old | 0
primiparous | 0
healthy | 0
uneventful pregnancy | -280
spontaneous labour | 0
normal vaginal delivery | 0
right medio-lateral episiotomy | 0
discharged home | 24
general weakness | 48
severe pain | 48
swelling at the episiotomy site | 48
tachycardia | 48
normal blood pressure | 48
ecchymosis | 48
induration | 48
severe tenderness | 48
no crepitus | 48
elevated white blood count | 48
elevated C-reactive protein | 48
intravenous fluids | 48
broad-spectrum antibiotics | 48
urgent exploration of the episiotomy site | 48
no obvious hematoma | 48
no pus collection | 48
viable tissues | 48
culture swabs collected | 48
surgical drain sited | 48
episiotomy wound edges approximated | 48
clinical picture deteriorated | 72
tachycardia | 72
hypotension | 72
transferred to intensive care unit | 72
further rise in CRP | 72
further rise in WBC | 72
pelvic CT scan | 72
bulky uterus | 72
pelvic ascites | 72
no evidence of tissue fluid or gas collection | 72
surgical consultation | 72
laparoscopy | 96
no evidence of uterine rupture | 96
no pelvic hematoma | 96
ascitic fluid drained | 96
culture swabs obtained | 96
perineal re-exploration | 96
unviable tissue | 96
extensive tissue debridement | 96
healthy viable tissues reached | 96
wound left open | 96
iodine-soaked pack applied | 96
antibiotics adjusted | 96
clinical condition improved | 120
repeated debridements | 120
V-Y advancement fascial flap | 168
wound closure | 168
discharged in good condition | 240
followed up in outpatient department | 240
recovered completely | 720
pregnant again | 720
regular antenatal care | 720
elective cesarean section | 752
Hailey-Hailey disease | -672
exacerbated by pregnancy | 48
exacerbated by trauma | 48
exacerbated by infection | 48
acantholysis | 96
dyskeratosis | 96
epidermal hyperplasia | 96
polymicrobial infection | 96
E. coli | 96
Enterococcus faecalis | 96
Bacteroides fragilis | 96