65 years old | 0
female | 0
diabetes | -7200
oral hypoglycemic agents | -7200
admitted to the hospital | 0
right flank pain | 0
fever | 0
blood pressure 80/50 mmHg | 0
temperature 39 °C | 0
pulse 130 beats/minute | 0
respiration rate 20 breaths/minute | 0
knocking tenderness on the right flank area | 0
WBC count 23,400/μL | 0
hemoglobin 9.7 g/dL | 0
platelet count 97,000/μL | 0
C-reactive protein 21.97 mg/dL | 0
blood urea nitrogen 35.3 mg/dL | 0
creatinine 2.21 mg/dL | 0
sodium 142 mEq/L | 0
potassium 3.7 mEq/L | 0
total protein 4.8 g/dL | 0
albumin 2.4 g/dL | 0
lactate dehydrogenase 472 U/L | 0
HbA1c 9.8% | 0
prothrombin time 17.5 seconds | 0
activated partial thromboplastin time 52.8 seconds | 0
antithrombin III 70.5% | 0
fibrin degradation products 49.2 μg/mL | 0
fibrinogen 429.3 mg/dL | 0
urinalysis specific gravity 1.028 | 0
urinalysis pH 5.0 | 0
urinalysis protein traces | 0
urinalysis WBCs 10-19 per high power field | 0
urinalysis RBCs 0-1 per high power field | 0
sinus tachycardia | 0
KUB nonspecific | 0
contrast-enhanced abdominal CT scan | 0
focal wedge-shaped perfusion defect in the upper pole of right kidney | 0
Escherichia coli isolated from blood and urine cultures | 0
intravenous ceftriaxone 2 g per day | 0
drowsy | 120
blood pressure 80/60 mmHg | 120
fever | 120
chest X-ray increased haziness on both lower lung fields | 120
WBC count 27,800/μL | 120
platelet count 26,000/μL | 120
creatinine 0.8 mg/dL | 120
chest CT scan | 120
passive atelectasis in both lungs | 120
no evidence of pneumonia | 120
echocardiography mildly decreased cardiac wall motion | 120
left ventricular dysfunction | 120
ejection fraction 47% | 120
no evidence of thrombus in all cardiac chambers | 120
diuretics and inotropes administered | 120
antibiotics changed to piperacillin sodium 4 g and tazobactam 0.5 g every 8 hours | 120
clinical course improved | 168
sudden onset of severe right flank pain | 312
tenderness | 312
urinalysis WBCs 1-4 per high power field | 312
urinalysis RBCs 5-9 per high power field | 312
lactate dehydrogenase 1768 U/L | 312
abdominal CT scan | 312
large perfusion defect in the upper to mid portion of the right kidney | 312
intravascular filling defect in the right renal artery | 312
prothrombin time 12.3 seconds | 312
activated partial thromboplastin time 23.8 seconds | 312
antithrombin III 84.7% | 312
fibrin degradation products 19.5 μg/mL | 312
fibrinogen >500 mg/dL | 312
factor assay V 81% | 312
proteins C and S normal | 312
lupus anticoagulant Ab not found | 312
flank pain resolved | 384
hematuria disappeared | 384
follow-up abdominal CT scan | 384
perfusion defect in the right kidney partially regressed | 384
size of right renal artery thrombus partially regressed | 384
discharged | 528