47 years old | 0
male | 0
primary school director | 0
goiter | 0
euthyroidism | 0
admitted to the hospital | 0
fever | -168
chills | -168
myalgias | -168
mucocutaneous jaundice | -96
yellowish diarrhea | -96
abdominal pain | -96
altered | 0
dehydrated | 0
conscious | 0
temperature 38°C | 0
blood pressure 90/70 mm Hg | 0
oxygen saturation 98% | 0
jaundice | 0
liver normal size | 0
spleen normal size | 0
white blood cells 29 000/mm3 | 0
neutrophils 91% | 0
hemoglobin 8.7 g/dL | 0
platelet counts 30 000/mm3 | 0
serum creatinine 76 mg/L | 0
urea 1.38 g/L | 0
alanine aminotransferase 140 IU/L | 0
aspartate aminotransferases 180 IU/L | 0
alkaline phosphatase 194 IU/L | 0
total bilirubin 425 mg/L | 0
prothrombin level 95% | 0
lumbar puncture | 0
clear cerebrospinal fluid | 0
cytochemical normal | 0
chest radiograph unremarkable | 0
abdominopelvic ultrasound | 0
normal-sized liver | 0
non-dilated bile ducts | 0
low abundance fluid effusion | 0
treated with ceftriaxone + ciprofloxacin + metronidazole + parenteral rehydration | 0
blood pressure 60/40 mm Hg | 72
hematemesis | 72
abdominal pain | 72
nausea | 72
tense and bloated abdomen | 72
depressible to palpation | 72
preserved transit | 72
null diuresis | 72
renal insufficiency | 72
urea 3.31 g/L | 72
creatinine 106 mg/L | 72
hyponatremia 115 mEq/L | 72
hemoglobin 6.7 g/dL | 72
procalcitonin 111 ng/mL | 72
creatine phosphokinase 833 IU/L | 72
lactate dehydrogenase 955 IU/L | 72
lipaemia 273 IU/L | 72
amylasemia 429 IU/L | 72
electrocardiography normal | 72
echocardiography normal | 72
abdominal CT angiography | 72
enlarged pancreas | 72
necrosis flow | 72
liquid digestive distension | 72
densification of the mesenteric fat | 72
intraperitoneal effusion | 72
transferred to medical resuscitation service | 72
noradrenaline | 72
vascular filling | 72
blood transfusions | 72
extrarenal purification sessions | 72
Inexium | 72
antibiotic therapy maintained | 72
gradual improvement | 120
diuresis initiated | 120
colors return | 120
kidney and liver tests correct | 408
blood cultures negative | 408
HBsAg negative | 408
anti-HAV IgM negative | 408
anti-HCV antibodies negative | 408
HIV serology negative | 408
SARS-CoV-2 viral RNA negative | 408
MAT serology positive | 408
Leptospira biflexa positive | 408
discharged | 408
follow-up | 480
no complication | 480