47 years old | 0
nulliparous | 0
female | 0
admitted to the hospital | 0
increasing abdominal girth | -336
fever | -48
no previous significant medical or surgical history | 0
nonsmoker | 0
stable relationship | 0
no history of sexually transmitted disease | 0
no intra-uterine copper device | 0
no previous gynecological problems | 0
temperature 38.5 C | 0
pulse 113 beats per minute | 0
blood pressure 76/46 mmHg | 0
pale | 0
clammy | 0
cachectic | 0
abdomen grossly distended | 0
abdomen tense | 0
large mass on the right side | 0
abdomen tender | 0
bowel sound not audible | 0
large umbilical hernia | 0
hemoglobin 7.8 g/dl | 0
WBC 21.7 | 0
CRP 205 | 0
clear lung fields on chest X-ray | 0
extensive intra-abdominal fluid on abdominal X-ray | 0
large ovarian mass on CT | 0
large ascites on CT | 0
left ureter obstructed | 0
malignant ovarian mass with superimposed infection | 0
started on cefuroxime | 0
started on Metronidazole | 0
laparotomy | 0
six liters of pus aspirated | 0
large cystic mass from right adnexa | 0
edematous tubes | 0
five liters of thick pus drained | 0
necrosis in cavity wall | 0
large uterus with multiple fibroids | 0
subtotal hysterectomy | 0
left ovary removed | 0
hernial sac excised | 0
hernia repaired | 0
no bowel perforation | 0
appendix normal | 0
abdominal washout with saline | 0
two drains inserted | 0
mass closure of abdomen | 0
estimated blood loss one liter | 0
admitted to intensive care | 0
ventilatory support | 0
inotropic cardiac support | 0
six units of blood transfusion | 24
tracheostomy | 48
pus culture grew Bacteroids fragilis | 24
no other bacteria grew | 24
antibiotics changed to Tazocine | 24
inflammatory markers rising | 24
became apyrexial | 24
remained on antibiotics for 10 days | 240
histology confirmed multiple fibroids | 240
right ovarian cyst wall showed marked inflammation | 240
endometriosis identified on ovary surface | 240
endometriotic cyst confirmed in left ovary | 240
started to improve | 96
CRP 33 | 96
discharged home | 336