71 years old | 0
female | 0
admitted to the hospital | 0
unconscious state | -24
stroke | -24
hypertension | -24
ischaemic heart disease | -24
peripheral vascular disease | -24
septic shock | -48
elevated erythrocyte sedimentation rate | -48
elevated C-reactive protein | -48
yeast in blood culture | -48
caspofungin | -48
died | 48
history of hypertension | -336
history of ischaemic heart disease | -336
history of peripheral vascular disease | -336
lower limb ischaemia | -336
hospitalized for lower limb ischaemia | -336
discharged | -336
Candida parapsilosis | -336
turquoise blue colonies on CHROMagar Candida | -336
identified as C. parapsilosis by VITEK 2 yeast identification system | -336
sequencing of ITS region of rDNA | -336
Lodderomyces elongisporus | -336
long ellipsoidal-shaped ascospores | -336
Internally transcribed spacer region of ribosomal DNA | -336
sequencing of ITS region of rDNA | -336
ascospores on acetate ascospore agar | -336
antifungal susceptibility | -336
MIC values | -336
amphotericin B | -336
0.012 | -336
fluconazole | -336
0.125 | -336
voriconazole | -336
0.004 | -336
posaconazole | -336
0.003 | -336
itraconazole | -336
0.008 | -336
flucytosine | -336
0.064 | -336
caspofungin | -336
0.064 | -336
micafungin | -336
0.003 | -336
unusual yeast in the absence of any known risk factors | -336
inoculation of the yeast from the skin or translocation from the gastrointestinal tract | -336
L. elongisporus is a recognized bloodstream pathogen | -336
little is known about its virulence attributes or its environmental niche | -336
global prevalence | -336
isolated from patients in distant geographic regions | -336
Mexico | -336
Malaysia | -336
China | -336
Australia | -336
Middle East | -336
Japan | -336
Spain | -336
Korea | -336
COPD | -336
ESRD | -336
endocarditis | -336
osteomyelitis | -336
brain embolic lesions | -336
intravenous drug user | -336
blue-green colonies on CHROMagar | -336
ITS region sequence analysis | -336
Candida metappsilosis | -336
C. orthopsilosis | -336
C. parapsilosis | -336
turquoise blue colonies on CHROMagar Candida | -336
identified as C. parapsilosis by VITEK 2 yeast identification system | -336
PCR sequencing of ITS region of rDNA | -336
L. elongisporus | -336
MALDI-TOF MS | -336
sequence analysis of ITS region and D1–D2 domains of rDNA | -336
trauma | -336
thoracoabdominal aortic replacement complicated with aortoesophageal fistula | -336
catheter | -336
dark green colonies Candida agar medium | -336
identified as C. parapsilosis by VITEK 2 system | -336
sequence analysis of ITS region and D1–D2 domains of rDNA | -336
COPD | -336
diabetes | -336
ESRD | -336
sequencing ITS region of rDNA | -336
turquoise blue colony on CHROMagar | -336
Candida medium | -336
VITEK 2 YST ID | -336
API 20C AUX | -336
MALDI-TOF MS | -336
score value | -336
1.79 | -336
lung cancer | -336
receiving immunosuppressive agents | -336
vascular catheter | -336
turquoise blue colony on CHROMagar | -336
identified as C. parapsilosis in VITEK 2 yeast identification system | -336
PCR sequencing of ITS region of rDNA | -336
hypertension | -336
ischaemic heart disease | -336
peripheral vascular disease | -336
caspofungin | -336
fluconazole | -336
voriconazole | -336
posaconazole | -336
itraconazole | -336
flucytosine | -336
caspofungin | -336
micafungin | -336
amphotericin B | -336
5-FC | -336
FL | -336
IT | -336
KE | -336
VO | -336
POS | -336
ISA | -336
CS | -336
AND | -336
MYC | -336
Lockhart 2008 | -336
BMD | -336
CLSI | -336
Tay 2009 | -336
Etest | -336
Daveson 2012 | -336
NA | -336
Hatanaka 2016 | -336
BMD | -336
CLSI | -336
Ahmad 2013 | -336
Etest | -336
Taj-Aldeen 2014 | -336
BMD | -336
CLSI | -336
Fernández-Ruiz 2017 | -336
BMD | -336
CLSI | -336
Lee 2018 | -336
ATB Fungus 3 | -336
uncommon yeast pathogens | -336
misidentified as a result of limitations of the currently available commercial yeast identification systems | -336
VITEK 2 | -336
C. parapsilosis complex | -336
C. parapsilosis | -336
C. orthopsilosis | -336
C. metapsilosis | -336
L. elongisporus | -336
multiplex PCR assay | -336
380 C. parapsilosis complex isolates | -336
retrospective characterization | -336
Mycology Reference Laboratory culture collection | -336
previously speciated by VITEK 2 | -336
three L. elongisporus isolates | -336
Kw2486/06 | -336
sputum of a cancer patient | -336
Kw554/08 | -336
catheter tip of a patient with fungaemia | -336
Kw3047/14 | -336
bloodstream of a cancer patient | -336
matrix-assisted laser desorption/ionization time-of-flight mass spectrometry | -336
identification of L. elongisporus | -336
rare yeast species | -336
exhibit reduced susceptibility to one or more commonly used antifungal agents | -336
prolonged survival of seriously ill patients | -336
intensive care units | -336
administration of multiple broad-spectrum antibiotics | -336
life support systems | -336
extended use of intravascular catheters | -336
selection pressure created by prophylactic and therapeutic use of antifungal agents | -336
colonization and invasive infection | -336
delay in accurate identification | -336
lack of experience in the management of such rare yeast infections | -336
higher mortality rates | -336