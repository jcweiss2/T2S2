53 years old | 0
female | 0
admitted to the hospital | 0
necrotizing fasciitis | 0
unconscious | 0
septic shock | 0
high temperature | 0
myalgia | 0
breathing difficulties | 0
respiratory failure | -672
mild hypertension | -672
obesity | -672
heavy smoker | -672
large necrotic area of skin and soft tissue | 0
purulent discharge | 0
palpable right axillary lymph nodes | 0
tachypneic | 0
heart rate of 115 bpm | 0
blood pressure of 80/50 mmHg | 0
leukocytosis | 0
increased erythrocyte sedimentation rate | 0
increased C-reactive protein | 0
low hemoglobin level | 0
increased serum creatine kinase | 0
resuscitated with intravenous fluids | 0
imaging of the breast, chest, and abdomen | 0
blood samples for blood culture | 0
treated with intravenous broad-spectrum antibiotics | 0
cefazolin | 0
gentamycin | 0
surgical debridement | 24
segmental partial mastectomy | 24
subtotal excision of both the outer quadrants of the right breast | 24
nipple and areola spared | 24
intraoperative wound tissue and exudate collected for microbiological examination | 24
area of 13×27 cm of excised breast tissue sent for histopathological examination | 24
histopathological examination described breast tissue with fibrosis, fat necrosis, chronic inflammation, and hemorrhage | 24
intubated | 24
stable vital signs | 24
hyperbaric oxygen therapy commenced | 96
extubated | 120
microbiology culture identified Staphylococcus aureus | 120
microbiology culture identified Klebsiella pneumoniae | 120
microbiology culture identified Acinetobacter baumanii | 120
Staphylococcus epidermidis isolated by blood culture | 120
intravenous antibiotic regimen changed to vancomycin | 120
intravenous antibiotic regimen changed to meropenem | 120
wounds managed with negative pressure wound therapy dressings | 120
foam dressings changed every 48 hours | 120
wounds appeared clean, healing with pink granulation tissue present, and reduced in size | 432
breast defect surgically repaired using a nipple and areola centralization technique | 432
defects in the right chest and flank continued to be managed with NPWT dressings | 432
discharged from the hospital with a portable NPWT device for home use | 744
CT scan of the soft tissues and breast performed every 14 days | 744
wounds had healed successfully | 1200
breast shape and volume retained with a good cosmetic effect | 1200