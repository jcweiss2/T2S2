54 years old | 0
male | 0
admitted to the hospital | 0
gastroesophageal reflux disease | -672
degenerative disc disease | -672
subacute onset of subjective fevers | -336
chills | -336
arthritis of his right knee | -336
arthritis of his left wrist | -336
erythema | -336
pain | -336
swelling | -336
visited a walk-in clinic | -336
prescribed naproxen | -336
temperature was 37.1°C | 0
pulse was 80 beats per minute | 0
blood pressure was 109/62 mm Hg | 0
respiratory rate was 24 breaths per minute | 0
oxygen saturation was 97% on room air | 0
grade III to VI early diastolic murmur | 0
faint crackles to the lung bases | 0
mild swelling and pain to his right knee | 0
mild swelling and pain to his left wrist | 0
no erythema | 0
no rash on his skin or mucosal surfaces | 0
diffuse bilateral B-lines | 0
pulmonary edema | 0
aortic regurgitation | 0
neutrophil-dominant leukocytosis | 0
hemoglobin of 126 g/L | 0
platelets of 164 × 10^9/L | 0
creatinine of 137 μmol/L | 0
C-reactive protein was 209 mg/L | 0
liver enzymes were within normal limits | 0
pulmonary edema on chest radiography | 0
complete heart block with a ventricular escape rate on electrocardiography | 0
bicuspid aortic valve | 0
severe aortic insufficiency | 0
aortic root abscess | 0
moderate mitral insufficiency | 0
fistula from the right ventricle to the aortic root | 0
blood cultures grew Neisseria gonorrhoeae | 0
gonococcal endocarditis | 0
empiric administration of intravenous ceftriaxone | 0
empiric administration of vancomycin | 0
stopped vancomycin | 24
prescribed oral azithromycin | 24
continued ceftriaxone | 24
admitted to the cardiac intensive care unit | 24
modified Bentall procedure | 48
surgical aortic valve replacement | 48
insertion of a bioprosthetic valve | 48
aortic root repair | 48
venous–arterial extracorporeal membrane oxygenation | 48
inotropic support | 48
temporary transvenous pacing | 48
aortic valve tissue gram stain and culture were negative for bacteria | 72
16S rRNA gene sequencing of aortic valve tissue confirmed the presence of N. gonorrhoeae | 72
NG-MAST of the porA and tbpB genes | 72
valvular pathology showed an active purulent process with neutrophilic infiltration | 72
acute tubular necrosis | 168
continuous renal replacement therapy | 168
implantation of a dual-chamber permanent pacemaker | 336
continued administration of ceftriaxone for 28 days | 336
transitioned from continuous renal replacement therapy to intermediate hemodialysis | 672
discharged home | 720
kidney function improved | 1440
stopped hemodialysis | 1440
nephrology follow-up | 2640