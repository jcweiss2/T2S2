55 years old | 0
male | 0
nonalcoholic steatohepatitis | -672
alpha 1 antitrypsin deficiency | -672
orthotopic liver transplant | 0
incarcerated inguinal hernia | 0
hernia repair | 0
cytomegalovirus viremia | 0
valganciclovir treatment | 0
discharged | 0
mycophenolate mofetil | 0
tacrolimus | 0
prednisone | 0
encephalopathy | 336
increasing home oxygen requirements | 336
admitted to hospital | 336
required 4L nasal cannula | 336
oxygen saturation >92% | 336
sparse speech | 336
disorientation | 336
nonfocal neurologic examination | 336
white blood cell count 9.3 × 10^9/L | 336
creatinine 2.12 mg/dL | 336
blood urea nitrogen 53 mg/dL | 336
arterial ammonia 204 µmol/L | 336
induction dosing of intravenous ganciclovir | 336
empiric antibiotic coverage with vancomycin | 336
meropenem | 336
micafungin | 336
intravenous micronutrient supplementation for B1, B6, and levocarnitine | 336
lumbar puncture | 336
encapsulated yeast suspicious for Cryptococcus | 336
liposomal amphotericin B | 336
flucytosine | 336
continuous renal replacement therapy (CRRT) | 336
rifaximin | 336
zinc | 336
lactulose | 336
ammonia level climbed to 692 µmol/L | 360
neurological deterioration | 360
mechanical ventilation | 360
empiric intravenous doxycycline | 360
urine and bronchial aspirate obtained for Mycoplasma and Ureaplasma PCR | 360
ammonia levels fell to <100 µmol/L | 384
Cryptococcal serum and cerebrospinal fluid (CSF) antigen titers positive | 384
cultures from bronchoalveolar lavage, CSF, and blood revealed cryptococcal growth | 384
repeat lumbar punctures | 384
opening pressures greater than 45 cmH2O | 384
large volume drainage every 48 hours | 384
thrombocytopenia | 384
mental status transiently improved | 408
unable to wean from mechanical ventilation | 408
tracheostomy | 408
persistent hydrocephalus | 432
oliguric renal failure | 432
progressive splenic infarcts with necrosis | 432
splenectomy | 432
sepsis | 432
duodenal leak | 432
renal failure | 432
failure to thrive | 432
moved to comfort care in hospice | 456
urea cycle disorder screening studies | 456
low urine orotic level | 456
normal serum citrulline and arginine level | 456