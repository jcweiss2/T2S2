23 years old | 0
female | 0
pregnant | 0
36th week of gestation | 0
admitted to the emergency room | 0
high-grade fever | -168
abnormal movements of eyes and limbs | -168
fever onset | -168
abnormal movements onset | -167
no history of drug or toxin intake | 0
no significant past medical history | 0
restless | 0
sick | 0
blood pressure 90/50 mm Hg | 0
pulse rate 120 beats/minute | 0
respiratory rate 32 breaths/minute | 0
oxygen saturation 96% on room air | 0
bilateral basal crepitations | 0
cigarette burn eschar | 0
conscious | 0
oriented to time, place and person | 0
conjugate, chaotic, multidirectional eye movements | 0
myoclonic jerks | 0
normal tone | 0
normal power | 0
normal deep tendon reflexes | 0
no features of parkinsonism | 0
no features of cerebellar dysfunction | 0
elevated leukocyte count | 0
thrombocytopenia | 0
deranged renal function | 0
deranged hepatic function | 0
normal serum electrolyte levels | 0
emergency cesarean section | 0
intensive care admission | 0
treated with injectable azithromycin | 0
supportive management | 0
diagnosis of scrub typhus confirmed by IgM ELISA | 0
vasculitis markers negative | 0
autoimmune and paraneoplastic antibody profile nonrevelatory | 0
serology for HIV, hepatitis B, and hepatitis C negative | 0
VDRL test negative | 0
brain MRI with contrast normal | 0
cerebrospinal fluid examination normal | 0
electroencephalography normal | 0
PET-CT of the whole body normal | 0
OMS resolved over two weeks | 336
no specific treatment or immunotherapy | 336 
opsoclonus-myoclonus syndrome | -168 
discharged | 336