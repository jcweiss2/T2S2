61 years old | 0
male | 0
admitted to the hospital | 0
dyspnoea | 0
NYHA class IV | 0
anasarca | 0
electrocardiogram demonstrates ventricular fibrillation | 0
ventricular fibrillation | -144
internal cardioverter defibrillator interrogation | 0
type 2 amiodarone-induced thyrotoxicosis | -336
discontinuation of amiodarone | -336
initiation of thiamazole therapy | -336
normal thyroid function tests | -336
trans-oesophageal echocardiogram | 480
no evidence of intracardiac thrombi | 480
external defibrillations | 480
re-initiation of oral amiodarone | 480
discontinuation of amiodarone | 672
acute kidney injury | 1008
anuria | 1008
admission to the intensive care unit | 1008
initiation of continuous veno-venous haemodialysis | 1008
exacerbation of chronic driveline infection | 1024
shared decision for best supportive care | 1024
death | 1104
septic shock | 1104
multi-organ failure | 1104
left ventricular assist device implantation | -6048
dilated cardiomyopathy | -6048
heart failure | -6048
morbid obesity | -3024
chronic driveline infection | -6048
absent arterial pulse | 0
normal capillary refill time | 0
normal core temperature | 0
unremarkable neurologic exam | 0
elevated serum creatinine | 0
elevated N-terminal prohormone of brain natriuretic peptide | 0
elevated serum lactate level | 0
global akinesia of all cardiac chambers | 0
profound dilation of the right ventricle | 0
faint movements of the tricuspid valve leaflets | 0
initiation of intravenous furosemide | 0
external defibrillation | 0
multiple unsuccessful attempts to restore normal rhythm | 480
initiation of oral amiodarone | 480
multiple unsuccessful defibrillations | 672
end-stage renal failure | 1008
sepsis | 1104