27 years old | 0
Hispanic | 0
male | 0
admitted to the hospital | 0
fevers | -120
chills | -120
intermittent epigastric pain | -120
pain started acutely | -120
eating dinner | -120
burning pain | -120
non-radiating pain | -120
pain lasted 20 minutes | -120
pain recurred | -120
subjective fevers | -48
subjective chills | -48
vomiting | -48
denies diarrhea | -48
denies sick contacts | -48
denies recent travel | -48
denies dysuria | -48
denies hematuria | -48
denies chest pain | -48
denies shortness of breath | -48
tachycardic | 0
afebrile | 0
normotensive | 0
diaphoretic | 0
mildly jaundiced | 0
sclera icteric | 0
lungs clear | 0
cardiac exam negative | 0
extremities normal | 0
no edema | 0
no rash | 0
mildly tender in epigastrium | 0
abdomen soft | 0
abdomen non-distended | 0
no rebound tenderness | 0
no involuntary guarding | 0
no Rovsing’s sign | 0
no Obturator sign | 0
no Murphy’s sign | 0
leukocytosis | 0
toxic granulations | 0
neutrophilic predominance | 0
thrombocytopenic | 0
elevated D-dimer | 0
elevated fibrinogen | 0
elevated total bilirubin | 0
elevated alkaline phosphatase | 0
normal chest radiograph | 0
normal electrocardiogram | 0
treated for severe sepsis | 0
treated for septic shock | 0
received normal saline | 0
received broad-spectrum antibiotics | 0
vital signs normalized | 12
feeling better | 12
abdominal ultrasound | 12
liver normal | 12
no intra- or extra-hepatic ductal dilatation | 12
kidneys normal | 12
aorta normal | 12
spleen normal | 12
pancreas normal | 12
gallbladder wall thickened | 12
no stones | 12
no sludge | 12
no peri-cholecystic fluid | 12
surgical consult | 12
possible acute cholecystitis | 12
possible cholangitis | 12
admitted to medical intensive care unit | 24
infectious workup | 24
tested for influenza | 24
tested for viral hepatitis | 24
tested for HIV | 24
tested for malaria | 24
tested for tularemia | 24
blood cultures grew E. coli | 48
antibiotics tailored | 48
CT of abdomen and pelvis | 72
dilated and thick walled retrocecal appendix | 72
adjacent inflammation | 72
free fluid | 72
inflammation of gallbladder wall | 72
laproscopic appendectomy | 96
procedure without complications | 96
intravenous antibiotics continued | 96
discharged | 144
elevated white blood cell count | 144
elevated total bilirubin | 144
antibiotics discontinued | 144
follow-up in surgery clinic | 168
feeling better | 168
minimal pain | 168
staples removed | 168
lost to follow up | 168
pylephlebitis diagnosed | 72
pylephlebitis treated | 72
anticoagulation not used | 72