52 years old | 0
male | 0
admitted to intensive care unit | 0
high grade fever | 0
shortness of breath | 0
hypotension |4 0
urosepsis | 0
poor oral intake | -672
significant weight loss | -672
no cough | -672
no expectoration | -672
no nausea | -672
no vomiting | -672
no dysuria | -672
no bleeding | -672
no loose bowel movements | -672
no alteration of higher mental functions | -672
drinking unpasteurized camel milk | -672
hypertension | -672
diabetes | -672
single | -672
denies sexual activities | -672
military service | -672
no past history of sexually transmitted diseases | -672
no blood transfusion | -672
no homosexuality | -672
no travel outside the country | -672
moderate distress | 0
febrile (38.1°C) | 0
decreased breath sounds bilaterally | 0
blood pressure 100/50 mmHg | 0
visible carotid pulsations | 0
no bruits | 0
non-elevated jugular venous pressure | 0
normal heart sounds | 0
soft abdomen | 0
non-tender abdomen | 0
no hepatosplenomegaly | 0
no pain on deep palpation | 0
hemoglobin 85 g/liter | 0
total leucocyte count 6200/mm3 | 0
normal platelet count (1.6 × 109/liter) | 0
C reactive protein 222 mg/L | 0
no malaria parasites | 0
internal hemorrhoids | 0
gastritis | 0
negative Helicobacter pylori stain | 0
CT scan no mediastinal lymphadenopathy | 0
CT scan no hilar lymphadenopathy | 0
CT scan no axillary lymphadenopathy | 0
3 cm right pleural effusion | 0
1.4 cm left pleural effusion | 0
minor pericardial effusion | 0
no focal changes in liver | 0
no focal changes in pancreas | 0
no focal changes in spleen | 0
no focal changes in kidneys | 0
no focal changes in adrenals | 0
no retroperitoneal lymphadenopathy | 0
no intraperitoneal lymphadenopathy | 0
minor free abdominal fluid | 0
lesser pelvic fluid | 0
non-typhoidal Salmonella Group D in blood | 0
non-typhoidal Salmonella Group D in urine | 0
sensitivity to piperacillin/tazobactam | 0
sensitivity to ciprofloxacin | 0
sensitivity to ampicillin | 0
resistance to cefuroxime | 0
resistance to gentamicin | 0
resistance to trimethoprim/sulfamethoxazole | 0
investigation for malignancy | 0
investigation for tuberculosis | 0
investigation for HIV | 0
positive ELISA | 0
positive Western blot | 0
HIV diagnosis | 0
negative cytology for malignancy | 0
negative sputum smears | 0
negative fluorescence microscopy for acid-fast bacilli | 0
treated with ciprofloxacin | 0
switched to piperacillin/tazobactam | 72
treatment duration 7 days | 168
negative urine culture | 168
recovered without renal complications | 168
