76 years old | 0
male | 0
admitted to the hospital | 0
fatigue | -720
anorexia | -720
dyspnea | -720
hypertension | 0
type two diabetes | 0
smoking | 0
alcoholism | 0
temperature 37.8 degrees Celsius | 0
heart rate 56 beats per minute | 0
blood pressure 132/53 mmHg | 0
respiratory rate 40 per minute | 0
oxygen saturation 94% on room air | 0
bilateral pulmonary crackles | 0
white blood cell count of 35,000/μL | 0
creatinine of 1.38 mg/dL | 0
troponin-I of 0.128 ug/L | 0
pulmonary edema | 0
first degree AV block | 0
left bundle branch block | 0
treated with ceftriaxone | 0
treated with furosemide | 0
treated with supplemental oxygen | 0
worsening dyspnea | 24
third degree heart block | 24
transvenous pacing | 24
aortic valve endocarditis | 24
transferred to the coronary care unit | 48
transesophageal-echocardiography | 48
native aortic valve endocarditis | 48
vegetation and abscess | 48
fistula into left ventricular outflow tract | 48
small shunt into the right atrium | 48
mitral-aortic continuity involvement | 48
large vegetation | 48
gram negative rods in blood cultures | 120
Capnocytophaga canimorsus identified | 144
sensitive to ceftriaxone | 144
sensitive to ampicillin | 144
sensitive to ciprofloxacin | 144
dog exposure | 144
severe dog bites | -2160
cardiac surgery | 240
aortic valve replacement | 240
mitral valve repair | 240
closure of a Sinus of Valsalva aneurysm | 240
pathology of the aortic valve | 240
negative gram-stain | 240
negative bacterial culture | 240
post-operative blood cultures negative | 240
discharged | 480
antimicrobial treatment | 0 
planned duration of antimicrobial treatment six weeks | 0