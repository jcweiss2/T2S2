57 years old | 0
female | 0
intractable low back pain | -8760
severely impaired mobility | -8760
lumbar laminectomy and fusion | -8760
posterior spinal instrumentation | -8760
motor strength 4/5 in lower limbs | -8760
decreased sensation in bilateral dermatomes | -8760
adjacent segment disease | -8760
revision surgery | 0
posterior laminectomies | 0
posterior spinal fusion | 0
bilateral transpedicular instrumentation | 0
hemovac drain placement | 0
severe headache | 48
somnolence | 48
left hemiparesia | 48
intraparenchymal hemorrhage in right parietal lobe | 48
subarachnoid hemorrhage | 48
bilateral symmetrical cerebellar hemorrhages | 48
pneumocephalus | 48
hemovac drain removal | 48
antiedema treatment | 48
antiepileptic treatment | 48
neurological improvement | 72
in-patient rehabilitation | 72
cognitive impairment | 120
residual dysphagia | 120
neurogenic bladder | 120
aspiration pneumonia | 2160
sepsis | 2160
death | 2160