61 years old | 0
    male | 0
    arterial hypertension | -8760
    severe heart failure | -8760
    left ventricular ejection fraction of 30% | -8760
    carvedilol | -8760
    ivabradine | -8760
    losartan | -8760
    stage IIIB chronic renal failure | -8760
    urinary symptoms | -8760
    fever | -8760
    diaphoresis | -8760
    low back pain | -8760
    hypotension | -8760
    dyspnea | -8760
    increased acute phase reactants | -8760
    sepsis | -8760
    hospitalization in intensive care unit | -8760
    alterations in calcium | -8760
    severe hyperparathyroidism | -8760
    functional adenoma in the lower left parathyroid | -8760
    surgery for hyperparathyroidism | -8760
    chest x-ray lesions | -8760
    admitted for excisional biopsy | 0
    thin patient | 0
    chronic disease | 0
    deformity in the neck | 0
    severe dorsal kyphoscoliosis | 0
    secondary asymmetry of the right ribcage | 0
    decreased intercostal spaces | 0
    increased dyspnea | 0
    NYHA class III | 0
    blood pressure 120/70 mm Hg | 0
    heart rate 100 bpm | 0
    breathing frequency 16 bpm | 0
    no cyanosis | 0
    jugular engorgement at 90° | 0
    no neck masses | 0
    tachycardic rhythmic heart | 0
    no murmurs or gallop | 0
    decreased breath sounds | 0
    abdomen without ascites or masses | 0
    edema grade II | 0
    no chest wall lesions | 0
    mild anemia | 0
    moderate restrictive ventilatory pattern | 0
    no post-bronchodilator changes | 0
    DLCO 109% | 0
    chronic kidney disease stable | 0
    thoracic CT lesions | 0
    decision for surgical resection | 0
    hospitalized in ICU pre-surgically | 0
    intravenous levosimendan | 0
    red blood cell transfusion | 0
    thoracoscopic resection | 0
    partial resection of ribs | 0
    hemodynamic instability | 24
    vasoactive support with norepinephrine | 24
    prolonged mechanical ventilation | 24
    tracheostomy | 24
    vasoactive drugs removed | 168
    invasive ventilatory support removed | 168
    tracheostomy removed | 168
    physical rehabilitation | 168
    respiratory rehabilitation | 168
    ossifying lipoma diagnosis | 168
    mature adipose tissue | 168
    thin bone trabeculae | 168
    no medullary stroma | 168
    no recurrence of lesions | 168
    no chemotherapeutic treatment | 168
    frequent medical controls | 168
<|eot_id|>
