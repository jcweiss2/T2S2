40 years old|0
    woman|0
    placenta previa totalis|0
    Cesarean section|0
    first baby delivered by Cesarean section|-87600
    myomectomy|-78744
    myoma in the low portion of uterus|-78744
    preoperative laboratory tests normal|0
    invasive arterial blood pressure monitoring|0
    anesthesia induced with thiopental sodium 250 mg|0
    anesthesia induced with succinylcholine 66 mg|0
    intubation|0
    anesthesia maintained with sevoflurane 1.2 vol%|0
    anesthesia maintained with nitrous oxide 50%|0
    volume-controlled ventilation with 50% oxygen|0
    electrocardiogram monitoring|0
    bispectral index monitoring|0
    pulse oximetry monitoring|0
    end-tidal carbon dioxide partial pressure 30-35 mmHg|0
    atracurium 25 mg injected intravenously|0
    baby delivered|9
    Apgar score 8 at 1 minute|9
    Apgar score 9 at 5 minutes|9
    no complications with the fetus|9
    placenta removed|9
    bleeding observed in the uterus|9
    methyl ergonovine 0.2 mg injected intravenously|9
    central venous catheter inserted|9
    packed RBCs administered|9
    vital signs stable|9
    systolic blood pressure 110B120 mmHg|9
    diastolic blood pressure 70B80 mmHg|9
    heart rate 75B85 beatsBmin|9
    bispectral index 50B65|9
    uterine suture completed|100
    EtCO2 partial pressure dropped abruptly|100
    systolic blood pressure dropped abruptly|100
    SpO2 90%|100
    ventricular fibrillation|100
    operation stopped|100
    chest compression started|100
    additional help requested|100
    defibrillation attempted with 200 Joule|100
    epinephrine injected|100
    atropine injected|100
    bicarbonate injected|100
    chest compression continued|100
    normal sinus rhythm not returned|100
    systolic blood pressure maintained 60B100 mmHg|100
    manual ventilation with 100% oxygen|100
    arterial oxygen saturation 86%|100
    arterial blood gas analysis pH 7.32|100
    arterial blood gas analysis PaCO2 35 mmHg|100
    arterial blood gas analysis PaO2 56 mmHg|100
    arterial blood gas analysis HCO3- 18.0 mmolB|100
    arterial blood gas analysis SaO2 86.0%|100
    blood-like secretion exited endotracheal tube|100
    EtCO2 partial pressure apnea|100
    bispectral index maintained above 40|100
    cardiac compression attempted for 40 minutes|100
    defibrillation performed three times|100
    epinephrine 60 mg used|100
    atropine 5 mg used|100
    bicarbonate 120 mEq used|100
    calcium chloride 1200 mg used|100
    heart rhythm not returned|100
    CPR not stopped|100
    endotracheal tube secretion flow|100
    corrugating tube exchanged five times|100
    EtCO2 partial pressure monitoring stopped|100
    tube continuously suctioned|100
    manual ventilation maintained with 100% oxygen|100
    CPR continued for 50 minutes|100
    normal sinus rhythm returned|250
    blood pressure 90B50 mmHg|250
    heart rate 110 beatsBmin|250
    mannitol 20% 100 ml injected|250
    lasix 20 mg injected|250
    methylprednisolone 500 mg injected|250
    obstetricians re-stitched wound|250
    no urine output during CPR|250
    urine output exceeding 200 mlBhour after ROSC|250
    no uterine bleeding observed|250
    hysterectomy not performed|250
    vaginal bleeding developed|310
    heart rate increased to 120B130 beatsBmin|310
    hysterectomy performed|310
    transesophageal echocardiography probe inserted|310
    thrombus in heart not found|310
    global hypokinesia in left ventricle|310
    platelet count 39000|310
    prothrombin time 28.6 sec|310
    activated partial thrombin time 129.1 sec|310
    fibrinogen 60 mgBdl|310
    d-dimer >20 µgBml|310
    disseminated intravascular coagulation suspected|310
    whole blood 3 units transfused|310
    packed cells 10 units transfused|310
    platelets 20 units transfused|310
    fresh frozen plasma 10 units transfused|310
    total anesthesia time 8 hours 40 minutes|310
    transferred to intensive care unit|310
    chest radiography pulmonary edema|310
    transfusion and fluid therapy|310
    suspected DIC by amniotic fluid embolism|310
    recovered to drowsy state 2 hours postoperation|330
    responded to pain stimulation|330
    pulmonary edema slight improvement 6 hours postoperation|390
    transthoracic echocardiography no regional wall motion abnormality|390
    ventilator breathing|390
    alert mental state 16 hours postoperation|460
    extubation performed|460
    vital signs stable|460
    arterial blood gas analysis pH 7.605|460
    arterial blood gas analysis PaCO2 25.3 mmHg|460
    arterial blood gas analysis PaO2 98.5 mmHg|460
    arterial blood gas analysis HCO3- 24.6 mmolB|460
    arterial blood gas analysis SaO2 98.4%|460
    hemoglobin 9.9 gBdl|460
    platelet 108000|460
    PTB16.6 sec|460
    aPTT 48.5 sec|460
    fibrinogen 263 mgBdl|460
    d-dimer 4.51 µgBml|460
    sudden loss of consciousness 30 minutes post extubation|490
    cardiac arrest developed|490
    defibrillation performed|490
    mental state recovered|490
    heart rhythm recovered|490
    tachyarrhythmia 7 hours post extubation|520
    cardiac arrest developed|520
    condition deteriorated 5 days postoperation|120
    multi-organ failure|120
    ECMO support|120
    continuous renal replacement therapy|120
    died 6 days postoperation|144
    