22 years old|0
White|0
G2P1001 woman|0
presented to a county hospital|0
28 1/7 weeks of gestation|0
cerebrovascular accident tenderness|0
malaise|0
polysubstance abuse|0
methicillin-sensitive Staphylococcus aureus bacteremia (MSSA)|0
hepatitis C virus|0
undetectable viral load|0
endocarditis|-8760
admitted a year ago|-8760
treated with 6 weeks of IV antibiotics|-8760
planned for surgical management but was lost to follow-up|-8760
COVID-19 pneumonia|0
pyelonephritis|0
MSSA bacteremia|0
thrombocytopenia|0
admitted to the intensive care unit (ICU)|0
respiratory failure|0
intubated|0
transesophageal echocardiogram|0
severe tricuspid valve (TV) regurgitation|0
large TV vegetations (2 × 1 cm)|0
flail TV leaflets|0
severe valve malcoaptation|0
received betamethasone for fetal lung maturation|0
transferred to a tertiary care hospital|0
cardiothoracic surgery team recommended medical management with IV antibiotics|0
plan to consider valve surgery after delivery|0
patient's condition improved with antibiotic treatment|0
extubated|0
transferred to the maternal-fetal medicine (MFM) unit|0
29 3/7 weeks of gestation|-168
fetal monitoring|0
Subutex initiation|0
continuation of IV antibiotics|0
infectious diseases (ID) team consulted|0
recommended continuation of IV cefazolin|0
29 6/7 weeks of gestation|72
tachypneic|72
tachycardic|72
required increasing oxygen supplementation|72
computed tomography angiogram|72
new septic emboli throughout the lungs bilaterally|72
small pericardial effusion|72
multidisciplinary discussion|72
AngioVac procedure recommended|72
preprocedure echocardiogram|168
ejection fraction of 60%|168
moderate TV regurgitation|168
continued presence of mobile vegetation on the TV|168
AngioVac procedure performed|264
30 2/7 weeks of gestation|264
general anesthesia|264
continuous fetal monitoring|264
obstetrician present|264
neonatal ICU (NICU) on standby|264
placed in supine position with leftward tilt|264
Foley catheter placed|264
external fetal heart monitor placed|264
access obtained to both femoral veins|264
access obtained to right internal jugular vein|264
intracardiac echocardiogram directed to right atrium|264
intracardiac echocardiography identified vegetations on posterior and anterior leaflets of TV|264
vegetations along eustachian valve|264
AngioVac cannula introduced through right internal jugular vein|264
directed to right atrium under fluoroscopic guidance|264
ultrasound guidance directed toward vegetations|264
venous bypass circuit activated|264
multiple passes made until most vegetations (80%) were debulked|264
vegetations grew S aureus|264
procedure uncomplicated and well tolerated|264
postoperative echocardiogram|264
ejection fraction of 57%|264
continued presence of mobile vegetations on TV|264
flail TV|264
severe TV regurgitation|264
postoperative blood cultures negative|408
1 week after procedure|408
32 5/7 weeks of gestation|1032
nonreassuring fetal heart tracing of uncertain etiology|1032
delivered via uncomplicated primary low transverse CD|1032
fetal malpresentation|1032
biophysical profile of 4/8|1032
live-born male infant|1032
Apgar scores of 9 and 9|1032
placental pathology|1032
3-vessel cord|1032
no evidence of funisitis or chorioamnionitis|1032
scattered perivillous fibrin deposition|1032
calcification|1032
neonate admitted to NICU|1032
respiratory distress syndrome|1032
prematurity|1032
prolonged course due to nutritional needs|1032
discharged on day 35 of life|1032
postpartum course complicated by preeclampsia with severe features|1032
received magnesium|1032
started on long-acting nifedipine|1032
improvement|1032
transferred back to cardiothoracic surgery|1848
postpartum day 7|1848
repeat echocardiogram|1848
severe TV regurgitation|1848
TV vegetations|1848
flair leaflet|1848
Chiari network in right atrium|1848
dilated right atrium|1848
normal ventricular function|1848
patent foramen ovale|1848
blood cultures showed no growth|1848
TV replacement with porcine valve|2304
postpartum day 16|2304
primary closure of patent foramen ovale|2304
completed antibiotics course|2304
discharged on postpartum day 24|2304
