58 years old | 0
    male | 0
    presented to the Emergency Department | 0
    three-day history of fever | -72
    three-day history of worsening perineal erythema | -72
    three-day history of pain | -72
    mild seasonal allergies | 0
    very good functional status | 0
    inguinal herniorrhaphy three years prior | -26280
    fexofenadine | 0
    pseudoephedrine | 0
    not in acute distress | 0
    significant perineal cellulitis | 0
    significant pain | 0
    preoperative chest X-ray with no infiltrates | 0
    preoperative chest X-ray with no pulmonary edema | 0
    preoperative chest X-ray with no cardiomegaly | 0
    computed tomography demonstrated extensive inflammation of the perineum and scrotum | 0
    computed tomography demonstrated subcutaneous air | 0
    diagnosis of Fournier's gangrene | 0
    normotensive | 0
    tachycardic (heart rate 110 – 120 beats / minute) | 0
    no cardiac murmurs | 0
    electrocardiogram without ST, T-wave changes | 0
    no third heart sound | 0
    no peripheral edema | 0
    no jugular venous distention | 0
    clear lungs on auscultation bilaterally | 0
    baseline SpO2 98% on room air | 0
    hemoglobin 14.9 g/dL | 0
    hematocrit 44% | 0
    white blood cell count 12.7 × 10³/mL | 0
    platelet count 146,000/mL | 0
    sodium 135 mmol/L | 0
    potassium 4.3 mmol/L | 0
    chloride 99 mmol/L | 0
    HCO3 26 mmol/L | 0
    blood urea nitrogen 16 mg/dL | 0
    creatinine 1.14 mg/dL | 0
    without nourishment for >8 hours preoperatively | 0
    emergency surgical debridement of Fournier's gangrene | 0
    premedicated with midazolam 2 mg IV | 0
    anesthesia induced with propofol 200 mg IV | 0
    anesthesia induced with fentanyl 100 mcg IV | 0
    no central venous pressure monitor placed | 0
    laryngeal mask airway (LMA, size number 4) placed without difficulty | 0
    anesthesia maintained with sevoflurane 2–3% | 0
    received fentanyl 500 mcg intraoperatively | 0
    received dilaudid 1 mg intraoperatively | 0
    remained hemodynamically stable | 0
    tachypneic (respiratory rate 35 breaths/minute) | 0
    surgical blood loss ~200 mL | 0
    procedure uneventful | 0
    sevoflurane discontinued | 0
    able to follow commands | 0
    forcefully bit down on the LMA before removal | 0
    laryngospasm noted after LMA removal | 0
    concurrent tachycardia | 0
    concurrent hypertension | 0
    positive pressure via face mask unsuccessful | 0
    administered propofol IV | 0
    administered succinylcholine IV | 0
    orotracheal intubation with 7.5 ETT | 0
    bilateral rales on auscultation | 0
    pink frothy secretions suctioned | 0
    brief episode of tachycardia (120–130 beats per minute) | 0
    brief episode of hypertension (170–180/90–100 mmHg) | 0
    SpO2 85–88% despite FiO2 100% | 0
    ABG pH 7.27 | 0
    ABG PaCO2 59 mmHg | 0
    ABG PaO2 46 mmHg | 0
    ABG HCO3 16 mmol/L | 0
    ABG base excess –1.9 | 0
    ABG oxygen saturation 75% | 0
    ABG lactate 1.27 mmol/L | 0
    SIMV at 12 cycles/minute | 0
    tidal volume 750 mL | 0
    pressure support 10 cm H2O | 0
    PEEP 10 cm H2O | 0
    PEEP increased to 12 cm H2O | 0
    SpO2 >90% | 0
    peak and plateau pressures minimally elevated | 0
    ability to generate negative pressure adequate (>–25 cm H2O) | 0
    transferred to ICU | 24
    continued on SIMV | 24
    tidal volume 580 mL | 24
    FiO2 100% | 24
    pressure support 15 cm H2O | 24
    PEEP 12 cm H2O | 24
    initial ICU ABG pH 7.6 | 24
    initial ICU ABG PaCO2 25 mmHg | 24
    initial ICU ABG PaO2 165 mmHg | 24
    initial ICU ABG HCO3 27 mmol/L | 24
    initial ICU ABG SpO2 99% | 24
    ventilator adjustments made | 24
    ICU admission chest radiograph with bilateral patchy infiltrates | 24
    ICU admission chest radiograph with no pneumothoraces | 24
    ICU admission chest radiograph with no effusions | 24
    ICU admission chest radiograph with normal heart size | 24
    FiO2 weaned to 40% over 12 hours | 36
    ABG pH 7.45 | 36
    ABG PCO2 41 mmHg | 36
    ABG PaO2 78 mmHg | 36
    ABG HCO3 28 mmol/L | 36
    ABG base excess 3.8 | 36
    ABG oxygen saturation 96% | 36
    positive fluid balance during first few days | 72
    negative fluid balance thereafter | 72
    arterial line with pulse wave variability | 72
    planned re-debridement on postoperative day 2 | 48
    not extubated until postoperative day 3 | 72
    acute shortness of breath after extubation | 72
    ABG pH 7.49 | 72
    ABG PCO2 39 mmHg | 72
    ABG PaO2 62 mmHg | 72
    ABG HCO3 29 mmol/L | 72
    ABG SpO2 93% | 72
    placed on CPAP 10 cm H2O | 72
    chest radiogram improvement | 72
    patchy infiltrates persisted | 72
    administered furosemide 40 mg IV | 72
    improvement in oxygenation | 72
    improvement in shortness of breath | 72
    improvement in roentgenographic examination | 72
    received furosemide 20 mg IV two additional doses over 24 hours | 96
    weaned off oxygen on postoperative day 6 | 144
    chest radiogram near complete resolution | 144
    discharged on postoperative day seven | 168
    doing well at three-month follow-up | 2160
    uneventful skin grafting | 2160
    no general anesthesia-related complications | 2160
    