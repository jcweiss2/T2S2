73 years old | 0
male | 0
found unconscious | -1
brought to emergency department | 0
empty bottle of Supracide insecticide found | -1
suicide note found | -1
past medical history unremarkable | 0
no history of hypertension | 0
no history of diabetes | 0
body weight 45 kg | 0
comatose | 0
Glasgow coma scale score 3 | 0
pinpoint pupils | 0
blood pressure 120/100 mm Hg | 0
pulse rate 108 per minute | 0
respiration rate 24 per minute | 0
body temperature 36°C | 0
salivation increased | 0
rales increased | 0
intubated | 0
mechanical ventilation started | 0
activated charcoal given | 0
atropine given | 0
pralidoxime infusion started | 0
arterial pH 7.220 | 0
PCO2 36.7 mm Hg | 0
PO2 59.9 mm Hg | 0
bicarbonate 14.7 mmol/L | 0
serum lactate 7.8 mmol/L | 0
blood urea nitrogen 18 mg/dl | 0
serum creatinine 1.2 mg/dl | 0
plasma cholinesterase level <200 units/L | 0
blood pressure dropped to 70/40 mm Hg | 6
norepinephrine infusion started | 6
urine output decreased to 25 ml/hr | 6
blood gas analysis pH 7.154 | 6
PCO2 20.8 mm Hg | 6
PO2 323 mm Hg | 6
bicarbonate 7.1 mmol/L | 6
CRRT initiated | 6
CVVHDF started | 6
norepinephrine requirement decreased | 26
patient's condition deteriorated | 24
died on the fourth day | 96
plasma cholinesterase levels measured | 24
prefilter plasma cholinesterase levels <200 U/L | 24
postfilter plasma cholinesterase levels 358 U/L | 7
postfilter plasma cholinesterase levels 689 U/L | 24