74 years old | 0
male | 0
end-stage renal disease | 0
admitted to hospital | 0
spring | 0
syncope during hemodialysis session | -24
returned from cottage in eastern Ontario | -24
fever (38.6°C) | 24
tachycardia (101 beats/min) | 24
confused | 24
no nuchal rigidity | 24
no jaundice | 24
no cardiorespiratory abnormalities | 24
no lymphadenopathy | 24
no hepatosplenomegaly | 24
no abdominal tenderness | 24
mild anemia | 24
slight elevation in aspartate transaminase | 24
working diagnosis of sepsis | 24
started on intravenous piperacillin–tazobactam | 24
started on intravenous vancomycin | 24
clinical status deteriorated over following 4 days | 120
high-grade fevers (up to 40.1°C) | 120
decreasing level of consciousness | 120
hypotensive | 120
transferred to intensive care unit | 120
vasopressor support | 120
intubation | 120
anti-infective drugs changed to acyclovir | 120
anti-infective drugs changed to ampicillin | 120
anti-infective drugs changed to ceftriaxone | 120
anti-infective drugs changed to vancomycin | 120
anemia | 120
thrombocytopenia | 120
transaminitis | 120
marked hyperferritinemia | 120
suspicion of hemophagocytic lymphohistiocytosis | 120
magnetic resonance imaging of brain normal | 120
tick discovered attached to left calf | 120
Ixodes scapularis confirmed | 120
peripheral blood smear showed morulae within granulocytes | 120
added oral doxycycline | 120
concern for HLH | 120
bone marrow aspiration and biopsy showed hemophagocytosis | 120
blood cultures negative | 120
urine culture negative | 120
serological testing for hepatitis B negative | 120
serological testing for hepatitis C negative | 120
serological testing for HIV negative | 120
serological testing for Epstein–Barr virus negative | 120
serological testing for cytomegalovirus negative | 120
PCR tests of cerebrospinal fluid for herpes simplex virus negative | 120
PCR tests of cerebrospinal fluid for varicella zoster negative | 120
PCR tests of cerebrospinal fluid for enterovirus negative | 120
PCR tests of cerebrospinal fluid for adenovirus negative | 120
requested CSF cell count, glucose, and protein not completed | 120
ordered serology and molecular testing for tick-borne pathogens | 120
positive for Anaplasma phagocytophilum (PCR) | 120
positive for Borrelia burgdorferi (Western blot and ELISA) | 120
positive for Powassan virus (serology) | 120
diagnosed with severe human granulocytic anaplasmosis | 120
diagnosed with secondary HLH | 120
diagnosed with Lyme disease | 120
diagnosed with Powassan virus | 120
completed 10-day course of doxycycline | 120
completed 3-week course of ceftriaxone | 120
clinical improvement with antimicrobials | 120
did not start other treatments for HLH | 120
discharged home | 1320
seen in follow-up 3 months after presentation | 2280
clinically well | 2280
complete resolution of hematologic derangements | 2280
