39 years old | 0
female | 0
partial pancreaticoduodenectomy | -2190
periampullary neuroendocrine tumor | -2190
locoregional extension | -2190
metastatic lymph nodes | -2190
histopathology | -2190
neuroendocrine tumor | -2190
gastrin | -2190
Ki 67 5% | -2190
Grade 2 | -2190
liver metastases | -1092
lanreotide | -1092
sunitinib | -546
intolerance | -274
extreme fatigue | -274
muscle weakness | -274
delirium | -274
peptide receptor radiotherapy | -274
moon face | 0
hirsutism | 0
severe proximal weakness | 0
anemia | 0
hyperglycemia | 0
severe hypokalemia | 0
elevated 24-h urinary free cortisol | 0
elevated morning serum cortisol | 0
elevated plasmatic ACTH | 0
SCS | 0
EAS | 0
ketoconazole | 0
acute upper gastrointestinal bleeding | 0
hemodynamic instability | 0
subendocardial ischemia | 0
atrial fibrillation | 0
hemodynamic support | 0
Forrest Ib gastric ulcer | 0
endoscopic treatment | 0
intravenous fluconazole | 0
mental state improvement | 48
decreased morning cortisol | 48
dose titration | 48
increased liver transaminases | 120
decreased fluconazole dose | 120
cortisolemia decrease | 168
bilateral adrenalectomy | 360
hypokalemia | 360
metabolic alkalosis | 360
acetazolamide | 360
spironolactone | 360
amiloride | 360
thrombocytopenia | 360
platelet transfusions | 360
intravenous Gamma globulin | 360
bone marrow biopsy | 360
hypocellularity | 360
Eltrombopag | 360
platelet count improvement | 360
hemodynamic stability | 432
lower cortisol levels | 432
successful bilateral adrenalectomy | 432
replacement doses of hydrocortisone | 432
fludrocortisone | 432
lanreotide 120 LAR | 432
sepsis | 720
emphysematous cystitis | 720
disseminated Herpes Zoster infection | 720
antibiotics | 720
intravenous acyclovir | 720
chemoembolization | 720
liver metastases decrease | 720
rehabilitation therapy program | 17520
good general health | 17520
active life | 17520