9 years old | 0
female | 0
admitted to the hospital | 0
low-grade fever | -24
sore throat | -24
swelling of the neck | -24
dysphagia | -24
born at a rural hospital in Yemen | -9 years
received Bacillus Calmette-Guérin vaccination | -9 years
received hepatitis B vaccination | -9 years
no other vaccinations | -9 years
no known previous medical problems | 0
close contact with other sick patients | -48
brother died due to acute febrile illness | -48
febrile | 0
tachycardia | 0
average respiratory rate | 0
normal blood pressure | 0
weight 22 kg | 0
swelling of the right side of the neck | 0
inflamed pharyngotonsillar area | 0
white patches with enlarged tonsils | 0
lungs clear to auscultation | 0
hemoglobin 13.5 g/dL | 0
white blood cell count 11,700 cells/mm3 | 0
platelet count 95,000/mm3 | 0
elevated blood urea nitrogen | 0
elevated creatinine | 0
throat swab Gram stain showed gram-positive bacilli | 0
throat swab culture showed C. diphtheriae | 0
elevated troponin T level | 0
elevated creatine kinase-MB level | 0
elevated pro-brain natriuretic peptide | 0
started on DAT | 24
started on penicillin G | 24
started on ceftriaxone | 24
developed abdominal pain | 72
vomiting | 72
mild ascetic fluid collection | 72
increased blood urea nitrogen | 72
increased creatinine | 72
elevated creatine kinase-MB level | 72
contacted CDC regarding re-dosing of DAT | 72
recommended re-dosing of DAT | 72
condition continued to worsen | 120
developed generalized edema | 216
hypotension | 216
diminished urine output | 216
declared dead | 216
acute myocarditis | 216
cardiogenic shock | 216