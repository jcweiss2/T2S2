62 years old | 0
male | 0
admitted to the hospital | 0
ankle twisting injury | -72
undisplaced fracture medial malleolus | -72
below knee ankle plaster | -72
elevation | -72
analgesic with proteolytic | -72
itching | -36
pain | -36
swelling | -36
erythema | -36
fever | -36
progressive swelling | -36
crepitus | -36
blisters | -36
serous discharge | -36
discoloration of tissue | -36
necrosis | -36
foul smell | -36
slab removal | -36
clinical diagnosis of necrotizing fasciitis | -36
laboratory risk indicator for NF score | -36
erythrocyte sedimentation rate | -36
C-reactive protein | -36
white blood cells | -36
hemoglobin | -36
platelet | -36
Na | -36
creatinine kinase | -36
urea | -36
alanine transaminase | -36
total bilirubin | -36
albumin | -36
creatinine | -36
blood sugar | -36
serology for human immunodeficiency virus | -36
hepatitis B | -36
blood culture | -36
glycated hemoglobin | -36
anti-nucleosome antibody | -36
anti-dsDNA | -36
referral to tertiary care center | -24
incision in the skin | -24
local anesthetic agent infiltration | -24
lack of bleeding | -24
dishwater-colored fluid | -24
tissue dissection | -24
positive finger probe test | -24
Pseudomonas aeruginosa | -24
tissue biopsy | -24
gas gangrene | -24
piperazillin-tazobactam | -24
meropenem | -24
teicoplanin | -24
clindamycin | -24
above knee amputation | -168
debridement | -168
septic shock | -168
acute renal failure | -480
death | -480
limb cleaning | -72
plaster material | -72
gypsum | -72
cotton bandage | -72
thermogenic effect | -72
inadequate wrap | -72
soft roll | -72
Stockey net | -72
tap water | -72
plastic bucket | -72
culture for Pseudomonas | -72