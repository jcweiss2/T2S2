47 years old | 0
woman | 0
admitted to the emergency department | 0
fever | -96
left loin pain | -96
autosomal dominant polycystic kidney disease | 0
polycystic liver disease | 0
blood pressure 127/91 mmHg | 0
heart rate 133 beats/min | 0
respiratory rate 20/min | 0
body temperature 38.5 °C | 0
hard mass palpable at belly button on right abdomen | 0
no abdominal tenderness | 0
percussion pain in left kidney area | 0
leukocytosis 10.62 × 10^9/L | 0
platelet count 97 × 10^9/L | 0
C-reactive protein 214.5 mg/L | 0
serum creatinine 97.6 μmol/L | 0
plasma fibrinogen 6.63 g/L | 0
numerous white blood cells in urine | 0
computed tomography revealed multiple air pockets in left collecting system | 0
multiple hypodense cysts in bilateral kidneys | 0
multiple renal stones in left pelvis | 0
left hydronephrosis | 0
diagnosed with left type I EPN | 0
diagnosed with ADPKD | 0
oral antibiotic treatment (nitrofurantoin 100 mg q8 h) | 0
condition rapidly deteriorated | 24
insertion of double “J” stent on left side | 24
urine specimen collection for culture | 24
left collecting system full of pus | 24
culture yielded ESBL-positive Escherichia coli | 24
antibiotics changed to imipenem-cilastatin | 24
postoperative CT showed left D-J tube well positioned | 24
air spaces in left collecting system disappeared | 24
left hydronephrosis significantly better | 24
discharged | 432
readmitted | 1440
oral antibiotic treatment (nitrofurantoin 50 mg q8 h) | 1440
flexible ureteroscopy lithotripsy | 1440
urine cultures negative | 1440
surgery performed | 1440
shivering | 1440
blood pressure 60/40 mmHg | 1440
heart rate 133/min | 1440
temperature 41°C | 1440
white blood cell count 0.50 × 10^9/L | 1440
platelet count 117 × 10^9/L | 1440
severe hematuria | 1440
transferred to intensive care unit | 1440
intravenous antibiotics (meropenem 1.0 g q8 h) | 1440
right internal jugular vein punctured | 1440
norepinephrine prescribed | 1440
right radial artery punctured | 1440
fresh plasma transfusion 600 mL | 1440
blood cultures negative | 1440
general condition improved | 1440
transferred back to general ward | 1440
meropenem treatment continued | 1440
postoperative CT showed stones cleared in left renal pelvis | 1440
few stones remained in lower calyx | 1440
discharged | 1440
oral antibiotics (fosfomycin trometamol 3.0 g qod) | 1440
serum creatinine remained below 100 μmol/L | 1440
CT showed no stones in left renal pelvis | 1440
stones in lower calyx smaller and fewer | 1440
