30 years old | 0
male | 0
admitted to the emergency room | 0
mechanical ileus | 0
enterocutaneous fistula | 0
abdominal pain | 0
difficulty in defecation | 0
sudden changes in mental status | 0
stupor | 0
vomiting | 0
sepsis | 0
blood pressure 60/40 mmHg | 0
heart rate 140 beats/min | 0
MELAS syndrome | -6048
partial seizure | -6048
carbamazepine | -6048
valproic acid | -6048
mental retardation | -6048
cerebral infarction | -6048
lactic acidosis | -6048
white blood cells 2.9 × 10^3 /μl | 0
lactic acid 142.1 mg/dl | 0
aspartate transaminase 141.1 U/L | 0
alanine transaminase 124.7 U/L | 0
creatine kinase 353.0 U/L | 0
CK-MB 20.79 ng/ml | 0
blood urine nitrogen 36.7 mg/dl | 0
creatinine 1.10 mg/dl | 0
prothrombin time 17.7 s | 0
international normalized ratio 1.57 | 0
activated partial thromboplastin time 56.7 s | 0
metabolic acidosis | 0
pH 7.170 | 0
PaO2 129.5 mmHg | 0
PaCO2 36.8 mmHg | 0
base excess −15.2 mM/L | 0
HCO3- 13.6 mM/L | 0
lactate 131.7 mg/dl | 0
Wolff–Parkinson–White syndrome | 0
high sensitivity troponin-T 205 ng/L | 0
pro B-type natriuretic peptide 313.7 pg/ml | 0
hypoglycemia 55.1 mg/dl | 0
dobutamine | -1
norepinephrine | -1
drowsy-to-stupor mental status | 0
cardiopulmonary resuscitation not performed | 0
emergency total colectomy | 0
terminal ileostomy | 0
TIVA | 0
propofol | 0
remifentanil | 0
dexmedetomidine | 0
anesthesia induction | 0
propofol infusion | 0
dexmedetomidine infusion | 5
remifentanil infusion | 5
rocuronium | 5
endotracheal intubation | 5
mechanical ventilation | 5
fluid management | 5
hypotension | 80
epinephrine | 80
vasopressin | 80
dexmedetomidine stopped | 180
remifentanil stopped | 205
sugammadex | 210
extubation | 212
discharged to intensive care unit | 210
cardiac arrest | 720
death | 720
sepsis persisted | 720
condition worsened | 720