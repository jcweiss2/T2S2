67 years old | 0
male | 0
admitted to the hospital | 0
sudden onset confusion | 0
dysarthria | 0
tested positive for SARS-CoV-2 | -336
symptoms of sore throat | -336
headache | -336
fever | -336
body aches | -336
diarrhea | -336
initial symptoms improved | -168
symptomatically hypoxic | 0
oxygen saturation of 75% on room air | 0
oxygen saturation improved to 95% | 0
lymphocytopenia | 0
thrombocytopenia | 0
borderline lactic acidosis | 0
mixed respiratory and metabolic acidosis | 0
bilateral airspace opacities | 0
generalized seizure | 12
cardiac arrest | 12
resuscitation | 12
heparin anticoagulation initiated | 12
vasopressors initiated | 12
mechanical ventilation initiated | 12
ventilator set to airway-pressure-release-ventilation mode | 12
switched to pressure-control mode | 24
focal region or wedge-shaped low attenuation in the left temporal region | 24
diffuse subpleural pneumonitis | 24
regions of ground-glass opacities | 24
consolidation | 24
paraseptal emphysema | 24
acute bilateral pulmonary emboli | 24
evidence of right ventricular dysfunction | 24
increasing vasopressor requirements | 120
increasing oxygen demands | 120
unchanged chest radiograph | 120
comfort care measures initiated | 120
terminally extubated | 120
died | 120 
hypercoagulability | -336
hyper-tension | 0
dyslipidemia | 0
prothrombin time-international normalized ratio | 0
sequential organ failure assessment score | 0
SIC score calculated to be 5 | 0
D-dimer | 0
prothrombin time | 0
complete blood count | 0 
white blood cell count | 0
hemoglobin | 0
hematocrit | 0
platelets | 0
absolute lymphocytes | 0
lactic acid | 0
creatinine | 0
albumin | 0
troponin I | 0
troponin T | 0
NT-proBNP | 0
PaO2/FiO2 | 0 
INR | 0