45 years old | 0
male | 0
referred to our hospital | 0
admitted to our hospital | 0
general malaise | 0
fever | 0
2-week history of purpura | -336
pancytopenia | 0
leukopenia | 0
anemia | 0
thrombocytopenia | 0
computed tomography showed diffusely increased bone marrow concentration | 0
no liver enlargement | 0
no splenic enlargement | 0
bone marrow aspiration unsuccessful | 0
bone marrow biopsy | 0
acute panmyelosis with myelofibrosis | 0
induction therapy started | -192
idarubicin hydrochloride | -192
cytosine arabinoside | -192
cefozopran treatment started | -336
left cheek cellulitis | -576
cellulitis failed to respond to cefozopran | -576
switched to meropenem/vancomycin | -648
blood cell recovery | -672
improved cellulitis | -672
antibiotic therapy switched to levofloxacin | -672
bone marrow aspiration failed | -672
peripheral blood cell count within normal limits | -672
Wilm's tumor 1 mRNA count decreased | -672
hematological complete remission | -672
consolidation therapy started | -672
febrile neutropenia | -504
switched levofloxacin to cefozopran | -504
sustained hyperthermia | -552
blood culture test performed | -552
indwelling central venous catheter removed | -552
chest radiograph showed pneumonia | -576
switched to meropenem and amikacin | -576
transferred to ICU | -576
intubation | -600
blood culture revealed S. maltophilia | -600
sputum culture revealed S. maltophilia | -600
SMX-TMP administered | -600
levofloxacin administered | -600
ceftazidime administered | -600
minocycline administered | -600
hematic tracheal aspirates reported | -624
intravenous granulocyte-colony stimulating factor administered | -624
neutropenia resolved | -648
ventilator condition deteriorated | -648
airway pressure-release ventilation initiated | -672
intermittent prone positioning initiated | -672
respiratory failure | -672
PaO2/FiO2 ratio 69.5 | -672
FiO2 0.85 | -672
PaCO2 40 mmHg | -672
respiratory rate 20 | -672
PEEP 14 | -672
PIP 27 cmH2O | -672
chest CT showed massive consolidation | -672
opacities around lung fields | -672
use of catecholamines reduced | -672
met ARDS criteria | -672
severe ARDS | -672
bronchoalveolar lavage cell counts | -672
blood culture negative | -672
sputum culture negative | -672
VV ECMO initiated | -816
ventilator settings lowered | -816
right lung collapsed | -816
left lung partially collapsed | -816
VV ECMO-dependent | -816
tracheotomy performed | -840
partially awakened | -840
lungs gradually opened | -840
regained spontaneous breathing | -840
active mobilization of bronchial secretions | -840
weaned off VV ECMO | -888
mechanical ventilation support | -888
bilateral pulmonary infiltration improved | -888
biphasic positive airway pressure weaned | -1056
oxygen supplementation discontinued | -3144
discharged from hospital | -3480
chest CT showed improved pneumonia | -3480
additional consolidation chemotherapy postponed | -3480
regained functional status | -3480
subsequent consolidation chemotherapy | -3480
allogenic hematopoietic stem cell transplantation | -3480
complete remission | -3480
