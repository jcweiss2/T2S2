39 years old | 0
male | 0
PEG tube dependence (replaced 6 months prior) | -4320
high grade fever of 103F | -24
recurrent episodes of coffee ground emesis | -24
intubated | 0
diffused crackles throughout the lung fields | 0
mild epigastric distention | 0
left lower quadrant tenderness | 0
PEG tube in place | 0
loose external bumper | 0
clean insertion site | 0
unable to twirl PEG tube | 0
unable to retract PEG tube | 0
unable to advance PEG tube | 0
normal sphincter tone | 0
hemoccult negative stool | 0
hemodynamically unstable | 0
low blood pressure | 0
norepinephrine | 0
mechanical ventilation | 0
100% fraction of inspired oxygen | 0
white blood cells 26,000 k/ul | 0
hemoglobin 12.9 g/dl | 0
granulocyte 80.1% | 0
sodium 157 mmol/l | 0
potassium 2.9 mmol/L | 0
chloride 116 mmol/L | 0
bicarbonate 31 mmol/l | 0
BUN 50 mg/dl |&lt;!&gt;!
