66 years old | 0
female | 0
admitted to the hospital | 0
crown tumor | -672
clear-cell carcinoma | -672
computed tomography (CT) | -672
right renal tumor | -672
lung metastases | -672
bone metastases | -672
metastatic right renal cell carcinoma | -672
cT1bN0M1 | -672
laparoscopic right renal resection | -672
sunitinib | -504
axitinib | -168
nivolumab | 0
pazopanib | 0
IMDC intermediate risk | 0
serum uric acid level | 0
normal serum uric acid level | 0
discharged | 240
CTCAE v4.0 grade 2 fatigue | 48
CTCAE v4.0 grade 2 nausea | 48
grade 1 diarrhea | 48
temperature of 40.5°C | 48
blood pressure of 132/48 mm Hg | 48
heart rate of 120 beats per minute | 48
no abdominal pain | 48
lung metastasis decreased | 48
CTCAE grade 2 acute kidney injury | 48
disseminated intravascular coagulation | 48
hydration | 48
thrombomodulin alpha | 48
broad-spectrum antibiotics meropenem | 48
hyperphosphatemia | 72
hyperuricemia | 72
hypocalcemia | 72
acute renal failure | 72
tumor lysis syndrome (TLS) | 72
intensive care unit | 72
renal replacement therapy | 96
poor prognosis | 96
palliative care | 120
death | 120