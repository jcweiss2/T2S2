42 years old | 0
male | 0
admitted to the hospital | 0
high-grade fever | -504
chills | -504
productive cough | -504
weight loss | -336
diarrhea | -336
right middle zone consolidation | -504
Klebsiella pneumoniae | -504
levofloxacin | -504
amikacin | -504
metronidazole | -504
fluconazole | -504
empiric anti-tuberculosis therapy | -504
recurrent upper respiratory tract infections | -7200
pneumonia | -6048
pulmonary tuberculosis | -6048
pulmonary tuberculosis | -4320
monthly episodes of watery diarrhea | -4320
fever | 0
tachycardia | 0
tachypnea | 0
blood pressure 110/60 | 0
bilateral crepitations | 0
PaO2 58 mm Hg | 0
admitted to the intensive care unit | 0
right middle and lower zone consolidation | 0
non-resolving pneumonia | 0
meropenem | 0
levofloxacin | 0
endotracheal intubation | 24
bilateral alveolar shadows | 120
PaO2/FiO2 59/1 | 120
noradrenaline | 120
targocid | 120
colistin | 120
amphotericin-B | 120
trimethoprim-cotrimoxazole | 120
primary immune deficiency | 120
CVID | 120
intravenous immunoglobulin | 168
hypogammaglobulinemia | 168
afebrile | 192
reduced FiO2 requirements | 192
tracheostomy | 744
decannulation | 768
clearing of alveolar shadows | 768
residual bronchiectasis | 768
ambulatory | 2160
discharge | 2160
follow-up | 2160
replacement IVIG | 2160
chest physiotherapy | 2160