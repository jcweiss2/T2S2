57 years old | 0
female | 0
type 2 diabetes | 0
poorly controlled | 0
HbA1c 148 mmol/mol | 0
lower back pain | 0
no trauma | 0
history of right hallux apical neuropathic ulcer | -120
complicated by osteomyelitis | -120
non-healing wound following left forefoot amputation | -288
left fifth toe ulcer | -408
peripheral vascular disease | 0
peripheral neuropathy | 0
diabetic retinopathy | 0
diabetic nephropathy | 0
atrial fibrillation | 0
hypertension | 0
WHO performance status score 2 | 0
Metformin MR 1 g twice-daily | 0
Lantus 18 units at night | 0
aspirin 75 mg once-daily | 0
bisoprolol 7.5 mg once-daily | 0
cholecalciferol 20 000 units once week | 0
ramipril 5 mg once-daily | 0
rivaroxaban 20 mg once-daily | 0
acutely confused | 0
septic | 0
no headache | 0
no respiratory symptoms | 0
no urinary symptoms | 0
no gastrointestinal symptoms | 0
BP 102/84 mmHg | 0
heart rate 110/min | 0
temperature 33.7°C | 0
normal heart sounds | 0
no added murmurs | 0
clear chest | 0
unremarkable abdominal examination | 0
soft tissue infection | 0
capillary refill time 3 s | 0
biphasic Doppler signals | 0
lumbar vertebral tenderness | 0
bilateral lower limb weakness | 0
absent reflexes | 0
acute renal failure | 0
profound metabolic acidosis | 0
oliguria | 0
pH 7.13 | 0
pCO2 4.2 kPa | 0
lactate 14.6 mmol/L | 0
bicarbonate 10.3 mmol/L | 0
base excess -18.9 mmol/L | 0
normal confusion screen | 0
negative chest radiograph | 0
negative urine cultures | 0
no acute intracranial haemorrhage | 0
no collection | 0
no infarct | 0
collapsible inferior vena cava | 0
poorly filled right ventricle | 0
significant volume depletion | 0
no abdominal free fluid | 0
no abdominal aortic aneurysm | 0
diffusely diseased arteries | 0
calcified plaques | 0
no haemodynamically significant stenosis | 0
biphasic spectral waveforms | 0
mixed growth | 0
Pseudomonas sp. | 0
yeast | 0
negative right foot wound swabs | 0
previous foot ulcer swabs | -408
mixed anaerobes | -408
S. aureus | -408
Pseudomonas sp. | -408
Beta haemolytic group B Streptococcus | 0
severely impaired systolic function | 0
Visual EF 25-30% | 0
unremarkable abdominal imaging | 0
severe osteomyelitis | 24
L3/L4 discitis | 24
L4/L5 discitis | 24
adjacent vertebral end-plate oedema | 24
posterior epidural collection | 24
canal compression | 24
T12 to L4 | 24
ciprofloxacin | 24
gentamicin | 24
meropenem | 48
ceftriaxone | 72
improved inflammatory markers | 168
persistent lower limb neurology | 168
further signs of sepsis | 1920
death | 1920
septicaemia | 1920
epidural abscess | 1920
diabetic foot ulcer | 1920