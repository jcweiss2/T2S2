73 years old | 0
man | 0
brought to the Emergency Department | 0
altered mental status | -72
weak | -672
lethargic | -672
agitated | 0
confused | 0
not oriented to person | 0
not oriented to place | 0
not oriented to time | 0
febrile | 0
101.5°F | 0
tachycardic | 0
pulse 115/min | 0
regular rate | 0
regular rhythm | 0
hypotensive | 0
blood pressure 85/60 mm Hg | 0
respiratory rate 20/min | 0
oxygen saturation 99% | 0
multiple stage 3 to 4 draining ulcers | 0
left lower extremity | 0
bilateral lower-extremity +2 pitting edema | 0
no tenderness | 0
no ecchymosis | 0
no external signs of trauma | 0
leukocytosis | 0
13,000/µL | 0
bandemia 27% | 0
dehydration | 0
elevated lactate 47 mg/dL | 0
urinary tract infection | 0
urine output decreased | 0
150 ml in 5 h | 0
infection | 0
cellulitis | 0
decubitus ulcers | 0
sepsis criteria | 0
4-liter bolus of normal saline | 0
maintenance rate 250 ml/h | 0
broad-spectrum IV antibiotics | 0
hypotensive persisted | 0
vasopressors initiated | 0
norepinephrine | 0
normal cardiac markers | 0
normal EKG | 0
normal sinus rhythm | 0
tachycardia | 0
echocardiography ejection fraction 55% | 0
mild diastolic dysfunction | 0
central venous pressure 8 cmH2O | 0
cardiogenic shock ruled out | 0
transferred to intensive care unit | 0
surgical debridement | 0
infected decubitus ulcer | 0
initial blood cultures | 0
wound cultures | 0
Streptococcus agalactiae | 0
urine culture | 0
Citrobacter amalonaticus | 0
WBC count trended down | 0
lactic acid normalized | 0
Doppler studies | 0
right lower-extremity occluding thrombus | 0
popliteal vein | 0
superficial femoral vein | 0
weight-based unfractionated heparin | 0
adjusted daily | 0
coagulation profile | 0
cell counts measured daily | 0
PT measured daily | 0
INR measured daily | 0
aPTT measured daily | 0
anti-Factor Xa activity measured daily | 0
fibrinogen 220 mg/dL | 0
fibrinogen degradation product 35 mg/dL | 0
D-dimer 300 ng/mL | 0
DIC ruled out | 0
altered consciousness persisted | 0
lab values stable | 0
hemoglobin drop | 72
13.4 g/dL to 6.1 g/dL | 72
heparin discontinued | 72
coagulopathy reversed | 72
2 units fresh frozen plasma | 72
4 units packed red blood cells | 72
hemoglobin steady | 72
no overt bleeding | 72
no occult bleeding | 72
fecal occult blood tests negative | 72
CT abdomen and pelvis | 72
retroperitoneal hematoma | 72
expansion left iliopsoas musculature | 72
left common iliac arteries | 72
left external iliac arteries | 72
no increase in size of hematoma | 72
serial CT scans | 72
inferior vena cava filter | 72
no angiography | 72
no surgical intervention | 72
hemoglobin stable | 72
died | 168
multi-organ failure | 168
