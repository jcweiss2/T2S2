29 years old | 0
    male | 0
    regular consumer of alcohol | 0
    heavy consumer of alcohol | 0
    lumberjack | 0
    fever | -336
    cough | -336
    confused state | 0
    septic shock | 0
    neck stiffness | 0
    bilateral upper limbs power normal | 0
    bilateral lower limbs power normal | 0
    normal tone | 0
    normal reflexes | 0
    normal heart sounds | 0
    no murmur | 0
    bilateral lung crepitations | 0
    fluid resuscitation | 0
    vasopresssor required | 0
    mechanical ventilator | 0
    admitted to intensive care unit | 0
    anaemia | 0
    thrombocytopenia | 0
    normal total white cells | 0
    normal renal function | 0
    splenic microabscesses | 0
    bilateral lung fields consolidation | 0
    normal computed tomography of the brain | 0
    no signs of inflammation in cerebrospinal fluid | 0
    no signs of infection in cerebrospinal fluid | 0
    Burkholderia pseudomallei blood culture | 0
    ventilator associated pneumonia | 72
    multidrug-resistant Acinetobacter baumanii respiratory tract infection | 192
    bacteraemic with Burkholderia pseudomallei | 288
    left side hemiplegia | 600
    pansystolic murmur | 600
    right corona radiata infarct | 600
    high parietal petechia haemorrhage | 600
    thickened mitral valve | 600
    vegetation on posterior mitral valve leaflet | 600
    moderate eccentric mitral regurgitation | 600
    sepsis-induced supraventricular tachycardia | 168
    persistent high-grade temperature | 96
    leukopenia | 96
    oral trimethoprim-sulfamethoxazole started | 168
    IV ceftazidime | 0
    IV C-penicillin | 0
    IV imipenem | 96
    IV ampicilin-sulbactam | 336
    IV gentamicin | 168
    oral co-trimoxazole continued | 2016
    discharged | 2016
    minimal residual left sided weakness | 2016
    Modified Rankin Score of 2 | 2016
    activities of daily living independently | 2016
    intact cognitive function | 2016
    transferred to cardiac referral centre | 2016
    vegetation on mitral valve resolved | 6048
    residual moderate mitral regurgitation | 6048
    left ventricular ejection fraction 66.5% | 6048
    Modified Rankin Score of 2 at nine months | 6048
    cerebral infarct | 600
    haemorrhages | 600
    septic emboli to the brain | 600
    disseminated melioidosis | 0
    infective endocarditis | 600
    cerebral infarct complication | 600
    haemorrhages complication | 600
    blood culture no growth | 576
    blood culture no growth | 624
    blood culture no growth | 648
    blood culture Burkholderia pseudomallei | 144
    blood culture Burkholderia pseudomallei | 288
    multidrug-resistant Acinetobacter baumanii respiratory tract | 264
    fluid resuscitation | 0
    vasopresssor highest dose 0.27 mcg/kg/min | 96
    ventilator support high setting | 336
    IV noradrenaline | 0
    IV ceftazidime | 0
    IV C-penicillin | 0
    IV imipenem | 96
    oral trimethoprim-sulfamethoxazole | 168
    IV ampicilin-sulbactam | 336
    IV gentamicin | 168
    IV ceftazidime continued | 1008
    oral co-trimoxazole monotherapy | 2016
    discharged after 12 weeks | 2016
    transferred to cardiac referral centre | 2016
    follow-up at nine months | 6048
    echocardiogram resolved vegetation | 6048
    residual moderate mitral regurgitation | 6048
    left ventricular ejection fraction 66.5% | 6048
    Modified Rankin Score of 2 | 6048
    no known medical illness | 0
    missing from work | -96
    bilateral lung crepitations | 0
    bilateral lung fields consolidation | 0
    normal heart sounds | 0
    no murmur | 0
    normal computed tomography of the brain | 0
    no signs of inflammation in cerebrospinal fluid | 0
    no signs of infection in cerebrospinal fluid | 0
    Burkholderia pseudomallei confirmed by PCR | 0
    gentamicin-susceptible isolate | 0
    positive blood cultures on Day 6 | 144
    positive blood cultures on Day 12 | 288
    blood culture no growth on Day 24 | 576
    blood culture no growth on Day 26 | 624
    blood culture no growth on Day 27 | 648
    left-sided hemiparesis | 600
    pansystolic murmur | 600
    right corona radiata infarct | 600
    high parietal petechia haemorrhage | 600
    thickened mitral valve | 600
    vegetation on posterior mitral valve leaflet | 600
    moderate eccentric mitral regurgitation | 600
    septic embolus suspected | 600
    prolapsed mitral valve | 600
    cerebral infarct | 600
    haemorrhages | 600
    intensive phase therapy extended to 6 weeks | 1008
    IV ceftazidime continued | 1008
    IV gentamicin for 14 days | 168
    concurrent oral co-trimoxazole | 168
    eradication phase therapy | 2016
    activities of daily living independently | 2016
    intact cognitive function | 2016
    transferred to cardiac referral centre | 2016
    follow-up at nine months | 6048
    echocardiogram resolved vegetation | 6048
    residual moderate mitral regurgitation | 6048
    left ventricular ejection fraction 66.5% | 6048
    Modified Rankin Score of 2 | 6048
    no medical illness | 0
    alcohol consumption | 0
    fever duration 2 weeks | -336
    cough duration 2 weeks | -336
    missing from work | -96
    brought to hospital | 0
    septic shock secondary to pneumonia | 0
    blood culture Burkholderia pseudomallei | 0
    started IV ceftazidime and IV C-penicillin | 0
    ventilator associated pneumonia | 72
    multidrug-resistant Acinetobacter baumanii | 192
    bacteraemic on Day 6 | 144
    bacteraemic on Day 12 | 288
    blood culture no growth on Day 24 | 576
    blood culture no growth on Day 26 | 624
    blood culture no growth on Day 27 | 648
    left side hemiplegia | 600
    pansystolic murmur | 600
    echocardiography | 600
    computed tomography of the brain | 600
    started IV gentamicin | 168
    completed intensive phase antibiotics | 504
    discharged from hospital | 2016
    last follow-up visit | 6048
    cerebral infarct | 600
    haemorrhages | 600
    septic emboli | 600
    infective endocarditis | 600
    mitral valve vegetation | 600
    gentamicin-susceptible strain | 0
    IV ceftazidime and gentamicin combination | 168
    oral co-trimoxazole continuation | 2016
    residual left sided weakness | 2016
    Modified Rankin Score of 2 | 2016
    activities of daily living | 2016
    intact cognitive function | 2016
    transferred to cardiac centre | 2016
    follow-up at nine months | 6048
    resolved vegetation | 6048
    residual mitral regurgitation | 6048
    left ventricular ejection fraction 66.5% | 6048
    Modified Rankin Score of 2 | 6048
    no known medical illness | 0
    regular alcohol consumer | 0
    heavy alcohol consumer | 0
    lumberjack occupation | 0
    fever for 2 weeks | -336
    cough for 2 weeks | -336
    missing from work | -96
    confused state | 0
    septic shock | 0
    neck stiffness | 0
    normal limbs power | 0
    normal tone | 0
    normal reflexes | 0
    normal heart sounds | 0
    no murmur | 0
    bilateral lung crepitations | 0
    fluid resuscitation | 0
    vasopresssor | 0
    mechanical ventilator | 0
    ICU admission | 0
    anaemia | 0
    thrombocytopenia | 0
    normal white cells | 0
    normal renal function | 0
    splenic microabscesses | 0
    bilateral lung consolidation | 0
    normal CT brain | 0
    no inflammation in CSF | 0
    no infection in CSF | 0
    B. pseudomallei blood culture | 0
    ventilator-associated pneumonia | 72
    MDR A. baumanii | 192
    bacteraemia Day 6 | 144
    bacteraemia Day 12 | 288
    no growth Day 24 | 576
    no growth Day 26 | 624
    no growth Day 27 | 648
    left hemiplegia | 600
    pansystolic murmur | 600
    CT brain infarct | 600
    CT brain haemorrhage | 600
    echocardiogram vegetation | 600
    mitral regurgitation | 600
    supraventricular tachycardia | 168
    high temperature | 96
    leukopenia | 96
    started co-trimoxazole | 168
    IV imipenem | 96
    IV ampicilin-sulbactam | 336
    IV gentamicin | 168
    extended ceftazidime | 1008
    co-trimoxazole monotherapy | 2016
    discharged | 2016
    residual weakness | 2016
    Modified Rankin 2 | 2016
    daily activities independent | 2016
    intact cognition | 2016
    transferred | 2016
    follow-up 9 months | 6048
    resolved vegetation | 6048
    residual regurgitation | 6048
    LVEF 66.5% | 6048
    Modified Rankin 2 | 6048
    cerebral infarct | 600
    haemorrhages | 600
    septic emboli | 600
    infective endocarditis | 600
    mitral vegetation | 600
    gentamicin susceptibility | 0
    ceftazidime and gentamicin | 168
    co-trimoxazole continued | 2016
    residual weakness | 2016
    Rankin 2 | 2016
    activities independent | 2016
    intact cognition | 2016
    transfer to cardiac centre | 2016
    follow-up | 6048
    resolved vegetation | 6048
    residual regurgitation | 6048
    LVEF 66.5% | 6048
    Rankin 2 | 6048
    no medical history | 0
    alcohol use | 0
    lumberjack | 0
    fever 2 weeks | -336
    cough 2 weeks | -336
    missing work | -96
    confusion | 0
    septic shock | 0
    neck stiffness | 0
    normal limbs | 0
    normal tone | 0
    normal reflexes | 0
    heart sounds normal | 0
    no murmur | 0
    lung crepitations | 0
    fluid resuscitation | 0
    vasopresssor | 0
    ventilator | 0
    ICU | 0
    anaemia | 0
    thrombocytopenia | 0
    normal WBC | 0
    normal renal | 0
    splenic abscesses | 0
    lung consolidation | 0
    CT brain normal | 0
    CSF no inflammation | 0
    CSF no infection | 0
    B. pseudomallei culture | 0
    ventilator pneumonia | 72
    MDR A. baumanii | 192
    bacteraemia Day 6 | 144
    bacteraemia Day 12 | 288
    no growth Day 24 | 576
    no growth Day 26 | 624
    no growth Day 27 | 648
    hemiplegia | 600
    murmur | 600
    CT infarct | 600
    CT haemorrhage | 600
    echocardiogram vegetation | 600
    regurgitation | 600
    tachycardia | 168
    high temp | 96
    leukopenia | 96
    co-trimoxazole start | 168
    imipenem | 96
    ampicilin-sulbactam | 336
    gentamicin | 168
    extended ceftazidime | 1008
    co-trimoxazole mono | 2016
    discharge | 2016
    weakness residual | 2016
    Rankin 2 | 2016
    activities independent | 2016
    cognition intact | 2016
    transfer | 2016
    follow-up 9 months | 6048
    vegetation resolved | 6048
    regurgitation residual | 6048
    LVEF 66.5% | 6048
    Rankin 2 | 6048
    cerebral infarct | 600
    haemorrhages | 600
    emboli | 600
    endocarditis | 600
    mitral vegetation | 600
    gentamicin use | 168
    co-trimoxazole | 2016
    residual weakness | 2016
    Rankin 2 | 2016
    activities | 2016
    cognition | 2016
    transfer | 2016
    follow-up | 6048
    resolved vegetation | 6048
    regurgitation | 6048
    LVEF | 6048
    Rankin 2 | 6048
    no medical issues | 0
    alcohol regular | 0
    alcohol heavy | 0
    lumberjack | 0
    fever 2 weeks | -336
    cough 2 weeks | -336
    missing work days | -96
    confusion | 0
    septic shock | 0
    neck stiffness | 0
    limb power normal | 0
    tone normal | 0
    reflexes normal | 0
    heart normal | 0
    no murmur | 0
    lung sounds | 0
    fluid given | 0
    vasopresssor | 0
    ventilator | 0
    ICU | 0
    anaemia | 0
    thrombocytopenia | 0
    WBC normal | 0
    renal normal | 0
    spleen abscesses | 0
    lung consolidation | 0
    CT brain normal | 0
    CSF normal | 0
    B. pseudomallei positive | 0
    ventilator pneumonia | 72
    MDR A. baumanii | 192
    blood culture Day 6 | 144
    blood culture Day 12 | 288
    no growth Day 24 | 576
    no growth Day 26 | 624
    no growth Day 27 | 648
    hemiplegia | 600
    murmur | 600
    CT infarct | 600
    CT haemorrhage | 600
    echo vegetation | 600
    regurgitation | 600
    tachycardia | 168
    high temperature | 96
    leukopenia | 96
    co-trimoxazole start | 168
    imipenem | 96
    ampicilin-sulbactam | 336
    gentamicin | 168
    ceftazidime extended | 1008
    co-trimoxazole alone | 2016
    discharge | 2016
    weakness | 2016
    Rankin 2 | 2016
    daily activities | 2016
    cognition intact | 2016
    transfer | 2016
    follow-up | 6048
    vegetation gone | 6048
    regurgitation remains | 6048
    LVEF 66.5% | 6048
    Rankin 2 | 6048
    cerebral infarct | 600
    haemorrhages | 600
    emboli | 600
    endocarditis | 600
    vegetation | 600
    gentamicin | 168
    co-trimoxazole continued | 2016
    weakness | 2016
    Rankin 2 | 2016
    activities | 2016
    cognition | 2016
    transfer | 2016
    follow-up | 6048
    resolved | 6048
    regurgitation | 6048
    LVEF | 6048
    Rankin | 6048
    no medical problems | 0
    alcohol | 0
    job | 0
    fever | -336
    cough | -336
    missing | -96
    confused | 0
    septic shock | 0
    neck stiff | 0
    limbs normal | 0
    tone | 0
    reflexes | 0
    heart | 0
    no murmur | 0
    lungs | 0
    fluids | 0
    vasopresssor | 0
    ventilator | 0
    ICU | 0
    anaemia | 0
    low platelets | 0
    WBC | 0
    kidneys | 0
    spleen abscess | 0
    lung consolidation | 0
    CT brain | 0
    CSF | 0
    B. pseudomallei | 0
    ventilator pneumonia | 72
    MDR A.