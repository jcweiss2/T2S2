42 years old | 0
female | 0
Thai | 0
motorcycle accident | -12
left knee pain | -12
drowsiness | -12
subdural hematoma | -12
multiple shallow abrasion wounds | -12
pain at the lateral tibial plateau | -12
limited range of left knee motion | -12
combined tibial plateau fracture | -12
tibial tubercle avulsion | -12
long leg slab | -12
white blood cell count 19,490 /μL | -12
hematocrit 26.7% | -12
hemoglobin 8.6 g/dL | -12
polymorphonuclear neutrophils 85.5% | -12
lymphocytes 6.0% | -12
eosinophils 0.2% | -12
monocytes 8.2% | -12
platelets 336,000/μL | -12
admitted to intensive care unit | 0
close clinical observation | 0
open reduction and internal fixation | 120
locking plate | 120
cloudy fluid collection | 120
Staphylococcus aureus | 120
intravenous ceftriaxone | 120
intravenous clindamycin | 120
fever | 168
redness around the surgical wound | 168
sepsis investigation | 168
chest radiograph | 168
urine sample | 168
erythrocyte sedimentation rate more than 140 mm/h | 168
C-reactive protein more than 19.2 mg/dL | 168
irrigation and debridement | 192
necrotic tissue removal | 192
necrotic tissue culture | 192
Staphylococcus aureus | 192
hemoculture negative | 192
intravenous ceftriaxone and clindamycin | 192
oral Augmentin | 312
inflammatory markers disappeared | 432
able to walk without aid | 432
union of the left tibial plateau | 1056
plain radiograph | 1056