53 years old | 0
    male | 0
    admitted to the Emergency Department | 0
    sudden loss of vision in left eye | -120
    feeling unwell | -120
    shortness of breath | -120
    generalized body pains | -120
    fever | -120
    chills | -120
    denied headache | 0
    denied extremity weakness or numbness | 0
    denied chest pain | 0
    denied cough | 0
    denied abdominal pain | 0
    denied nausea | 0
    denied vomiting | 0
    chronic obstructive lung disease | -175200
    exploratory laparotomy | -105120
    gunshot wound | -105120
    tobacco smoking | 0
    active illicit IV drug use | 0
    temperature 36.8ºC | 0
    heart rate 92 bpm | 0
    blood pressure 91/55 mmHg | 0
    respiratory rate 18 breaths/min | 0
    oxygen saturation 92% | 0
    moderate respiratory distress | 0
    diffuse bilateral rhonchi | 0
    regular heart rate | 0
    regular rhythm | 0
    ejection murmur in tricuspid area | 0
    soft abdomen | 0
    nontender abdomen | 0
    left eye endophthalmitis | 0
    increasingly short of breath | 0
    hypotensive | 0
    intubated | 0
    fluid resuscitation | 0
    vasopressor therapy | 0
    vitreous tap | 0
    intravitreal vancomycin injection | 0
    intravitreal ceftazidime injection | 0
    empiric IV vancomycin | 0
    empiric IV cefepime | 0
    empiric moxifloxacin eye drops | 0
    elevated white blood cell count 28000/mm³ | 0
    hemoglobin 8.4 g/dL | 0
    platelet count 210000/mm³ | 0
    creatinine 1.45 mg/dL | 0
    urine drug screen positive for benzodiazepine | 0
    urine drug screen positive for opiates | 0
    blood cultures obtained | 0
    HIV nonreactive | 0
    chest X-ray left upper lobe reticulonodular infiltrates | 0
    chest X-ray prominent pulmonary arteries | 0
    chest X-ray coarse left basilar markings | 0
    chest X-ray coarse right upper lung zone markings | 0
    CT thorax multiple scattered cystic-like opacities | 0
    CT thorax consolidation | 0
    CT thorax suspicious for multifocal pneumonia | 0
    CT orbit minimal edema left preseptal soft tissues | 0
    CT orbit thickening left sclera | 0
    CT orbit intraconal fat stranding | 0
    CT orbit suspicious for preseptal cellulitis | 0
    CT orbit suspicious for postseptal cellulitis | 0
    transthoracic echocardiogram large vegetation tricuspid valve | 0
    transthoracic echocardiogram small vegetation septal leaflet | 0
    blood cultures positive for Serratia marcescens | 24
    switched to meropenem | 24
    switched to gentamicin | 24
    vancomycin continued | 24
    cardiothoracic surgeon consulted | 24
    tricuspid valve replacement | 48
    left upper lung abscess drainage | 48
    tricuspid valve vegetation | 48
    severe tricuspid regurgitation | 48
    Epic porcine tissue valve placed | 48
    tricuspid valve culture Serratia marcescens | 48
    lung abscess culture Serratia marcescens | 48
    dark red blood from nasogastric tube | 72
    low hemoglobin | 72
    suspected gastrointestinal bleeding | 72
    esophagogastroduodenoscopy esophagitis | 72
    clotted blood in stomach fundus | 72
    ischemic ulcers | 72
    septic emboli | 72
    hemoclips placed | 72
    critically ill in ICU | 96
    vitreous culture left eye Serratia marcescens | 96
    stable left eye | 96
    no hypopyon | 96
    switched to ciprofloxacin | 96
    discontinued vancomycin | 96
    continued meropenem | 96
    continued gentamicin | 96
    negative follow-up blood cultures | 192
    S. marcescens susceptible to ciprofloxacin | 192
    switched to IV ciprofloxacin | 192
    persistent chemosis | 192
    cloudy anterior chamber | 192
    possible infection progression | 192
    repeat CT orbit minimal preseptal swelling | 192
    repeat intravitreal ceftazidime | 192
    B-scan ultrasound increased vitreous debris | 336
    posterior hyaloid detachment | 336
    retinal detachment | 336
    small loculations | 336
    pars plana vitrectomy | 360
    subconjunctival pus | 360
    360-degree conjunctival peritomy | 360
    hazy lens | 360
    lens removed | 360
    sclera erosion | 360
    purulent intraocular drainage | 360
    vitreous biopsy | 360
    anterior chamber paracentesis | 360
    iris membrane removed | 360
    intravitreal vancomycin injection | 360
    intravitreal ceftazidime injection | 360
    posterior perforation | 360
    left eye enucleation | 456
    vitreous culture Serratia marcescens | 456
    left eye culture Serratia marcescens | 456
    continued meropenem | 0
    continued oral ciprofloxacin | 0
    discharged to nursing home | 840
    Staphylococcus aureus bacteremia | 4368
    continued IV drug use | 4368
    