45 years old | 0
male | 0
farmer | 0
admitted to the hospital | 0
shortness of breath | 0
altered sensorium | 0
inability to speak | 0
weakness of bilateral lower limbs | 0
snake bite | -48
swelling of the left leg | -48
anasarca | -48
anti-snake venom | -48
non-diabetic | 0
no history of hypertension | 0
no history of tuberculosis | 0
no history of chronic disease | 0
no melaena | 0
no bleeding manifestations | 0
history of smoking | 0
intake of alcohol | 0
minimally conscious | 0
reduced alertness | 0
non-cooperative | 0
disoriented | 0
blood pressure 106/60 mmHg | 0
cardiac rate 102 beats per minute | 0
respiratory rate 20 breaths per minute | 0
body temperature 37.2°C | 0
SpO2 91% | 0
bilateral crepitations | 0
pitting edema over the left foot | 0
non-tender | 0
raised temperature | 0
non-distinct impressions of two rows of teeth | 0
hemoglobin level 15 g/dl | 0
total leukocyte count 24.37×10^9/L | 0
neutrophils 89% | 0
lymphocytes 6% | 0
platelet count 19,000 per cubic millimeter | 0
blood urea 122 mg/dl | 0
serum creatinine 5.01 mg/dl | 0
serum sodium 117 mEq/L | 0
serum potassium 5.1 mEq/L | 0
no deep vein thrombosis | 0
bilateral mildly raised renal cortical echo-genicity | 0
coagulation profile normal | 0
PT 12.7 s | 0
INR 1.03 | 0
serum procalcitonin level 0.27 ng/ml | 0
normal left ventricular function | 0
bilateral multiple B lines | 0
interstitial pulmonary edema | 0
intubation | 0
transferred to ICU | 0
provisional diagnosis of snake bite with cellulitis | 0
sepsis | 0
acute kidney injury | 0
disseminated intravascular coagulation | 0
dual-antibiotic treatment | 0
piperacillin plus tazobactam | 0
clindamycin | 0
magnesium sulphate dressing | 0
random donor platelets | 0
continuous renal replacement therapy | 24
metoclopramide | 0
calcium polystyrene sulfonate | 0
glucose-insulin drip | 0
pantoprazole | 0
vitamin K | 0
magnesium sulphate | 0
conjugated estrogen | 0
condition worsened | 48
no reduction in swelling | 48
body temperature 37.8-38.9°C | 48
persistence of bilateral chest crepitations | 48
normal blood glucose levels | 48
total leukocyte count 31.65×10^9/L | 168
neutrophil 91% | 168
lymphocyte 7% | 168
Klebsiella pneumoniae | 192
tigecycline | 192
loading dose 100 mg | 192
maintenance dose 50 mg every 12 h | 192
improvement in condition | 216
reduction in swelling | 216
sharp fall in serum procalcitonin level | 216
normal body temperature | 216
hypoglycemic episode | 240
severe palpitations | 240
tremors | 240
sweating | 240
blood glucose level 47 mg/dl | 240
dextrose infusion | 240
relief of symptoms | 240
blood glucose level 83 mg/dl | 240
hypoglycemic episode | 264
blood glucose level 49 mg/dl | 264
hyperventilating | 264
profuse sweating | 264
palpitations | 264
dextrose infusion | 264
blood glucose level 86 mg/dl | 264
tigecycline stopped | 360
meropenem | 360
clindamycin | 360
polymyxin B | 360
no hypoglycemic episodes | 360
blood glucose levels below normal | 360
gradual rise in blood glucose levels | 408
condition improved | 456
reduction of swelling | 456
CRRT stopped | 456
serum creatinine normal | 456
urea levels normal | 456
electrolyte levels normal | 456
signs of sepsis reappeared | 648
Enterobacter spp. | 696
doxycycline | 696
minocycline | 696
tetracycline | 696
tigecycline | 696
loading dose 100 mg | 696
maintenance dose 50 mg every 12 h | 696
hypoglycemic attacks | 720
sweating | 720
palpitations | 720
blood glucose level 25 mg/dl | 720
dextrose infusion | 720
tigecycline discontinued | 744
minocycline | 744
cefoperazone plus sulbactam | 744
no hypoglycemic episodes | 744
blood glucose levels below normal | 744
gradual rise in blood glucose levels | 768
condition improved | 912
reduction of swelling | 912
reversal of sepsis | 912
discharged from ICU | 912