40 years old | 0
male | 0
admitted to the hospital | 0
severe diffuse abdominal pain | -8
abdominal bloating | -8
diarrhea | -8
nausea | -8
ruptured diverticulum | -120 months
acute diverticulitis | -24 months
acute diverticulitis | -12 months
mild periodic discomfort | -1 month
fever | 0
abdominal distension | 0
tenderness | 0
abdominal tenderness on deep palpation | 0
no stool in the vault | 0
temperature 38.8°C | 0
heart rate 120 beats/min | 0
normal blood pressure | 0
normal oxygen saturation | 0
hemoglobin 15.9 g/dl | 0
WBC 19.120 | 0
CRP 270.6 mg/l | 0
CPK 543 U/l | 0
GLU 125 mg/dl | 0
LDH 481 U/l | 0
fibrinogen 4.4 g/l | 0
Na 141 mEq/l | 0
K 5.2 mEq/l | 0
stenosis of the sigmoid colon | 0
marked dilation of the descending colon | 0
marked dilation of the transverse colon | 0
marked dilation of the ascending colon | 0
marked dilation of the cecum | 0
deterioration | 8
signs of sepsis | 8
multiorgan failure | 8
severe dyspnea | 8
metabolic acidosis | 8
intubation | 8
CRP 318 mg/l | 8
CPK 543 U/l | 8
fibrinogen 6 g/l | 8
creatinine 2.2 mg/dl | 8
PT 28.20 s | 8
INR 2.56 | 8
D-dimer 2,223.2 μg/l | 8
Na 133 mEq/l | 8
K 5.4 mmol/l | 8
P 5.4 mg% | 8
toxic megacolon | 8
surgical assessment | 8
emergency laparotomy | 8
extensive necrotic colon | 8
total colectomy | 8
protective loop ileostomy | 8
transfer to intensive care unit | 8
extubation | 20
transfer to ward | 20
discharge | 240
histological examination | 240
resolving necrotic colon | 240
no malignancy | 240
loop ileostomy reversal | 2160
good health | 4320