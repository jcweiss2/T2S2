56 years old | 0
male | 0
intermittent chest tightness | -168
shortness of breath | -168
chest tightness | -168
tremor of the hands | -24
loss of appetite | -24
general malaise | -24
loss of consciousness | -24
no history of alcohol consumption | 0
no history of drug abuse | 0
no history of high-risk behaviors causing PLA | 0
denies hypertension | 0
denies diabetes | 0
denies heart diseases | 0
no family history of hypertension | 0
no family history of diabetes | 0
no family history of heart diseases | 0
abdomen soft with right upper quadrant tenderness | 0
no rebound pain | 0
no muscle tension | 0
body temperature 39.2 °C | 0
blood pressure 98/56 mmHg | 0
heart rate 84 beats per min | 0
respiratory rate 26 breaths per min | 0
white blood cell count 22.22×109/L | 0
neutrophil percentage 91.7% | 0
platelet count 26 × 109/L | 0
pH 7.28 | 0
PCO2 27 mmHg | 0
PO2 64 mmHg | 0
HCO3- 12.7 mmol/L | 0
BE -12.5 mmol/L | 0
C-reactive protein level > 90 mg/L | 0
interleukin 6 > 5000 pg/mL | 0
procalcitonin > 100 ng/mL | 0
myoglobin > 2000 ug/L | 0
cranial CT showing thickened nasopharynx soft tissue | 0
thoracic CT showing bilateral pneumonia | 0
thoracic CT showing lung air sac in right lung apex | 0
thoracic CT showing multiple nodules in bilateral lungs | 0
thoracic CT showing bilateral pleural effusion | 0
abdominal and pelvic CT showing foci in right lobe of liver | 0
abdominal and pelvic CT showing mixed density in segment IV of liver | 0
needle-like high-density shadow in liver | 0
brown drainage from gastric tube | 0
history of eating fish before onset | 0
PLA caused by fishbone puncture | 0
severe pneumonia | 0
acute respiratory failure | 0
septic shock | 0
anti-inflammatory rescue therapy | 0
electrolyte correction | 0
nutritional support | 0
recurrent fever | 0
no significant decreases in inflammatory index | 0
repeat abdominal CT showing combined density | 0
laparoscopic exploration | 0
dense adhesions between pylorus and hepatic hilum | 0
liver swollen at ligamentum teres root | 0
fishbone found during operation | 0
abscess cavity incised | 0
white pus drained | 0
drainage tube placed | 0
small amount of reddish drainage fluid | 0
inflammatory indexes decreased | 120
symptoms and discomfort disappeared | 120
drainage tube removed | 120
discharged | 120
unremarkable follow-up at 2 weeks | 336
unremarkable follow-up at 2 months | 1440
