53 years old | 0
African American | 0
female | 0
coronary artery disease | 0
end-stage renal disease | 0
cervical carcinoma | 0
right atrial thrombus | 0
presented to emergency department | 0
bleeding profusely from rectum | 0
placement of two self-expanding nasal tampons | -24
transfusion of two units PRBCs | -24
MTP started | 0
administration of 2g tranexamic acid | 0
taken to operating room | 12
surgical efforts failed to control bleeding | 12
pelvic radiation therapy | -672
total colectomy | 12
proctoscopy | 12
massive blood from lower rectum/anal canal | 12
balloon tamponade with Penrose drain and Foley catheter | 12
TEG results: normal R time | 12
decreased alpha angle | 12
decreased maximum amplitude | 12
coagulopathy secondary to fibrinogen deficiency | 12
coagulopathy secondary to platelet deficiency | 12
administration of FFP | 12
administration of cryoprecipitate | 12
administration of platelets | 12
concern for apixaban-related coagulopathy | 12
consultation with interventional radiology | 18
transfer to SICU | 18
assembly of rapid transfuser devices | 18
insertion of wide-bore central venous catheter | 18
continued MTP | 18
goal MAP 50-60 mmHg | 18
administration of norepinephrine | 18
administration of vasopressin | 18
intermittent epinephrine boluses | 18
guided by vital signs | 18
guided by bedside echocardiography | 18
guided by serial TEG | 18
guided by serum lactate | 18
guided by base deficit | 18
blood loss >14L in 90 minutes | 18
identification of fistula between right common iliac and rectum | 24
placement of covered stent | 24
bleeding stopped | 24
administration of 60 units PRBC | 24
administration of 23 units FFP | 24
administration of 20 packs platelets | 24
administration of 6 units cryoprecipitate | 24
administration of 2g TXA | 24
administration of 30L crystalloid | 24
administration of 2L albumin | 24
serial FoCUS | 24
hypothermia improved | 24
serum lactate improved | 24
base deficit improved | 24
minimal ventilatory support | 24
closure of abdomen | 96
successful extubation | 96
transfer to floor | 96
no lung injury | 120
no volume overload | 120
no coagulopathy | 120
no cardiomyopathy | 120
