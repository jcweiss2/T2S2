66 years old | 0
female | 0
Hashimoto’s disease | -1920
pulmonary embolism | -1920
recurrent fever | 0
suspected connective tissue disease | 0
fever persisted | 0
admitted to the hospital | 0
antibiotic therapy | 0
pneumonia | 0
urinary tract inflammation | 0
human immunodeficiency virus excluded | 0
hepatitis C virus excluded | 0
cytomegalovirus excluded | 0
toxoplasmosis excluded | 0
Lyme disease excluded | 0
tuberculosis excluded | 0
bone marrow biopsy | 0
no evidence of proliferative disease | 0
diagnosis of SLE | 0
methylprednisolone 80 mg/day | 0
shortness of breath | 24
progressive decrease in blood pressure | 24
elevated procalcitonin serum concentration | 24
transferred to the Intensive Care Unit | 24
severe infection with risk of septic shock | 24
empirical antibiotic treatment | 24
glucocorticosteroid therapy | 24
atrial fibrillation | 24
amiodarone | 24
sinus rhythm | 24
re-hospitalized in the rheumatology department | 168
immunoglobulins infusions | 168
flaccid four-limb weakness | 168
dominant weakness of the left upper limb | 168
right lower limb weakness | 168
brain imaging by magnetic resonance imaging | 168
no abnormalities found | 168
episode of unconsciousness | 168
left eye turning | 168
hypotension | 168
transthoracic echocardiography | 168
computed tomography of coronary arteries | 168
no significant deviations found | 168
electroencephalography recording | 168
no irritation changes typical for epilepsy | 168
electromyography | 168
generalized axonal damage of peripheral nerve motor fibers | 168
F wave disturbance from the right median nerve | 168
limit values of conduction in sensory fibers of the right ulnar nerve | 168
depletion of exercise recording | 168
increased percentage of polyphasia | 168
critical illness polyneuropathy suspected | 168
follow-up EMG | 672
intensification of the lesions | 672
acute axonal polyneuropathy | 672
significant predominance of lesions in the nerves of the lower extremities | 672
acute denervation | 672
methotrexate 15 mg/week | 672
hydroxychloroquine planned | 672
low molecular weight heparin | 672
transferred to the department of rehabilitation | 672
generalized weakness of trunk and limb muscle strength | 672
tetraparesis | 672
left upper limb dominance | 672
global paresis of the lower limbs | 672
abolition of tendon reflexes in the limbs | 672
lower limb allodynia | 672
pregabalin | 672
comprehensive improvement program | 672
gradual verticalization | 672
increase of muscular strength | 672
isometric exercises | 672
learning to change position in the bed | 672
coordination exercises | 672
improvement in muscle strength | 672
functional status improvement | 672
independent bed position changes | 1512
walker-assisted walking | 1512
next cycle of rehabilitation | 2520
gait improvement | 2520
high support walking | 2520
stairs walking | 2520
rising after a fall | 2520
left shoulder strengthening | 2520
range of mobility improvement | 2520
significant functional improvement | 2520
discharge | 3024
short distance walking | 3024
two-wheel support walking | 3024
Barthel Index improvement | 3024
