67 years old | 0
African-American | 0
male | 0
admitted to the hospital | 0
achy, non-radiating pain in chest | -72
acute left foot pain | -72
fatigue | -72
malaise | -72
nausea | 0
vomiting | 0
sweating | 0
ESRD | -6480
hemodialysis | -2628
non-ischemic heart failure | -0
pericardial effusion | -0
low-grade follicular cell lymphoma | -0
stroke | -0
DVT | -0
pulmonary embolism | -0
paroxysmal atrial fibrillation | -0
COPD | -0
hepatitis C infection | -0
chronic anemia | -0
medication non-adherence | -0
multiple dialysis catheter placements | -0
AV fistula creation | -0
atrial flutter ablation | -0
hernia repair | -0
elevated troponin | 0
WBC count | 0
neutrophils | 0
ECG | 0
nuclear stress test | 72
LV ejection fraction | 72
perfusion defect | 72
ischemic changes | 72
low-grade fever | 24
blood cultures | 24
gram-positive rods | 24
diphtheroid | 24
endocarditis | 0
transthoracic echocardiogram | 0
mitral valve vegetation | 0
severe mitral annular calcification | 0
moderate mitral regurgitation | 0
mild mitral stenosis | 0
aortic valve leaflets | 0
mild to moderate tricuspid regurgitation | 0
vancomycin | 0
femoral permcath replacement | 0
Corynebacterium jeikeium | 0
resistant to penicillin | 0
resistant to ceftriaxone | 0
resistant to meropenem | 0
sensitive to vancomycin | 0
repeated blood cultures | 72
positive for diphtheroid | 72
new femoral permcath | 216
discharged | 216
Corynebacterium jeikeium endocarditis | 216
vancomycin | 216
dialysis session | 216
recovered | 432
dialysis catheter malfunction | 432
no follow-up | 432