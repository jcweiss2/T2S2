18 years old | 0
male | 0
shortness of breath | -8
severe right-sided chest pain | -8
fever | -336
sore throat | -336
dysphagia | -336
fatigue | -336
admitted to hospital | -144
Penicillin V | -144
discharged after 24 h observation | -144
IM confirmed | 0
EBV specific antibodies detected | 0
right chest pain | 0
tenderness |,0
dyspnoeic | 0
respiratory rate of 30 breaths per minute | 0
peripheral oxygen saturations of 94% | 0
temperature 37.4°C | 0
pulse rate 120 beats per minute | 0
blood pressure 100/70 mmHg | 0
bilateral symmetrical tonsillar swelling | 0
white exudate | 0
bilateral cervical lymphadenopathy | 0
leucocytosis | 0
elevated C-reactive protein | 0
elevated liver enzymes | 0
computed tomography imaging | 0
extensive pneumomediastinum | 0
mediastinal fat stranding | 0
pockets of fluid in the anterior mediastinum | 0
small right pleural effusion | 0
inflammatory consolidation in the right lung | 0
reactive lymph nodes | 0
splenomegaly | 0
enlarged lymphoid tissue in the posterior nasopharynx | 0
no evidence of oesophageal perforation | 0
no peritonsillar abscess | 0
no retropharyngeal abscess | 0
IV opioid analgesia | 0
fluid resuscitation | 0
amoxicillin | 0
clavulanic acid | 0
cardiothoracic surgery consultation | 0
deterioration | 4
increased chest pain | 4
worsening physiology | 4
antibiotics changed to IV Piperacillin | 4
tazobactam | 4
clindamycin | 4
video-assisted thoracoscopic surgery | 4
drainage and decortication of right pleural empyema | 4
drainage of multiple mediastinal abscesses | 4
debridement of mediastinal necrotic tissue | 4
insertion of right-sided intercostal drain | 4
Fusobacterium necrophorum detected | 4
Dialister pneumosintes detected | 4
Peptostreptococcus anaerobius detected | 4
admitted to intensive care unit | 4
22-day period in hospital | 528
14 days of intensive care | 336
discharged home well | 528
