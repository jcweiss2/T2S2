65 years old | 0
female | 0
rheumatic valve disease | -8760
surgical mitral valve repair | -8760
percutaneous exchange of the mitral valve | -240
dyspnea on the slightest effort | -720
paroxysmal nocturnal dyspnea | -720
orthopnea | -720
dry cough | -720
fever | -720
treated for dengue fever | -960
admitted to the hospital | 0
paroxysmal atrial flutter | 240
decreased level of consciousness | 240
anisocoric pupils | 240
referred to the intensive care unit | 240
drowsy | 240
pale | 240
hydrated | 240
acyanotic | 240
afebrile | 240
arterial blood pressure 122/73 mm Hg | 240
heart rate 96 beats per minute | 240
respiratory rate 14 breaths per minute | 240
heart auscultation normal | 240
murmurs absent | 240
respiratory auscultation normal | 240
abdomen examination normal | 240
mild edema in the lower limbs | 240
hemoglobin 8.5 g/dL | 240
hematocrit 25% | 240
white blood cells 16,200/mm3 | 240
platelets 192,000/mm3 | 240
mild anisocytosis and microcytosis | 240
urea 67 mg/dL | 240
creatinine 2.39 mg/dL | 240
sodium 132 mmol/L | 240
potassium 3.6 mmol/L | 240
C reactive protein 11.2 mg/dL | 240
APACHE II score 22 | 240
SAPS III score 64 | 240
dental evaluation indicated precarious dentition | 240
blood culture samples collected | 240
empirical treatment with ceftriaxone associated with gentamicin | 240
transesophageal echocardiogram | 240
vegetation in the ventricular face of the anterior mitral valve leaflet | 240
sensitive conduction aphasia | 480
mild right central paralysis | 480
ischemic stroke suspected | 480
brain tomography | 480
hypodense left insular lobe | 480
mechanical thrombectomy indicated | 480
arteriogram | 480
failed partial filling of the parietal branch of the left middle cerebral artery | 480
worsened level of consciousness | 720
hemodynamic instability | 720
need for hemodialysis | 720
orotracheal intubation | 720
vasoactive drugs initiated | 720
brain edema in the posterior circulation region | 720
hypodensity in the left thalamus | 720
septic shock | 720
refractory to therapeutic measures | 720
death | 720
Haemophilus parainfluenzae grew in the four blood culture samples | 720
blood culture conducted in diffusion discs | 720
microorganism sensitive to all the tested B-lactamic compounds | 720