69 years old | 0
woman | 0
stabbed herself in the abdomen with a kitchen knife | 0
suicidal intent | 0
admitted to emergency department | 0
blood pressure could not be measured | 0
pulseless electrical activity | 0
body temperature 35.0 °C | 0
oxygen saturation 99% | 0
Glasgow Coma Scale score of 3 | 0
agonal respiration | 0
5 cm wound on upper abdomen | 0
intra-abdominal fluid collection | 0
emergency thoracotomy | 0
aortic cross-clamping | 0
open cardiac massage | 0
aorta clamped for 15 min | 0
epinephrine administered thrice | 0
temporary return of spontaneous circulation | 0
hemodynamically unstable | 0
laparotomy performed | 0
injuries to common hepatic artery | 0
injuries to splenic artery | 0
injuries to pancreas | 0
injuries to spleen | 0
injuries to liver | 0
ligation of injured arteries | 0
left gastric artery not identified | 0
branch arising directly from aorta injured | 0
ligation on branch | 0
distal pancreatectomy | 0
splenectomy | 0
liver sutured | 0
norepinephrine administered | 0
second-look surgery | 24
no active bleeding | 24
no ischemic change | 24
hospital day 3 | 72
no vasopressor requirement | 72
abdominal wall closure | 72
regular examinations | 72
enhanced CT scan on hospital day 4 | 96
disruption of celiac artery | 96
gastroduodenal artery arising from superior mesenteric artery | 96
right gastric arteries not observed | 96
left gastroepiploic arteries not observed | 96
right gastroepiploic arteries not observed | 96
short gastric arteries not observed | 96
gastroscopy on hospital day 9 | 216
patchy mucosal necrosis on gastric upper body | 216
conservative treatment administered | 216
no significant change after 2 weeks | 216
hospital day 23 | 552
fever 39 °C | 552
pain in the stomach | 552
white blood cell count 34,000/mm³ | 552
C reactive protein 13.4 mg/dL | 552
CT scan demonstrating air in gastric wall | 552
intra-abdominal free air | 552
gastric necrosis suspected | 552
gastroscopy revealing extensive mucosal necrosis | 552
emergency surgery | 552
necrosis of stomach | 552
total gastrectomy | 552
Roux-en-Y reconstruction | 552
histological findings of stomach | 552
diffuse necrotic changes | 552
inflammatory cell infiltrations | 552
no evidence of invasive fungal infection | 552
leakage on duodenal stump | 696
continuous tube drainage | 696
consciousness became clear | 696
rehabilitation in bed | 696
sepsis due to Pseudomonas aeruginosa infection | 1680
disseminated intravascular coagulation | 1680
general condition gradually deteriorated | 1680
died 70 days after admission | 1680
