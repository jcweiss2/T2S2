2 years old | 0
male | 0
admitted to the hospital | 0
collapse | -1
unresponsive | -1
persistently alerted level of conscious | 0
normal vital signs | 0
dual heart sounds | 0
clear chest | 0
soft and nontender abdomen | 0
generalized poor tone | 0
no neurological deficits | 0
no significant medical or antenatal history | 0
no regular medications | 0
not recently been unwell | 0
commenced on intravenous ceftriaxone | 0
commenced on aciclovir | 0
mild neutrophilia | 0
hypokalaemia | 0
metabolic acidosis | 0
level of consciousness improved | 12
transferred to tertiary center | 12
dysmetria | 12
dysphagia | 12
deranged coagulation profile | 12
international-normalized ratio of 1.7 | 12
activated-partial thromboplastin time of 62 | 12
fibrinogen level of 0.9 | 12
blood cultures taken | 12
infectious serology taken | 12
autoimmune and vasculitic screen taken | 12
lumbar puncture taken | 12
possible bite mark on the lip | 12
serum samples for snake venom-specific enzyme immunoassay taken | 12
acute respiratory distress | 24
transferred to pediatric intensive care unit | 24
encephalopathic | 24
intubated | 24
ventilated | 24
given cryoprecipitate | 24
continued on aciclovir | 24
continued on ceftriaxone | 24
commenced on methylprednisolone | 24
echocardiogram performed | 24
echocardiogram normal | 24
MRI with contrast of the brain | 48
multiple supra and infratentorial anterior and posterior circulation infarcts | 48
no associated hemorrhage | 48
managed conservatively | 72
antibiotics ceased | 72
antivirals ceased | 72
corticosteroids ceased | 72
extubated | 72
specialized testing of blood sample returned positive result for Eastern Brown snake venom | 72
returned to pediatrics ward | 72
dysmetria resolved | 96
dysphagia resolved | 96
discharged | 96
received ongoing rehabilitation | 96
received physical therapy | 96
received occupational therapy | 96
made a good recovery | 168
meeting all developmental milestones | -672 
bite by an Australian Eastern Brown snake | -1