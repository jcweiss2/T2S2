68 years old | 0
male | 0
transferred from another institution | 0
progressively worsening tachypnea | -720
increased fraction of inspired oxygen (FIO2) requirements | -720
endotracheal intubation | -720
initiation of mechanical ventilation | -720
morbid obesity | 0
systemic arterial hypertension | 0
diabetes mellitus | 0
chronic lung disease | 0
heavy smoking history | 0
ramipril | 0
amlodipine | 0
metformin | 0
metoprolol | 0
no recent or remote exposure to corticosteroids therapy | 0
no recent or remote exposure to immunosuppressive agents | 0
blood pressure 86/52 mm Hg | 0
mean arterial pressure 63 | 0
heart rate 104 beats/min | 0
respiratory rate 24 breaths/min | 0
temperature 37 °C | 0
bilateral rales | 0
wheezing | 0
white blood cell (WBC) count 16.4 × 103/mm3 | 0
alanine aminotransferase (ALT) level 119 U/L | 0
lactate dehydrogenase (LDH) level 488 U/L | 0
blood urea nitrogen (BUN) level 36 mg/DL | 0
creatinine level within normal limits | 0
cardiac enzymes within normal limits | 0
coagulation profile within normal limits | 0
HIV test negative | 0
arterial blood gas (ABG) pH 7.24 | 0
pCO2 level 69 mm Hg | 0
PaO2 level 67 mm Hg | 0
initial chest X-ray bilateral increased interstitial markings | 0
left retrocardiac consolidation | 0
chest computed tomography (CT) bilateral ground-glass opacities | 0
no evidence of pulmonary embolism | 0
venous Doppler ultrasound no evidence of deep venous thrombosis | 0
electrocardiogram (ECG) sinus tachycardia | 0
no ST-segment abnormalities | 0
no T-wave abnormalities | 0
transthoracic echocardiogram (TTE) normal left ventricular ejection fraction | 0
normal right ventricular systolic function | 0
no evidence of pulmonary hypertension | 0
admitted to intensive care unit (ICU) | 0
empiric intravenous antimicrobial therapy vancomycin | 0
empiric intravenous antimicrobial therapy cefepime | 0
empiric intravenous antimicrobial therapy azithromycin | 0
vasopressors norepinephrine continuous infusion | 0
presumptive septic shock | 0
severe community-acquired pneumonia (CAP) | 0
blood cultures negative | 0
respiratory cultures negative | 0
Legionella urinary antigen negative | 0
Streptococcus pneumoniae urinary antigen negative | 0
serum cryptococcal antigen negative | 0
antimicrobials discontinued after 7 days | 168
procalcitonin level 0.25 ng/mL | 0
(1-3)-β-D-glucan assay 32 pg/mL | 0
increased FIO2/PEEP requirements | 0
ARDS | 0
decreased PaO2/FIO2 ratio | 0
worsening bilateral infiltrates on CXR | 0
increased vasopressors requirements | 0
acute kidney injury | 0
optimal sedation achieved | 0
analgesia achieved | 0
fentanyl continuous infusion | 0
propofol continuous infusion | 0
neuromuscular blocking agent (cisatracurium) infusion initiated | 0
epoprostenol added | 0
extracorporeal membrane oxygenation (ECMO) therapy deemed inappropriate | 0
plateau pressures < 35 cm H2O | 0
BAL positive for Pneumocystis jirovecii DNA | 0
CMV antigenemia negative | 0
serum immunoglobulin levels within normal limits | 0
complement component 3 (C3) diminished | 0
complement component 4 (C4) diminished | 0
CH50 levels diminished | 0
repeated HIV test non-reactive | 0
T-lymphocytes cell count (CD4) 97 cells/µL | 0
absolute lymphocytes cell count 377 × 103/µL | 0
intravenous antimicrobial therapy trimethoprim-sulfamethoxazole initiated | 0
steroids methylprednisone initiated | 0
repeated chest CT diffuse ground-glass opacities | 0
severe pneumomediastinum | 0
pneumopericardium | 0
bilateral pneumothorax | 0
clinical condition worsening | 0
withdrawal of artificial life support | 336
patient expired | 336
