Here is the table of events and timestamps:

age 43 | 0
female | 0
history of difficult-to-manage bronchial asthma | 0
hospitalized in the last 8 months | 0
asthmatic crisis | 0
24-hour history of dry cough | -24
progressive dyspnea | -24
psychomotor agitation | -24
audible wheezing | -24
salbutamol and ipratropium bromide | -24
diaphoretic | -24
tachycardic | -24
dyspneic | -24
supraclavicular retractions | -24
respiratory rate of 30 breaths/minute | -24
ambient oxygen saturation 87% | -24
auscultation with abolished vesicular murmur in both lung fields | -24
Glasgow coma scale (GCS) 12/15 | -24
arterial blood gases (ABG) analysis | -24
respiratory acidosis | -24
hypoxemia | -24
invasive ventilatory support | -24
midazolam | -24
propofol | -24
hydrocortisone 100 mg IV every 8 hours | -24
magnesium sulfate | -24
antibiotics (piperacillin tazobactam and clarithromycin) | -24
sepsis and/or shock | -24
multiple organ failure | -24
metabolic variables such as hyperglycemia | -24
duration of mechanical ventilation | -24
deep sedation | -24
neuromuscular blocking agents (NMB) | -48
cisatracurium | -48
ventilatory weaning | -48
dexmedetomidine | -48
improvement in ABG | -48
GCS 15/15 | -48
weakness of the neck flexor muscles | -48
facial paresis | -48
could not move all 4 limbs | -48
muscular strength 1/5 in lower limbs | -48
muscular strength 2/5 in upper limbs | -48
flaccid hyporeflexia | -48
preserved sensitivity | -48
brain and cervical MRI | -48
cerebrospinal fluid study | -48
EMG | -48
signs of denervation and irritability | -48
myopathic pattern | -48
polyneuropathic compromise | -48
axonal pattern in conduction velocity | -48
diagnosis of ICUAW | -48
physiotherapy and comprehensive rehabilitation | -48
ventilator was withdrawn | -10
MRC score of 55 points | -10
normal ABG control | -10
symptomatic resolution | -10
symptomatic resolution was achieved | -10