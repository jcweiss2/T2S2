42 years old | 0
male | 0
admitted to the hospital | 0
acute kidney injury | 0
dyspnea | 0
swelling in the face | -8760
swelling in the upper arms | -8760
HAE suspected | 0
C4 level low | 0
C1-INH level low | 0
high doses of androgen therapy | -672
Danazol | -672
kidney injury worsened | -168
chronic kidney disease | -168
kidney transplant surgery | 0
hemodialysis | -168
C1-INH level low | -7
FFP administered | -1
surgery | 0
anesthesia induced | 0
intubation | 0
mechanical ventilation | 0
surgery ended | 4
neuromuscular blockade reversed | 4
extubation | 4
immunosuppressants administered | 4
ganciclovir administered | 4
prostaglandin E1 administered | 4
vital signs stable | 4
urine output | 4
hemoglobin level | 5
coagulation tests | 5
dyspnea | 24
abdominal discomfort | 24
hypotension | 24
tachycardia | 24
loss of consciousness | 24
intubation | 24
mechanical ventilation | 24
norepinephrine administered | 24
dobutamine administered | 24
abdominal distension | 24
massive serosanguineous fluids | 24
generalized edema | 24
low urine output | 24
low hemoglobin level | 24
coagulopathy | 24
DIC diagnosed | 24
transfusion | 24
CRRT | 24
second-look operation | 48
no anastomosis leakage | 48
normal blood flow to kidney | 48
severe generalized edema | 48
hypoalbuminemia | 48
C1-INH level increased | 48
albumin administered | 48
danazol administered | 48
FFP transfusions | 48
pulmonary edema | 96
pneumonia | 96
rejection of transplanted kidney | 96
severe hypotension | 96
death | 120