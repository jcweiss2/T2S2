78 years old | 0
    male | 0
    admitted to the Department of Ophthalmology | 0
    current smoker | 0
    hypertension | -26304
    hyperlipidemia | -26304
    nifedipine | -26304
    candesartan | -26304
    atorvastatin | -26304
    doxazosin | -26304
    sarpogrelate | -26304
    levofloxacin eye drops started | 0
    cataract surgery | 0
    fever | 72
    dyspnea | 72
    no change in surgical sites | 72
    cefcapene pivoxil | 72
    hypoxia | 72
    oliguria | 72
    neutrophilia | 72
    elevation of C-reactive protein | 72
    impairment of liver function | 72
    impairment of kidney function | 72
    chest X-ray showed bilateral non-segmental consolidation | 72
    CT showed bilateral non-segmental consolidation | 72
    thickening of the bronchovascular bundles | 72
    pleural effusion | 72
    no abnormal findings in electrocardiogram | 72
    no abnormal findings in ultrasound cardiography | 72
    differential diagnosis considered | 72
    continuous hemodiafiltration | 72
    tazobactam/piperacillin started | 72
    ventilatory support | 72
    renal function improved | 72
    respiratory failure prolonged | 72
    fever prolonged | 72
    meropenem started | 72
    increase in airway pressure | 72
    wheezes developed | 72
    corticosteroid treatment | 72
    microbial examinations negative | 72
    autoantibody tests negative | 72
    bronchoalveolar lavage fluid obtained | 240
    lymphocytes increased | 240
    eosinophils increased | 240
    diagnosis of drug-induced lung injury | 240
    nicardipine hydrochloride stopped | 240
    sivelestat sodium stopped | 240
    levofloxacin injection started | 240
    respiratory condition worsened | 240
    liver dysfunction re-emerged | 240
    levofloxacin injections stopped | 240
    steroid therapy administered | 240
    respiratory failure improved | 240
    liver dysfunction improved | 240
    fever continued | 240
    levofloxacin eye drops continued | 240
    levofloxacin eye drops discontinued | 240
    fever resolved | 528
    respiratory failure resolved | 528
    extubated | 528
    drug lymphocyte stimulation test positive for levofloxacin | 528
    discharged | 1368
    steroid therapy continued | 1368
    no recurrence | 1368
