47 years old | 0
female | 0
26-pack-year history of cigarette smoking | 0
10-year history of consumption of more than 1 glass of alcohol per day | 0
untreated chronic psoriasis vulgaris | 0
found unconscious | 0
previously treated with meropenem | -48
intravenous infusion of 1 g meropenem every 12 hours for 2 days | -48
interhospital transfer to OMFS Clinic | 0
evaluation and treatment of extensive infection of occipital excoriated psoriatic plaque |6 0
normal temperature | 0
tachypnea | 0
tachycardia | 0
hypotension | 0
tumefaction in the right area of face and neck | 0
bilateral palpebral microabscesses | 0
large occipital psoriatic plaque | 0
massive crepitations in the occipital and posterior cervical regions | 0
emergency surgery | 1
wide posterior cervical incision | 1
right submandibular incision | 1
extensive necrosis | 1
wide excision | 1
sterile dressing | 1
extensive washing with oxygenated water and povidone-iodine solution | 1
postoperative contrast-enhanced computed tomography scan | 1
empirical antibiotic therapy | 1
limited right lateral cervical and supraclavicular necrectomy | 72
leukocytosis | 72
fever 38.8°C | 72
bacteriological wound drainage and drug sensitivity testing | 144
Staphylococcus epidermidis | 144
Klebsiella sp. | 144
Acinetobacter sp. | 144
sensitivity limited to colistin | 144
treatment with colistin | 144
previous antibiotics continued | 144
entire face became edematous | 168
necrectomy of the entire epicranial galea | 168
necrectomy of the right temporal fascia | 168
clean wounds with granulation tissue | 1080
denuded skull bone | 1080
plastic reconstruction with flaps and grafts | 1080
transferred to Plastic Surgery Department | 1080
discharged | 1824
no hyperbaric oxygen therapy | 0
