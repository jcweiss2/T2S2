36 years old | 0
male | 0
no pathological history of interest | 0
admitted to the outpatient clinic | 0
swallowing difficulties | -72
plain chest radiography with a water soluble contrast swallow | -72
PPI therapy | -72
six food elimination diet | -72
noncompliant for follow-up | -72
presented to the emergency department | 0
swallowing complaints | 0
EFBI | 0
plain chest radiography with a water soluble contrast swallow | 0
gastroscopy | 0
food bolus impaction | 0
subcutaneous emphysema | 0
thoracic computer tomography | 0
pneumomediastinum | 0
esophageal perforation | 0
febrile | 0
chest pain | 0
no emphysema | 0
auscultatory bilateral soft rough breathing sounds | 0
hemodynamically stable | 0
blood pressure 140/90mmHg | 0
arterial pulse 85bpm | 0
oxygen saturation 98% | 0
increased inflammatory markers | 0
mild eosinophilia | 0
plain chest radiography with a water soluble contrast swallow | 0
esophageal stricture | 0
esophageal food bolus impaction | 0
esophageal perforation | 0
transhiatal esophagectomy | 24
cervical esophagostomy | 24
pyloromyotomy | 24
feeding jejunostomy | 24
histologic examination | 24
eosinophilic esophagitis | 24
eosinophilic gastritis | 24
postoperative period | 24
nutritional support | 24
imagistic control | 24
blood tests survey | 24
control contrast study | 48
jejunostomy tube | 48
Nutrison Advanced Peptisorb | 48
abdominal discomfort | 48
discharged | 240
hypoalbuminemia | 720
poor enteral nutrition | 720
cervical esophagogastrostomy | 8760
gastric pull-up | 8760
postoperative period | 8760
anastomotic integrity | 8784
contrast imaging study | 8784
clear fluids | 8784
oral administration | 8784
enteral tube feeding | 8784
full fluid consistency | 8784
discharged | 8928
follow-up | 17520
correct oral nutrition | 17520
no episodes of swallowing disorders | 17520
no dysphagia | 17520
no EFBI | 17520
no malabsorption syndrome | 17520