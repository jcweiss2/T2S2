49 years old | 0
female | 0
upper respiratory tract infection | -48
rhinorrhea | -48
cough | -48
fever | -48
lethargy | -48
fatigue | -48
loss of appetite | -48
dehydrated | -48
reduced urine output | -48
syncopal attack | -72
nausea | -72
vomiting | -72
admitted to hospital | 0
no detectable pulse | 0
no measurable blood pressure | 0
blueish extremities | 0
brief intermittent episodes of syncope | 0
fully awake and mentally coherent | 0
intravenous Ringer’s solution | 0
hypotension | 0
hemoconcentration | 0
hypoalbuminemia | 0
generalized edema | 0
increased white blood cell count | 0
neutrophilia | 0
elevated creatinine | 0
elevated serum glutamic oxaloacetic transaminase | 0
elevated creatinine kinase | 0
elevated C-reactive protein | 0
low albumin | 0
fasciotomy | 5
pleural effusions | 24
retropharyngeal edema | 24
necrotic areas in leg muscles | 48
elevated creatine kinase | 96
anemia | 120
transfusion | 120
discharged from hospital | 720
rehabilitation | 720
orthopedic support for walking | 720
weakness | 720
reduced quality of life | 720
frequent upper respiratory tract infections | 720
monoclonal gammopathy | 0
IgG-kappa paraprotein | 0
low IgG | 0
low IgA | 0
normal IgM | 0
low mannose-binding lectin | 0
family history of monoclonal gammopathy | 0
family history of cardiovascular disease | 0
family history of cancer | 0
family history of diabetes | 0
intravenous immunoglobulin | 120
terbutaline | 720
theophylline | 720
appendicitis | -604800
sepsis | -604800
urinary tract infections | -604800
cystitis | -604800
pyelonephritis | -604800
premature birth | -1411200
toxemia | -1411200
Rhesus incompatibility | -1411200
exchange transfusion | -1411200
increased blood glucose during pregnancy | -1411200
fasciotomy #2 | 24
furosemide | 12
IVIG treatment | 120
SAG | 264
normal complement levels | 8760
low mannose-binding lectin | 8760
normal lectin activation pathway | 8760
normal alternative activation pathway | 8760
normal classic activation pathway | 8760