74 years old | 0
female | 0
ulcerative colitis | -17280
colectomy | -17280
ileostomy | -17280
hypertension | -17280
presented to the emergency department | 0
fatigue | 0
myalgia | 0
confusion | 0
temperature of 100°F | 0
blood pressure of 108/60 mmHg | 0
heart rate of 106 bpm | 0
respiratory rate of 20 breaths per minute | 0
disoriented to the surrounding environment | 0
unremarkable neurologic examination | 0
normal S1 and S2 without murmurs | 0
decreased breath sounds on lung bases | 0
sodium of 128 mEq/L | 0
creatinine of 1.21 mg/dL | 0
elevated lactate at 3.0 mEq/L | 0
urinary tract infection | 0
white blood cell count of 8.8 k/cmm | 0
hemoglobin of 15.1 g/dL | 0
platelet count of 131 k/cmm | 0
unremarkable CT of the brain | 0
unremarkable chest X-ray | 0
resuscitated with intravenous fluid | 0
started on IV ceftriaxone | 0
admitted for treatment of sepsis | 0
discharged after 3 days | 72
improvement of mentation to baseline | 72
resolution of acute kidney injury | 72
resolution of hyponatremia | 72
resolution of lactic acidosis | 72
returned to the ED | 72
significant weakness | 72
inability to ambulate | 72
elevated temperature of 103°F | 72
heart rate of 115 bpm | 72
blood pressure of 90/65 mmHg | 72
respiratory rate of 24 breaths per minute | 72
normal mental status | 72
white blood cell count of 3.31 k/cmm | 72
hemoglobin of 13.2 g/dL | 72
platelet count of 60 k/cmm | 72
lactic acid of 5.4 mEq/L | 72
AST of 237 U/L | 72
ALT of 189 U/L | 72
alkaline phosphatase of 146 U/L | 72
right middle lobe infiltrates | 72
started on vancomycin | 72
started on piperacillin-tazobactam | 72
admitted to the medical floor | 72
developed worsening respiratory status | 96
requiring noninvasive mechanical ventilation | 96
transferred to the medical intensive care unit | 96
bilateral pleural effusions | 96
thoracentesis | 96
removal of 750cc of exudative fluid | 96
progressively hypoxemic | 96
bilateral interstitial infiltrates consistent with ARDS | 96
required intubation | 96
fever persisted | 96
continuous decline in her state | 96
negative blood cultures | 96
negative sputum cultures | 96
negative urine cultures | 96
negative stool cultures | 96
white blood cell count of 1.4 k/cmm | 96
hemoglobin of 8.5 g/dL | 96
platelet count of 45 k/cmm | 96
worsening kidney function tests | 96
creatinine of 2.1 mg/dL | 96
BUN of 65 mg/dL | 96
worsening liver transaminases | 96
jaundice worsened | 96
coagulopathy | 96
elevated INR at 8 | 96
acute liver injury | 96
normal Factor V activity | 96
normal Factor VIII activity | 96
ruled out DIC | 96
unremarkable abdominal ultrasound | 96
unremarkable MRI of the liver | 96
unremarkable MRI of the pancreas | 96
elevated LDH at 1367 U/L | 96
elevated triglycerides at 808 mg/dL | 96
fibrinogen of 240 mg/dL | 96
elevated ferritin at 40,000 ng/mL | 96
suspected secondary HLH | 96
bone marrow biopsy | 96
normocellular marrow with myeloid predominance | 96
mild granulocyte atypia | 96
increased histiocytes | 96
CD163 immunostaining showed increased histiocytes | 96
hemophagocytosis consistent with HLH | 96
started on dexamethasone | 96
started on etoposide | 96
improvement of clinical status | 96
improvement of cell counts | 96
improvement of liver functions | 96
negative viral serologies | 96
negative HIV | 96
negative CMV | 96
negative HSV type 1 | 96
negative HSV type 2 | 96
negative EBV | 96
negative hepatitis B virus | 96
negative hepatitis C virus | 96
negative antinuclear antibody | 96
negative double-stranded DNA antibody | 96
negative rheumatoid factor | 96
negative autoimmune hepatitis workup | 96
ruled out hereditary hemochromatosis | 96
diagnosed with HLH | 96
met 5 out of 8 HLH-2004 criteria | 96
fever | 96
cytopenia of 2 cell lines | 96
elevated ferritin >500 ng/mL | 96
elevated fasting triglyceride >265 mg/dL | 96
hemophagocytosis in bone marrow | 96
improved respiratory status | 96
weaned off mechanical ventilation | 96
normalization of liver enzymes | 96
readmitted to the hospital | 672
persistent confusion | 672
diagnosed with HLH with central nervous system involvement | 672
worsening cognitive impairment | 672
increased protein level on cerebrospinal fluid | 672
pleocytosis on cerebrospinal fluid | 672
started on intrathecal methotrexate | 672
no improvement in symptoms | 672
changed goals of care to comfort care | 672
passed away | 792
