2.5 years old | 0
male | 0
Pearson syndrome | 0
myelodysplasia | 0
impaired immunity | 0
admitted to the hospital | 0
history of Pearson syndrome | -8760
filgrastim therapy | -8760
bone marrow aspirate | -144
blast cells | -144
monosomy 7 | -144
scraped his left first toe | -336
erythematous scabbed lesion | -336
treated with clindamycin | -336
progressive swelling and erythema | -168
hospitalization | -168
intravenous vancomycin | -168
absolute neutrophil count 6895 | 0
did not improve | 48
cefepime | 48
magnetic resonance imaging | 48
osteomyelitis | 48
sepsis of the first metatarso-pharyngeal joint | 48
voriconazole | 48
ambisome | 48
Orthopedics consultation | 48
aspiration of the first metatarsal | 48
serosanguinous fluid | 48
Fusarium species | 48
suppurative arthritis | 48
invasive fungal disease | 48
severe hypotension | 72
transfer to pediatric intensive care unit | 72
restoration of perfusion | 72
intravenous fluids | 72
dobutamine | 72
blood cultures negative | 72
computed tomography scan | 72
no evidence of fungal dissemination | 72
stabilized | 96
edema and erythema did not improve | 96
biopsy of the first metatarsal | 120
washout of the joint | 120
culture negative for fusarium | 120
fungal elements in bone tissue | 120
voriconazole discontinued | 120
amphotericin B continued | 120
caspofungin | 120
minimal clinical improvement | 240
repeat MRI | 240
progression of bone destruction | 240
joint space widening | 240
partial foot amputation | 360
eradication of osteomyelitis | 360
bone marrow transplant | 360
monosomy 7 | 360
monocytic leukemia | 360
orthopedic surgeons | 360
partial amputation | 360
wide surgical excision | 360
foot instability | 360
future ambulation | 360
Gomori methenamine silver stain | 360
Periodic acid-Schiff stain | 360
fungal hyphae | 360
yeast-like structures | 360
osteomyelitis | 360
abscess formation | 360
caspofungin discontinued | 362
amphotericin B discontinued | 367
bone marrow transplantation | 367
no evidence of recurrent infection | 744
viral respiratory illness | 744
respiratory failure | 744
renal failure | 744
underlying metabolic disorder | 744
death | 744