40 years old | 0
male | 0
admitted to the hospital | 0
resuscitation for cardiac arrest | 0
ventricular fibrillation | 0
Graves’ disease | -120
paroxysmal atrial flutter | -120
atrial fibrillation | 0
ventricular extra systoles | 0
q-waves in anterior leads | 0
elevated troponin-T | 0
elevated creatine kinase | 0
cardiomegaly | 0
dilatation of left ventricle | 0
ejection fractions 25-30% | 0
hypofunction of right ventricle | 0
inferoseptal akinesia | 0
normal coronary arteries | 0
cardiac magnetic resonance imaging | 0
late gadolinium enhancement | 0
Cardiac-Resynchronization-Therapy-Defibrillator device | 24
anticoagulants | 24
antiarrhythmics | 24
statin | 24
heart failure therapy | 24
muscle weakness | -8760
elevated total CK | -8760
proximal weakness of all extremities | 0
progressive muscular weakness | 8760
repetitive supraventricular arrhythmias | 8760
repetitive ventricular arrhythmias | 8760
elevated cardiac enzymes | 8760
serological tests for myositis-specific autoantibodies | 8760
whole-body positron-emission-tomography computed-tomography | 8760
pulmonary function tests | 8760
muscle biopsy | 8760
fiber variability | 8760
cell necrosis | 8760
immune-mediated necrotizing myopathy | 8760
Prednisolone | 8760
improved physical performance | 8760
methotrexate | 10920
tapered prednisolone | 10920
continued clinical improvement | 10920
stable LVEF | 10920
worsening of muscle weakness | 12744
dyspnea | 12744
rising total CK | 12744
pulmonary congestion | 12744
diuretics | 12744
increased methotrexate | 12744
transitory improvement | 12744
cardiogenic shock | 18144
decompensated severe biventricular failure | 18144
inotropic support | 18144
amiodarone | 18144
upregulation of CRT pace | 18144
glucocorticoids | 18144
biventricular hypofunction | 18144
dilatation of left ventricle | 18144
LVEF 10-15% | 18144
nonviable perfusion defect | 18144
myocardial biopsy | 18144
mild to moderate hypertrophy | 18144
maturing replacement fibrosis | 18144
alcian-positive matrix | 18144
endothelial proliferation | 18144
inflammatory cells | 18144
cyclosporine | 18960
mycophenolate mofetil | 18960
prednisolone | 18960
stable peripheral muscle function | 18960
no cardiac improvement | 18960
AMA testing | 20304
AMA positive | 20304
rituximab therapy | 20640
no cardiac improvement | 20640
severe chronic renal impairment | 20976
liver failure | 20976
not a candidate for heart transplantation | 20976
cardiogenic shock | 21216
septic shock | 21216
death | 21216