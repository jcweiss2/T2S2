75 years old | 0
male | 0
Type 2 diabetes mellitus | 0
hypertension | 0
chronic thrombocytopenia | 0
chronic kidney injury | 0
admitted to the hospital | 0
ruptured AAA | -29 months
resection of AAA | -29 months
placement of aortobifemoral bypass graft | -29 months
postoperative renal failure | -29 months
dialysis | -29 months
rigors | -48 hours
dysuria | -48 hours
polyuria | -48 hours
burning micturition | -48 hours
fever | -24 hours
weakness | -24 hours
lethargy | -24 hours
cough denied | 0
chest pain denied | 0
palpitations denied | 0
nausea denied | 0
vomiting denied | 0
constipation denied | 0
blood pressure 70/35 mmHg | 0
blood pressure 90/48 mmHg | 0
temperature 101 degrees Fahrenheit | 0
heart rate 90/min | 0
respiratory rate 20/min | 0
white blood cell count 18,000 | 0
lactic acid 4.1 | 0
20 percent bands | 0
platelet count 20,000 | 0
urinalysis with white blood cells | 0
urinalysis with red blood cells | 0
moderate leukocyte esterase | 0
diffuse abdominal tenderness | 0
peri-umbilical tenderness | 0
severe sepsis | 0
urinary tract infection | 0
high anion gap metabolic acidosis | 0
lactic acidosis | 0
Eggerthella lenta septicemia | 0
Escherichia coli ESBL-positive urinary tract infection | 0
IV antibiotics with etrapenem | 0
abdominal CT with contrast | 0
induration with inflammatory changes around the aortobifemoral bypass graft | 0
stranding around the aorta near the iliac components | 0
air bubble between the components | 0
aortoenteric fistula | 0
graft replacement surgery recommended | 0
graft replacement surgery refused | 0
treatment with IV antibiotics | 0
repeated blood cultures negative | 24 hours
discharged home on antibiotics | 24 hours