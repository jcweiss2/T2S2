72 years old | 0
male | 0
immunocompetent | 0
admitted to the hospital | 0
severe high fever | -72
gastrointestinal symptoms | -72
genitourinary symptoms | -72
diagnosed with acute prostatitis | -72
started on systemic antibiotic therapy | -72
gentamycin 240 mg per 24 h i.v. | -72
urine culture collected | -72
ampicillin-resistant K. pneumoniae isolated | -72
floaters in the right eye | -48
loss of vision | -48
referred to a local ophthalmologist | -48
intraocular inflammation | -45
topical therapy with cycloplegics and corticosteroid eye drops | -45
little benefit | -42
presented to the Eye Hospital | -42
endogenous endophthalmitis suspected | -42
best corrected visual acuity (BCVA) in the right eye was hand motion | -42
intraocular pressure was 12 mmHg | -42
dilated slit lamp eye examination | -42
marked exudation in the anterior chamber | -42
poorly dilated, round pupil | -42
fibrin on the anterior lens capsule | -42
opaque fundus view | -42
right eye ultrasound | -42
vitreous chamber with hyper-reflective signal compatible with abscess or hemorrhage | -42
underwent an urgent and complete pars plana vitrectomy (PPV) | -42
vitreous biopsy | -42
intravitreal injection of vancomycin 1 mg/0.1 ml + ceftazidime 2 mg/0.1 ml | -42
intraoperatively, the retina appeared moderately ischemic | -42
signs of vasculitis | -42
area of infiltrated retina temporal to the central fovea | -42
vitreous samples underwent Gram staining and microbiological cultures | -42
growth of K. pneumoniae | -42
inflammation slowly started to subside | -39
microbiological examinations showed that this strain of K. pneumoniae was resistant to ampicillin | -39
sensitive to all other tested antibiotics | -39
targeted injection of ceftazidime intravitreally | -39
developed fever | -39
sepsis suspected | -39
transferred to the infectious disease department | -39
examined daily by an ophthalmologist | -36
re-deterioration of the vision | -36
referred to the emergency eye clinic | -36
ophthalmoscopy examination | -36
opacities in the vitreous | -36
retinal detachment temporal to the central fovea | -36
moderate cataract | -36
underwent phacoemulsification with in-the-bag intraocular lens (IOL) implantation | -36
posterior capsulotomy | -36
PPV | -36
intraoperative retinal examination | -36
vitreous cavity highly infiltrated with dense inflammatory cells and fibrin | -36
temporal to the fovea was a large retinal necrotic area | -36
no laser photocoagulation nor cryotherapy performed | -36
silicone oil chosen | -36
large barrage around the extensive necrotic area deemed unnecessary | -36
postoperative followup | 0
scar tissue developed in the location of the necrotic retina | 0
retina was flat | 0
inflammation completely disappeared | 0
BCVA improved to 0.2 on the Snellen chart | 0
10-month followup period | 240
retina remained attached and without new changes | 240
silicone oil removed | 240
intraoperatively, laser photocoagulation around the edges of retinal defects performed | 240
visual function improved | 240
retina remained attached | 240
optical coherence tomography scan | 240
regular foveal contour despite the large temporal retinal defect | 240
final BCVA stabilized to 0.3 after 3 months | 360