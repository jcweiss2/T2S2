48 years old | 0
female | 0
admitted to the emergency room | 0
shortness of breath | -3
headache | -3
nausea | -3
increased blood pressure | -3
painless loss of vision | 0.17
heart rate of 104/min | 0
BP of 220/120 mm of Hg | 0
basal crepitations | 0
drowsy but arousable | 0
normal pupillary reflex | 0
normal extra-ocular movements | 0
normal fundoscopy | 0
no light perception | 0
no signs of meningeal irritation | 0
normal hemoglobin | 0
mild leukocytosis | 0
elevated C-reactive protein | 0
normal ESR | 0
normal liver function tests | 0
normal renal function tests | 0
normal coagulation profile | 0
normal autoantibodies | 0
normal neoplastic markers | 0
increased protein level in cerebrospinal fluid | 0
pulmonary edema | 0
normal arterial blood gas analysis | 0
bilateral occipital, parietal and subcortical white matter T2/FLAIR hyperintensities | 0
PRES | 0
nitroglycerin infusion | 0
furosemide | 0
calcium channel blockers | 0
telmisartan | 0
normal lipid profile | 0
normal thyroid profile | 0
diffuse theta/delta slowing | 0
bilateral temporal–occipital epileptiform discharges | 0
normal electrocardiogram | 0
normal echocardiogram | 0
normal ultrasound abdomen | 0
normal renal artery doppler | 0
normal neck vessel doppler | 0
reduced shortness of breath | 120
regaining vision completely | 120
BP of 160/90 mmHg | 96
Telmisartan 40 mg once daily | 96
Cilnidipine 10 mg BID | 96
Hydrochlorothiazide 12.5 mg once daily | 96
Metoprolol 25 mg BID | 96
paradoxical BP increase | 96
elevated urine metanephrine | 96
elevated plasma metanephrine | 96
irregularly marginated, locally infiltrative retroperitoneal mass | 96
paraganglioma | 96
Phenoxybenzamine | 96
surgical resection of the tumor | 168
biopsy confirmed neuroendocrine tumor | 168
discharged in a stable condition | 168
normal BP | 168