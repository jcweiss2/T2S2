41 years old | 0
    man | 0
    presented with pain in the right lower posterior teeth | -168
    swelling in the oral region | -168
    swelling in the maxillofacial region | -168
    swelling in the head and neck regions | -168
    difficulty in breathing | -48
    difficulty in swallowing | -48
    pain in the right lower posterior teeth | -168
    placed a cigarette butt dipped in pesticide "Miehailin" into dental cavity | -168
    no significant improvement in dental pain | -144
    visited a local community clinic | -144
    removed the cigarette butt | -144
    received infusion of anti-inflammatory drugs | -144
    odontogenic infections gradually became aggravated | -120
    spread to floor of the mouth | -120
    spread to submandibular space | -120
    spread to neck | -120
    spread to chest | -120
    spread to waist | -120
    spread to back | -120
    spread to temporal areas | -120
    difficulty in breathing | -48
    difficulty in swallowing | -48
    difficulty in eating | -48
    transferred to our hospital for follow-up treatment | 0
    emergency admission | 0
    mentally exhausted | 0
    poor diet | 0
    poor sleep | 0
    weight loss of approximately 2.5 kg | 0
    healthy history | 0
    no specific diseases | 0
    acutely painful face | 0
    extensive swelling in bilateral temporal region | 0
    extensive swelling in oral region | 0
    extensive swelling in maxillofacial region | 0
    extensive swelling in neck region | 0
    extensive swelling in chest region | 0
    extensive swelling in waist region | 0
    extensive swelling in back region | 0
    pneumatosis in bilateral temporal region | 0
    pneumatosis in oral region | 0
    pneumatosis in maxillofacial region | 0
    pneumatosis in neck region | 0
    pneumatosis in chest region | 0
    pneumatosis in waist region | 0
    pneumatosis in back region | 0
    skin redness | 0
    high temperature | 0
    submandibular space pulsation when touched | 0
    neck region pulsation when touched | 0
    purulent fluid (black, thin, with bubbles, foul odor) | 0
    mouth opening less than 1 cm | 0
    leukocyte count 13.53 × 109/L | 0
    neutrophil ratio 88.40% | 0
    hypersensitive C-reactive protein > 180 mg/L | 0
    procalcitonin 9.8 ng/mL | 0
    potassium 5.65 mmol/L | 0
    sodium 136.4 mmol/L | 0
    chlorine 101.9 mmol/L | 0
    calcium 1.91 mmol/L | 0
    magnesium 0.93 mmol/L | 0
    alanine aminotransferase 19 U/L | 0
    glutamic oxaloacetic aminotransferase 23 U/L | 0
    creatinine 94 µmol/L | 0
    urea 19.1 mmol/L | 0
    platelet count 41.0 × 109/L | 0
    D-dimer 1184 ng/mL | 0
    blood culture positive for Streptococcus viridans | 0
    sensitive to penicillin antibiotics | 0
    extensive swelling in soft tissues bilaterally in oral region | 0
    extensive swelling in soft tissues bilaterally in maxillofacial region | 0
    extensive swelling in soft tissues bilaterally in temporal region | 0
    extensive swelling in soft tissues bilaterally in cervical region | 0
    extensive swelling in soft tissues bilaterally in parapharyngeal space | 0
    extensive swelling in soft tissues bilaterally in chest region | 0
    extensive swelling in soft tissues bilaterally in back region | 0
    extensive swelling in soft tissues bilaterally in mediastinum | 0
    extensive swelling in soft tissues bilaterally in posterior abdominal wall region | 0
    upper respiratory tract narrowed slightly | 0
    bilateral lung pneumothorax | 0
    bilateral pleural effusion | 0
    bilateral pericardial effusion | 0
    left lung pneumothorax (20%-30% compression) | 0
    pulmonary infection in both lungs | 0
    severe multi-space infections bilaterally in oral region | 0
    severe multi-space infections bilaterally in maxillofacial region | 0
    severe multi-space infections bilaterally in head and neck regions | 0
    secondary infections in thorax | 0
    secondary infections in back | 0
    secondary infections in waist | 0
    mediastinal abscess | 0
    bilateral pneumothorax | 0
    bilateral pulmonary infection | 0
    purulent pleural effusion | 0
    pericardial effusion | 0
    secondary thrombocytopenia | 0
    transferred to ICU | 0
    consultations with multiple departments | 0
    abscess incision and drainage in oral region | 0
    abscess incision and drainage in maxillofacial region | 0
    abscess incision and drainage in head and neck regions | 0
    thoracic puncture | 0
    pericardial puncture | 0
    catheter drainage | 0
    pneumothorax management | 0
    management of back infections | 0
    management of waist infections | 0
    anesthesia and respiratory management | 0
    platelet transfusion | 0
    blood transfusion | 0
    intensive care | 0
    antimicrobial administration (Norvancomycin hydrochloride) | 0
    nutritional support | 0
    water, electrolyte, and acid-base stability management | 0
    platelets decreased to 22.00 × 109/L | 24
    alanine aminotransferase 186 U/L | 24
    glutamic oxalate aminotransferase 450 U/L | 24
    cholinesterase 968 U/L | 24
    urea 21.3 mmol/L | 24
    creatinine 153 µmol/L | 24
    potassium 4.77 mmol/L | 24
    sodium 148.8 mmol/L | 24
    chlorine 114.6 mmol/L | 24
    calcium 1.38 mmol/L | 24
    alanine aminotransferase increased to 168 U/L | 48
    glutamic oxalate aminotransferase increased to 1025 U/L | 48
    cholinesterase increased to 814 U/L | 48
    urea increased to 34.44 mmol/L | 48
    creatinine increased to 259 µmol/L | 48
    septic shock | 72
    sudden respiratory arrest | 72
    sudden cardiac arrest | 72
    cardiopulmonary resuscitation | 72
    death | 72
    acute hepatic insufficiency | 72
    acute renal insufficiency | 72
    acute multiple organ failure | 72
    septic shock | 72
    severe multi-space infections bilaterally in oral region | 72
    severe multi-space infections bilaterally in maxillofacial region | 72
    severe multi-space infections bilaterally in head and neck regions | 72
    secondary infections in thorax | 72
    secondary infections in back | 72
    secondary infections in waist | 72
    mediastinal abscess | 72
    bilateral pneumothorax | 72
    bilateral pulmonary infection | 72
    purulent pleural effusion | 72
    pericardial effusion | 72
    secondary thrombocytopenia | 72

<|eot_id|>