49 years old | 0
male | 0
admitted to the hospital | 0
fever | 0
chills | 0
diarrhea | 0
highest temperature was 40 °C | -72
history of acute pancreatitis | -2628
history of fatty liver | -2628
liver cirrhosis | -30
mild ascites | -30
esophageal variceal ligation | -16
drunk wine 0.5 kg/day | -8760
intermittently seditious | 0
confused | 0
disoriented | 0
skin was yellowish | 0
shifting dullness was positive | 0
lower limb edema was moderate | 0
body temperature was 38.7 °C | 0
heart rate was 100 beats per minute | 0
blood pressure was 100/54 mmHg | 0
WBC was 6.0 × 10^9/L | 0
neutrophilic granulocyte percentage was 68.5% | 0
hemoglobin was 69 g/L | 0
total bilirubin was 126.8 μmol/L | 0
direct bilirubin was 61.5 μmol/L | 0
alanine aminotransferase was 37.39 U/L | 0
aspartate aminotransferase was 54.7 U/L | 0
γ-glutamyl transpeptidase was 72.05 U/L | 0
albumin was 29 g/L | 0
blood urea nitrogen was 9.77 mmol/L | 0
creatinine was 67.8 μmol/L | 0
prothrombin time was 30.7 s | 0
INR was 2.90 | 0
procalcitonin was 25.24 ng/mL | 0
PaO2 was 79 mmHg | 0
FiO2 was 29.0% | 0
pneumonia | 0
hydrothorax | 0
liver cirrhosis | 0
splenomegaly | 0
cholecystitis | 0
ascites | 0
right renal calculus | 0
ACLF grade 1 | 0
Child-Pugh score was 12 | 0
MELD score was 25.4 | 0
treated with ademetionine | 0
treated with L-Ornithine-L-Aspartate | 0
treated with montmorillonite powder | 0
treated with bifidobacterium lactobacillus tripterygium | 0
treated with ceftriaxone sodium | 0
febrile | 24
temperature was up to 38.5 °C | 24
BP was 59/23 mmHg | 24
heart rate was 110 beats per minute | 24
oliguria | 24
septic shock | 24
blood culture findings revealed epidermal staphylococcus and gram-positive bacteria | 24
WBC was 9.9 × 10^9/L | 24
GR% was 84.4% | 24
Hb was 63 g/L | 24
TBIL was 138.6 μmol/L | 24
DBIL was 85.5 μmol/L | 24
AST was 40.51 U/L | 24
γ-GGT was 63.38 U/L | 24
BUN was 15.76 mmol/L | 24
Cr was 143.56 μmol/L | 24
PT was 33.6 s | 24
INR was 3.25 | 24
AKI stage 2 | 24
ACLF grade 2 | 24
red blood cells were transfused | 24
dopamine was infused | 24
meropenem was infused | 24
terlipressin was infused | 24
hematemesis | 28
esomeprazole was infused | 28
somatostatin was infused | 28
human albumin was infused | 28
BP was 86/57 mmHg | 48
heart rate was 110 beats per minute | 48
body temperature was 37 °C | 48
WBC was 5.4 × 10^9/L | 48
GR% was 78.4% | 48
Hb was 94 g/L | 48
TBIL was 155.9 μmol/L | 48
DBIL was 90.4 μmol/L | 48
AST was 32.52 U/L | 48
γ-GGT was 52.3 U/L | 48
BUN was 10.27 mmol/L | 48
Cr was 42.04 μmol/L | 48
GR% improved | 120
C-reaction protein improved | 120
procalcitonin improved | 120
Cr improved | 120
urine volume improved | 120
fecal occult blood test was negative | 312
WBC was 11.1 × 10^9/L | 312
GR% was 65.5% | 312
Hb was 84 g/L | 312
Cr was 54.56 μmol/L | 312
C-reaction protein was 16.5 mg/L | 312
procalcitonin was 0.03 ng/mL | 312
no ACLF | 312
discharged | 312
mild distension of abdomen | 504
mild lower limb edema | 504
Hb was 87 g/L | 504
TBIL was 77.4 μmol/L | 504
DBIL was 40.9 μmol/L | 504
AST was 54.77 U/L | 504
ALT was 28.05 U/L | 504
γ-GGT was 61.07 U/L | 504
ALB was 30.6 g/L | 504
BUN was 5.36 mmol/L | 504
Cr was 36.79 μmol/L | 504
PT was 19.7 s | 504
INR was 1.67 | 504
furosemide was prescribed | 504
spironolactone was prescribed | 504