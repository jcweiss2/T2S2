75 years old | 0
female | 0
multiple left renal calculi | -672
right upper ureteric calculus | -672
abdominal X-ray | -672
sonography | -672
PCNL | -24
severe bleeding | -24
percutaneous nephrostomy drainage tube placement | -24
transfer to hospital | -24
hemodynamically unstable condition | 0
resuscitation | 0
blood transfusion | 0
acute kidney injury | 0
serum urea 105 mg/dL | 0
serum creatinine 5.77 mg/dL | 0
noncontrast CT abdomen | 0
PNDT in renal vein | 0
suspected renal vein thrombosis | 0
hemodialysis | 24
bilateral urinary diversion | 24
cystoscopy | 48
right-sided double-J stent placement | 48
left-sided percutaneous nephrostomy | 48
sepsis | 0
improvement of condition | 72
CT renal angiography | 96
dynamic renal scan | 168
confirmation of PNDT in renal vein | 168
renal vein thrombosis | 168
no uptake in left kidney | 168
planning for left nephrectomy | 168
laparoscopic left simple nephrectomy with thrombectomy | 192
dense adhesions | 192
two renal arteries | 192
PNDT in renal vein with thrombus | 192
clipping of renal arteries | 192
clipping of renal vein | 192
removal of PNDT | 192
operative time 125 min | 192
evaluation of specimen | 192
direct tract from renal cortex into renal vein | 192
intra-abdominal drain removal | 216
discharge | 216
planning for right ureteroscopic lithotripsy | 216