5 years old | 0
male | 0
presented with fever | -1464
presented with night sweats | -1464
presented with weight loss | -1464
presented with cough | -1464
bilateral anterior cervical lymph nodes enlargement | 0
peripheral cyanosis in digits | 0
hemoglobin concentration: 128 g/L | 0
white blood cell count: 9.12×109/L | 0
platelet count: 329×109/L | 0
normal liver enzymes | 0
normal serum bilirubin | 0
normal creatinine | 0
normal blood urea nitrogen | 0
blood culture: no bacterial growth | 0
chest X-ray: bilateral airway narrowing | 0
neck CT scan: multiple bilateral anterior cervical lymphadenopathy | 0
neck CT scan: supraclavicular lymphadenopathy | 0
neck CT scan: infraclavicular lymphadenopathy | 0
neck CT scan: mass effect | 0
neck CT scan: largest lymph node 20 × 15 mm | 0
neck CT scan: cystic degeneration suggestive of central necrosis | 0
neck CT scan: thyroid gland heterogenous density | 0
chest CT scan: bilateral nodular and micronodular lung densities | 0
chest CT scan: hilar lymphadenopathy | 0
abdominal CT scan: mild hepatomegaly | 0
abdominal CT scan: paraaortic lymph node enlargement | 0
clinical impression: tuberculosis or Hodgkin’s lymphoma | 0
excisional biopsy of cervical lymph node | 0
bone marrow trephine biopsy | 0
histopathological examination: malignant thyroid glands | 0
histopathological examination: papillary growth | 0
histopathological examination: nuclear clearing | 0
histopathological examination: nuclear grooves | 0
histopathological examination: residual rim of lymph node tissue | 0
bone marrow biopsy: negative for metastasis | 0
diagnosis of metastatic papillary thyroid carcinoma | 0
clinical stage-I disease | 0
total thyroidectomy | 0
cervical lymph nodes excision | 0
radioactive iodine therapy | 0
complete remission | 0
developed respiratory symptoms | 4320
CT scan: multiple bilateral pulmonary nodules | 4320
multiple admissions to ICU for unstable vital signs | 4320
died of septicemia by methicillin-resistant Staphylococcus aureus | 4416
blood culture: no bacterial growth |$ 
