77 years old | 0
male | 0
admitted to the hospital | 0
syncope | 0
hypertension | -672
hyperlipidemia | -672
uncontrolled diabetes mellitus type two | -672
diabetic foot ulcers | -672
osteomyelitis | -672
peripheral vascular disease | -672
coronary artery disease | -672
pacemaker/defibrillator implantation | -6120
systolic heart failure | -6120
ischemic cardiomyopathy | -6120
dizziness | -72
dyspnea | -72
fevers | -72
elevated blood glucose | -72
lethargy | -72
rigors | -72
chills | -72
malaise | -72
elevated troponin | 0
elevated NT-proBNP | 0
leukocytosis | 0
wide complex tachycardia | 0
tachypnea | 0
hypertension | 0
cardioversion | 0
 Levophed initiation | 0
empiric antibiotic therapy | 0
agonal breathing | 0
intubation | 0
transfer to ICU | 0
hypotension | 0
dopamine initiation | 0
cardiac catheterization | 0
PCI | 0
stent deployment | 0
pseudoaneurysm identification | 0
IABP insertion | 0
persistent ventricular tachycardia | 0
lidocaine infusion | 0
amiodarone infusion | 0
MSSA positive blood cultures | 48
elevated liver function tests | 48
elevated creatinine | 48
IABP removal | 48
vancomycin transition to linezolid | 48
Levophed titration | 48
extubation | 72
BiPAP initiation | 72
volume overload | 72
monitored diuresis | 72
IV amiodarone transition to oral | 72
Infectious Disease Service consultation | 72
cefazolin and rifampin initiation | 72
leukocytosis resolution | 96
defervesce | 96
ventricular tachycardia episodes | 96
AICD discharges | 96
pacemaker interrogation | 96
lidocaine infusion resumption | 96
mexiletine initiation | 120
amiodarone continuation | 120
TEE recommendation | 120
transcutaneous pacer pads placement | 120
palliative care consideration | 120
Diuril initiation | 120
Precedex discontinuation | 120
lidocaine drip transition to amiodarone | 144
mexiletine continuation | 144
amiodarone infusion continuation | 144
TTE | 144
dilated left ventricle | 144
segmental wall motion abnormalities | 144
LVEF 35% | 144
moderate concentric left ventricular hypertrophy | 144
left atrial enlargement | 144
mitral annular calcification | 144
mild mitral regurgitation | 144
TEE | 168
fibrinous lead vegetations | 168
probable abscess | 168
lateral wall of the right atrium | 168
4.0×4.4×3.9 cm abscess | 168
lucent core | 168
encasing the lead | 168
gentamicin initiation | 168
tertiary care transfer proposal | 168
transfer decline | 192
lidocaine and amiodarone drips discontinuation | 192
mexiletine and amiodarone continuation | 192
defibrillator and detection functions inhibition | 192
pacemaker function intact | 192
antibiotic treatment continuation | 192
discharge home with hospice | 216