63 years old | 0
female | 0
chronic hepatitis B-related cirrhosis | -8760
Child-Pugh class A | -8760
oral antiviral treatment with entecavir | -8760
type II Diabetic mellitus | -8760
hypertension | -8760
HCC | -720
AJCC/TNM stage II | -720
BCLC stage B | -720
transarterial chemoembolization | -720
TACE | -720
follow-up contrast-enhanced CT | -30
poorly enhanced nodules | -30
RFA | 0
ultrasound-guided RFA | 0
general anesthesia | 0
fever | 6
chills | 6
dyspnea | 6
abdominal pain | 6
body temperature increased | 6
heart rate increased | 6
blood pressure decreased | 6
WBC increased | 6
neutrophil predominant | 6
hyperlactatemia | 6
CRP increased | 6
AST increased | 6
ALT increased | 6
total bilirubin increased | 6
albumin decreased | 6
INR increased | 6
Cr increased | 6
Ammonia increased | 6
abdominal ultrasound | 6
hyperechoic change | 6
air formation | 6
contrast-enhanced CT | 6
necrotic changes | 6
air component | 6
intra-tumoral abscess formation | 6
septic shock | 6
oxygen supplement | 6
aggressive fluid resuscitation | 6
empirical antibiotic | 6
intravenous Flomoxef | 6
ultrasound-guided aspiration | 6
pus discharge | 6
pus culture | 6
packed red blood cell transfusion | 6
fresh frozen plasma transfusion | 6
anemia correction | 6
coagulopathy correction | 6
C. perfringens infection | 78
liver abscess | 78
blood culture | 78
drug sensitivity test | 78
Flomoxef susceptible | 78
abscess aspiration | 78
antibiotics completion | 78
infection control | 78
discharged | 720
stable condition | 720
follow-up contrast-enhanced CT | 2160
complete ablation | 2160
no local tumor recurrence | 2160