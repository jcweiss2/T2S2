48 years old | 0
man | 0
presented to the Emergency Room | 0
headache | 0
subarachnoid hemorrhage | 0
untreated hypertension | 0
no smoking history | 0
no family history of thrombotic disease | 0
admitted to hospital | 0
surgical titanium clipping for left intracranial aneurysms | 0
surgery completed without complications | 0
transferred from ICU to general ward | 72
receiving rehabilitation (walking and brain training) | 72
high grade fever | 120
chills | 120
nausea | 120
ceftriaxone initiated | 120
vancomycin initiated | 120
possible meningitis | 120
hypotensive | 144
tachycardia | 144
temperature 37.4°C | 144
blood pressure 62/52 mmHg | 144
heart rate 110/min | 144
respiratory rate 26 breaths/min | 144
oxygen saturation 68% at 3 L/min supplemental oxygen | 144
cold limbs | 144
cyanosis | 144
tachypnea | 144
leukocytosis (WBC 20,900/μL) | 144
elevated AST (103 U/L) | 144
elevated ALT (106 U/L) | 144
elevated serum creatinine (3.71 mg/dL) | 144
elevated C-reactive protein (29.33 mg/dL) | 144
normal protein C level | 144
pyuria | 144
bacteriuria | 144
acute focal bacterial nephritis | 144
septic shock due to nephritis | 144
intravenous fluid resuscitation | 144
meropenem (1 g 12h) | 144
vancomycin (1 g q24h) | 144
metronidazole (500 mg q8h) | 144
norepinephrine | 144
vasopressin | 144
methylprednisolone 200 mg/day | 144
recombinant thrombomodulin for DIC | 144
continuous hemodiafiltration | 144
Enterobacter aerogenes in blood cultures | 168
sensitive to meropenem and piperacillin/tazpbactum | 168
high-grade fever | 168
DIC | 168
platelet transfusion | 168
extensive purpura | 168
purpura fulminans due to infection | 168
skin purpura and necrosis | 168
skin biopsy necrosis and bullae | 168
thrombosis | 168
planned limb amputation | 168
hypotension improved temporarily | 216
low platelet levels improved temporarily | 216
high-grade persistent fever | 216
chills | 216
changed all devices (central venous catheter, arterial line, vascular access) | 216
two sets of blood cultures | 216
persistent bacteremia with Enterobacter aerogenes | 216
transfusion dependent | 216
progressing anemia | 216
low platelet levels | 216
received 100 units of platelets | 216
received 10 units of red blood cells | 216
condition progressively worsened | 456
died | 456
autopsy multiple abscesses and thrombosis in lung, intestinal tract, kidney | 456
