29 years old | 0
male | 0
admitted to the hospital | 0
severe dysphonia | 0
dyspnea | 0
15 kg weight loss in 6 months | -4320
recurrent fever | 0
coughing | -336
fever | -336
leg pain | -336
elevated lactate dehydrogenase (298 U/L) | -336
elevated C-reactive protein (11.5 mg/dL) | -336
elevated uric acid (8.7 mg/dL) | -336
elevated d-dimer (1.58 mg/dL) | -336
discharged | -336
symptomatic treatment | -336
suspected viral infection | -336
no imaging diagnostics | -336
elevated LDH (444 U/L) | 0
elevated uric acid (8 mg/dL) | 0
elevated CRP (27.7 mg/dL) | 0
cervical lymphadenopathy | 0
supraclavicular lymphadenopathy | 0
left vocal cord paresis | 0
FDG-PET/MRI | 0
FDG uptake in left hemithorax | 0
FDG uptake in mediastinum | 0
FDG uptake in supraclavicular lymph nodes | 0
infradiaphragmal lymph nodes |0
intrapulmonary masses | 0
cervical lymph node removal | 0
diffuse proliferation of centroblastic lymphoid cells | 0
high proliferative activity (80% Ki-67 positivity) | 0
CD20 positive | 0
Pax5 positive | 0
Bcl6 positive | 0
MUM-1 positive | 0
CD5 negative | 0
CD23 negative | 0
Cyclin D1 negative | 0
CD30 negative | 0
EBV negative | 0
diffuse large B-cell lymphoma diagnosis | 0
stage IVB DLBCL | 0
bone marrow biopsy no infiltration | 0
dexamethasone prephase | 0
rapid regression of dyspnea | 0
rapid regression of dysphonia | 0
Rituximab-CHOP regimen | 0
Rituximab 375 mg/m2 | 0
doxorubicin 50% reduction | 0
cyclophosphamide 50% reduction | 0
vincristine 2 mg | 0
vincristine 1 mg | 0
prednisolone 100 mg | 0
cotrimoxazole prophylaxis | 0
valaciclovir prophylaxis | 0
posaconazole prophylaxis | 0
ciprofloxacin prophylaxis | 0
PEGylated granulocyte colony-stimulating factor | 0
outpatient cycles 2-6 | 0
additional rituximab doses | 0
PET/MRI complete remission | 0
mediastinal lymphadenopathy | 8760
hilar lymphadenopathy | 8760
thoracoscopy biopsy | 8760
chronic inflammation | 8760
no neoplasia | 8760
biopsy-proven complete remission | 8760
Nijmegen breakage syndrome diagnosis | -262080
stage IV nodular sclerosis cHL | -17520
CR after 4 cycles of chemotherapy | -17520
liver failure | -17520
kidney failure | -17520
fungal sepsis | -17520
restored liver function | -17520
restored kidney function | -17520
selective IgG4 deficiency | -262080
previous genotoxic chemotherapy | -17520
secondary malignancies risk | 0
life-threatening infections absence | 0
individualized regimen | 0
extended prophylaxis | 0
monitoring | 0
functional imaging without DNA damage | 0
aggressive therapy | 0
standard immunochemotherapy | 0
second complete remission | 0
