49 years old|0
    morbidly obese|0
    African American|0
    man|0
    end-stage renal disease|0
    peritoneal dialysis (PD)|0
    hypertension|0
    admitted to the hospital|0
    nausea|-96
    nonbilious nonbloody emesis|-96
    severe diffuse abdominal pain|-96
    symptoms reported to outpatient PD nurse|-48
    cloudy white fluid|-48
    peritoneal fluid sent for evaluation|-48
    culture sent for evaluation|-48
    started on 1 g intraperitoneal cefazolin|-48
    started on 1 g intraperitoneal ceftazidime|-48
    fever (101.5 °F) measured on home thermometer|-24
    PD for 2 years|0
    no prior similar episode|0
    oliguric at baseline|0
    not using sterile aseptic technique during last week|0
    using dish towels to wipe hands before accessing transfer set|0
    using dish towels to wipe hands after accessing transfer set|0
    afebrile on admission|0
    blood pressure 95/72 mmHg|0
    heart rate 88 bpm|0
    respiratory rate 20 breaths/min|0
    acute distress secondary to abdominal pain|0
    distended abdomen|0
    tender to light palpation|0
    positive fluid wave|0
    dull to percussion|0
    leukocytosis 13,700|0
    potassium 3.3 mmol/L|0
    anion gap 25|0
    peritoneal fluid total white blood cell count 93,557|-48
    neutrophil predominance 80%|-48
    organism identified as Acinetobacter pittii on hospital day 1|24
    susceptibilities pending|24
    started on intraperitoneal ceftazidime|24
    started on intraperitoneal gentamicin|24
    susceptibilities returned on hospital day 2|48
    sensitive to ceftazidime (4 μg/mL)|48
    blood culture results showed no growth on day 5|120
    continued on intraperitoneal ceftazidime 1.5 g as last fill for 21 days|0
    persistence of cloudy effluent as an outpatient|0
    treatment extended to 28 days|0
    readmitted to the hospital for fever on day 34|816
    readmitted to the hospital for abdominal pain on day 34|816
    peritoneal fluid cell count elevated to 43,245/μL|816
    80% neutrophils|816
    cultures growing same organism|816
    initially treated with dual therapy of vancomycin and gentamicin|816
    subsequently placed on intravenous ceftazidime|816
    blood cultures in second hospital stay showed no growth|816
    improvement in abdominal pain|816
    decreasing intraperitoneal white blood cell count|816
    PD catheter removed|816
    hemodialysis (HD) initiated via tunneled HD catheter|816
    discharged with 2-week course of ciprofloxacin|816
    plan for HD until kidney transplant becomes available|816
    asymptomatic upon completion of therapy|816
    no growth in blood cultures|816
    no prior similar episode|0
    oliguric at baseline|0
    not using sterile aseptic technique during last week|0
    using dish towels to wipe hands before accessing transfer set|0
    using dish towels to wipe hands after accessing transfer set|0
    afebrile on admission|0
    blood pressure 95/72 mmHg|0
    heart rate 88 bpm|0
    respiratory rate 20 breaths/min|0
    acute distress secondary to abdominal pain|0
    distended abdomen|0
    tender to light palpation|0
    positive fluid wave|0
    dull to percussion|0
    leukocytosis 13,700|0
    potassium 3.3 mmol/L|0
    anion gap 25|0
    peritoneal fluid total white blood cell count 93,557|-48
    neutrophil predominance 80%|-48
    organism identified as Acinetobacter pittii on hospital day 1|24
    susceptibilities pending|24
    started on intraperitoneal ceftazidime|24
    started on intraperitoneal gentamicin|24
    susceptibilities returned on hospital day 2|48
    sensitive to ceftazidime (4 μg/mL)|48
    blood culture results showed no growth on day 5|120
    continued on intraperitoneal ceftazidime 1.5 g as last fill for 21 days|0
    persistence of cloudy effluent as an outpatient|0
    treatment extended to 28 days|0
    readmitted to the hospital for fever on day 34|816
    readmitted to the hospital for abdominal pain on day 34|816
    peritoneal fluid cell count elevated to 43,245/μL|816
    80% neutrophils|816
    cultures growing same organism|816
    initially treated with dual therapy of vancomycin and gentamicin|816
    subsequently placed on intravenous ceftazidime|816
    blood cultures in second hospital stay showed no growth|816
    improvement in abdominal pain|816
    decreasing intraperitoneal white blood cell count|816
    PD catheter removed|816
    hemodialysis (HD) initiated via tunneled HD catheter|816
    discharged with 2-week course of ciprofloxacin|816
    plan for HD until kidney transplant becomes available|816
    asymptomatic upon completion of therapy|816
    no growth in blood cultures|816
    no prior similar episode|0
    oliguric at baseline|0
    not using sterile aseptic technique during last week|0
    using dish towels to wipe hands before accessing transfer set|0
    using dish towels to wipe hands after accessing transfer set|0
    afebrile on admission|0
    blood pressure 95/72 mmHg|0
    heart rate 88 bpm|0
    respiratory rate 20 breaths/min|0
    acute distress secondary to abdominal pain|0
    distended abdomen|0
    tender to light palpation|0
    positive fluid wave|0
    dull to percussion|0
    leukocytosis 13,700|0
    potassium 3.3 mmol/L|0
    anion gap 25|0
    peritoneal fluid total white blood cell count 93,557|-48
    neutrophil predominance 80%|-48
    organism identified as Acinetobacter pittii on hospital day 1|24
    susceptibilities pending|24
    started on intraperitoneal ceftazidime|24
    started on intraperitoneal gentamicin|24
    susceptibilities returned on hospital day 2|48
    sensitive to ceftazidime (4 μg/mL)|48
    blood culture results showed no growth on day 5|120
    continued on intraperitoneal ceftazidime 1.5 g as last fill for 21 days|0
    persistence of cloudy effluent as an outpatient|0
    treatment extended to 28 days|0
    readmitted to the hospital for fever on day 34|816
    readmitted to the hospital for abdominal pain on day 34|816
    peritoneal fluid cell count elevated to 43,245/μL|816
    80% neutrophils|816
    cultures growing same organism|816
    initially treated with dual therapy of vancomycin and gentamicin|816
    subsequently placed on intravenous ceftazidime|816
    blood cultures in second hospital stay showed no growth|816
    improvement in abdominal pain|816
    decreasing intraperitoneal white blood cell count|816
    PD catheter removed|816
    hemodialysis (HD) initiated via tunneled HD catheter|816
    discharged with 2-week course of ciprofloxacin|816
    plan for HD until kidney transplant becomes available|816
    asymptomatic upon completion of therapy|816
    no growth in blood cultures|816
    no prior similar episode|0
    oliguric at baseline|0
    not using sterile aseptic technique during last week|0
    using dish towels to wipe hands before accessing transfer set|0
    using dish towels to wipe hands after accessing transfer set|0
    afebrile on admission|0
    blood pressure 95/72 mmHg|0
    heart rate 88 bpm|0
    respiratory rate 20 breaths/min|0
    acute distress secondary to abdominal pain|0
    distended abdomen|0
    tender to light palpation|0
    positive fluid wave|0
    dull to percussion|0
    leukocytosis 13,700|0
    potassium 3.3 mmol/L|0
    anion gap 25|0
    peritoneal fluid total white blood cell count 93,557|-48
    neutrophil predominance 80%|-48
    organism identified as Acinetobacter pittii on hospital day 1|24
    susceptibilities pending|24
    started on intraperitoneal ceftazidime|24
    started on intraperitoneal gentamicin|24
    susceptibilities returned on hospital day 2|48
    sensitive to ceftazidime (4 μg/mL)|48
    blood culture results showed no growth on day 5|120
    continued on intraperitoneal ceftazidime 1.5 g as last fill for 21 days|0
    persistence of cloudy effluent as an outpatient|0
    treatment extended to 28 days|0
    readmitted to the hospital for fever on day 34|816
    readmitted to the hospital for abdominal pain on day 34|816
    peritoneal fluid cell count elevated to 43,245/μL|816
    80% neutrophils|816
    cultures growing same organism|816
    initially treated with dual therapy of vancomycin and gentamicin|816
    subsequently placed on intravenous ceftazidime|816
    blood cultures in second hospital stay showed no growth|816
    improvement in abdominal pain|816
    decreasing intraperitoneal white blood cell count|816
    PD catheter removed|816
    hemodialysis (HD) initiated via tunneled HD catheter|816
    discharged with 2-week course of ciprofloxacin|816
    plan for HD until kidney transplant becomes available|816
    asymptomatic upon completion of therapy|816
    no growth in blood cultures|816
    no prior similar episode|0
    oliguric at baseline|0
    not using sterile aseptic technique during last week|0
    using dish towels to wipe hands before accessing transfer set|0
    using dish towels to wipe hands after accessing transfer set|0
    afebrile on admission|0
    blood pressure 95/72 mmHg|0
    heart rate 88 bpm|0
    respiratory rate 20 breaths/min|0
    acute distress secondary to abdominal pain|0
    distended abdomen|0
    tender to light palpation|0
    positive fluid wave|0
    dull to percussion|0
    leukocytosis 13,700|0
    potassium 3.3 mmol/L|0
    anion gap 25|0
    peritoneal fluid total white blood cell count 93,557|-48
    neutrophil predominance 80%|-48
    organism identified as Acinetobacter pittii on hospital day 1|24
    susceptibilities pending|24
    started on intraperitoneal ceftazidime|24
    started on intraperitoneal gentamicin|24
    susceptibilities returned on hospital day 2|48
    sensitive to ceftazidime (4 μg/mL)|48
    blood culture results showed no growth on day 5|120
    continued on intraperitoneal ceftazidime 1.5 g as last fill for 21 days|0
    persistence of cloudy effluent as an outpatient|0
    treatment extended to 28 days|0
    readmitted to the hospital for fever on day 34|816
    readmitted to the hospital for abdominal pain on day 34|816
    peritoneal fluid cell count elevated to 43,245/μL|816
    80% neutrophils|816
    cultures growing same organism|816
    initially treated with dual therapy of vancomycin and gentamicin|816
    subsequently placed on intravenous ceftazidime|816
    blood cultures in second hospital stay showed no growth|816
    improvement in abdominal pain|816
    decreasing intraperitoneal white blood cell count|816
    PD catheter removed|816
    hemodialysis (HD) initiated via tunneled HD catheter|816
    discharged with 2-week course of ciprofloxacin|816
    plan for HD until kidney transplant becomes available|816
    asymptomatic upon completion of therapy|816
    no growth in blood cultures|816
    no prior similar episode|0
    oliguric at baseline|0
    not using sterile aseptic technique during last week|0
    using dish towels to wipe hands before accessing transfer set|0
    using dish towels to wipe hands after accessing transfer set|0
    afebrile on admission|0
    blood pressure 95/72 mmHg|0
    heart rate 88 bpm|0
    respiratory rate 20 breaths/min|0
    acute distress secondary to abdominal pain|0
    distended abdomen|0
    tender to light palpation|0
    positive fluid wave|0
    dull to percussion|0
    leukocytosis 13,700|0
    potassium 3.3 mmol/L|0
    anion gap 25|0
    peritoneal fluid total white blood cell count 93,557|-48
    neutrophil predominance 80%|-48
    organism identified as Acinetobacter pittii on hospital day 1|24
    susceptibilities pending|24
    started on intraperitoneal ceftazidime|24
    started on intraperitoneal gentamicin|24
    susceptibilities returned on hospital day 2|48
    sensitive to ceftazidime (4 μg/mL)|48
    blood culture results showed no growth on day 5|120
    continued on intraperitoneal ceftazidime 1.5 g as last fill for 21 days|0
    persistence of cloudy effluent as an outpatient|0
    treatment extended to 28 days|0
    readmitted to the hospital for fever on day 34|816
    readmitted to the hospital for abdominal pain on day 34|816
    peritoneal fluid cell count elevated to 43,245/μL|816
    80% neutrophils|816
    cultures growing same organism|816
    initially treated with dual therapy of vancomycin and gentamicin|816
    subsequently placed on intravenous ceftazidime|816
    blood cultures in second hospital stay showed no growth|816
    improvement in abdominal pain|816
    decreasing intraperitoneal white blood cell count|816
    PD catheter removed|816
    hemodialysis (HD) initiated via tunneled HD catheter|816
    discharged with 2-week course of ciprofloxacin|816
    plan for HD until kidney transplant becomes available|816
    asymptomatic upon completion of therapy|816
    no growth in blood cultures|816
    no prior similar episode|0
    oliguric at baseline|0
    not using sterile aseptic technique during last week|0
    using dish towels to wipe hands before accessing transfer set|0
    using dish towels to wipe hands after accessing transfer set|0
    afebrile on admission|0
    blood pressure 95/72 mmHg|0
    heart rate 88 bpm|0
    respiratory rate 20 breaths/min|0
    acute distress secondary to abdominal pain|0
    distended abdomen|0
    tender to light palpation|0
    positive fluid wave|0
    dull to percussion|0
    leukocytosis 13,700|0
    potassium 3.3 mmol/L|0
    anion gap 25|0
    peritoneal fluid total white blood cell count 93,557|-48
    neutrophil predominance 80%|-48
    organism identified as Acinetobacter pittii on hospital day 1|24
    susceptibilities pending|24
    started on intraperitoneal ceftazidime|24
    started on intraperitoneal gentamicin|24
    susceptibilities returned on hospital day 2|48
    sensitive to ceftazidime (4 μg/mL)|48
    blood culture results showed no growth on day 5|120
    continued on intraperitoneal ceftazidime 1.5 g as last fill for 21 days|0
    persistence of cloudy effluent as an outpatient|0
    treatment extended to 28 days|0
    readmitted to the hospital for fever on day 34|816
    readmitted to the hospital for abdominal pain on day 34|816
    peritoneal fluid cell count elevated to 43,245/μL|816
    80% neutrophils|816
    cultures growing same organism|816
    initially treated with dual therapy of vancomycin and gentamicin|816
    subsequently placed on intravenous ceftazidime|816
    blood cultures in second hospital stay showed no growth|816
    improvement in abdominal pain|816
    decreasing intraperitoneal white blood cell count|816
    PD catheter removed|816
    hemodialysis (HD) initiated via tunneled HD catheter|816
    discharged with 2-week course of ciprofloxacin|816
    plan for HD until kidney transplant becomes available|816
    asymptomatic upon completion of therapy|816
    no growth in blood cultures|816
    no prior similar episode|0
    oliguric at baseline|0
    not using sterile aseptic technique during last week|0
    using dish towels to wipe hands before accessing transfer set|0
    using dish towels to wipe hands after accessing transfer set|0
    afebrile on admission|0
    blood pressure 95/72 mmHg|0
    heart rate 88 bpm|0
    respiratory rate 20 breaths/min|0
    acute distress secondary to abdominal pain|0
    distended abdomen|0
    tender to light palpation|0
    positive fluid wave|0
    dull to percussion|0
    leukocytosis 13,700|0
    potassium 3.3 mmol/L|0
    anion gap 25|0
    peritoneal fluid total white blood cell count 93,557|-48
    neutrophil predominance 80%|-48
    organism identified as Acinetobacter pittii on hospital day 1|24
    susceptibilities pending|24
    started on intraperitoneal ceftazidime|24
    started on intraperitoneal gentamicin|24
    susceptibilities returned on hospital day 2|48
    sensitive to ceftazidime (4 μg