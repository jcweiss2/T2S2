65 years old | 0
male | 0
hypertension | 0
depression | 0
fevers | -168
malaise | -168
chest x-ray | -168
COVID swab | -168
admitted to ambulatory respiratory care unit | -24
referred to emergency department | -24
found to be in shock | 0
admitted to medical intensive care unit | 24
cardiac biomarkers peak | 12
able to be fully weaned from vasopressor support | 12
transferred to cardiac intensive care unit | 24
transferred out of cardiac intensive care unit to general cardiology service | 72
coronary angiogram | 96
cardiac magnetic resonance imaging | 120
myopericarditis | 120
anaplasma polymerase chain reaction testing | 144
discharged | 144
follow-up 2 weeks | 336
followed up with infectious disease | 336
stopped antibiotics | 336
repeat cardiac magnetic resonance imaging | 336
follow-up 4 weeks | 672
followed up with heart failure | 672
back to baseline functional status | 672
electrocardiogram | 672
ambulatory rhythm monitoring | 672
dental work | -24
ill-appearing | 0
temperature 97.7 Fahrenheit | 0
heart rate 63 beats per minute | 0
blood pressure 74/44 mm of mercury | 0
respiratory rate 20 breaths per minute | 0
oxygen saturation 99% on room air | 0
crackles at the right lung base | 0
II out of VI holosystolic murmur at the cardiac apex | 0
AST 89 IU/L | 0
ALT 103 IU/L | 0
proBNP of 16 093 pg/mL | 0
Troponin-T of 0.79 ng/mL | 0
CRP > 300 mg/L | 0
creatinine 2.6 mg/dL | 0
lactate 3.4 mmol/L | 0
atrial fibrillation | 0
non-specific intraventricular conduction delay | 0
minimal ST elevation in the lateral leads | 0
amlodipine | 0
losartan | 0
lamotrigine | 0
vancomycin | 0
ceftriaxone | 0
doxycycline | 0
unfractionated heparin | 0
apixaban | 120
fever abated | 12
blood pressure stabilized | 12
vasopressors weaned | 12
renal function improved | 12
cardiac biomarkers peaked | 12
peak troponin-T 1.24 | 12
CK-MB 57 | 12
coronary angiography | 96
obstructive coronary artery disease | 96
LVEF 54% | 120
dilated right ventricle | 120
moderate-to-severe RV systolic dysfunction | 120
tricuspid annular plane systolic excursion 1.3 cm | 120
leftward interventricular septal shift in systole and diastole | 120
mild to moderate tricuspid regurgitation | 120
no significant left-sided valvular disease | 120
no pericardial effusion | 120
Lyme IgG serology positive | 120
western blot negative for three of three different IgM bands | 120
positive for only one of 10 different IgG bands | 120
anaplasma serologies positive for IgM | 144
anaplasma serologies negative for IgG | 144
anaplasma phagocytophilum DNA detected | 144
mixed shock | 0
vasodilation | 0
hypovolaemia | 0
RV dysfunction | 0
myopericarditis | 120
conduction system disease | 0
atrial fibrillation | 0
sinus rhythm | 672
no conduction abnormalities | 672
no recurrent atrial fibrillation | 672
no episodes of high-grade heart block | 672
LVEF of 59% | 672
normal RV size and systolic function | 672
resolution of the pericardial effusion | 672
normal T2 signal intensity | 672