45 years old | 0
male | 0
admitted to the hospital | 0
epigastric pain | -72
abdominal tenderness | 0
elevated serum creatinine | 0
elevated blood urea | 0
abdominal CT scan with contrast | 0
chest X-ray | 0
fentanyl | 0
paracetamol | 0
fever | -96
non-productive cough | -96
dyspnea | -96
lymphopenia | -96
nasopharyngeal swab | -96
oropharyngeal swab | -96
COVID-19 diagnosis | -96
airborne isolation | -96
wheezes | -192
respiratory rate of 33 per minute | -192
heart rate of 115 beats per minute | -192
oxygen saturation 94% | -192
bilateral infiltrates | -192
elevated c-reactive protein | -192
elevated liver enzyme | -192
elevated urea | -192
elevated creatinine | -192
intubation | -192
hydroxychloroquine | -192
azithromycin | -192
tocilizumab | -192
methylprednisolone | -192
extubation | -288
discharge | 840
newly diagnosed with hypertension | 0
chronic kidney disease | 0
acute kidney injury | 0
kidney ultrasound | 0
hydration | 0
improvement of respiratory symptoms | -288
improvement of abdominal pain | -288