21 years old | 0
man | 0
evaluated in the Emergency Department | 0
rapidly progressive shortness of breath | -120
fever | -120
sore throat | -120
empiric treatment with vancomycin | 0
empiric treatment with piperacillin-tazobactam | 0
empiric treatment with azithromycin | 0
endotracheal intubation | 0
worsening hypoxemic respiratory failure | 0
acute respiratory distress syndrome | 0
CT imaging demonstrated bilateral pulmonary infiltrates | 0
CT imaging demonstrated thrombophlebitis of the left internal jugular vein | 0
blood cultures drawn on admission | 0
blood cultures grew Fusobacterium necrophorum | 0
blood cultures grew Granulicatella | 0
clinical diagnosis of septic thrombophlebitis | 0
clinical diagnosis of Lemierre syndrome | 0
antibiotics narrowed to piperacillin-tazobactam | 72
febrile | 0
worsening hypoxemia | 0
high positive end-expiratory pressure titration | 0
neuromuscular blockade | 0
vancomycin restarted | 168
repeated sampling of the respiratory system for cultures | 0
routine culture of sputum | 24
sputum culture identified normal respiratory flora | 24
BAL specimens obtained | 72
BAL specimens obtained | 168
BAL specimens revealed no growth | 72
BAL specimens revealed no growth | 168
persistent leukocytosis | 0
developed empyemas | 168
developed bilateral pneumothoraces | 168
surgical chest tube insertions | 168
bacterial culture performed on pleural fluid | 168
pleural fluid grew Mycoplasma hominis | 168
azithromycin therapy restarted | 168
fevers subsided | 216
clinically improved | 408
liberated from mechanical ventilation | 408
discharged from the hospital | 480
blood samples collected | 0
respiratory samples collected | 0
bacterial DNA sequencing performed | 0
plasma biomarkers measured | 0
endotracheal aspirates drawn | 0
endotracheal aspirates drawn | 72
endotracheal aspirates drawn | 168
sequencing of the 16S rRNA gene | 0
sequencing on the Illumina MiSeq platform | 0
analysis using custom mothur-based pipelines | 0
Fusobacterium dominated respiratory aspirates | 0
Mycoplasma taxa present | 0
repeat 16S sequencing performed | 168
Mycoplasma increased in abundance | 168
Fusobacterium decreased in abundance | 168
whole metagenome sequencing performed | 0
detection of Mycoplasma hominis | 0
detection of Fusobacterium necrophorum | 0
plasma biomarkers RAGE elevated | 0
plasma biomarkers IL-6 elevated | 0
plasma biomarkers procalcitonin elevated | 0
RAGE persistently elevated | 168
IL-6 persistently elevated | 168
procalcitonin persistently elevated | 168
RAGE decreased | 336
IL-6 decreased | 336
procalcitonin decreased | 336
negative procalcitonin levels | 240
