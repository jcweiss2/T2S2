83 years old | 0
male | 0
admitted to the hospital | 0
disorientation | 0
weakness | 0
cough | -24
prostate cancer | -672
GnRH agonist treatment | -672
fatigue | -216
itching | -216
cold intolerance | -216
whole-body edema | -216
bicalutamide | -168
silodosin | -168
antihistamine | -168
tuberculosis | -10000
transection of the left upper lobe | -10000
Hashimoto's disease in family | -10000
pale | 0
depressed level of consciousness | 0
Glasgow Coma Scale of 9 | 0
low blood pressure | 0
bradycardia | 0
hypothermia | 0
respiratory rate | 0
oxygen saturation | 0
distant heart sounds | 0
decreased breath sounds | 0
sparse hair | 0
thinning of the outer eyebrows | 0
macroglossia | 0
hoarse voice | 0
thickened skin | 0
hyperkeratosis | 0
pitting edema | 0
elevated aspartate transaminase | 0
elevated creatine kinase | 0
elevated brain natriuretic peptide | 0
sinus bradycardia | 0
low voltage in the limb and chest leads | 0
cardiomegaly | 0
normal cardiac structure and function | 0
catecholamine infusion | 0
improved hemodynamics | 24
withdrawal of catecholamine infusion | 48
deteriorated consciousness | 48
coma | 48
endotracheal intubation | 48
shock state | 48
thyroid hormone replacement | 48
levothyroxine | 48
levotriiodothyronin | 48
nasogastric tube | 48
improved general condition | 120
withdrawal hypothermia | 120
discontinued catecholamine infusion | 144
sedative agent | 168
recombinant human thrombomodulin | 168
disseminated intravascular coagulation | 168
regained full consciousness | 264
discharged from intensive-care unit | 264
extubation | 360
noninvasive positive pressure ventilation | 360
relapse of hypercapnia | 360
whole-body computed tomography | 360
acute pancreatitis | 360
elevated elastase 1 level | 360
tube feeding | 360
respiratory rehabilitation | 360
improved respiratory state | 432
ceased noninvasive positive pressure ventilation | 432
massive abdominal pain | 504
peripancreatic effusion | 504
elevated white blood cells | 504
elevated C-reactive protein | 504
broad-spectrum antibiotics | 504
septic shock | 504
death | 840
autopsy | 840
necrotic changes in the pancreatic parenchyma | 840
extensive necrotic and purulent lesions | 840
disseminated abscesses | 840
Hashimoto's thyroiditis | 840
reduction in prostate cancer | 840