68 years old | 0
male | 0
admitted to the hospital | 0
arterial hypertension | -672
dyslipidemia | -672
fever | -72
wheezing | -72
Atorvastatin | -672
Candesartan | -672
SARS-CoV-2 positive | 0
bilateral interstitial pneumonia | 0
high-resolution computed tomography | 0
blood pressure 117/74 mmHg | 0
heart rate 83 bpm | 0
peripheral oxygen saturation 79% | 0
sinus rhythm | 0
narrow QRS complex | 0
normal atrioventricular conduction | 0
no ST-T segment abnormalities | 0
Azithromycin | 0
Methylprednisolone | 0
Remdesivir | 0
Enoxaparin | 0
Insulin Lispro | 0
High Flow Nasal Cannula | 0
antihypertensive therapy discontinued | 0
statin therapy discontinued | 0
clinical status improved | 96
HRCT performed | 96
reduction of severity score | 96
sudden worsening of dyspnea | 672
increased heart rate | 672
ST-T segment morphological alterations | 672
BP 154/75 mmHg | 672
HR 85 bpm | 672
SpO2 97% | 672
ST-elevation myocardial infarction | 672
Acetylsalicylic acid | 672
Ticagrelor | 672
Bisoprolol | 672
Atorvastatin | 672
hypokinesis in the mid-apical anterior segment | 672
no evidence of intra-cardiac thrombi | 672
percutaneous coronary intervention | 675
critical stenosis of left anterior descending artery | 675
percutaneous transluminal coronary angioplasty | 675
drug eluting stent | 675
left hemiplegia | 687
National Institutes of Health Stroke Scale score 7 | 687
acute right frontal ischemic lesion | 687
fibrinolysis not performed | 687
discharged | 720
no clinical evidence of residual neurologic deficit | 744