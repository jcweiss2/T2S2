1½ years old | 0
male | 0
admitted to the hospital | 0
fever | -360
loose motions | -360
cough | -240
cold | -240
productive cough | -240
post-tussive vomiting | -240
breathlessness | -240
measles | -1095
incomplete immunization | -1095
OPV vaccine | -1095
BCG vaccine | -1095
lethargy | 0
pallor | 0
dusky | 0
shallow respiration | 0
bounding pulse | 0
low blood pressure | 0
depressed anterior fontanel | 0
dry tongue | 0
altered sensorium | 0
generalized hypotonia | 0
sluggish reflexes | 0
flexed plantar | 0
lost skin turgor | 0
malnourished | 0
protein energy malnutrition | 0
diarrhea with severe dehydration | 0
respiratory infection | 0
pallor | 0
hemoglobin 11g% | 0
leukocytosis | 0
thrombocytopenia | 0
normal liver function | 0
normal renal function | 0
negative Widal test | 0
normal X-ray chest | 0
IV fluids | 0
Inj. Cefotaxime | 0
Inj. Amikacin | 0
Inj. Calcium gluconate | 0
IV IgG | 0
ventilator | 0
Inj. Metronidazole | 96
reduced hemoglobin | 504
persistent leukocytosis | 504
low total protein | 504
low albumin | 504
another stool sample sent | 168
no Campylobacter species | 168
V. vulnificus growth | 168
sensitive to amikacin | 168
resistant to amoxicillin-clavulanic acid | 168
resistant to cefotaxime | 168
resistant to nalidixic acid | 168
resistant to co-trimoxazole | 168
resistant to tetracycline | 168
resistant to norfloxacin | 168
Klebsiella pneumoniae | 168
Acinetobacter species | 168
Inj. Imipenem | 168
Inj. Ciprofloxacin | 168
Inj. Promethazine | 168
nebulization | 168
transferred to ward | 720
Inj. Amikacin | 720
discharged | 744
stable condition | 744