19 years old | 0
male | 0
admitted to the hospital | 0
fever | -168
body ache | -168
throat pain | -168
decreased oral intake | -168
low systolic/diastolic | 0
infusing 1500 ml of normal saline | 0
broad-spectrum antibiotic | 0
inotropic support | 0
noradrenaline | 0
dengue test | 0
typhoid test | 0
malaria test | 0
leptospira test | 0
negative test results | 0
deranged KFT | 0
deranged LFT | 0
pancytopenia | 0
coagulation disturbance | 0
organomegaly | 0
hepatospenomegaly | 0
clinical hematology consultation | 0
HLH suspected | 0
further investigations | 0
hematological parameters sent | 0
coagulation parameters sent | 0
serum triglyceride sent | 0
serum fibrinogen level sent | 0
serum Ferritin sent | 0
KFT repeated | 0
LFT repeated | 0
bone marrow biopsy | 0
intubated | 0
IV methylprednisolone pulse | 0
TPE started | 0
lactate dehydrogenase | 0
fibrinogen | 0
ferritin | 0
fasting triglyceride | 0
LFT deranged | 0
KFT deranged | 0
coagulation profile deranged | 0
hemophagocytosis in bone marrow | 0
TPE procedures | 24
TPE using COM.TEC | 24
written consent | 24
benefits and risks explained | 24
standard TPE procedure | 24
plasma volume exchanges | 24
FFP used | 24
peripheral femoral line | 24
aseptic precautions | 24
organ function improved | 72
extubated | 72
Hb% improved | 72
absolute neutrophil count improved | 72
platelet count improved | 72
prothrombin time/international normalized ratio improved | 72
fibrinogen improved | 72
fasting triglyceride improved | 72
serum ferritin improved | 72
blood transfusion | 72
packed red cells | 72
FFP | 72
single donor platelet concentrates | 72
cryoprecipitate | 72
discharged | 384
hematological parameters normal | 384
biochemical parameters normal | 384
coagulation parameters normal | 384