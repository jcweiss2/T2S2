32 years old | 0
female | 0
no significant past medical history | 0
no known allergies | 0
dental abscess | -120
treated with amoxicillin/clavulanate | -120
odynophagia | -72
painful left submandibular oedema | -72
severe upper airway respiratory distress | -72
trismus | -72
extension of inflammatory signs to anterior cervical region | -72
stable vitals | -72
oxygen saturation 97% | -72
no fever | -72
leukocytosis | -72
C-reactive protein 33.36 mg/dL | -72
cervical and thoracic CT scan | -72
diffuse thickening of soft tissues | -72
phlegmon and emphysema | -72
abscess extension to submandibular, parapharyngeal and retrosternal spaces | -72
left internal jugular vein thrombosis | -72
transferred to tertiary referral centre | -48
evaluated by Maxillofacial Surgery | -48
fibreoptic nasotracheal intubation | -24
surgical drainage of abscesses | 0
admitted to Intensive Care Unit | 0
airway management | 0
daily bedside drainage of submandibular region | 0
intravenous corticosteroids | 0
empiric antibiotic therapy with ceftriaxone and metronidazole | 0
extension of vein thrombosis to brachiocephalic vein | 48
intravenous non-fractioned heparin | 48
Gram staining demonstrated polymicrobial flora | 48
abscess cultures grew Streptococcus anginosus | 72
blood cultures were sterile | 72
HIV 1/2 antibodies/antigen assay was negative | 72
all serum immunoglobulins were normal | 72
clinical and imaging improvement | 192
successful extubation | 192
transferred to infirmary for postoperative care | 192
CT reevaluation demonstrated persistence of left internal jugular vein thrombosis | 240
favourable clinical progress | 240
defervescence | 240
neck tenderness resolution | 240
recovered without sequelae | 240
discharged | 600
anticoagulation with enoxaparin | 600