39 years old | 0
man | 0
presented to the emergency department | -168
isolated episode of fever | -168
axillary temperature: 39°C | -168
diffuse myalgia | -168
pleuritic type precordial chest pain | -144
progressive dyspnea | -144
diabetes mellitus type 1 | 0
insulin treatment | 0
apyrexial | 0
dyspneic at rest | 0
respiratory rate of 24/min | 0
blood pressure of 160/90 mmHg | 0
pulse rate of 130 beats per minute | 0
distended jugular veins | 0
pericardial friction rub | 0
heart sounds not muffled | 0
pulmonary auscultation diminished sounds in bases | 0
abdominal examination unremarkable | 0
sinus tachycardia | 0
normal amplitude QRS complexes | 0
concaved ST elevation | 0
concordant T waves in DII, DIII, V4, V5, V6 leads | 0
reciprocal ST depression | 0
PR elevation in lead aVR | 0
PR depression in lead DII | 0
massively enlarged globular cardiac shadow | 0
left pleural effusion | 0
white-blood-cell count of 10,800/μl | 0
83% segmented cells | 0
9% lymphocytes | 0
hemoglobin of 10.5 g/dl | 0
platelet count of 182,000/μl | 0
CRP was 192 U/l | 0
normal renal function tests | 0
normal liver function tests | 0
NT-proBNP levels was 1155 pg/ml | 0
admitted to the intensive care unit | 0
arterial line placed | 0
pulsus paradoxus observed | 0
echocardiogram demonstrated good left ventricular function | 24
ejection fraction of 78% | 24
no valve dysfunctions | 24
massive pericardial effusion | 24
right ventricular systolic collapse | 24
cardiac tamponade | 24
pericardiocentesis performed | 24
aspiration of 160 ml purulent fluid | 24
pericardial fluid 500,000 nucleated cells/μl | 24
80% segmented cells | 24
8% lymphocytes | 24
2% eosinophils | 24
1000 red blood cells/μl | 24
lactate dehydrogenase of 19,523 U/l | 24
triglycerides of 90 mg/dl | 24
glucose of 36 mg/dl | 24
protein of 5.9 g/dl | 24
pH of 6.0 | 24
direct microbiological analysis revealed gram-positive cocci | 24
no acid-fast bacilli present | 24
vancomycin started | 24
rapid HIV test positive | 24
follow-up echocardiogram showed fluid reaccumulation | 48
right ventricular collapse | 48
urgent surgical approach indicated | 48
drain placed in pericardial sac | 48
bacterial culture set up | 48
fungal culture set up | 48
tuberculous culture set up | 48
Methicilin-sensitive S. aureus in two samples | 48
high ADA levels >200 U/l | 48
episodes of fever | 120
continuous drainage of purulent fluid | 120
tuberculostatic drugs initiated | 120
HIV positive | 120
CD4 count 28 cells/μl | 120
HIV viral load 347,609 copies/mm3 | 120
pericardial biopsy non-specific inflammation | 120
culture negative | 120
thoracic drain placed for pleural effusion | 120
no empyema | 120
chest CT no pulmonary parenchymal lesion | 120
no lymphadenopathy | 120
abdominal CT normal | 120
tuberculosis treatment | 168
fluid aspect reduced | 168
pericardial drain removed | 168
pericardial fluid cultures negative for fungal | 168
tuberculous cultures negative | 168
cytology for malignant cells negative | 168
corticosteroids not prescribed | 168
echocardiogram no fluid reaccumulation | 168
constrictive pericarditis patterns | 168
rifampin prescribed | 168
isoniazid prescribed | 168
pyrazinamide prescribed | 168
ethambutol prescribed | 168
elective pericardiectomy considered | 168
