42 years old | 0
male | 0
hypertension | -120
shortness of breath | -120
subjective fever | -120
chills | -120
cough | -120
generalized bone pain | -120
intermittent headache | -120
watery diarrhea | -120
anorexia | -120
home temperature recording of 105 °F | -120
admitted to the hospital | 0
dyspneic | 0
unable to speak in full sentences | 0
breath sounds were equal | 0
symmetrical chest wall expansion | 0
regular rhythm | 0
strong and symmetrical peripheral pulses | 0
alert and oriented | 0
no focal neurological deficits | 0
chest X-ray | 0
scattered bilateral airspace opacities | 0
sodium: 120 mEq/L | 0
potassium: 4 mEq/L | 0
blood urea nitrogen: 21 mg/dL | 0
creatinine: 1.1 mg/dL | 0
white blood cell: 13 900/µL | 0
neutrophil %: 89.4 | 0
lymphocyte %: 5.5 | 0
hemoglobin: 13.3 g/dL | 0
platelets: 250 000/µL | 0
D-dimer: 2.74 | 0
C-reactive protein: 29.32 mg/dL | 0
ferritin: 826.30 ng/mL | 0
lactate dehydrogenase: 1883 U/L | 0
interleukin-6: 224.35 pg/mL | 0
troponin <0.019 ng/mL | 0
RT-PCR nasopharyngeal swab returned positive for COVID | 0
nonrebreather mask | 0
nasal cannula | 0
ceftriaxone | 0
azithromycin | 0
hydroxychloroquine | 0
tocilizumab | 0
remdesivir | 0
severe hypoxia | 48
oxygen saturation to the 60s | 48
intubated | 48
hypotension | 48
vasopressor therapy | 48
lactate remained below 2.5 | 48
serum creatinine remained below 0.8 mg/dL | 48
troponinemia worsened | 48
heparin drip | 48
fluctuating hypoxia | 48
sedatives | 48
paralytics | 48
febrile | 48
pressor support | 48
duplex study | 72
no deep vein thrombosis | 72
transthoracic echocardiography | 72
no intracavitary thrombus | 72
diminished pupillary reflexes | 144
mid-dilated pupils | 144
no corneal or oculocephalic reflexes | 144
computed tomography head | 144
large ischemic infarcts | 144
bilateral occipital | 144
left parietal | 144
right temporal | 144
right frontal lobes | 144
downward herniation | 144
CT chest with angiography | 144
extensive multifocal dense ground-glass opacities | 144
no PE | 144
pronounced dead | 168