19 years old | 0
male | 0
head injury | -1
sound gun trauma | -1
increased intracranial pressures | -1
cerebellar damage | -1
admitted to ICU | 0
unconscious | 0
intubated | 0
Glasgow coma score 3E | 0
skin incision | 0
soft tissue defects | 0
light and corneal reflexes negative | 0
no spontaneous breathing | 0
heart rate 56 beats/min | 0
blood pressure 80/40 mmHg | 0
body temperature below 36°C | 0
central venous pressure 1 cm H2O | 0
brain CT | 0
bone fragments in right temporal region | 0
hemorrhagic contusion area | 0
edema in right frontotemporal area | 0
mechanical ventilation | 0
low blood pressure | 0
central venous pressure | 0
crystalloid fluid administration | 0
dopamine infusion | 0
mannitol therapy | 0
furosemide administration | 0
metoclopramide HCl administration | 0
famotidine administration | 0
acetylcysteine administration | 0
normal blood biochemistry values | 0
toxicological evaluation | 0
no emergency operation | 0
noradrenaline infusion | 24
nutritional status assessment | 24
enteral feeding | 24
eye opening and closing | 48
blinking | 48
light and corneal reflex positive | 48
no spontaneous limb movement | 48
no response to pain stimuli | 48
percutaneous tracheotomy | 120
LIS diagnosis | 168
vertical eye movements | 168
quadriplegia | 168
brain CT repeated | 168
minimal pressure in pons and mesencephalon | 168
partial compression in fourth ventricle | 168
hyperdense area in cerebellum | 168
MRI planned | 168
antibiotic treatment | 168
pulmonary edema | 168
acute respiratory distress syndrome | 168
ventilation modes adjusted | 168
melena | 408
decrease in Hb and htc | 408
blood and blood product replacement | 408
omeprazole administration | 408
death | 864
multiorgan failure | 864
postmortem macroscopic examination | 864
ischemia in cerebellum | 864
vertebrobasilar artery system normal | 864