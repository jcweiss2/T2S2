4 years old | 0
female | 0
developmental delay | -8760
myelomeningocele | -8760
hydrocephalus | -8760
neurogenic bladder | -8760
recurrent urinary tract infections | -8760
admitted to hospital for urosepsis | -720
hemolytic uremic syndrome | -720
chronic renal failure | -720
discharged on peritoneal dialysis | -720
seizure-like activity | -48
fever | -48
distended abdomen | -48
tachycardic | -48
tachypneic | -48
normal oxygen saturations on room air | -48
given lorazepam | -48
given fosphenytoin | -48
given antibiotics | -48
transferred to facility | -48
chest x-ray performed | -24
enlarged cardiac silhouette | -24
suspicious for tamponade | -24
transthoracic echocardiogram performed | -12
moderate circumferential pericardial effusion | -12
diastolic right atrial collapse | -12
tamponade physiology | -12
taken to catheterization laboratory | 0
endotracheal intubation | 0
6-French pigtail catheter placed | 0
220 ml of serosanguineous fluid drained | 0
patient stabilized | 24
pericardial drainage minimal | 48
decision to discontinue drain | 48
attempted removal of drain | 48
patient became unresponsive | 48
decreased respiratory rate | 48
bradycardia | 48
chest compressions initiated | 48
patient ventilated via bag mask | 48
patient started breathing spontaneously | 48
palpable pulse | 48
bedside chest x-ray performed | 48
transferred to operating room | 72
TTE-guided withdrawal of drain | 72
patient became profoundly hypotensive | 72
bradycardic | 72
external cardiac compressions initiated | 72
0.35 flex guidewire passed into catheter | 72
catheter and wire advanced back into chest | 72
patient stabilized hemodynamically | 72
decision to remove catheter under direct visualization | 72
sternotomy performed | 72
catheter found to course around pulmonary artery and aorta | 72
traction on catheter resulted in complete occlusion of main pulmonary artery | 72
severe reduction in pulmonary blood flow | 72
abrupt fall in end-tidal carbon dioxide | 72
drain surgically removed | 72
patient recovered in pediatric intensive care unit | 120