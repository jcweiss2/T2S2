50 years old | 0
female | 0
celiac disease | 0
iron deficiency anemia | 0
hypothyroidism | 0
admitted to the medical ward | 0
chronic febrile illness | 0
drenching night sweats | 0
fungal esophagitis | 0
antifungal medication | 0
frequent nausea | 0
no vomiting episodes | 0
normal bowel motion | 0
CT scan | 0
incidental tumor finding | 0
liver lesions | 0
mild pericardial effusion | 0
echocardiogram | 0
normal ejection fraction | 0
liver lesion biopsy | 0
GIST diagnosis | 0
referred to medical oncologist | 0
imatinib 400 mg daily | -2160
generalized fatigability | -2160
symptomatic anemia | -2160
bleeding tumor | -2160
multiple transfusions | -2160
follow-up CT scan | -2160
tumor progression | -2160
started sunitinib | -2160
hospital stay | 0
echocardiography | 0
persistent tachycardia | 0
small pericardial effusion | 0
high ejection fraction | 0
presented to emergency department | 24
generalized abdominal pain | 24
multiple vomiting episodes | 24
no bowel motion | 24
tachycardic | 24
tachypneic | 24
nasal cannula oxygenation | 24
generalized abdominal tenderness | 24
guarding | 24
rigid abdomen | 24
significant rise in lactate level | 24
unremarkable laboratory test | 24
sinus tachycardia | 24
CT scan abdomen | 24
ischemic jejunal loops | 24
pneumoperitoneum | 24
emergency laparotomy | 24
turbid intraperitoneal fluid | 24
large mid-jejunal mass | 24
adherent mass | 24
bowel perforation | 24
edematous bowel | 24
mass resection | 24
small bowel resection | 24
side-to-side anastomosis | 24
hypotension episodes | 24
intraoperative pericardial window | 24
200 mL serous fluid drained | 24
intraperitoneal drains inserted | 24
extubated | 24
transferred to ICU | 24
adjuvant Regorafenib | 24
adjuvant Pazopanib | 24
unsuccessful chemotherapy | 24
liver metastasis | 24
obstructive phenomena | 24
PTC required | 24
passed away | 24
histopathological examination | 24
GIST 12x11x9cm | 24
mitotic rate 11 MF/50 HPF | 24
negative mesenteric lymph node | 24
CD117 immunoreactive | 24
DOG1 immunoreactive | 24
high-grade anaplastic areas | 24
