60 years old | 0
male | 0
admitted to the hospital | 0
diffuse itchy skin | -168
eczema-like symptoms | -168
vitiligo | -6720
anemia | -6720
occupational exposures | -6720
smoker | -6720
alcohol use | -6720
dermatitis | -504
topical nystatin | -504
nummular eczema | -168
topical hydrocortisone | -168
cetirizine | -168
naproxen | -168
oral prednisone | -168
unremitting itching | -168
edematous nasal mucosal | -168
posterior oropharyngeal erythema | -168
maculopapular erythematous rash | -168
topical triamcinolone | -168
hydroxyzine | -168
persistent intense pruritus | -84
lesions on face, chest, and abdomen | -84
sarcoidosis | -84
lichen planus | -84
disseminated lupus erythematosus | -84
lymphoma | -84
syphilis | -84
punch biopsies | -84
CTCL | -84
CD3+ | -84
CD4+ | -84
CD8+ | -84
CD4:CD8 ratio > 2:1 | -84
loss of CD7 lymphocyte staining | -84
CD20 | -84
CD30+ | -84
Treponema pallidum stain | -84
T-cell gene rearrangement | -84
atypical lymphoid epidermal infiltrate | -84
irregular nuclear contour | -84
dermal/epidermal junction | -84
inflammatory dermal infiltrate | -84
CT/PET scan | -56
moderately avid and enlarged bilateral axillary, inguinal, and supraclavicular lymph nodes | -56
pathology from lymph node biopsy | -56
CTCL | -56
tumor staging | -56
IVA2 | -56
T4N3M0B0 | -56
doxepin | -56
warfarin | -56
second opinion | -28
Cleveland Clinic Oncology | -28
clobetasol | -28
desonide | -28
oral bexarotene | -28
gabapentin | -28
bilateral foot pain and swelling | -12
lower extremity duplex | -12
extreme pain | 0
open skin wounds | 0
yellow-green fluids | 0
large eschar | 0
foul-smelling fluid | 0
excoriating wounds | 0
broad-spectrum antibiotics | 0
CT chest/abdomen/pelvis | 0
axillary adenopathy | 0
enlarged bilateral inguinal and external iliac chain lymph nodes | 0
subcutaneous lesions | 0
skin cultures | 0
MRSA | 0
Diphtheroid | 0
left inguinal lymph node excision | 48
left anterior abdominal wall biopsy | 48
debridement of chest wall eschar | 48
large cell transformation | 48
romidepsin | 48
COVID-19 | 48
discharge to SNF | 336
diffuse large lesions | 672
purulent foul-smelling discharge | 672
excruciating pain | 672
infected skin lesions | 672
admission to ED | 672
aggressive pain management | 672
broad-spectrum antibiotic therapy | 672
romidepsin held | 672
extensive excisional debridement | 696
necrotic tissue | 696
MRSA | 696
group B Streptococcus bacteremia | 696
T4N3M0B1 | 696
mechanical ventilation | 696
surgical ICU | 696
critically hypotensive | 720
decreased urine output | 720
leukocytosis | 720
group G streptococcus | 720
MRSA bacteremia | 720
spontaneous breathing trial | 720
code status changed to DNR | 816
comfort care only | 816
extubated | 816
expired | 864