62 years old | 0
female | 0
admitted to the hospital | 0
history of UC | -12
5-aminosalicylic acid | -12
acute severe flare of UC | -168
infliximab | -168
computed tomography | -168
perinuclear anti-neutrophilic cytoplasmic antibody | -168
antinuclear antibody | -168
breast carcinoma | -36
family history of UC | -12
fever | 0
cough | 0
vomiting | 0
diarrhea | 0
generalized weakness | 0
confusion | 0
lethargy | 0
low Glasgow coma scale | 0
mild neck stiffness | 0
elevated C-reactive protein | 0
stable hemoglobin | 0
negative Coronavirus disease 2019 | 0
lower respiratory tract infection | 0
piperacillin/tazobactam | 0
admitted to the intensive care unit | 0
positive blood cultures for L. monocytogenes | 24
listeriosis | 24
bacterial meningitis | 24
lumbar puncture | 24
grossly cloudy cerebrospinal fluid | 24
elevated white blood cell count | 24
low cerebrospinal fluid glucose | 24
raised cerebrospinal fluid protein | 24
discharged from intensive care unit | 168
flare of colitis | 744
Mayo 3 endoscopic appearance | 744
vedolizumab | 744
colectomy | 912
subtotal colectomy | 912
unremarkable post-surgical course | 936