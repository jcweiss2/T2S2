81 years old | 0
man | 0
admitted to a primary hospital | 0
lower abdominal pain | 0
bloody diarrhea | 0
no specific past medical history | 0
abdominal computed tomography | 0
thickness of the descending colon wall | 0
intravenous hydration | 0
antibiotic therapy | 0
cefotiam | 0
levofloxacin | 0
ischemic colitis | 0
hospital day 2 | 48
follow-up abdominal computed tomography | 48
ascites | 48
thickness of the entire colon wall | 48
hospital day 4 | 96
transferred to our hospital | 96
renal dysfunction | 96
convulsion | 96
first aid station | 96
patient's consciousness was slightly clouded | 96
temperature 38.0°C | 96
blood pressure 140/92 mm Hg | 96
heart rate 95/min | 96
skin was cold and moist | 96
abdomen was distended | 96
abdomen was tympanic | 96
generalized tenderness | 96
severe inflammation | 96
anemia | 96
low platelet count | 96
blood gas analysis | 96
hypoxemia | 96
metabolic acidosis | 96
low CO2 level | 96
tachypnea | 96
colonoscopy | 96
diffuse mucosal edema | 96
ulcer formation | 96
bleeding from the rectum to the ascending colon | 96
no evidence of free air | 96
whole colon wall was markedly thickened | 96
huge ascites | 96
gradually, patient's vital signs deteriorated | 96
blood pressure 60/40 mm Hg | 96
heart rate 115/min | 96
severe disturbance of consciousness | 96
generalized cyanosis | 96
necrotic ischemic colitis | 96
septic shock | 96
emergency surgery | 96
operative findings | 96
large amount of ascites | 96
colon wall was markedly edematous and sclerotic | 96
inflammation of the transverse colon | 96
necrosis | 96
extended right hemicolectomy | 96
ileostomy | 96
resected specimen | 96
hemorrhagic necrosis of the transverse colon | 96
pathological findings | 96
mucosal hemorrhagic necrosis | 96
submucosal edema | 96
venous dilatation | 96
congestion of blood | 96
ischemic colitis | 96
stool culture | 96
O157 | 96
verotoxin | 96
hemorrhagic colitis | 96
HUS | 96
acute encephalopathy | 96
O157 infection | 96
after the operation | 96
treated in the intensive care unit | 96
ventilation | 96
delayed emergence from anesthesia | 96
encephalopathy | 96
poor oxygenation | 96
intensive care | 96
HUS improved | 96
encephalopathy improved | 96
no dialysis | 96
discharged | 792
