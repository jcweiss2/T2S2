45 years old | 0
    female | 0
    admitted to the hospital | 0
    shortness of breath | -48
    malaise | -1440
    lethargy | -1440
    slow speech | -1440
    edema of the face | -1440
    edema of the extremities | -1440
    progressive weight gain | -1440
    no history of medical illness | -1440
    no drug history | -1440
    temperature 36°C | 0
    blood pressure 90/52 mmHg | 0
    heart rate 74 beats/min | 0
    BMI 32.6 kg/m² (obese) | 0
    hypothermic | 0
    pulsus paradoxus | 0
    facial edema | 0
    coarse hair | 0
    dry skin | 0
    engorged jugular vein | 0
    mild pallor | 0
    non-pitting edema of the extremities | 0
    oxygen saturation 84% | 0
    cardiac apical impulse not visible | 0
    apex beat not felt | 0
    soft and distant heart sounds | 0
    bilateral basal rales | 0
    mild hepatomegaly | 0
    delayed relaxation of deep reflexes | 0
    chest radiogram cardiomegaly with globular enlargement | 0
    electrocardiogram low voltage pattern with electrical alternans | 0
    echocardiogram massive pericardial effusion | 0
    early diastolic RV collapse | 0
    swinging motion of heart | 0
    prominent respiratory alteration of RV dimension | 0
    right atrial and RV collapse during diastole | 0
    pericardial effusion all around | 0
    small cardiac chambers | 0
    predominant diastolic heart failure | 0
    right ventricular diastolic collapse | 0
    diagnosis of large pericardial effusion | 0
    diagnosis of cardiac tamponade | 0
    pericardiocentesis procedure | 0
    450 ml pericardial fluid tapped | 0
    pericardial fluid yellowish golden | 0
    oxygen saturation increased to 94% | 0
    post-pericardiocentesis chest radiogram reduced cardiomegaly | 24
    post-pericardiocentesis echocardiogram minimal pericardial effusion | 24
    thyroid function test high TSH | 24
    thyroid function test low T3 | 24
    thyroid function test low T4 | 24
    treated with thyroxine 100 μg daily | 24
    thyroxine increased to 200 μg daily | 336
    discharged after 2 weeks | 336
    follow-up echocardiogram after 3 months | 2160
    near total resolution of pericardial effusion | 2160
    symptoms and signs disappeared | 2160
    Hb 11.5 g% | 0
    ESR 24 | 0
    total leukocyte count 9850 mm³ | 0
    platelet count 2.1 lac | 0
    BUL 24 mg% | 0
    serum creatinine 1.1 mg% | 0
    LFT normal | 0
    TSH 84 mU/ml | 0
    T3 26.2 ng/dl | 0
    T4 0.56 μg/dl | 0
    total cholesterol 317 mg/dl | 0
    HDL-C 52 mg/dl | 0
    triglyceride 214 mg/dl | 0
    serum sodium 136 mEq/l | 0
    serum potassium 4.2 mEq/l | 0
    HIV negative | 0
    HbSAg negative | 0
    pericardial fluid lymphocytes 8–10/mm³ | 0
    pericardial fluid proteins 4.7 g% | 0
    pericardial fluid sugar 80 mg% | 0
    pericardial fluid cholesterol 192 mg% | 0
    no organisms grown on culture | 0

<|eot_id|>

