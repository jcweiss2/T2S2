38 years old | 0
male | 0
agammaglobulinaemia | 0
non-compliance with monthly immunoglobulin administration | -672
presented to emergency department | 0
worsening dyspnoea | -24
productive cough | -24
recent fever | -24
tachycardic | 0
tachypnoeic | 0
febrile | 0
body temperature 38.7°C | 0
blood pressure 78/51 mmHg | 0
oxygen saturation 85% | 0
placed on non-rebreather mask | 0
aggressive fluid resuscitation | 0
chest X-ray infiltrates left lower lobe | 0
mild left pleural effusion | 0
community-acquired pneumonia diagnosis | 0
septic shock diagnosis | 0
ceftriaxone initiation | 0
clarithromycin initiation | 0
arterial oxygen pressure 65 mmHg | 0
persistent hypoxaemia | 0
worsening respiratory distress | 0
transferred to ICU | 0
sedated | 0
intubated | 0
ventilated | 0
chest X-ray increasing left pleural effusion | 0
chest tube insertion | 0
drained empyema | 0
persistent hypotension | 0
norepinephrine initiation | 0
haemodynamic stability restored | 0
urine output improving | 0
CT scan thorax homogeneous density air bronchogram left upper lobe | 48
lingula involvement | 48
left lower lobe involvement | 48
Gram stain sputum Gram-negative bacilli | 48
aerobic blood cultures Gram-negative coccobacilli | 48
identified as A. calcoaceticus | 48
sensitive to ceftazidime | 48
sensitive to cefepime | 48
sensitive to colistin | 48
sensitive to tigecycline | 48
sensitive to meropenem | 48
sensitive to piperacillin | 48
sensitive to cotrimoxazole | 48
sensitive to ciprofloxacin | 48
negative influenza viruses A and B | 48
negative pneumococcus urinary antigen | 48
negative Legionella urinary antigen | 48
intravenous immunoglobulins administered | 24
C-reactive protein peak 271 mg/L | 48
procalcitonin peak 16.22 ng/mL | 48
colistin initiation | 48
cefepime initiation | 48
pressors stopped | 72
weaned off mechanical ventilation | 72
extubated | 72
imaging minimal left pleural effusion | 72
chest tube removed | 72
ciprofloxacin initiation | 72
discharged | 336
ciprofloxacin continued for 2 weeks | 336
clinical stability maintained | 336
