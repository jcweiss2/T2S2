78 years old | 0
    male | 0
    admitted to the intensive care unit | 0
    acute respiratory distress | 0
    acute diastolic decompensation | 0
    started on 50% oxygen via mask | 0
    nothing by mouth | 0
    enoxaparin | 0
    amiodarone | 0
    digoxin | 0
    respiratory failure | 0
    intubated | 0
    mild leukocytosis | 0
    hemoglobin 9.1 g/dL | 0
    hematocrit 27.6% | 0
    platelet 468.0 K/uL | 0
    serum chemistries within normal limits | 0
    urine cultures | 0
    sputum cultures | 0
    three sets of blood cultures | 0
    treated empirically for septic shock | 0
    intravenous vancomycin | 0
    cefepime | 0
    clindamycin | 0
    computed tomography demonstrated persistent esophageal leakage of contrast | 0
    bronchopulmonary fistula | 0
    blood cultures positive for A. israelii | 0
    esophageal rupture | - (prior to admission)
    COPD | - (prior to admission)
    atrial fibrillation | - (prior to admission)
    Clostridium difficile infection | - (prior to admission)
    empyema with mediastinitis | - (prior to admission)
    esophageal repair | - (prior to admission)
    gastrostomy tube insertion | - (prior to admission)
    sudden onset respiratory distress | - (en route to facility)
    chest pain | - (en route to facility)
    back pain | - (en route to facility)
    hypotension | - (en route to facility)
    tachycardia | - (en route to facility)
    decreased bilateral air entry | 0
    dullness to percussion of the right lung | 0
    respiratory distress | - (en route to facility)
    septic shock | 0
    surgical debulking | - (prior to admission)
    relapse | - (future potential event)
    penicillin therapy | - (future treatment)
    surgical resection | - (future potential event)
    oral penicillin therapy | - (future treatment)
    <|eot_id|>
    78 years old | 0
male | 0
admitted to the intensive care unit | 0
acute respiratory distress | 0
acute diastolic decompensation | 0
started on 50% oxygen via mask | 0
nothing by mouth | 0
enoxaparin | 0
amiodarone | 0
digoxin | 0
respiratory failure | 0
intubated | 0
mild leukocytosis | 0
hemoglobin 9.1 g/dL | 0
hematocrit 27.6% | 0
platelet 468.0 K/uL | 0
serum chemistries within normal limits | 0
urine cultures | 0
sputum cultures | 0
three sets of blood cultures | 0
treated empirically for septic shock |3 0
intravenous vancomycin | 0
cefepime | 0
clindamycin | 0
computed tomography demonstrated persistent esophageal leakage of contrast | 0
bronchopulmonary fistula | 0
blood cultures positive for A. israelii | 0
esophageal rupture | - (prior to admission)
COPD | - (prior to admission)
atrial fibrillation | - (prior to admission)
Clostridium difficile infection | - (prior to admission)
empyema with mediastinitis | - (prior to admission)
esophageal repair | - (prior to admission)
gastrostomy tube insertion | - (prior to admission)
sudden onset respiratory distress | - (en route to facility)
chest pain | - (en route to facility)
back pain | - (en route to facility)
hypotension | - (en route to facility)
tachycardia | - (en route to facility)
decreased bilateral air entry | 0
dullness to percussion of the right lung | 0
respiratory distress | - (en route to facility)
septic shock | 0
surgical debulking | - (prior to admission)
relapse | - (future potential event)
penicillin therapy | - (future treatment)
surgical resection | - (future potential event)
oral penicillin therapy | - (future treatment)