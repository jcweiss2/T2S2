40 years old | 0
male | 0
admitted to the hospital | 0
multiple gunshots to the chest, abdomen, and pelvis | -1
resuscitative thoracotomy | 0
emergent exploratory laparotomy | 0
splenectomy | 0
direct repair of enterotomies | 0
gastrotomy | 0
traumatic IVC injury | 0
abdominal packing | 0
temporary abdominal closure | 0
mass transfusion protocol | 0
transferred to the surgical trauma intensive care unit | 0
high sanguineous output from abdominal wound | 7
hemodynamically unstable | 7
noticeable hemoperitoneum | 7
increasing drain output | 7
vascular surgery consulted | 7
multidisciplinary team meeting | 7
decision to proceed with IVC venogram | 7
IVC venogram with possible repair | 7
activated semihybrid circulatory dynamics laboratory | 7.34
ultrasound-guided access of the right femoral vein | 7.52
8F sheath placed | 7.52
IVC venogram obtained | 7.52
substantial blush within the suprarenal IVC | 7.52
IVUS probe advanced into the IVC | 7.52
measurements taken at the proximal and distal sites of the IVC injury | 7.52
Gore TAG 28.5-mm × 3.3-cm endograft cuff deployed | 7.52
completion venogram obtained | 7.52
tilting of the first cuff with an incomplete seal | 7.52
second Gore TAG endograft cuff deployed | 7.52
complete seal obtained | 7.52
access site closed | 7.52
coagulation panel ordered | 9.34
returned to the trauma intensive care unit | 9.34
abdominal washout | 24
follow-up computed tomography scan | 336
no stent graft migration or extravasation | 336
discharged home | 168
prescription for daily 75 mg clopidogrel and 81 mg aspirin | 168
follow-up at 30 days | 720