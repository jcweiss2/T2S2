39 years old | 0
    female | 0
    ingested ∼500 caffeine tablets | 0
    dissolved in water | 0
    caffeine overdose | 0
    generalized tonic–clonic seizure | -60
    treated by emergency medical service | -60
    three episodes of broad complex tachycardia | -60
    cardiopulmonary resuscitation | -60
    defibrillations | -60
    epinephrine | -60
    amiodarone | -60
    intubated | 0
    sinus rhythm | 0
    blood pressure 62/33 mmHg | 0
    heart rate 140/min | 0
    activated charcoal administered | 0
    multiple ventricular extrasystoles | 0
    intravenous magnesium | 0
    intravenous calcium | 0
    hypotension | 0
    received 9 L crystalloids | 0
    repeated epinephrine boluses | 0
    continuous epinephrine infusion | 0
    lactic acidosis | 0
    intravenous sodium bicarbonate | 0
    haemodialysis initiated | 300
    cardiovascular instability | 300
    lactic acidosis persisted | 300
    epinephrine replaced by dobutamine | 300
    hypotension-induced acute renal failure | 336
    rhabdomyolysis-induced acute renal failure | 336
    creatine kinase max 69 885 U/L | 336
    aspartate transaminase max 1908 U/L | 336
    volume overload | 336
    persistent haemodynamic instability | 336
    chronic venoBvenous haemodiafiltration initiated | 336
    haemodialysis therapy recommenced | 504
    pulmonary failure | 504
    tricuspid endocarditis | 504
    line sepsis | 504
    renal function improved | 504
    haemodialysis therapy stopped | 504
    caffeine serum concentration 2.95 mmol/L | 0
    survived caffeine overdose | 0
    lethal dose caffeine | 0
    serum caffeine concentrations measured | 0
    toxic effects central nervous system | 0
    adrenergic effects | 0
    tachyarrhythmias | 0
    vasodilation | 0
    hypotension persisted | 0
    hypokalaemia | 0
    leucocytosis | 0
    glycogenolysis | 0
    lipolysis | 0
    lactic acidosis caused by shock-induced tissue hypoxia | 0
    rhabdomyolysis | 0
    caffeine demethylated to paraxanthine | 0
    theobromine | 0
    theophylline | 0
    hepatic cytochrome P450 CYP1A2 system involved | 0
    plasma protein binding of caffeine 36% | 0
    caffeine removed by haemodialysis | 0
    disequilibrium syndrome risk | 0
    toxin removal principle | 0
    line sepsis risk | 0
    tricuspid endocarditis risk | 0
    haemodialysis advocated for severe caffeine intoxication | 0
    clinical course complications | 0
    repeated haemodialysis sessions benefit | 0

<|eot_id|>