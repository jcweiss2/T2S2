72 years old | 0
woman | 0
history of bilateral breast cancers | 0
unusual occipital neck mass | 0
presented to the emergency department | 0
complained of shortness of breath | 0
haemoglobin of 4.2 g/dl | 0
cyst developed after minor trauma in 1967 | -168
mass started to grow over the past few years | -24000
mass periodically drain | -24000
mass scab over | -24000
mass drain again | -24000
mass began to bleed | -24000
portion of the mass fallen out | -120
mass bled more profusely | -120
developed severe diffuse swelling in arms | -240
developed severe diffuse swelling in legs | -240
developed severe diffuse swelling in trunk | -240
afebrile | 0
haemodynamically stable | 0
hypertensive to 170/70 mmHg | 0
oxygen saturation of 100% on 4-l nasal cannula | 0
clear lung sounds | 0
severe upper extremity pitting oedema | 0
severe lower extremity pitting oedema | 0
baseball-sized malodorous occipital mass | 0
mass soft to touch | 0
thick oozing purulent drainage | 0
white blood cell count of 8.3*103/μl | 0
haemoglobin of 4.7 g/dl | 0
albumin of 2.9 g/dl | 0
INR of 1.6 | 0
B-type natriuretic peptide level of 666 pg/ml | 0
chest X-ray showed mild interstitial oedema | 0
severe anaemia | 0
recurrent bleeding from the neck mass | 0
cause of shortness of breath | 0
primary differential for anasarca included nephrotic syndrome | 0
primary differential for anasarca included cirrhosis | 0
primary differential for anasarca included liver metastases | 0
mass suspicious for malignancy | 0
CT pan-scan ordered | 0
patient not able to tolerate CT pan-scan | 0
remained in the emergency department for more than 24 h | 24
transfused three units of packed red blood cells | 0
became febrile to 101.2 °F | 24
became tachycardic to 110 bpm | 24
fever ascribed to transfusion reaction | 24
acetaminophen ordered | 24
temperature increased to 102 °F | 24
heart rate increased to 120 bpm | 24
tachypnoeic to 30 breaths per minute | 24
hypertensive to 200/60 mmHg | 24
lactate level of 2.7 mEq/l | 24
white blood cell count of 24.3*103/μl | 24
6% band forms | 24
blood cultures grew E. coli | 24
started on vancomycin | 24
started on piperacillin–tazobactam | 24
creatinine doubled from 0.72 mg/dl to 1.46 mg/dL | 24
INR of 2.4 | 24
platelet count fell from 127*103/μl to 86*103/μl | 24
fibrinogen of 224 mg/dl | 24
d-dimer level of 4668 ng/ml | 24
disseminated intravascular coagulation secondary to severe sepsis | 24
breathing became increasingly laboured | 24
placed on bilevel non-invasive positive pressure ventilation | 24
transferred to medical intensive care unit | 24
hypotensive to 80/40 mmHg | 24
vasopressors initiated | 24
urinalysis notable for pyuria with greater than 180 white blood cells per hpf | 24
intubated | 24
sedated | 24
pan-CT scan performed | 24
obstructing left distal ureteric stone measuring up to 1.6 cm | 24
proximal dilation | 24
hydronephrosis | 24
taken to operating room for extraction and stenting | 24
weaned from vasopressors | 24
could not be extubated for a day | 24
chest X-ray showed increasing pulmonary oedema | 24
became oliguric | 24
creatinine elevated to 6.4 mg/dl | 24
urgently dialyzed | 24
stabilized | 24
transferred back to general medicine service after ten days | 240
discharged from the hospital on day 28 | 672
required haemodialysis for several months | 2160
kidney function recovered | 2160
neck mass excised | 2160
pathology showed benign haemangioma | 2160
infected haematoma | 2160
abscess formation | 2160
severe sepsis due to urinary tract infection | 24
urinary tract infection caused by obstructing ureteric stone | 24
