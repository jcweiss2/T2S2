67 years old | 0
female | 0
hypertension | 0
type 2 diabetes mellitus | 0
dyslipidemia | 0
abdominal pain | -72
bleeding diarrhoea | -72
nausea | -72
admitted to emergency department | 0
blood pressure 95/71 mmHg | 0
temperature 36.3 °C | 0
oxygen saturation 92% | 0
diffuse abdominal painful | 0
leucocytes count 7.3 × 10^3 μL | 0
haemoglobin 12.6 g/dL | 0
platelet count 96 × 10^3 μL | 0
serum creatinine 1.45 mg/dL | 0
serum sodium 132 mmol/L | 0
serum potassium 4.5 mmol/L | 0
diagnosed of acute gastroenteritis | 0
treated with fluids | 0
treated with proton pump inhibitor | 0
treated with antiemetics | 0
treated with intravenous antibiotic therapy | 0
anuria | 0
unfavourable evolution on blood test | 0
abdominal CT scan | 24
proctitis | 24
cortical hypoperfusion of both kidneys | 24
admitted to intensive care unit | 72
neurological failure | 72
bradipsiquia | 72
anuria | 72
worsen of blood test analysis | 72
haemoglobin 11.2 g/dL | 72
haptoglobin < 6.63 mg/dL | 72
lactate dehydrogenase 1125 U/L | 72
elevated schistocytes count on blood smear | 72
negative direct antiglobulin test | 72
diagnosed of microangiopathic haemolytic anemia | 72
thrombocytopenia | 72
diagnosed of TMA | 72
treated with urgent plasma exchange | 72
treated with methylprednisolone | 72
haemodialysis | 72
ADAMTS13 test | 96
normal ADAMTS13 levels | 96
maintenance of plasma exchange | 96
complement c3 levels on low limit of normal range | 96
isolation of verotoxin 2-secreting Escherichia Coli | 120
discontinuation of plasma exchange | 120
favourable clinical evolution | 120
progressive improvement of neurological symptoms | 120
transferred to ward | 120
recovery of diuresis | 336
renal biopsy | 336
histological changes compatible with thrombotic microangiopathic involvement | 336
anaemia increased | 144
red-cell transfusion | 144
platelet transfusion | 72
discharged | 672