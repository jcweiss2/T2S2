3 years old | 0
female | 0
admitted to the hospital | 0
fever | -72
respiratory distress | -72
family history of secondary parental consanguinity | 0
sibling died from fever | -6300
cousin died due to unknown cause | -13140
ampicillin-sulbactam treatment | 0
azithromycin treatment | 0
COVID-19 PCR negative | 0
low consciousness level | 0
confusion | 0
high blood pressure | 0
crackles in both lungs | 0
deep tendon reflexes normoactive | 0
light reflex normal | 0
COVID-19 PCR positive | 168
hydroxychloroquine treatment | 168
favipiravir treatment | 168
intubated | 72
ventilated | 72
hemoglobin level 6.5 g/dl | 72
white blood cell count 16 160/mm3 | 72
platelet count 503 000/mm3 | 72
blood urea nitrogen 44 mg/dl | 72
creatinine 0.8 mg/dl | 72
AST 65 U/l | 72
ALT 57 U/l | 72
total bilirubin 0.68 mg/dl | 72
sedimentation rate 60 mm/hour | 72
D-dimer 5820 µg/l | 72
thorax computerized tomography (CT) showed bilateral effusion and atelectasis | 72
pleural effusion resolved | 168
marked consolidation areas and ground glass opacities | 168
teicoplanin treatment | 168
cefotaxime treatment | 168
amlodipine treatment | 96
esmolol infusion | 96
furosemide infusion | 96
albumin transfusion | 96
peripheral blood smear showed 64% polymorphonuclear leukocytes | 120
bone marrow aspiration | 120
normocellular bone marrow | 120
renal Doppler ultrasound | 120
left ventricular hypertrophy | 120
mitral insufficiency | 120
azithromycin stopped | 120
cefotaxime tapered to meropenem | 120
intravenous immunoglobulin (IVIG) | 168
erythrocyte transfusions | 168
anuric | 240
thrombocytopenia | 240
microangiopathic hemolytic anemia | 240
HUS diagnosis | 240
schistocytes | 240
ADAMTS-13 activity level normal | 240
disseminated intravascular coagulation ruled out | 240
plasmapheresis | 240
hemodialysis | 240
extubated | 336
urine output increased | 336
LDH values decreased | 336
blood pressure reduced | 336
platelet count increased | 336
oral antihypertensive medication | 336
asymptomatic | 672
hemodynamic parameters normalized | 672
discharged | 672
oral antihypertensive treatment discontinued | 840
control CT | 1008
sequelae pleuroparenchymal shrinkage | 1008
faintly circumscribed, slightly ground glass densities | 1008