24 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
severe headache | -72 | 0 | Factual
projectile vomiting | -72 | 0 | Factual
no fever | -72 | 0 | Negated
no convulsions | -72 | 0 | Negated
no focal neurological deficit | -72 | 0 | Negated
symptomatic treatment outside | -72 | 0 | Factual
no relief | -72 | 0 | Factual
admission to hospital | 0 | 0 | Factual
provisional diagnosis of metabolic encephalopathy | 0 | 0 | Possible
symptomatic treatment | 0 | 0 | Factual
altered sensorium | 0 | 24 | Factual
Glasgow Coma Scale-9 | 0 | 24 | Factual
high-grade fever | 0 | 24 | Factual
chills | 0 | 24 | Factual
transfer to intensive care unit | 0 | 24 | Factual
dyselectrolytemia | 0 | 24 | Factual
low serum phosphate | 0 | 24 | Factual
neutrophilic leukocytosis | 0 | 24 | Factual
cerebrospinal fluid sent for evaluation | 0 | 24 | Factual
empirical treatment with ceftriaxone | 0 | 24 | Factual
Gram stain of CSF | 0 | 24 | Factual
polymorphs and lymphocytes in CSF | 0 | 24 | Factual
Gram-positive bacilli in CSF | 0 | 24 | Factual
culture of CSF | 0 | 24 | Factual
Listeria monocytogenes in CSF | 0 | 24 | Factual
blood culture at admission | 0 | 0 | Factual
Gram-positive bacilli in blood culture | 0 | 0 | Factual
Listeria monocytogenes in blood culture | 0 | 24 | Factual
switch to meropenem | 24 | 24 | Factual
clinical improvement | 24 | 48 | Factual
microbiological improvement | 24 | 48 | Factual
discharge | 48 | 48 | Factual