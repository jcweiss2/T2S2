numbness and weakness in lower extremities | -720
numbness and weakness progressed to hands and neck | -720
presumptive diagnosis of Guillain-Barré syndrome (GBS) | -720
admission to community hospital | 0
lumbar puncture | 0
albuminocytologic dissociation in cerebrospinal fluid | 0
brain magnetic resonance imaging (MRI) scan | 0
small vessel ischemic changes | 0
intravenous immunoglobulin (IVIG) treatment | 0
worsening pancytopenia | 120
encephalopathy | 120
transfer to specialist center | 120
hypotensive | 120
unresponsive to verbal stimuli | 120
minimally responsive to painful stimuli | 120
Glasgow Coma Scale (GCS) score of 6 | 120
anasarcic | 120
flaccid paralysis of all four extremities | 120
malnourished and septic state | 120
calcium of 6.7 mg/dL | 120
hemoglobin of 9.4 g/dL | 120
white cell count of 2.1×10^9/L | 120
phosphorus of 1.1 mg/dL | 120
creatinine <0.2 mg/dL | 120
albumin <1.5 gm/dL | 120
lactate of 4 mmol/L | 120
nutritional risk screening (NRS-2002) score of 5 | 120
malnutrition universal screening (MUST) score of 5 | 120
intubated | 120
resuscitated with intravenous fluids | 120
intravenous infusion of norepinephrine | 120
meropenem treatment | 120
vancomycin treatment | 120
anidulafungin treatment | 120
empirical treatment with high-dose intravenous thiamine | 120
electroencephalogram (EEG) | 168
diffuse slow waves | 168
severe metabolic encephalopathy | 168
brain magnetic resonance imaging (MRI) scan | 216
hyperintensity of bilateral medial thalamus | 216
Wernicke’s encephalopathy | 216
serum thiamine level of 104 nmol/L | 216
improved mental status | 288
able to understand simple commands | 288
discontinuation of norepinephrine | 288
discontinuation of antimicrobial treatment | 288
extubated | 360
electromyography (EMG) | 504
severe sensorimotor polyneuropathy | 504
transferred out of intensive care unit (ICU) | 1008
discharge | 1008 
thiamine supplementation | 0