39 years old | 0
businessman | 0
male | 0
admitted to ICU | 0
history of acute onset severe abdominal pain | 0
vomiting | 0
binge drinking | -24
chronic alcoholic | -8760
history of irregularly treated hypertension | -8760
normal baseline creatinine values | -8760
no history of chest pain | 0
conscious | 0
restless | 0
distended and tender abdomen | 0
in shock | 0
high total leukocyte count | 0
serum creatinine 4 mg/dl | 0
lipase 1500 IU/L | 0
normal ECG | 0
normal TTE | 0
SAP | 0
septic shock | 0
acute kidney injury | 0
raised intra-abdominal pressure | 0
treated with broad-spectrum antibiotics | 0
treated with anti-fungals | 0
treated with vasopressor | 0
treated with inotropes | 0
mechanical ventilation | 0
tracheostomy | 0
enteral nutrition | 0
renal replacement therapy | 0
multiple percutaneous drainages | 0
necrosectomy | 0
calcification of mitral leaflet | 1008
calcification of myocardium | 1008
grade I diastolic dysfunction of left ventricle | 1008
ring calcification around left ventricle | 1008
non-specific ST-T changes | 1008
normal cardiac enzyme markers | 1008
normal serum calcium | 0
normal phosphorus levels | 0
initiation of left ventricular wall calcification | 504
multi-drug-resistant complicated intra-abdominal infection | 1200
septic shock | 1200
death | 1200