55 years old | 0
male | 0
farmer | 0
admitted to the hospital | 0
repeated fever | -168
tick bite | -240
chills | -168
fatigue | -168
fever without an obvious cause | -168
body temperature normalized | -120
fever recurred | -120
no history of smoking | 0
no history of allergy | 0
no abnormalities in personal history | 0
no abnormalities in marital history | 0
no abnormalities in familial history | 0
temperature 40°C | 0
respiratory rate 20 breaths/minute | 0
blood pressure 116/65 mmHg | 0
no ecchymosis | 0
no bleeding points | 0
slightly coarse sounds in both lungs | 0
no obvious dry and wet rales | 0
heart rhythm regular | 0
pain in the liver on percussion | 0
palpable lymph node enlargement | 0
total white blood cell count 3.1 × 10^9/L | 0
neutrophil count 2.48 × 10^9/L | 0
hemoglobin 138 g/L | 0
platelet count 112 × 10^9/L | 0
C-reactive protein 66.7 mg/L | 0
negative for hepatitis B surface antigen | 0
urinalysis normal | 0
chest computed tomography revealed mild inflammation in both lungs | 0
chest computed tomography revealed emphysema | 0
diagnosed with sepsis | -48
diagnosed with pneumonia | -48
piperacillin 4.5 g every 8 hours for 2 days | -48
no significant improvement | -24
treatment changed to Tienam injection 1.0 every 8 hours for 2 days | -24
no observable improvement | 0
admitted to Lishui People’s Hospital | 0
delirious | 0
responded suspiciously to bending of his neck | 0
white blood cell count 3.5 × 10^9/L | 0
red blood cell count 4.38 × 10^12/L | 0
hemoglobin 132 g/L | 0
platelet count 61 × 10^9/L | 0
erythrocyte sedimentation rate 17 mm/hour | 0
prothrombin time 13.1 s | 0
d-dimer 4546 µg/L | 0
total protein 53.4 g/L | 0
alanine aminotransferase 285 U/L | 0
aspartate aminotransferase 235 U/L | 0
total bile acids 30.9 µmol/L | 0
C-reactive protein 130.8 mg/L | 0
no blood plasmodia detected | 0
serologically negative for human immunodeficiency virus | 0
serologically negative for hepatitis C | 0
serologically negative for anti-Epstein–Barr virus IgG | 0
serologically negative for syphilis | 0
serologically negative for pneumonia antibody | 0
Widal test negative | 0
Weil–Felix test negative | 0
urinalysis revealed weakly positive signal for urinary microalbumin | 0
cerebrospinal fluid transparency clear | 0
Pandy’s test revealed weak positivity for chloride | 0
Pandy’s test revealed weak positivity for total protein | 0
Pandy’s test revealed weak positivity for IgG | 0
cerebrospinal fluid and blood culture sterile | 0
mild mitral valve and tricuspid valve reflux | 0
cardiac arrhythmia | 0
calcification in the left renal cortex and prostate | 0
hepatomegaly with echogenicity | 0
gallbladder wall thickening | 0
abdominal cavity effusion | 0
inflammation in both lungs | 0
multiple small nodules in the right and left lower lobes | 0
patchy fibrosis in the right middle lung lobe and upper lobes of both lungs | 0
emphysema | 0
hepatomegaly | 0
dilatation of intrahepatic lymphatic vessels | 0
gallbladder wall edema | 0
ascites | 0
enlarged lymph nodes in the abdominal cavity and retroperitoneum | 0
multiple low-density lesions in the spleen | 0
possible splenic infarction | 0
small cysts in caudate hepatic lobes | 0
small cyst in the left kidney | 0
calcification foci in the prostate | 0
bilateral pleural effusion | 0
NGS identified Q fever associated with Coxiella infection | 120
doxycycline hydrochloride enteric-coated capsules administered | 120
compound glycyrrhizin and reduced glutathione injection administered | 120
fever relieved | 144
chills relieved | 144
discharged from the hospital | 144
doxycycline anti-infection sustained | 144
compound glycyrrhizin/doxycycline treatment sustained | 144
no side effects of therapy reported | 144