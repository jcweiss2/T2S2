75 years old | 0
male | 0
admitted to the hospital | 0
acute ischemic stroke | 0
thrombotic occlusion of the M1 segment of the left A. cerebri media | 0
coronary angiography | -16
intervention for non-ST-elevation myocardial infarction | -16
right-sided hemiplegia | 0
mechanical thrombectomy | 0
aspiration pneumonia | 0
piperacillin/tazobactam | -7
recurrent sinus bradycardia | 0
intermittent ventricular escape rhythm | 0
third-degree sinoatrial block | 0
2-chamber pacemaker implantation | 0
povidone-iodine solution | 0
discharged to a neurological rehabilitation facility | 4
readmitted | 11
fever | 11
hyperthermic, reddened pacemaker incision site | 11
leucocytosis | 11
elevated C-reactive protein | 11
blood cultures | 11
ampicillin/sulbactam | 11
system extraction | 12
intraprocedural inspection of the pacemaker pocket | 12
old hematoma | 12
swab samples of pacemaker and pocket | 12
explanted leads | 12
transferred to intensive care unit | 12
persisting sinoatrial block | 12
transesophageal echocardiography (TEE) | 12
mobile vegetation from the right atrium to the superior vena cava | 12
ghosts | 12
device-associated endocarditis | 12
blood cultures positive for C. difficile | 14
pacemaker samples positive for C. difficile | 14
pocket swab cultures positive for C. difficile | 14
stool sample | 14
toxigenic C. difficile strains | 14
nontoxigenic isolate | 14
antimicrobial testing | 14
ribotyping | 14
minimum inhibitory concentration | 14
vancomycin | 14
metronidazole | 14
genotyping | 14
whole-genome sequencing | 14
clonality of the RT014 isolates | 14
mixed strain colonization | 14
detailed medical history | 14
no signs of previous C. difficile infection | 14
no contact with infectious diarrhea | 14
abdominal ultrasound | 14
no pathologies | 14
antibiotic treatment switched to intravenous vancomycin and oral metronidazole | 17
laboratory tests revealed normalization of leukocytes and C-reactive protein | 20
oral antibiotic therapy switched from metronidazole to vancomycin | 20
repeated blood cultures and stool samples during therapy remained negative | 23
transferred back to the rehabilitation facility | 23
intravenous vancomycin continued for a total of 30 days | 23
oral vancomycin administered for a total of 42 days | 23
tapering regime | 23
readmitted for pacemaker reimplantation | 50
TEE revealed complete elimination of vegetations | 50
repeated blood cultures and skin swabs of the groin, axilla, rump, and pacemaker pocket were negative for C. difficile | 50
colonoscopy showed no signs of intestinal inflammation | 50
noninflamed sigmoid diverticula | 50
toxigenic C. difficile was again isolated from follow-up stool samples | 50
genotyping revealed a different toxigenic RT005 | 50
reinfection | 50
reimplantation of the pacemaker was performed on the contralateral side | 53
released to a rehabilitation facility | 53
oral vancomycin tapering regime for another 50 days | 53
follow-up visit 2 months after reimplantation | 105
normal pacemaker function with no sign of infection | 105