28 years old | 0
    male | 0
    presented to the Emergency Department via Emergency Medical Services | 0
    found unresponsive | -24
    hypothermic | 0
    hypoxic | 0
    core body temperature of 32.7°C | 0
    required 3 L of supplemental oxygen per nasal cannula | 0
    blood pressure 116/42 mmHg | 0
    heart rate 90 beats per minute | 0
    pupils equal and reactive to light | 0
    non-icteric sclera | 0
    dry oral mucous membranes | 0
    regular heart rate and rhythm | 0
    no murmurs | 0
    no jugular venous distension | 0
    no edema of the lower extremities | 0
    intact radial and dorsal pedal pulses | 0
    Kussmaul breathing | 0
    clear to auscultation bilaterally | 0
    soft and nontender abdomen | 0
    multiple tattoos | 0
    no rashes | 0
    no lesions | 0
    obtunded | 0
    arousable | 0
    able to follow commands | 0
    arterial blood gas pH 6.85 | 0
    carbon dioxide 14.0 kPa | 0
    oxygen 164.0 kPa | 0
    bicarbonate 2.3 mmol/L | 0
    base excess −29.6 mmol/L | 0
    potassium 9.0 mmol/L | 0
    ECG suspicious for STEMI | 0
    consulted Cardiology | 0
    initial ECG irregular rhythm without consistent p-wave to QRS complexes | 0
    rSR’ with down-sloping S-wave | 0
    inverted T-waves | 0
    hyperkalemia | 0
    treated with calcium carbonate | 0
    treated with insulin therapy | 0
    diabetic ketoacidosis | 0
    repeat ECG showed improvement | 24
    sodium 115 mmol/L | 0
    potassium 9.0 mmol/L | 0
    chloride 76 mmol/L | 0
    blood urea nitrogen 88 mmol/L | 0
    creatinine 4.8 mmol/dL | 0
    glucose 1375 mmol/L | 0
    calcium 7.9 mmol/L | 0
    alkaline phosphatase 112 μkat/L | 0
    bicarbonate <5.0 mmol/L | 0
    alanine aminotransferase 40 μkat/L | 0
    aspartate aminotransferase 26 μkat/L | 0
    albumin 3.5 g/L | 0
    total bilirubin 0.5 μmol/L | 0
    osmolality 330 mmol/kg | 0
    creatinine phosphokinase 176 units/L | 0
    troponin-I 0.596 μg/L | 0
    c-reactive protein 0.1 mg/L | 0
    glomerular filtration rate 15 mL/s | 0
    creatinine kinase-MB 5.3 μg/L | 0
    myoglobin 551 nmol/L | 0
    white blood cell count 29.4×109/L | 0
    hemoglobin 8.1 g/L | 0
    hematocrit 25% | 0
    mean corpuscular volume 86.8 fL | 0
    platelet count 301×109/L | 0
    intubated | 0
    central venous access placed | 0
    dialysis catheter placed | 0
    covered with Bair Hugger | 0
    covered with heated blankets | 0
    intravenous access started | 0
    aggressive volume resuscitation with 4 L normal saline | 0
    admitted to Intensive Care Unit | 0
    hyperosmolar coma | 0
    type I diabetes mellitus | 0
    insulin therapy non-compliance | -672
    alcohol use | -672
    diabetic ketoacidosis addressed with fluid resuscitation | 24
    initiated insulin infusion | 24
    consulted Nephrology | 24
    life-threatening electrolyte abnormalities | 24
    systemic inflammatory response syndrome | 24
    suspected sepsis | 24
    elevated prolactin level | 24
    placed on empiric antibiotic therapy with vancomycin | 24
    placed on empiric antibiotic therapy with meropenem | 24
    chest radiography confirmed left lower-lobe aspiration pneumonia | 72
    lactic acidosis | 72
    initial cardiac troponin-I 0.596 μg/L | 0
    subsequent cardiac troponin-I 19.1 μg/L | 72
    peak cardiac troponin-I 20.452 μg/L | 96
    on weight-based heparin infusion | 72
    on antiplatelet therapy | 72
    no significant cardiac history | 0
    presentation of DKA | 0
    profound hypovolemia | 0
    WHO fourth universal definition type-II myocardial infarction | 72
    preserved ejection fraction | 72
    absence of significant cardiac wall motion abnormalities | 72
    biochemically improved | 144
    clinically improved | 144
    eager for discharge | 144
    no documented seizures | 144
    no agonal nocturnal respirations after extubation | 144
    medical therapies optimized | 144
    discharged home | 144
    atorvastatin 80 mg P.O. QHS | 144
    aspirin 81 mg p.o. daily | 144
    metoprolol tartrate 12.5 mg p.o. BID | 144
    amlodipine 5 mg p.o. daily | 144
    Levemir 25 units subcutaneous qam | 144
    Levemir 10 units subcutaneous qpm | 144
    nov-Log subcutaneous carb count | 144
    subsequent Cardiology follow-up | 168
    history of syncope | -672
    continued isolated dizzy spells | -672
    prior Brugada-like ECG findings | -672
    high-risk diabetes | -672
    left heart catheterization | 168
    selective coronary angiogram | 168
    left ventriculo-gram | 168
    normal epicardial coronary arteries | 168
    ejection fraction of 65% | 168
    referred for electrophysiology consultation | 168
    no family history of sudden cardiac death | 0
    no proband-positive Brugada syndrome family history | 0
    Brugada pattern secondary to Brugada phenocopy | 0
    severe dehydration | -672
    severe electrolyte derangements | -672
    severe metabolic derangements | -672
    acute renal failure | 0
    sepsis | 0
    type-II myocardial infarction | 72
    EMS ECG interpreted as acute anterior myocardial infarction | -24
    ED ECG findings secondary to hyperkalemia | 0
    treated with calcium carbonate | 0
    treated with bicarbonate | 0
    treated with insulin infusion therapy | 0
    no cardiac resuscitation | 0
    no ventricular arrhythmias | 0
    subsequent ECGs demonstrated normalization of Brugada pattern | 72
    resolution of electrolyte derangements | 72
    resolution of metabolic derangements | 72
    no chest pain | 0
    no sudden cardiac death presentation | 0
    hyperacute T wave | 0
    right axis deviation | 0
    widened QRS duration | 0
    absence of P waves | 0
    consumption of ethyl alcohol | -672
    hyperglycemia | -672
    diabetic ketoacidosis | 0
    acidosis | 0
    no ventricular fibrillation | 0
    referred to Electrophysiology | 168
    no ICD implantation | 168
    no ventricular tachycardia identification | 168
    no experimental EP ablation of RVOT | 168
    no quinidine consideration | 168
    STEMI mimics | 0
    Brugada syndrome | 0
    Brugada phenocopy | 0
    hyperkalemia- and acidemia-induced Brugada pattern | 0
    no genetic testing | 168
    no provocative testing confirmation | 168
    