55 years old | 0
male | 0
non-smoker | 0
admitted to the hospital | 0
fever | 0
joint pain | 0
cold, painful extremities | 0
non-erosive RA | -2190
rheumatoid factor positive | -2190
anti-cyclic citrullinated peptide negative | -2190
methotrexate | -730
lcSSc overlap syndrome | -730
RP | -730
sclerodactyly | -730
telangiectasia | -730
sicca symptoms | -730
anti-nuclear antibodies positive | -730
anti-RNP (U1RNP) specificity | -730
cold digits | 0
small joint synovitis of the hands and feet | 0
raised white cell count | 0
neutrophil count | 0
C-reactive protein (CRP) 301 mg/L | 0
empirical intravenous antibiotics | 0
oral corticosteroids (prednisolone 20 mg od) | 0
continuous prostaglandin analog (iloprost) infusion | 0
body temperature spiked | 24
inflammatory markers rose | 24
antibiotic therapy broadened | 24
transesophageal echocardiogram | 24
no vegetations | 24
multiple sets of blood cultures returned negative | 24
computed tomography of the chest, abdomen, and pelvis | 24
no occult source of sepsis | 24
necrosis of the hands and feet | 168
therapeutic dose of low-molecular weight heparin | 168
clopidogrel | 168
iloprost infusion uptitrated | 168
magnetic resonance angiography | 168
no macrovascular occlusions | 168
intravenous methylprednisolone (500 mg) | 240
CRP fell to 153 mg/L | 240
wet gangrene of the lower limbs | 240
bilateral below-knee amputations | 240
postoperatively | 240
prednisolone 60 mg daily | 240
infusions of intravenous immunoglobulin (IVIG) | 240
demarcation of tissue gangrene | 288
no further progression of necrosis | 288
ulnar and radial pulses strong | 288
CRP fell rapidly | 288
antibiotics stopped | 288
mycophenolate mofetil (MMF) initiated | 288
negative tests for anti-centromere/anti-Scl70 antibodies | 288
negative tests for anti-neutrophil cytoplasmic antibody (ANCA) | 288
negative tests for antiphospholipid antibodies | 288
negative tests for cryoglobulins | 288
negative serology for viruses hepatitis B, C, and HIV | 288
lipid profile within normal limits | 288
plastic surgeon advised amputation at both elbows | 288
conservative management | 288
dry gangrene | 288
monthly IVIG | 4320
weaning dose of prednisolone | 4320
vasodilator therapy including sildenafil | 4320
MMF uptitrated to 1g BD | 4320
rivaroxaban added | 4320
discharged to rehabilitation | 4032
learned to use prostheses independently | 4032
auto-amputation of fifth digits | 8760
limited surgical resection of remaining necrotic digits | 10920
remains in remission on medical therapy | 10920
significant functional impairment | 10920
manages well | 10920