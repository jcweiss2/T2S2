47 years old | 0
male | 0
Japanese | 0
admitted to the hospital | 0
septic shock | 0
necrotising fasciitis of the axilla | 0
Group A streptococci detected in blood | 0
Group A streptococci detected in soft tissue | 0
hypertension | -672
amlodipine administered | -672
invasive positive-pressure ventilation performed | 0
penicillin G administered | 0
norepinephrine administered | 0
serial debridement performed | 1
serial debridement performed | 2
serial debridement performed | 3
intravenous norepinephrine tapered | 3
normal ECG findings | 24
complete atrioventricular block developed | 96
cardiac arrest | 96
cardiopulmonary resuscitation performed | 96
return of spontaneous circulation achieved | 96
epinephrine administered | 96
inverted T waves on leads I, aVL and precordial leads V5 and V6 | 96
ST depression on leads I, aVL and precordial leads V1–V6 | 96
first-degree atrioventricular block | 96
hypokinesia of the inferior wall | 96
temporary pacemaker insertion | 96
coronary angiography performed | 96
no significant stenosis in coronary arteries | 96
coronary spastic angina suspected | 96
provocative testing with ergonovine performed | 96
coronary spasm with ST segment elevation confirmed | 96
intracoronary administration of isosorbide nitrate | 96
coronary spasm relieved | 96
nifedipine administered | 96
no recurrence of coronary spasm or atrioventricular block | 120
temporary pacing discontinued | 144
negative blood culture confirmed | 216
extubation | 216
transferred from intensive care unit to general ward | 240
discharged | 1176
no further complaints of chest pain | 1176
no changes on cardiac monitoring | 1176
no recurrence of symptoms at 3 months | 3264