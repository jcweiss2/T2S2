63 years old | 0
male | 0
admitted to hospital | 0
fever | -72
mental obtundation | -72
right-sided otitis media | 0
purulent discharge | 0
Glasgow Coma Scale score 4 | 0
temperature 36.8° C | 0
pulse 124 | 0
respiration 20 | 0
blood pressure 137/79 mmHg | 0
mild divergent strabismus | 0
eye deviation to the left | 0
deep tendon reflexes symmetric and enhanced | 0
Babinski's sign negative | 0
leukocyte count 18.5 × 10^9/L | 0
neutrophils 91% | 0
monocytes 7% | 0
lymphocytes 3% | 0
red blood cell count 4.7 × 10^12/L | 0
hemoglobin 143 g/L | 0
platelets 172 × 10^9/L | 0
erythrocyte sedimentation rate 80 per h | 0
C-reactive protein 75.5 mg/L | 0
fibrinogen 4.13 g/L | 0
prothrombin and partial-thromboplastin times normal | 0
serum concentration of lactate 6.0 mmol/L | 0
magnesium 0.5 mmol/L | 0
phosphorus 0.43 mmol/L | 0
total bilirubin normal | 0
aminotransferases normal | 0
lactate dehydrogenase normal | 0
glucose normal | 0
alkaline phosphatase normal | 0
serum protein electrophoresis normal | 0
sodium 134 mmol/L | 0
potassium 3.0 mmol/L | 0
chloride 97 mmol/L | 0
urea nitrogen 5.0 mmol/L | 0
creatinine 88 μmol/L | 0
cerebrospinal fluid examination | 0
white cells 200,000 per cubic millimeter | 0
polymorphonuclear cells 95% | 0
CSF glucose 0.0 mmol/L | 0
total protein concentration 12.1 g/L | 0
lactate 15.9 mmol/L | 0
intravenous ceftriaxone 4 g per day | 0
dexamethasone 48 mg/day | 0
native and contrast-enhanced brain CT scans normal | 0
transcranial Doppler ultrasonography | 0
absent diastolic blood flow velocities | 0
mean arterial pressure 72 mmHg | 0
carbon-dioxide reactivity impaired | 0
breath holding index 0.80 | 0
bilateral increase in optic nerve sheath diameter | 0
mild therapeutic hypothermia | 0
norepinephrine support | 0
hypothermia induced | 0
continuous veno-venous hemofiltration | 0
marked reduction in optic nerve sheath diameter | 24
improvement of mean blood flow velocities | 24
patient became alert | 120
followed simple commands | 120
mild diffuse brain edema | 120
flaccid paraplegia | 120
areflexia | 120
sensory level at T8 | 120
loss of bladder control | 120
repeated lumbar puncture | 120
bloody-brown fluid | 120
magnetic resonance imaging of the spine | 120
scattered multiple hyperintensive lesions | 120
myelitis | 120
high-dose methylprednisolone | 120
total plasma exchange | 120
neurological deficit unchanged | 168
transferred to rehabilitation center | 1440
Glasgow Coma Scale score 15 | 1440
Glasgow Outcome Scale score 3 | 1440
Karnofsky performance score 60% | 1440
rehabilitation treatment unsuccessful | 2880
patient remained paraplegic | 2880
urinary incontinence | 2880