12 years old | 0
    male | 0
    Maori | 0
    presented to hospital | 0
    acute otitis media | -24
    perforation | -24
    neck swelling | -24
    neck pain | -24
    features of septic shock | 0
    urgent ICU admission | 0
    endotracheal intubation | 0
    computed tomography scan | 0
    retropharyngeal phlegmon | 0
    obstructive thrombi in left internal jugular vein | 0
    obstructive thrombi in parts of right internal jugular vein | 0
    pulmonary septic emboli | 0
    multiple pulmonary lesions | 0
    differential diagnosis of Lemierre’s syndrome | 0
    antibiotics started | 0
    cefotaxime | 0
    metronidazole | 0
    flucloxacillin | 0
    lincomycin | 0
    cultures from external ear canal | 0
    blood cultures | 0
    growth of MSSA | 0
    initial echocardiogram normal | 0
    infective endocarditis excluded | 0
    blood cultures positive for first 3 days | 0
    blood cultures clear of MSSA after 3 days | 72
    high-frequency ventilation | 24
    hypoxia | 24
    increase in mean airway pressure to 28 cm H2O | 24
    inspired oxygen fraction of 0.5 | 24
    worst oxygenation index 40 | 24
    repeat CT scan on day three | 72
    progression of jugular clots | 72
    progression of pulmonary emboli | 72
    progression of pulmonary cavitating lesions | 72
    increasing cardiovascular support | 72
    noradrenaline 0.3 µg/kg/min | 72
    adrenaline 0.05 µg/kg/min | 72
    vasopressin 1 U/h | 72
    adequate blood pressure | 72
    deterioration requiring escalation of cardiorespiratory support | 72
    attempt to minimize ventilation pressures | 72
    prevent further lung injury | 72
    prevent pulmonary air leaks | 72
    commenced on ECLS via femoral veno-arterial cannulation | 72
    ECLS cannulation | 72
    rest ventilation instituted | 72
    pressure control ventilation | 72
    peak inspiratory pressures of 15 cm H2O | 72
    positive end-expiratory pressure of 5 cm H2O | 72
    right-sided pneumothorax | 72
    drained pneumothorax | 72
    left-sided pneumothorax | 144
    hemoserous drain losses | 72
    total hemoserous drain losses 400 mL | 72
    no evidence for frank haemorrhage | 72
    inflammatory markers remained high | 72
    intermittently required inotropic support | 72
    ongoing systemic inflammation | 72
    CT imaging on day eight | 192
    abscess formation posterior to cervical vertebra one | 192
    osteomyelitis involving body of C1 | 192
    osteomyelitis involving dens of C2 | 192
    opacified left mastoid | 192
    decision to drain abscess posterior to C1 | 192
    cortical mastoidectomy | 192
    procedure performed in PICU in prone position | 192
    mastoid drilled out | 192
    retropharyngeal space not opened | 192
    heparin stopped | 192
    tranexamic acid given | 192
    bleeding around abscess well controlled | 192
    periosteal bleeding challenging to control | 192
    estimated blood loss 600–700 mL | 192
    peri-procedure red blood cells 1500 mL | 192
    peri-procedure pooled platelet 1100 mL | 192
    fibrinogen remained high | 192
    no cryoprecipitate required | 192
    no concentrated fibrinogen required | 192
    tranexamic acid 1800 mg | 192
    thrombelastogram showing hyperfibrinolysis | 192
    total blood during ECMO run 5700 mL | 192
    total platelets during ECMO run 3200 mL | 192
    total tranexamic acid during ECMO run 4600 mg | 192
    cultures from drained paravertebral abscess | 192
    growth of MSSA | 192
    cortical mastoidectomy destruction of malleus and incus | 192
    granulation tissue in attic | 192
    subtotal perforation | 192
    chronic middle ear process | 192
    posterior cervical muscle wound not primarily closed | 192
    negative pressure vacuum dressing | 192
    delayed primary closure | 192
    no requirement for repeat surgical drainage | 192
    CT imaging on day 13 | 312
    progression of lung abscesses | 312
    big abscess in right middle lobe | 312
    high risk of bronchopleural fistula | 312
    deferred drainage of abscess | 312
    improving pulmonary gas exchange | 312
    weaning from ECLS | 312
    successful decannulation | 384
    magnetic resonance imaging post decannulation | 384
    no further abscesses | 384
    invasive mechanical ventilation | 0
    mechanical ventilation until day 23 | 552
    post extubation respiratory support | 552
    non-invasive ventilation | 552
    high-flow nasal cannula oxygen | 552
    secondary pseudomonal sepsis | 552
    profound critical illness myopathy | 552
    CT imaging after extubation | 552
    pathological fractures of lateral masses of C1 | 552
    discharged from ICU | 1032
    follow-up imaging after ICU discharge | 1032
    improved lung fields | 1032
    improvement of cavitations | 1032
    resolution of fluid collections around C1 and C2 | 1032
    persistence of thrombi in jugular veins | 1032
    persistence of thrombi in venous sinuses | 1032
    intravenous flucloxacillin | 1032
    intravenous Bactrim | 1032
    oral Bactrim | 1032
    oral flucloxacillin | 1032
    continued for eight weeks | 1032
    planned for further four months | 1032
    CNS imaging done repeatedly | 0
    delineation of mastoid and C1 collections | 0
    screening for intracranial abscesses | 0
    small intracranial extradural collections | 0
    small scattered foci of haemorrhage in cerebellar hemispheres | 0
    MRI six months after discharge | 4032
    resolution of all abnormal findings | 4032
    small degree of gliosis in cerebellum | 4032
    osteomyelitis of C1 and C2 | 0
    fractures of lateral masses of C1 | 552
    halo-thoracic jacket applied | 552
    neurocognitive assessment | 4032
    normal motor outcome | 4032
    normal cognitive outcome | 4032
    normal behavioural outcome | 4032
    Pediatric Overall Performance Category Assessment PCPC=1 | 4032
    audiological assessment | 4032
    mild conductive loss on left | 4032
    bilateral sensorineural mid to high frequency loss | 4032
    discharged from hospital | 2880
    halo-thoracic jacket removal deferred | 2880
    consent obtained from parents | 0
    patient assented | 0
    