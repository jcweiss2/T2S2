35 years old | 0\
female | 0\
pregnant | 0\
admitted to the hospital | 0\
fever | -240\
cough | -240\
dyspnoea | -120\
aggravated dyspnoea | -120\
conscious of foetal movement | -560\
foetus had been active | -560\
recurrent fever | -240\
highest body temperature being 39.2 ℃ | -240\
decreased to normal after oral acetaminophen | -240\
accompanied by cough | -240\
yellow viscous sputum | -240\
chest distress | -240\
shortness of breath | -240\
without chills | -240\
cyanosis of the lip | 0\
thick breathing sounds in both lungs | 0\
dry and wet rales in the right lower lung | 0\
heart rate was regular | 0\
no noises were heard in the auscultation area of each valve | 0\
gestational and symmetric abdominal type | 0\
height of 166 cm | 0\
pre-pregnancy weight of 46.5 kg | 0\
body mass index of 16.87 | 0\
weight gain of 8.8 kg during pregnancy | 0\
uterine height was 34 cm | 0\
abdominal circumference was 89 cm | 0\
contractions were sporadic and weak | 0\
head presentation | 0\
foetal heart sounds were 142 beats/min | 0\
intrapelvic and extrapelvic measurements were normal | 0\
pH 7.472 | 0\
partial pressure of carbon dioxide 34.0 mmHg | 0\
partial pressure of oxygen 56 mmHg | 0\
sulfur dioxide 88.6% | 0\
C-reactive protein (CRP): 186.33 mg/L | 0\
erythrocyte sedimentation rate: 69.00 mm/h | 0\
procalcitonin (PCT): 2.24 ng/mL | 0\
White blood cell (WBC) 18.29 × 109/L | 0\
neutrophil % 90.10% | 0\
lymphocyte 0.97 × 109/L | 0\
Alkaline phosphatase 232 U/L | 0\
total bilirubin 23.1 μmol/L | 0\
albumin (ALB) 33.9 g/L | 0\
K+ 2.93 mmol/L | 0\
sodium 129 mmol/L | 0\
chloride 89 mmol/L | 0\
cardiac markers were normal | 0\
multiple plaques, miliary foci, nodular foci with partial consolidation and cavities in the upper and lower lobes of both lungs | 0\
single viable foetus | 0\
head presentation | 0\
oligohydramnios | 0\
no significant abnormalities in cardiac ultrasound and lower extremity vascular ultrasound | 0\
first menarche at the age of 15 | -7305\
menstrual cycle was regular | -7305\
last menstruation occurred on May 2, 2022 | -6720\
moderate menstrual volume and a normal colour | -6720\
no blood clots or painful menstruation | -6720\
married at an appropriate age | -7305\
spouse was healthy | -7305\
one pregnancy history | -7305\
full-term normal delivery of a female infant in 2006 | -7305\
weighing 3500 g and in good health | -7305\
Pregnancy combined with severe pneumonia novel coronavirus infection S. aureus infection type respiratory failure | 0\
late pregnancy with 34 + 4 wk G2P1 left occiput anterior | 0\
elderly second parturient women | 0\
maternal lower weight | 0\
oligohydramnion | 0\
premature live baby | 0\
electrolyte disturbance | 0\
hypoproteinaemia | 0\
cefoperazone sodium and sulbactam sodium for anti-infective therapy | 0\
10 mg dexamethasone to promote foetal lung maturation | 0\
oxyhemoglobin saturation continued to progressively decline | 12\
foetal heart sounds were 146 beats/min | 12\
caesarean section of the lower uterus | 12\
high-flow nasal cannula oxygen therapy | 12\
oxyhemoglobin saturation increased to 95%-98% | 24\
assisted ventilation by endotracheal intubation with a ventilator | 24\
empirical antibiotic therapy to prevent infection by intravenous drip of meropenem and vancomycin | 24\
symptomatic treatment of fluid and ALB infusion | 24\
irrigation solution was collected and tested for metagenomic next-generation sequencing (mNGS) by bedside tracheoscopy | 24\
S. aureus combined with novel coronavirus infection | 24\
no acid-fast bacilli in the sputum tuberculosis smear | 24\
tubercle bacillus-polymerase chain reaction (TB-PCR) and nontuberculosis mycobacterium-PCR were negative | 24\
galactomannan experiments were normal | 24\
intravenous drip of 1 g every 12 h (q12h) vancomycin and 1 g q8h meropenem | 24\
anticoagulant therapy | 24\
treatments to relieve the cough and reduce the amount of sputum | 24\
other symptomatic treatment | 24\
transitioned from assisted ventilation by the invasive ventilator to nasal tube oxygen with a flow rate of 3-4 L/min | 48\
multiple areas of inflammation in both lungs | 96\
mildly enlarged mediastinal lymph nodes | 96\
a small amount of bilateral pleural effusion | 96\
CRP was 38.54 mg/L | 96\
WBC count was 8.25 × 109/L | 96\
PCT was 0.129 ng/mL | 96\
potassium was 4.04 mmol/L | 96\
D-dimer was 2.44 mg/L | 96\
TB-PCR was negative | 96\
inflammatory lesions | 216\
pleural effusion had been absorbed | 216\
antibiotics were adjusted to sitafloxacin 50 mg twice daily | 216\
condition was stable | 264\
discharged from the hospital | 264\
multiple lung inflammation was absorbed slightly | 264\
multiple lung inflammation was apparently absorbed | 744