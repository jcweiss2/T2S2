24 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
pregnancy | 0 | 0 | Factual
abdominal pain | -120 | 0 | Factual
abdominal distension | -120 | 0 | Factual
constipation | -120 | 0 | Factual
admitted to hospital | 0 | 0 | Factual
dehydrated | 0 | 0 | Factual
hypotension | 0 | 0 | Factual
tachycardia | 0 | 0 | Factual
tachypnea | 0 | 0 | Factual
asymmetrically distended abdomen | 0 | 0 | Factual
tenderness all over abdomen | 0 | 0 | Factual
empty rectum on digital examination | 0 | 0 | Factual
foetal viability assessed | 0 | 0 | Factual
vaginal examination not suggestive of threatened preterm labour | 0 | 0 | Factual
elevated white cell count | 0 | 0 | Factual
normal urine analysis | 0 | 0 | Factual
ultrasound scan of abdomen and pelvis | 0 | 0 | Factual
distended bowel loop | 0 | 0 | Factual
moderate amount of free fluid in peritoneal cavity | 0 | 0 | Factual
single viable foetus | 0 | 0 | Factual
abdominal X-ray | 0 | 0 | Factual
dilated large bowel | 0 | 0 | Factual
abnormal gas pattern | 0 | 0 | Factual
coffee bean appearance | 0 | 0 | Factual
sigmoidoscopy | 0 | 0 | Factual
twisted sigmoid colon | 0 | 0 | Factual
failure to negotiate obstruction | 0 | 0 | Factual
foetal distress | 0 | 0 | Factual
deceleration in heart rate | 0 | 0 | Factual
concomitant caesarean section | 0 | 0 | Factual
laparotomy | 0 | 0 | Factual
enormously distended sigmoid loop | 0 | 0 | Factual
ischemic and gangrenous changes | 0 | 0 | Factual
no signs of perforation | 0 | 0 | Factual
lower segment caesarean section | 0 | 0 | Factual
preterm infant | 0 | 0 | Factual
male infant | 0 | 0 | Factual
weight 750g | 0 | 0 | Factual
admitted to neonatal ICU | 0 | 24 | Factual
mechanical ventilation | 0 | 24 | Factual
gangrenous sigmoid colon resection | 0 | 0 | Factual
Hartmann’s procedure | 0 | 0 | Factual
end colostomy | 0 | 0 | Factual
closure of rectal stump | 0 | 0 | Factual
post-operative course uneventful | 0 | 216 | Factual
discharged home | 216 | 216 | Factual
reversal of Hartmann’s | 4320 | 4320 | Factual
bowel continuity restored | 4320 | 4320 | Factual
colo-rectal anastomosis | 4320 | 4320 | Factual
child discharged home | 720 | 720 | Factual