high-grade fever | -72
pleuritic right lower chest pain | -72
cough | -72
elevated temperature | 0
bibasilar crackles | 0
lower extremity edema | 0
grade 3 holosystolic apical murmur | 0
mitral valve regurgitation | 0
long-term venous access port | 0
anemia | 0
hemoglobin 12.1 g/dL | 0
white blood cell count 15.1×103/µL | 0
absolute neutrophil count 13.2×103/µL | 0
b-type natriuretic peptide 788 pg/mL | 0
congestive heart failure | 0
left bundle branch pattern | 0
Corynebacterium CDC group G bacteremia | 0
gram positive rods | 0
moderate mitral valve regurgitation | 0
thickened anterior mitral leaflet | 0
pulmonary artery systolic pressure 84 mmHg | 0
bacterial IE | 0
vancomycin therapy | 0
clindamycin therapy | 0
discharged to extended care facility | 120
readmitted to hospital | 192
hypoxia | 192
worsening vegetations on echocardiogram | 192
mitral valve replacement | 216
coronary artery bypass grafting | 216
post-op acute kidney injury | 240
acute respiratory failure | 240
mechanical ventilation | 240
vancomycin resistant enterococcus | 360
urinary tract infection | 360
daptomycin therapy | 360
worsening congestive heart failure | 432
fever spikes | 600
hypotension | 600
transesophageal echocardiography | 600
recurrent vegetations of the bioprosthetic mitral valve | 600
doxycycline therapy | 600
aztreonam therapy | 600
anidulafungin therapy | 600
bioprosthetic mitral valve replaced | 624
limb ischemia | 696
disseminated intravascular coagulation | 696
multi-organ failure | 696
patient expired | 696
diphtheroids in blood cultures | -720
pneumonia | -720
levofloxacin therapy | -720