64 years old|0
male|0
hepatitis C virus infection|0
alcohol-related cirrhosis|0
hepatocellular carcinoma|0
liver transplant|0
ABO-identical|0
cadaveric donor|0
cytomegalovirus-seronegative donor|0
toxoplasma-seropositive donor|0
cytomegalovirus-seropositive recipient|0
toxoplasma-seropositive recipient|0
body mass index 24.5 kg/m²|0
Child–Pugh score A6|0
MELD score 10|0
transfused 2 units concentrated red cells|0
transfused 4 units fresh frozen plasma|0
tacrolimus|0
corticosteroid|0
increase in aspartate aminotransferase|9
increase in alanine aminotransferase|9
acute cellular rejection|9
steroid pulse therapy|-16
regression of rejection|16
discharged|25
readmitted|31
skin rash|31
generalized maculopapular eruption|31
erythema|31
palm rash|31
fever|31
severe leukopenia (0.45 mil/mm³)|31
anemia|31
low hemoglobin|31
low blood pressure|31
watery diarrhea|31
skin biopsies consistent with GVHD|31
vacuolar degeneration of the basal layer|31
epidermal infiltration by lymphocytes|31
necrotic eosinophilic keratinocytes|31
spongiosis|31
basal cell hydropic changes|31
apoptotic keratinocytes|31
lymphocytic exocytosis|31
satellite-cell necrosis|31
subepidermal cleft formation (grade III)|31
hypoplastic bone marrow|31
aplasia|31
single-cell necrosis (apoptosis)|31
gastric mucosa gland abscesses|31
partial mucosal denudation|31
chimerism (day 32)|32
donor T-lymphocyte macrochimerism 3-4%|32
intravenous methylprednisolone|31
antithymocyte globulin|31
no improvement in skin rash|31
progressive worsening of clinical condition|36
pulmonary insufficiency|36
renal insufficiency|36
agranulocytosis|36
multi-organ failure|36
death|36
