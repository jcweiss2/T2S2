52 years old | 0 | 0 
male | 0 | 0 
admitted to the hospital | 0 | 0 
right upper quadrant pain | -168 | 0 
abdominal fullness and distention | -168 | 0 
abdominal pain worsened after meals | -168 | 0 
denies nausea | -168 | 0 
denies vomiting | -168 | 0 
denies stiffness | -168 | 0 
denies fever | -168 | 0 
no past medical history | 0 | 0 
no history of close contact with infected individuals | 0 | 0 
no recent travel | 0 | 0 
no abdominal trauma | 0 | 0 
hepatic abscess | -24 | 0 
treated with hepatic puncture and drainage | -24 | 0 
afebrile | 0 | 0 
pulse rate of 80 beats/minute | 0 | 0 
blood pressure of 118/73 mmHg | 0 | 0 
respiratory rate of 26 breaths/minute | 0 | 0 
leukocyte count of 16.4×10^9/L | 0 | 0 
neutrophil 94.5% | 0 | 0 
haemoglobin level of 85 g/L | 0 | 0 
platelet count of 240×10^9/L | 0 | 0 
procalcitonin level of 2.3 ng/mL | 0 | 0 
plasma fibrinogen level of 7.48 g/L | 0 | 0 
liver function tests slightly abnormal | 0 | 0 
serum glutamic oxalacetic transaminase level of 67 U/L | 0 | 0 
glutamic-pyruvic transaminase level of 83 U/L | 0 | 0 
cholinesterase level of 1360 U/L | 0 | 0 
total protein level of 50.8 g/L | 0 | 0 
albumin level of 21.5 g/L | 0 | 0 
blood urea nitrogen level of 10.8 mmol/L | 0 | 0 
creatinine level of 51.3 umol/L | 0 | 0 
negative for HIV | 0 | 0 
negative for syphilis | 0 | 0 
abdominal distension | 48 | 48 
mild bellyache | 48 | 48 
extreme thirst | 48 | 48 
right abdominal tenderness | 48 | 48 
no rebound or guarding | 48 | 48 
temperature of 36.8 °C | 48 | 48 
drainage catheter yield of 150 mL of fulvous fluid | 48 | 48 
abdominal and pelvic computed tomography scan | 48 | 48 
irregular, slightly low-density lesion in the right posterior hepatic lobe | 48 | 48 
gas density shadow inside the lesion | 48 | 48 
liquid density shadow and high-density drainage tube shadow around the lower margin of liver | 48 | 48 
round-like low-density lesion in the right lobe of the liver | 48 | 48 
appendix thickened to about 20 mm in diameter | 48 | 48 
structure of the ascending colon near the ileocecal region became disorganised | 48 | 48 
multiple gas accumulation and dilation in the bowel | 48 | 48 
air-fluid levels inside the abdomen | 48 | 48 
hepatic abscesses | 48 | 48 
ileus | 48 | 48 
mild ascites | 48 | 48 
appendicitis | 48 | 48 
liver cyst | 48 | 48 
abdominal infection | 48 | 48 
peritonitis | 48 | 48 
pre-shock | 72 | 72 
insufficient blood pressure of 93/59 mmHg | 72 | 72 
exploratory laparotomy | 72 | 72 
fulvous purulent exudate and necrotic tissue in the extraperitoneal space and abdominal cavity | 72 | 72 
partial postnecrotic defect in the peritoneum | 72 | 72 
massive epiploon adhesion in the right upper abdomen | 72 | 72 
two perforations | 72 | 72 
one perforation under the right side of the liver | 72 | 72 
one perforation in the right ascending colon | 72 | 72 
ileocecal resection | 72 | 72 
partial resection of the ascending colon | 72 | 72 
ileostomy | 72 | 72 
drainage of hepatic, abdominal and extraperitoneal abscesses | 72 | 72 
orotracheal intubation | 72 | 96 
hypotension | 72 | 96 
anemia | 72 | 96 
fever | 72 | 96 
transferred to the intensive care unit | 96 | 96 
noradrenaline to maintain blood pressure | 96 | 120 
ventilator to assist breathing | 96 | 120 
intravenous hydration to enlarge blood capacity | 96 | 120 
nutritional support therapy | 96 | 120 
blood transfusion | 96 | 120 
blood cultures and drainage fluids sent | 96 | 96 
empirically started on intravenous tigecycline and piperacillin/tazobactam | 96 | 120 
temperature went up to 39.3°C | 120 | 120 
pulse rate of 130 beats/minute | 120 | 120 
leukocyte count of 35.9×10^9/L | 120 | 120 
neutrophils 92.4% | 120 | 120 
procalcitonin level of 8.15 ng/mL | 120 | 120 
C-reactive protein level of 174 mg/L | 120 | 120 
anaerobic blood culture vials drawn postoperatively were reported to be positive | 144 | 144 
Gram stain revealed short Gram-positive bacillus without spores | 144 | 144 
positive culture broth was inoculated onto blood agar base medium | 144 | 144 
anaerobically incubated for three more days | 144 | 168 
colony from the agar plate was identified as E. lenta by matrix-assisted laser desorption/ionization time-of-flight mass spectrometry | 168 | 168 
plasma fibrinogen fell to 1.0 g/L | 168 | 168 
tigecycline was replaced by teicoplanin | 168 | 168 
piperacillin/tazobactam was discontinued | 168 | 168 
ertapenem was added to teicoplanin | 168 | 168 
cultures of the drainage fluid were obtained with the isolation of organism as Escherichia coli | 168 | 168 
Escherichia coli was susceptible to ertapenem | 168 | 168 
treated with ertapenem and teicoplanin | 168 | 240 
fever, leukocytosis, procalcitonin level and C-reactive protein level promptly improved | 168 | 240 
transferred to the general ward | 240 | 240 
administered ertapenem and teicoplanin for another 14 days | 240 | 384 
debridement, dressing change and symptomatic supportive treatment | 240 | 384 
repeated blood cultures after the introduction of antibiotics were negative | 240 | 384 
repeat CT revealed that the size of the hepatic abscess and the amount of ascites decreased | 384 | 384 
further 7-day course of intravenous ertapenem and teicoplanin | 384 | 432 
symptoms achieved further alleviation | 432 | 432 
discharged from the hospital | 432 | 432 
prescription for oral antibiotics (clindamycin) | 432 | 432 
remained well as an outpatient | 432 | 504 
no recurrence of fever | 504 | 504 
complete resolution of the abscess | 504 | 504 
six-week course of intravenous ertapenem | 504 | 504