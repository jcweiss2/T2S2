68 years old | 0
woman | 0
diagnosed with CLL/SLL | 0
inguinal lymph node biopsy | 0
bone marrow biopsy | 0
FCR therapy | 0
completed 6 cycles | 0
total thyroidectomy | 0
chronic lymphocytic thyroiditis | 0
Hurthle cell adenoma | 0
excision of basal cell carcinoma | 0
chest wall | 0
lost to follow-up | 0
cervical lymphadenopathy | 0
modified treatment with Rituxan and Bendamustine | 0
FISH peripheral blood | 0
mono-allelic deletion of 13q14.3 locus | 0
regression of cervical lymphadenopathy | 0
complete remission | 0
left axillary lymphadenopathy | 0
CT imaging demonstrated 3.5 cm left axillary lymph node | 0
enlarged retroperitoneal lymph nodes | 0
enlarged mesenteric lymph nodes | 0
planned to start on Gazyva and Venetoclax | 0
Venetoclax held | 0
Gazyva given | 0
completed 3 doses of Gazyva | 0
clinical improvement | 0
regression of mesenteric lymphadenopathy | 0
Venetoclax dose held | 0
presented to Emergency Department | 0
recurrent fever (39.2°C) | 0
weakness | 0
abdominal pain | 0
vomiting | 0
elevated alkaline phosphatase (961 U/L) | 0
AST 10 | 0
ALT 26 | 0
total bilirubin 1.4 | 0
negative hepatitis A, B, C serology | 0
negative ANA | 0
negative ASMA | 0
no duct dilatation | 0
no gallbladder thickening | 0
no peripancreatic ascites | 0
extensive splenomegaly | 0
splenic varicosities | 0
ascites | 0
porta hepatis lymphadenopathy | 0
CT abdomen and chest confirmed hepatosplenomegaly | 0
enlarged intra-abdominal lymph nodes | 0
pleural effusion | 0
liver biopsy performed | 0
periportal fibrosis | 0
histiocytic-predominant inflammation | 0
acute granulomatous hepatitis | 0
hemophagocytosis | 0
no steatosis | 0
no cholestasis | 0
no malignancy | 0
no infectious agents (AFB and fungus) | 0
peritoneal fluid sparse normal-appearing small lymphocytes | 0
negative for carcinoma | 0
bone marrow biopsy suggested | 0
declined by patient | 0
received blood transfusion | 0
consultations by gastroenterology | 0
consultations by infectious disease | 0
consultations by hematology/oncology | 0
treated for neutropenic fever | 0
hypotension (BP 85/57 mmHg) | 0
transferred to Intensive Care Unit | 15
septic shock | 15
remained on vasopressors | 15
low blood pressure | 15
increasing respiratory distress | 15
hypoxia | 15
died | 72
autopsy showed diffuse lymphadenopathy | 72
multi-organ involvement by large atypical cells | 72
Reed-Sternberg cells (positive for CD30, CD15, Pax 5, Bcl-2, EBV (EBER)) | 72
negative CD20, ALK, CD138, kappa/lambda in situ hybridization | 72
CD68 predominant granulomatous areas in liver | 72
negative CD30 and T cell markers (CD5) | 72
negative anaplastic large T cell (ALCL) | 72
negative histiocyte-rich T-cell lymphoma | 72
CD30/CD15 abnormal large neoplastic cells in abdominal lymph nodes | 72
CD30/CD15 abnormal large neoplastic cells in para-aortic lymph nodes | 72
CD30/CD15 abnormal large neoplastic cells in mesenteric lymph nodes | 72
CD30/CD15 abnormal large neoplastic cells in perihilar lymph nodes | 72
CD30/CD15 abnormal large neoplastic cells in bilateral lungs | 72
CD30/CD15 abnormal large neoplastic cells in liver | 72
CD30/CD15 abnormal large neoplastic cells in spleen | 72
CD30/CD15 abnormal large neoplastic cells in pancreatic surface | 72
CD30/CD15 abnormal large neoplastic cells in fallopian tubes | 72
CD30/CD15 abnormal large neoplastic cells in bone marrow | 72
final diagnosis of CLL with transformation to Hodgkin’s lymphoma | 72
cause of death: sepsis | 72
