4 years old|0
girl|0
developmental delay|0
myelomeningocele|0
hydrocephalus|0
neurogenic bladder|0
recurrent urinary tract infections|0
urosepsis|-1440
hemolytic uremic syndrome|-1440
chronic renal failure|0
peritoneal dialysis|0
seizure-like activity|-24
fever|-24
distress|0
tachycardic|0
tachypneic|0
distended abdomen|0
normal oxygen saturations|0
lorazepam|0
fosphenytoin|0
antibiotics|0
chest x-ray|0
enlarged cardiac silhouette|0
transthoracic echocardiogram|0
moderate circumferential pericardial effusion|0
diastolic right atrial collapse|0
tamponade physiology|0
intravenous induction|0
endotracheal intubation|0
6-French pigtail catheter|0
pericardial space|0
220 ml serosanguineous fluid drained|0
pericardial drainage minimal|48
decision to discontinue drain|48
attempted removal|48
unresponsive|48
decreased respiratory rate|48
bradycardia|48
chest compressions|48
bag mask ventilation|48
breathing spontaneously|48
palpable pulse|48
chest x-ray|48
transfer to operating room|48
TTE-guided withdrawal|48
general anesthesia|48
minimal effusion|48
another attempted removal|48
profoundly hypotensive|48
bradycardic|48
external cardiac compressions|48
0.35 flex guidewire|48
catheter advanced into chest|48
hemodynamic stabilization|48
drain encircling major vessel|48
surgical removal via sternotomy|48
catheter course anteriorly and superiorly over pulmonary artery and aorta|48
catheter course posteriorly and inferiorly under heart|48
pigtail adjacent to atrial appendage|48
traction on catheter|48
complete occlusion of main pulmonary artery|48
severe reduction in pulmonary blood flow|48
abrupt fall in end-tidal carbon dioxide|48
drain surgically removed|48
recovery in pediatric intensive care unit|48
