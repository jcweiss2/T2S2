36 years old | 0
male | 0
admitted to the hospital | 0
COVID-19 | 0
persistent fever | -168
dry cough | -168
coryzal symptoms | -72
intubated and ventilated | -24
type 1 respiratory failure | -24
lower/mid zone and multiple peripheral opacities | 0
positive SARS-CoV-2 PCR swab result | 48
proinflammatory process | 0
raised C-Reactive Protein (CRP) | 0
ferritin | 0
D-dimer | 0
lymphocytopaenia | 0
neutrophilia | 0
concurrent bacterial infection | 0
nasogastric tube placement | 0
enteral tube feeding | 0
estimated energy requirements | 0
Penn State protocol | 0
Mifflin-St.Jeor formula | 0
ESPEN recommendations | 0
high energy/protein feeds | 0
propofol | 0
sedation | 0
paralysis | 0
proning | 0
ventilatory support | 0
pulmonary embolism (PE) | 0
CT pulmonary angiogram | 0
non-occlusive right lower lobe segmental and subsegmental PE | 0
extensive COVID-19 pneumonitis | 0
early evidence of fibrotic change | 0
multiple antibiotic therapies | 0
elevated procalcitonin | 0
ventilating in the prone position | 0
metabolic and logistical impacts | 0
low volume feeding | 0
gastrointestinal symptoms | 0
cyclical phases of bowels | 0
constipation | 0
abdominal distension | 0
laxatives/enemas | 0
gastric aspirates | 0
prokinetics | 0
severe weight loss | 1248
deconditioning | 1248
reduced appetite | 1248
poor oral intake | 1248
modified texture diet | 1248
enteral tube feeding | 1250
oral nutritional supplements | 1250
discharged | 1312
vitamin D levels | 1008
insufficient levels | 1008
Pabrinex | 0
vitamin preparation | 0
refeeding syndrome | 0
electrolyte disturbances | 0
water-soluble vitamins | 0
micronutrients | 0
deficiencies | 0
Black, Asian and Minority Ethnic communities | 0
supplementary parenteral nutrition | 0
logistical challenges | 0
enhanced dietetic roles | 0
anthropometric measures | 0
physical assessments | 0
gastric residual volumes | 0
nasogastric tube (NGT) placement | 0
feed delivery | 0