76 years old | 0
female | 0
diagnosed with mesenteric ischemia | 0
scheduled for emergency laparotomy | 0
Mallampati Class 2 | 0
no restriction of mouth opening | 0
no anticipated difficulty in intubation | 0
flexion of the neck normal | 0
extension of the neck normal | 0
blood pressure 100/70 mmHg | 0
tachycardia |%0
tachypnea | 0
ASA Grade IV E | 0
hypertensive | 0
diabetic | 0
past history of coronary artery disease | -?
ongoing mesenteric ischemia | 0
severe sepsis syndrome | 0
acute respiratory distress syndrome | 0
low hemoglobin 7.6 g/dL | 0
mild hyponatremia 128 mmol/l | 0
consultation with patient's relatives | 0
general anesthesia | 0
rapid sequence induction | 0
intubation | 0
preoxygenated for 5 min | 0
Sellick's maneuver applied | 0
pentothal sodium 150 mg IV | 0
rocuronium 100 mg IV | 0
attempt to open mouth after 1 min | 60
teeth firmly approximated | 60
mouth could not be opened | 60
no peripheral nerve stimulator | 60
second attempt 1 min later | 120
failed to open mouth | 120
failure to intubate | 120
mask ventilation attempted | 120
continued Sellick's maneuver | 120
jaw locked | 120
airway obstruction | 120
attempted nasopharyngeal airway | 120
every attempt unsuccessful | 120
teeth firmly opposed | 120
blind nasal intubation attempted | 120
unsuccessful blind nasal intubation | 120
no anticipated difficult ventilation | 0
equipment not prepared | 0
fiberoptic bronchoscope not available | 0
ineffective ventilation | 120
oxygen saturation decreased to 92% | 120
decision for tracheostomy | 120
surgeon summoned | 120
tracheostomy performed | 120
patient desaturating | 120
hemodynamics deteriorating | 120
sustained cardiac arrest | 120
could not be revived | 120
attempt to pull jaw anteriorly | 120
no forward motion of TMJ | 120
mouth opened 1 cm | 120
no history of TMJ disorders | -?
malignant hyperthermia questioned | 0
masseter spasm questioned | 0
no triggering drugs received | 0
TMJ displacement | 120
patient demise | 120
