42 years old | 0
male | 0
admitted to the hospital | 0
severe shock | 0
febrile | 0
sedated with propofol | 0
invasive mechanical ventilation | 0
vasopressor and ionotropic support | 0
noradrenaline 0.5 μg/kg/min | 0
dobutamine 5 μg/kg/min | 0
systolic heart murmur | 0
abdomen soft | 0
no tenderness to deep palpation | 0
leukocytosis | 0
anemia | 0
prolonged international normalized ratio | 0
high prothrombin time | 0
acute kidney injury | 0
elevated aminotransferases | 0
hyperbilirubinemia | 0
elevated lactate dehydrogenase | 0
pro-calcitonin | 0
N-terminal pro b-type natriuretic peptide | 0
troponin | 0
metabolic acidemia | 0
high lactate levels | 0
left ventricle hypertrophy | 0
moderate-to-severe depression of global systolic function | 0
severe auricular dilatation | 0
thrombus in left auricular appendix | 0
native aortic valve vegetation | 0
severe septic shock | 0
multiple-organ dysfunction | 0
endocarditis | 0
empirical broad-spectrum antibiotics | 0
transferred to intensive care unit | 0
drug abuse history unknown | 0
negative for secondary causes of immunosuppression | 0
negative for syphilis | 0
blood cultures positive for Corynebacterium jeikeium | 0
initial clinical improvement | -216
severe hypotension | 216
vasopressor support re-introduced | 216
noradrenaline 1.9 μg/kg/min | 216
blood seen on nasogastric tube | 216
urgent upper endoscopy | 216
circumferential hemorrhagic mucosa | 216
fibropurulent plaques | 216
violaceus areas of elevated mucosa | 216
loss of vascular pattern | 216
pale mucosa | 216
hemorrhagic mucosa | 216
multiple erosions | 216
fibropurulent plaques | 216
biopsies consistent with extensive hemorrhagic necrosis | 216
acute kidney failure | 216
probable ischemic pancreatitis | 216
hepatitis | 216
contrast-enhanced abdominal computed tomography | -48
no alterations suggestive of intestinal ischemia | -48
no alterations suggestive of chronic liver disease | -48
died | 240
refractory multiple-organ dysfunction | 240