32 years old | 0
Gravida 2 Para 2 | 0
presented on postpartum day 7 | 0
uncomplicated late-term vaginal delivery | 0
fevers | 0
chills | 0
left distal lower extremity pain | 0
swelling | 0
swelling in the right knee | 0
denied recent injury | 0
unable to bear weight on the left side | 0
diffuse rash involving upper abdomen | 0
denied other postpartum complications | 0
continued breastfeeding | 0
history of stage IIa malignant peripheral nerve sheath tumor | -8760
in remission | -8760
treated 1-year prior | -8760
complete surgical excision | -8760
no chemotherapy | -8760
admitted in labor | 0
420/7 weeks gestation | 0
uncomplicated antepartum course | 0
group B streptococcus carrier screening negative | 0
small labial lacerations | 0
first-degree midline lacerations | 0
repaired at time of delivery | 0
minimal blood loss | 0
unremarkable postpartum course | 0
discharged home on postpartum day 1 | 24
reported fevers to 104°F at home | 144
temperature of 97.5°F | 0
heart rate of 68 bpm | 0
respiratory rate of 18 | 0
blood pressure of 107/69 | 0
mild distress | 0
moderate tight-like pain | 0
limited range of motion of left lower extremity | 0
focal area of erythema at left ankle | 0
exquisitely tender to palpation | 0
right knee swollen | 0
asymmetric in size | 0
peripheral pulses present | 0
nonperitoneal abdomen | 0
mildly tender uterus | 0
fundus firm at 4-cm below umbilicus | 0
faint maculopapular rash | 0
scant nonpurulent lochia | 0
leukocytosis 18,800 | 0
bandemia 23.7% | 0
lactate 1.6% | 0
urine culture with S. pyogenes | 0
orthopaedics consulted | 0
concern for compartment syndrome | 0
concern for necrotizing infection | 0
plain X-ray showed soft tissue edema | 0
no osseous abnormalities | 0
Doppler ultrasonography negative for deep vein thrombosis | 0
left ankle arthrocentesis | 0
normal appearing fluid | 0
heart rate 144 bpm | 2
temperature 102.6°F | 2
respiratory rate 20 | 2
MAP 66 | 2
SpO2 98% | 2
aggressive fluid resuscitation | 2
blood cultures obtained | 2
IV amoxicillin-sulbactam | 2
IV clindamycin | 2
suspicion for invasive GAS infection | 2
concern for TTS | 2
transfer to ICU | 2
CT of left lower extremity | 2
severe inflammation | 2
no abscess | 2
no necrotizing fasciitis | 2
severe pain | 2
left distal lower extremity fasciotomy | 2
no purulence | 2
no necrotic tissue | 2
normal appearing fascia | 2
edematous lateral compartment | 2
improvement in pain | 2
received albumin | 2
received norepinephrine | 2
received esmolol | 2
pressure support | 2
control of tachycardia | 2
received gentamicin for 48 hours | 2
endometritis coverage | 2
unclear source of infection | 2
tender uterus | 2
received therapeutic enoxaparin | 2
septic pelvic thrombophlebitis | 2
tachycardia resolved | 5
fevers resolved | 5
leukocytosis resolved | 5
stable for transfer out of ICU | 5
residual peroneal nerve palsy | 5
required reoperation on hospital day 8 | 192
concerns for myositis | 192
small area of purulence | 192
decreased contractility of anterior compartment | 192
no other abnormalities | 192
fever to 102.2°F on hospital day 13 | 312
new leukocytosis | 312
worsening pain in right knee | 312
arthrocentesis performed | 312
purulent fluid | 312
right knee arthroscopy | 312
synovectomy | 312
debridement | 312
inflamed proliferative synovium | 312
repeat right knee arthroscopic incision and drainage on hospital day 15 | 360
negative culture | 360
transitioned to IV penicillin G | 408
discharged on hospital day 19 | 456
continued treatment with IV penicillin | 456
additional 14 days of oral amoxicillin | 456
suspected endometritis | 456
no definite primary source | 456
cystitis less likely | 456
contamination with vaginal fluid | 456
continued physical and occupational therapy | 456
residual peroneal palsy | 456
no evidence of osteomyelitis | 456
chondromalacia of left patella | 456
ongoing pain | 456
diminished range of motion | 456
poor flexion | 456
poor wound healing | 456
consultation with outside orthopaedic facility | 456
multiple enlarged inguinal lymph nodes | 456
lymphadenopathy suspected reactive | 456
excisional biopsy of lymph node | 456
wound debridement | 456
lymph node biopsy negative for tumor | 456
reactive follicular hyperplasia | 456
blood cultures resolved | 456
resolution of GAS infection | 456
ongoing orthopaedic care | 456
physical therapy | 456
occupational therapy | 456
residual deficits | 456
malignant peripheral nerve sheath tumor in remission | -8760
