60 years old | 0
male | 0
homeless | 0
HIV positive | 0
CD4 count 604 | -744
HIV RNA PCR quantity 120,000 | -744
bilateral wrist pain | 0
left ankle swelling and pain | 0
pain 10/10 | 0
constant pain | 0
increased pain with movement | 0
no relief with ibuprofen | 0
history of gout attack | 0
denies intravenous drug abuse | 0
denies fever | 0
denies recent illness | 0
low grade fever 37.5 °C | 0
tachycardia 120 bpm | 0
non-toxic appearance | 0
no rashes | 0
limitation of active movement of bilateral wrists and left ankle | 0
warmth and tenderness to palpation in all 3 joints | 0
trace edema of the left ankle | 0
treated with colchicine | 0
treated with ibuprofen | 0
treated with hydrocodone/acetaminophen | 0
discharged home | 24
returned to ED with worsening pain | 72
returned to ED with erythema and swelling in left ankle | 72
returned to ED with new right ankle and left knee pain | 72
returned to ED with erythema and edema | 72
tachycardia 122 bpm | 72
labs obtained | 72
arthrocentesis of left knee performed | 72
treated with ketorolac | 72
peripheral WBC 9.4 | 72
uric acid 6.9 mg/dL | 72
joint aspirate WBC count 8.7 × 10^3 cells/μL | 72
no crystals | 72
discharged with nonsteroidal anti-inflammatory drugs | 96
discharged with rheumatology follow up | 96
diagnosis of inflammatory arthritis | 96
found unresponsive on a bench | 120
given naloxone without response | 120
hypertension 151/84 | 120
temperature 36.3°C | 120
tachycardia 138 bpm | 120
entire left lower extremity edema | 120
purpura throughout left leg and right ankle | 120
CT of left leg showed edema | 120
head CT negative | 120
acute renal failure with Cr 2.2 | 120
peripheral WBC 6.6 with 17% bands | 120
knee cultures growing gram negative coccobacilli | 120
taken to OR for washout | 120
admitted to intensive care unit | 120
intubated for airway protection | 120
blood and cerebral spinal fluid cultures grew N. meningitides | 120
required xigris and levophed for septic shock | 120
multiple surgical procedures for debridement/washouts | 120
multiple surgical procedures for I&Ds of bilateral lower extremities | 120
infected wounds from purpura fulminans | 120
wound vac management | 120
skin grafts to left lower extremity | 120
episode of acute renal failure due to urinary retention | 120
hydronephrosis | 120
urology consult | 120
taught to perform in-and-out catheterizations | 120
diagnosed with mild syndrome of inappropriate antidiuretic hormone | 120
placed on fluid restriction | 120
left-sided hearing loss due to meningitis | 120
developed right upper extremity deep vein thrombosis | 120
bridged from enoxaparin to warfarin | 120
treated for hospital-acquired urinary tract infections | 120
required multiple blood transfusions | 120
placed on nutritional supplementation for malnourishment | 120
neurology consult | 120
negative magnetic resonance image of the brain | 120
electroencephalography | 120
infectious disease consult | 120
treated with ceftriaxone | 120
treated with vancomycin and meropenem | 120
discharged to sub-acute rehabilitation facility | 1488