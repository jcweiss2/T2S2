79 years old | 0
gentleman | 0
spontaneous pneumomediastinum | 0
subcutaneous emphysema | 0
pneumonia | 0
no pre-existing lung disease | 0
presented | -96
increased shortness of breath | -96
pleuritic chest pain | -96
fevers | -96
non-productive cough | -96
Parkinson’s disease | 0
ischaemic heart disease | 0
hiatus hernia | 0
endoscopically investigated for dysphagia | 0
no firm diagnosis | 0
MEWS of 5 | 0
tachycardic (130 bpm) | 0
tachypnoeic (36 bpm) | 0
hypotensive (105/68 mmHg) | 0
febrile (39.0°C) | 0
oxygen saturations 92% on room air | 0
ABG pH 7.503 | 0
pCO2 3.60 | 0
pO2 7.66 | 0
SO2 92.5% | 0
lactate 3.0 | 0
reduced air entry in right upper zone | 0
right basal crepitations | 0
WBC count 1.6 | 0
CRP 320 | 0
AKI stage 1 | 0
creatinine 108 | 0
urea 13.3 | 0
sinus tachycardia | 0
right lower zone consolidation | 0
aspiration pneumonia | 0
AKI secondary to sepsis | 0
intravenous amoxicillin | 0
intravenous metronidazole | 0
intravenous fluids | 0
afebrile | 72
blood pressure 118/76 mmHg | 72
oxygen saturations 92% on 2L oxygen | 72
respiratory rate 20 bpm | 72
CRP 297 | 72
WBC 8.0 | 72
improved renal function | 72
tachycardic | 96
tachypnoeic | 96
increasing oxygen requirements at rest | 96
coarse crackles in right lower zone | 96
switched to piperacillin with tazobactam | 96
switched to clarithromycin | 96
subcutaneous emphysema in right hemithorax | 96
subcutaneous emphysema in right neck | 96
subcutaneous emphysema in right upper limb | 96
oxygen saturation 90% on 35% oxygen | 96
oxygen titrated upwards to >94% | 96
ABG Type 1 Respiratory Failure | 96
pCO2 4.09 | 96
pO2 6.88 | 96
sO2 89.9% | 96
stable blood pressure | 96
soft abdomen | 96
non-tender abdomen | 96
no external chest wall trauma | 96
chest x-ray showing subcutaneous emphysema | 96
suspected pneumomediastinum | 96
urgent CT scan | 96
bilateral consolidation | 96
subcutaneous emphysema of chest extending to neck | 96
extensive pneumomediastinum | 96
right 2–3 mm anterior pneumothorax | 96
no pre-existing lung disease | 96
pneumomediastinum secondary to pneumonia | 96
subcutaneous emphysema secondary to pneumonia | 96
subcutaneous emphysema descended into abdominal wall | 120
subcutaneous emphysema descended into lower limbs | 120
discussed with cardiothoracic surgery | 120
discussed with interventional radiology | 120
no interventions possible | 120
intensive care review | 120
invasive ventilation would worsen situation | 120
non-invasive ventilation would worsen situation | 120
treated with high-flow oxygen | 120
non-breathe mask | 120
clindamycin prescribed | 120
piperacillin with tazobactam continued | 120
clarithromycin continued | 120
clinically deteriorated | 120
maximum ward-based treatment | 120
guarded prognosis | 120
lack of response to treatment | 120
DNAR decision | 120
reviewed by palliative care team | 120
died of septic shock | 216
