65 years old | 0
female | 0
admitted to the hospital | 0
fever | 0
chills | 0
pain in left leg | 0
parkinsonism | -8760
diabetes mellitus | -8760
levodopa / carbidopa | -8760
rasagiline | -8760
ropinirole | -8760
trihexyphenidyl | -8760
amantadine | -8760
metformin | -8760
glipizide | -8760
cellulitis | 0
intravenous clindamycin | 0
intravenous benzylpenicillin | 0
high-temperature spikes | 72
tachycardia | 72
tachypnea | 72
hypotensive | 72
encephalopathic | 72
shifted to ICU | 72
intravenous linezolid | 72
intravenous piperacillin with tazobactam | 72
vancomycin not considered | 72
hemodynamics improved | 72
anti-parkinsonism drugs continued | 72
oral hypoglycemic agents stopped | 72
switched to insulin | 72
confused | 96
drowsy | 96
disoriented | 96
altered sensorium | 96
myoclonus | 96
tremors | 96
jerky movements | 96
no neck stiffness | 96
computed tomography of the brain | 96
cerebrospinal fluid analysis | 96
improving white blood cell counts | 96
better glycemic control | 96
sterile blood and pus cultures | 96
high temperature | 120
altered mental status | 120
myoclonus | 120
jerky movements | 120
tremors | 120
serotonin syndrome suspected | 120
linezolid stopped | 120
rasagiline stopped | 120
temperature settled | 128
heart rate normal | 144
sensorium improved | 144
tremors subsided | 144
shifted out of the ICU | 192
started walking with support | 240
discharged from the hospital | 240
anti-parkinsonism drugs | 240
rasagiline added | 240
regular follow-up with neurologist | 240
stable and asymptomatic for serotonin syndrome | 240