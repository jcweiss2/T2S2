20 years old | 0
male | 0
Caucasian | 0
admitted to the hospital | 0
abdominal pain | -144
watery diarrhoea | -144
nausea | -144
vomiting | -144
fever | -144
chills | -144
cough | -144
shortness of breath | -144
evaluated at outside ED | -144
prescribed oral ciprofloxacin | -144
prescribed metronidazole | -144
colitis | -144
tachycardic | 0
normotensive | 0
oxygen saturation 94% | 0
posterior oropharynx erythematous | 0
exudates | 0
enlarged cervical lymphadenopathy | 0
tender bilateral cervical lymphadenopathy | 0
left inguinal lymphadenopathy | 0
diffuse abdominal tenderness | 0
scleral injection | 0
mild conjunctivitis | 0
negative SARS-CoV-2 PCR | -144
negative rapid antigen test | 0
leukocytosis | 0
lymphopenia | 0
thrombocytopenia | 0
elevated C-reactive protein | 0
low fibrinogen level | 0
elevated D-Dimer | 0
infectious workup negative | 0
blood cultures negative | 0
urine cultures negative | 0
stool enteric panel negative | 0
respiratory viral panel negative | 0
computed tomography of abdomen and pelvis | 0
right-sided colitis | 0
right mesenteric lymphadenopathy | 0
mild hepatosplenomegaly | 0
normal chest X-ray | 0
started on piperacillin–tazobactam | 0
tachycardic | 24
intermittent fevers | 24
hypotension | 24
IV fluid boluses | 24
transferred to MICU | 24
started on IV norepinephrine | 24
mild respiratory distress | 24
oxygen saturation 85% | 24
nasal cannula | 24
bilateral pulmonary oedema | 24
elevated pro-brain natriuretic peptide | 24
elevated troponin T | 24
dilated cardiac chambers | 24
reduced left ventricular systolic function | 24
mild global hypokinesis | 24
normal right ventricular systolic function | 24
normal aortic root | 24
small pericardial effusion | 24
mild pulmonic regurgitation | 24
mild tricuspid regurgitation | 24
diagnosed with COVID-19 | -672
infectious disease team consulted | 24
diagnosis of MIS-C/MIS-A | 24
treated with IVIG | 24
treated with IV methylprednisolone | 24
heart rate normalized | 28
defervesced | 28
improvement in abdominal pain | 28
weaned off norepinephrine | 48
transferred out of MICU | 48
transitioned to oral prednisone | 120
tapered over 3 weeks | 240
started on IV furosemide | 120
started on angiotensin-converting enzyme inhibitor | 120
discharged on lisinopril | 120
discharged on carvedilol | 120
discharged on furosemide | 120
follow-up after 3 months | 744
complete resolution of symptoms | 744
scheduled for trans-thoracic echocardiogram | 744