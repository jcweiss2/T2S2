51 years old | 0
male | 0
admitted to the ICU | 0
bilateral nephrectomy | -48
invasive urothelial cancer | -48
hemodynamic monitoring | 0
high fever | 48
distributive shock | 48
c-reactive protein elevated | 48
septic shock | 48
antibiotics started | 48
Tazocin | 48
amikacin | 48
noradrenaline infusion | 48
continuous veno-venous hemofiltration | 48
increased noradrenaline infusion | 72
high fever persisted | 72
infectiologist and microbiologist consultation | 72
senior nephrologist-intensivist consultation | 72
bilateral resection of adrenal glands | -48
Addison’s disease | 72
hydrocortisone administered | 72
condition normalized | 84
antimicrobials stopped | 84
discharged | 96