24 years old | 0 | 0 
female | 0 | 0 
admitted to the hospital | 0 | 0 
severe headache | -72 | 0 
projectile vomiting | -72 | 0 
no fever | -72 | 0 
no convulsions | -72 | 0 
no focal neurological deficit | -72 | 0 
symptomatic treatment outside | -72 | 0 
no relief | -72 | 0 
provisional diagnosis of metabolic encephalopathy | 0 | 0 
symptomatic treatment | 0 | 0 
altered sensorium | 24 | 24 
Glasgow Coma Scale-9 | 24 | 24 
high-grade fever | 24 | 24 
chills | 24 | 24 
dyselectrolytemia | 24 | 24 
low serum phosphate | 24 | 24 
neutrophilic leukocytosis | 24 | 24 
cerebrospinal fluid sent for evaluation | 24 | 24 
empirically treated with ceftriaxone | 24 | 24 
Gram stain of CSF | 24 | 24 
Gram-positive bacilli in CSF | 24 | 24 
polymorphs in CSF | 24 | 24 
lymphocytes in CSF | 24 | 24 
culture of CSF | 24 | 48 
Listeria monocytogenes in CSF | 48 | 48 
blood culture | 0 | 24 
Gram-positive bacilli in blood culture | 0 | 24 
Listeria monocytogenes in blood culture | 24 | 24 
switched to meropenem | 48 | 48 
clinical improvement | 72 | 72 
microbiological improvement | 72 | 72 
discharged | 168 | 168