58 years old | 0
male | 0
admitted to the hospital | 0
shock | 0
diffuse ST-elevation at the electrocardiogram | 0
fever | -168
persistent cough | -168
nasopharyngeal swab test positive for SARS-CoV-2 | -48
fever decreased after 5 days of levofloxacin | 120
current smoker | 0
hypothyroidism | 0
chest X-ray | -2160
pneumological consultation | -2160
interstitial lung disease | -2160
high-resolution lung CT scan | -2160
right lung mass suspected for cancer | -2160
endobronchial ultrasound-guided transbronchial needle aspiration planned | -2160
severe hypotension | 0
asthenia | 0
emergency service called | 0
blood pressure 80/40 mmHg | 0
heart rate 110 bpm | 0
oxygen saturation 88% | 0
body temperature 37.5°C | 0
emergency coronary angiography | 0
absence of coronary artery disease | 0
normal left ventricular function |EOT_STREAM_EOF
high inflammatory markers | 0
increased liver enzymes | 0
normal troponin values | 0
respiratory alkalosis | 0
hyperlactatemia | 0
interstitial syndrome with bilateral B lines | 0
small sub-pleural consolidations | 0
bilateral pleural effusion | 0
diffuse pericardial effusion | 0
swinging heart | 0
inferior caval vein 2.2 cm | 0
no respiratory excursion | 0
left ventricular ejection fraction 50% | 0
blood pressure increased after fluid therapy | 0
pericardiocentesis not performed | 0
oxygen saturation deteriorated | 0
high flow oxygen therapy | 0
diagnosis of pericarditis | 0
corticosteroids started | 0
colchicine started | 0
heparin prophylaxis started | 0
high dose aspirin avoided | 0
empiric antibiotic therapy | 0
second nasopharyngeal swab negative for SARS-CoV-2 | 48
third nasopharyngeal swab negative for SARS-CoV-2 | 72
positive IgM and IgG antibodies for SARS-CoV-2 | 0
hemodynamically stable | 0
severe respiratory failure persisted | 0
total body CT | 0
locally advanced lung cancer | 0
subclavian artery and vein involvement | 0
thoracic lymph nodes involvement | 0
pleural effusion | 0
pericardial effusion | 0
histological examination confirmed lung adenocarcinoma | 0
oncologic evaluation | 0
moved to oncologic clinic | 168
died | 432
