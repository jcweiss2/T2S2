48 years old | 0
female | 0
obesity | 0
hypertension | 0
admitted to the hospital | 0
endoscopic sleeve gastroplasty | 0
no immediate procedural related complications | 0
general anesthesia | 0
endoscopic suturing system | 0
carbon dioxide insufflation | 0
full thickness U-shaped suture pattern | 0
five sutures | 0
antiemetics | 0
dipyrone | 0
omeprazole | 0
discharged | 24
abdominal pain | 72
emergency department visit | 72
readmitted to the hospital | 96
poor general health status | 96
signs of peritoneal irritation | 96
computed tomography | 96
fluid in the abdominal cavity | 96
laparoscopy | 96
biliary ascites | 96
gallbladder sutured to the gastric wall | 96
cholecystectomy | 96
review and lavage of the abdominal cavity | 96
admitted to the intensive care unit | 96
antibiotic therapy | 96
discharged | 480
weight loss | 4320
excellent general condition | 4320