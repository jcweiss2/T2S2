76 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
atrial fibrillation | -672 | 0 | Factual
rheumatic heart disease | -672 | 0 | Factual
congestive heart failure | -672 | 0 | Factual
preserved ejection fraction | -672 | 0 | Factual
digoxin | -672 | 0 | Factual
coumadin | -672 | 0 | Factual
generalized malaise | -168 | 0 | Factual
shortness of breath | -168 | 0 | Factual
lower extremity swelling | -168 | 0 | Factual
subjective fever | -168 | 0 | Factual
no chest pain | -168 | 0 | Negated
no orthopnea | -168 | 0 | Negated
no paroxysmal nocturnal dyspnea | -168 | 0 | Negated
blood pressure 79/54 mmHg | 0 | 0 | Factual
oral temperature 38.3°C | 0 | 0 | Factual
heart rate 55 beats/min | 0 | 0 | Factual
crackles up to the mid-lung fields bilaterally | 0 | 0 | Factual
irregularly irregular heart rhythm | 0 | 0 | Factual
2+ pitting edema up to the knees | 0 | 0 | Factual
congestion in the bilateral lower lung fields | 0 | 0 | Factual
cardiomegaly | 0 | 0 | Factual
sodium level 126 | 0 | 0 | Factual
potassium 5.2 | 0 | 0 | Factual
blood urea nitrogen 33 | 0 | 0 | Factual
creatinine 2.77 | 0 | 0 | Factual
white blood count 4.9 | 0 | 0 | Factual
INR 2.8 | 0 | 0 | Factual
signs of digoxin toxicity | 0 | 0 | Factual
peak troponin level 0.20 ng/mL | 0 | 0 | Factual
digoxin level 3.6 ng/mL | 0 | 0 | Factual
admitted to the Cardiac Intensive Care Unit | 0 | 0 | Factual
digoxin immune fab | 0 | 0 | Factual
ejection fraction 45% to 49% | 0 | 0 | Factual
possible vegetation on the mitral valve | 0 | 0 | Factual
severe eccentric mitral and tricuspid regurgitation | 0 | 0 | Factual
mitral valve vegetation measuring 1.2×0.7 cm | 0 | 0 | Factual
severe biatrial enlargement | 0 | 0 | Factual
left atrium volume 101.40 mL/m2 | 0 | 0 | Factual
right atrium volume 233.80 mL/m2 | 0 | 0 | Factual
blood cultures positive for Pasteurella multocida | 0 | 0 | Factual
ceftriaxone | 0 | 0 | Factual
septic emboli | 0 | 0 | Factual
owned 4 cats | -672 | 0 | Factual
evaluated for multi-valve replacement surgery | 0 | 0 | Factual
biopsy of the vegetation | 0 | 0 | Factual
condition stabilized | 0 | 168 | Factual
discharged to a skilled nursing facility | 168 | 168 | Factual
6-week course of ceftriaxone | 168 | 504 | Factual
readmitted for congestive heart failure exacerbation | 720 | 720 | Factual
hospice care | 720 | 720 | Factual