73 years old | 0
female | 0
admitted to the hospital | 0
left nasal obstruction | -480
left side facial pain | -480
headache | -480
history of COVID-19 infection | -720
home isolation treatment | -720
no steroid use | -720
black mucopurulent secretion | 0
oroantral ulcer | 0
fungal hyphae | 0
mucormycosis | 0
maxillary sinusitis | 0
oroantral fistula | 0
endoscopic surgical debridement | 0
inj. AmB 5 mg/kg/day | 0
bronchial asthma | 0
hypertension | 0
uncontrolled diabetes mellitus | 0
regular treatment | 0
normal airway examination | 0
total leucocyte count of 14,000/μL | 0
fasting blood sugar of 246 mg/dL | 0
HbA1c of 10.9% | 0
normal ECG | 0
normal CXR | 0
normal echocardiography | 0
normal PFT | 0
preoperative optimisation | 0
regular insulin | 0
nebulisation with budesonide | 0
nebulisation with salbutamol | 0
antifungal | 0
antibiotics | 0
control of blood sugar | 0
COVID-19 negative result | 0
RT-PCR test | 0
written informed consent | 0
inj. glycopyrrolate 0.2 mg | 0
inj. fentanyl 100 μg | 0
intravenous propofol | 0
vecuronium | 0
endotracheal tube | 0
oxygen | 0
nitrous oxide | 0
isoflurane | 0
controlled ventilation | 0
capnography | 0
neuromuscular monitoring | 0
urine output | 0
stable intraoperatively | 0
reversal of anaesthesia | 24
extubation | 24
postoperative ICU care | 24
inj. AmB | 24
monitoring of renal parameters | 24
monitoring of blood sugar | 24
discharge from ICU | -1 
Note: The time stamp for "discharge from ICU" is not mentioned in the text, so it is assumed to be after 24 hours.