60 years old | 0
male | 0
African descent | 0
gastroesophageal reflux disease | -7200
admitted to the hospital | 0
diffuse joint pain | -2160
joint swelling | -2160
diffuse rash | -2160
headaches | -2160
generalized weakness | -2160
subjective fevers | -2160
chills | -2160
profuse night sweats | -2160
unintentional 30-pound weight loss | -2160
pruritic rash | -2160
rash on face | -2160
rash on body | -2160
bilateral eye pain | -2160
eye swelling | -2160
double vision | -2160
mild vision blurriness | -2160
muscle weakness | -2160
dysphagia | -2160
diffuse alopecia | -2160
adjacent scarring | -2160
polymorphous rash | 0
hypopigmentation | 0
hyperpigmentation | 0
eczematous-like macules | 0
eczematous-like patches | 0
edematous joints | 0
tender joints | 0
symmetrical facial weakness | 0
decreased facial sensation | 0
proximal muscle weakness | 0
distal muscle weakness | 0
decreased muscle bulk | 0
increased muscle tone | 0
positive Babinski reflex | 0
hyperreflexive joint reflexes | 0
normocytic anemia | 0
thrombocytopenia | 0
elevated liver enzymes | 0
mild leukopenia | 0
unremarkable MRI scan | 0
unremarkable imaging | 0
mixed connective tissue disease | 0
dermatomyositis | 0
systemic lupus flare | 0
negative rheumatological panel | 0
perivascular dermatitis | 0
dermal mucin deposition | 0
negative infectious disease workup | 0
no signs of malignancy | 0
no monoclonal gammopathy | 0
mild muscle pain | 24
subcutaneous edema | 48
myositis | 48
focal myopathy | 72
denervation atrophy | 72
high-dose parenteral steroids | 72
immunosuppressive therapy | 72
oral hydroxychloroquine | 72
no clinical improvement | 120
worsening respiratory distress | 168
severe sepsis | 168
transferred to intensive care unit | 168
declined further escalation of care | 168
declined autopsy | 168
died | 168
gingival mucosal biopsy | 168
focal amyloid deposition | 168
novel mutation in gelsolin gene | 168
C>G1375 transversion | 168
proline 459 to arginine | 168
gelsolin domain 4 mutation | 168
widespread amyloidogenic protein deposition | 168
mucosal gingival involvement | 168
suspected liver involvement | 168
suspected heart involvement | 168
suspected kidney involvement | 168
gelsolin amyloid angiopathy | 168
nodular vascular amyloid deposition | 168
vascular amyloid staining | 168
amyloid deposits positive for Sulfated Alcian Blue | 168
atrophic myofibers | 168
systemic inflammatory syndrome | 168
multiorgan dysfunction | 168
novel mutation | 168
distinct clinical syndrome | 168
importance of considering rare diseases | 168
importance of considering atypical presentations | 168
amyloidosis consideration in multisystem pathology | 168
future research | 168
potential therapeutic targets | 168
decrease disease burden | 168
improve quality of life | 168