hypertension | 0
degenerative joint disease | 0
bilateral knee replacement | 0
substance abuse | 0
trauma to face and chest wall | 0
lightheadedness | 0
fatigue | 0
leukocytosis | 0
hemoglobin of 10.2 g | 0
venous lactic acid of 2.4 mol/l | 0
intramuscular and subpectoral hematoma in the right chest wall | 0
extrapleural extension into the chest | 0
acute right second through fifth anterior rib fractures | 0
bilateral lower lobe bronchopneumonia | 0
blood cultures obtained | 0
started on empiric antibiotics with intravenous piperacillin–tazobactam | 0
afebrile | 0
hypotensive with blood pressure of 60/40 mmHg | 0
admitted to the intensive care unit for suspected septic shock | 0
initiation of vasopressors | 0
antibiotics broadened to intravenous vancomycin, cefepime and metronidazole | 48
repeat blood, urine and sputum cultures obtained | 48
sputum cultures grew methicillin-resistant Staphylococcus aureus | 72
antibiotics narrowed to intravenous vancomycin | 96
left knee pain | 120
notable swelling on physical exam | 120
concern for infection of prosthetic knee joint | 120
sterile left knee aspiration | 120
synovial fluid was cloudy, amber colored | 120
white blood cells of 9.28 × 10^3/mcL | 120
calcium pyrophosphate crystals | 120
complete washout and debridement of the joint with retention of the prosthesis | 144
operative note described an infected knee with purulence | 144
antibiotic regimen transitioned to intravenous cefazolin | 168
cultures from the infected area grew C. bifermentans | 240
antibiotic regimen transitioned to intravenous ampicillin–sulbactam | 240
contrast computerized tomography scan of the abdomen | 240
human immunodeficiency virus screening | 240
discharged to a rehabilitation facility | 384
recovered full range of motion of his left knee | 744
no signs of lingering joint or systemic infection | 744
still taking Augmentin | 744
reported medication adherence | 744
had not yet opted to undergo colonoscopy | 744