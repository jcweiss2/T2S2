67 years old | 0
male | 0
admitted to the hospital | 0
SAP | 0
chronic pancreatitis | -672
diabetes | -672
consumed 5 liters of beer every day | -672
body temperature 36.6 | 0
blood pressure 172/94 mmHg | 0
heart rate 96 beats/min | 0
respiratory rate 21 breaths/min | 0
abdomen hard and flat with tenderness and defensiveness | 0
increased white blood cell count | 0
increased serum concentrations of C-reactive protein | 0
increased serum concentrations of amylase | 0
increased serum concentrations of lipase | 0
HbA1c 9.6% | 0
fluid resuscitation | 0
nafamostat mesylate | 0
antibiotics | 0
ICU | 0
abdominal pain improved | 12
inflammation improved | 12
high fever | 384
Candida albicans detected in blood | 384
Candida albicans detected in central venous catheter | 384
candidemia | 384
ophthalmologic examinations | 384
candida endophthalmitis | 384
exudative plaques consistent with fungal infection | 384
micafungin | 384
caspofungin | 384
fluconazole | 384
blood cultures evaluated weekly | 391
disappearance of C. albicans from bloodstream | 434
exudative plaques disappeared | 434
β-D glucan negative | 434
discharged | 2280
visual disturbance denied | 384 
no urinary tract infection | 384
no pneumonia | 384
no infected pancreatic fluid | 384