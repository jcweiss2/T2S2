66 years old | 0
male | 0
admitted to the Dermatology Clinic | 0
rash | -48
erythemato-violaceous macules and papules | -48
postblister erosions on the oral and nasal mucosa | -48
genital areas with deep fissures | -48
painful burning sensations | -48
prodromal flu-like symptoms | -48
fever | -48
fatigue | -48
malaise | -48
complicated diabetes mellitus type II | 0
chronic kidney disease Stage 5 | 0
chronic haemodialysis | 0
obstructive nephropathy | 0
right nephrostomy | 0
secondary renal hypertension | 0
mixed decompensate toxic cirrhosis | 0
hepatic encephalopathy | 0
insulin 10 UI b.i.d. | 0
amlodipine 5 mg q.d. | 0
carbamazepine 100 mg q.d. | 0
onset of illness | -48
hospitalized for haemodialysis | -48
itchy erythemato-papulous rash | -48
prodromal flu-like symptoms | -48
fever | -48
fatigue | -48
malaise | -48
extension of the rash | -24
appearance of purpuric elements | -24
flaccid blisters | -24
large areas of denudation | -24
preliminary diagnosis of drug-induced allergic vasculitis | -24
transferred to the Department of Dermatology | 0
malaise | 0
itchy rash | 0
erythemato-violaceous macules and papules | 0
flaccid blisters | 0
erosions | 0
denudation | 0
high blood pressure | 0
increased abdominal volume | 0
collateral venous circulation | 0
marked anemia | 0
leukocytosis | 0
neutrophilia | 0
thrombocytopenia | 0
inflammatory syndrome | 0
elevated ASLO titer | 0
elevated IgE | 0
nitrogen retention syndrome | 0
elevated blood sugar levels | 0
hydro-electrolyte imbalance | 0
abnormal liver function | 0
Gram stain and culture from genital secretion and skin lesions | 0
nasal swab | 0
bacterial supra-infection with Klebsiella pneumoniae | 0
diagnosis of toxic epidermal necrolysis | 0
drug reaction syndrome due to carbamazepine | 0
pulse-therapy with corticosteroid | 0
topical corticosteroids | 0
topical antiseptics | 0
antibiotics | 0
hydro-electrolyte rebalancing | 0
worsening condition of associated pathologies | 24
high blood sugar values | 24
worsening of nitrogenous retention | 24
low alkaline reserve | 24
hyponatremia | 24
hypokalemia | 24
episode of upper gastrointestinal hemorrhage | 24
transferred to an ICU | 24
treatment in the ICU | 24
satisfactory resolution of the muco-cutaneous aspects | 72
reduction in corticosteroids | 72
complete discontinuation of systemic corticosteroid | 120
resumption of dialysis | 120
electrolyte rebalancing | 120
normalization of renal function | 120
acid-basic balance | 120
discharged from the hospital | 360
advice to stop carbamazepine | 360
medically related drugs | 360