64 years old | 0
    male | 0
    history of chronic pancreatitis | 0
    pseudocysts | 0
    ascites | 0
    presented to outside hospital | 0
    increasing abdominal pain | 0
    hypoxic respiratory failure | 0
    hypotension | 0
    intubated | 0
    transferred to medical intensive care unit | 0
    treated for septic shock | 0
    infected pancreatic pseudocyst | 0
    severe necrotizing pancreatitis | 0
    CT imaging demonstrated 10.2 × 7.8 cm pseudocyst in head of pancreas | 0
    thrombosis in portal vein | 0
    thrombosis extending into splenic vein | 0
    thrombosis extending into superior mesenteric vein | 0
    diagnosed during previous admission | -168
    treated with anticoagulation | -168
    aggressive resuscitation | 0
    pseudocyst drainage by interventional radiology | 0
    complicated course | 0
    hematemesis | 0
    CT angiography demonstrated focus of arterial phase contrast media extravasation within pancreatic head pseudocyst | 0
    active hemorrhage from gastroduodenal artery | 0
    emergently brought to interventional radiology | 0
    therapeutic transcatheter embolization | 0
    conventional catheter angiogram of celiac artery showed occlusion of gastroduodenal artery | 0
    vasospasm | 0
    4-French catheter advanced into gastroduodenal artery | 0
    angiogram of proximal gastroduodenal artery demonstrated large bleeding pseudoaneurysm | 0
    extravasation into pseudocyst | 0
    microcatheter and guidewire advanced into pseudoaneurysm | 0
    2 mechanical detachable micro-coils deployed | 0
    post-coil embolization angiogram of celiac artery showed complete occlusion of gastroduodenal artery | 0
    no evidence of extravasation | 0
    post embolization superior mesenteric artery angiogram showed no active hemorrhage | 0
    clinical improvement over 6 weeks | 432
    discharged | 432
    anticoagulation for 6 months to treat superior mesenteric vein thrombosis | 432
    presented to outside hospital following fall | 2160
    hemothorax | 2160
    pneumothorax | 2160
    worsening ascites | 2160
    anasarca | 2160
    supratherapeutic INR of 4.9 | 2160
    transfused with 5 units of Fresh Frozen Plasma | 2160
    sudden cardiac arrest | 2160
    cardiopulmonary resuscitation | 2160
    2 rounds of epinephrine administration | 2160
    intubated | 2160
    transferred to institution | 2160
    two paracenteses performed | 2160
    8.5 L transudative fluid | 2160
    4.3 L transudative fluid | 2160
    portal venous hypertension | 2160
    CT angiography demonstrated persistent portal venous outflow obstruction | 2160
    chronic portal vein thrombosis extending into superior mesenteric vein | 2160
    referred to interventional radiology | 2160
    hepatic and portal vein venography | 2160
    core needle liver biopsy | 2160
    porto-systemic venous pressure measurement | 2160
    stent dilatation of portal vein and superior mesenteric vein | 2160
    right trans-jugular vein approach | 2160
    4-French catheter advanced into right hepatic vein | 2160
    two 19-gauge transvenous core needle liver biopsies obtained | 2160
    sheath needle used to puncture right hepatic vein into right portal vein branch | 2160
    4 French catheter advanced into portal vein | 2160
    portal vein venogram performed | 2160
    chronic occlusion of portal vein | 2160
    chronic occlusion of superior mesenteric vein | 2160
    reconstitution of portal vein in porta hepatis from collateral venous channels | 2160
    portal vein pressure measured as 20 Torr | 2160
    right hepatic vein pressure measured as 17 Torr | 2160
    portosystemic gradient of 3 Torr | 2160
    4 French catheter exchanged for long 4 French sheath | 2160
    4 French catheter advanced through hepatic parenchymal track into portal vein | 2160
    advanced through chronically occluded segment of portal vein and superior mesenteric vein | 2160
    superior mesenteric vein venogram performed | 2160
    4 cm long occlusion of central superior mesenteric vein | 2160
    occlusion extending into portal vein | 2160
    superior mesenteric vein pressure measured as 26 Torr | 2160
    superior mesenteric vein to systemic pressure gradient of 9 Torr | 2160
    pressure gradient across occlusion of 6 Torr | 2160
    10 mm self-expanding Nitinol stent deployed | 2160
    stent dilated with 8-mm angioplasty balloon | 2160
    post-stent dilatation superior mesenteric vein venogram demonstrated widely patent veins | 2160
    no residual stenosis | 2160
    no extravasation | 2160
    no thrombosis | 2160
    no dissection | 2160
    pressure measurements in superior mesenteric vein | 2160
    right hepatic vein | 2160
    right atrium of heart | 2160
    superior mesenteric vein pressure of 25 Torr | 2160
    right hepatic vein pressure of 23 Torr | 2160
    right atrial pressure of 19 Torr | 2160
    reduction of superior mesenteric vein to systemic pressure gradient from 9 to 2 Torr | 2160
    innumerable venous collateral channels pre-stent | 2160
    no venous collateral channels post-stent | 2160
    hepatopetal blood flow post-stent | 2160
    clinical symptom improvement | 2160
    discharged following day | 2184
    readmitted for lethargy | 2400
    hypotension | 2400
    recurrent ascites | 2400
    improved ascites | 2400
    superior mesenteric vein stent partially occluded | 2400
    anticoagulation resumed | 2400
    discharged 3 days later | 2424
    recovered remarkably | 2424
    asymptomatic at 3 months | 2424
    free of ascites at 3 months | 2424
    asymptomatic at 7 years | 2424
    free of ascites at 7 years | 2424
    duplex ultrasound at 3 months | 2424
    duplex ultrasound at 7 years | 2424
    widely patent superior mesenteric vein | 2424
    widely patent portal vein | 2424
    no ascites | 2424
    partial occlusion of SMV stent 1 week post-procedure | 2400
    anticoagulation resumed | 2400
    symptoms improved | 2400
    <|eot_id|>
    