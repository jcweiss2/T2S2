60 years old | 0
    male | 0
    vitiligo | 0
    anemia | 0
    presented to the emergency department | 0
    diffuse itchy skin | -504
    occupational exposures at a metal refinery | 0
    occupational exposures at a shipping dock | 0
    active pack-per-day smoker | 0
    35-year smoking history | 0
    drinks alcohol daily | 0
    denies illicit drug use | 0
    sexually active with multiple female partners | 0
    no significant family history | 0
    no travel outside the United States | 0
    dry circular rashes | 0
    widespread inguinal adenopathy | 0
    widespread axillary adenopathy | 0
    widespread supraclavicular adenopathy | 0
    normal complete blood count | 0
    normal comprehensive metabolic panel | 0
    normal lactate dehydrogenase | 0
    normal angiotensin-converting enzyme | 0
    negative human immunodeficiency virus serology | 0
    discharged | 0
    nummular eczema | 0
    topical hydrocortisone 2.5% | 0
    cetirizine 10 mg | 0
    naproxen 500 mg | 0
    oral prednisone taper | 0
    followed-up with PCP | -744
    unremitting itching | -744
    edematous nasal mucosal | -744
    posterior oropharyngeal erythema | -744
    maculopapular erythematous rash | -744
    topical triamcinolone 0.5% | -744
    hydroxyzine 10 mg | -744
    referred to Dermatology | -2184
    persistent intense pruritus | -2184
    lesions on face | -2184
    lesions on chest | -2184
    lesions on abdomen | -2184
    denies constitutional symptoms | -2184
    differential diagnosis included sarcoidosis | -2184
    differential diagnosis included lichen planus | -2184
    differential diagnosis included disseminated lupus erythematosus | -2184
    differential diagnosis included lymphoma | -2184
    differential diagnosis included syphilis | -2184
    punch biopsies performed | -2184
    morphologic findings consistent with CTCL | -2184
    immunophenotypic findings consistent with CTCL | -2184
    molecular findings consistent with CTCL | -2184
    CD3+ | -2184
    CD4+ | -2184
    CD8+ | -2184
    CD4:CD8 ratio > 2:1 | -2184
    significant loss of CD7 lymphocyte staining | -2184
    CD20 highlighted rare-scattered B lymphocytes | -2184
    CD30+ present in less than 5% of cells | -2184
    Treponema pallidum stain negative | -2184
    positive T-cell gene rearrangement studies | -2184
    atypical lymphoid epidermal infiltrate | -2184
    highly irregular nuclear contour | -2184
    splitting at the dermal/epidermal junction | -2184
    inflammatory dermal infiltrate | -2184
    small lymphocytes | -2184
    histiocytes | -2184
    eosinophils | -2184
    CT/positron emission tomography scan | -2184
    moderately avid bilateral axillary lymph nodes | -2184
    enlarged bilateral axillary lymph nodes | -2184
    enlarged inguinal lymph nodes | -2184
    enlarged supraclavicular lymph nodes | -2184
    ultrasound-guided left axillary lymph node biopsy | -2184
    pathology demonstrated CTCL | -2184
    tumor staging IVA2 | -2184
    T4N3M0B0 classification | -2184
    more than 80% cutaneous involvement | -2184
    clinically abnormal peripheral lymph nodes | -2184
    CD25 staining negative | -2184
    serology for HTLV-1 not obtained | -2184
    initiated doxepin 25 mg | -2184
    initiated warfarin 1 mg | -2184
    evaluated by Cleveland Clinic Oncology | -2184
    confirmed diagnosis | -2184
    added clobetasol 0.05% | -2184
    added desonide | -2184
    added oral bexarotene 200 mg/m2 | -2184
    added gabapentin 300 mg | -2184
    presented to ED with bilateral foot pain | -2184
    presented to ED with swelling | -2184
    bilateral lower extremity duplex negative | -2184
    discharged | -2184
    returned to ED with extreme pain | 0
    open skin wounds draining yellow-green fluids | 0
    large eschar draining foul-smelling fluid on chest | 0
    multiple excoriating wounds covering more than 70% of body | 0
    admitted for wound care | 0
    admitted for broad-spectrum antibiotics | 0
    CT chest/abdomen/pelvis showed axillary adenopathy | 0
    enlarged bilateral inguinal lymph nodes | 0
    enlarged external iliac chain lymph nodes | 0
    multiple subcutaneous lesions along ventral abdominal wall | 0
    staging T4N3M0B0 | 0
    skin cultures grew MRSA | 0
    skin cultures grew Diphtheroid | 0
    taken to operating room for left inguinal lymph node excision | 24
    left anterior abdominal wall biopsy | 24
    debridement of chest wall eschar | 24
    pathology showed MF with large cell transformation | 24
    discontinued bexarotene | 24
    initiated romidepsin 14 mg/m2 | 24
    COVID-related transfer denials | 0
    discharge to skilled nursing facility delayed | 336
    transferred to ED | 0
    admitted for excruciating pain | 0
    admitted for infected skin lesions | 0
    care-navigation team revealed discharge recommendation | 0
    transfer to burn ICU denied | 0
    aggressive pain management initiated | 0
    broad-spectrum antibiotic therapy initiated | 0
    romidepsin held | 0
    extensive excisional debridement | 48
    wound cultures positive for MRSA | 48
    blood cultures revealed group B Streptococcus bacteremia | 48
    staging T4N3M0B1 | 48
    post-operative mechanical ventilation | 48
    transferred to surgical ICU | 48
    condition deteriorated | 96
    critically hypotensive | 96
    decreased urine output | 96
    leukocytosis | 96
    repeat blood cultures positive for group G streptococcus | 96
    repeat blood cultures positive for MRSA bacteremia | 96
    failed spontaneous breathing trial | 144
    code status changed to do not resuscitate | 240
    patient extubated | 240
    patient expired | 336
