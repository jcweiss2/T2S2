85 years old | 0\
    male | 0\
    type 2 diabetes mellitus | 0\
    hypertension | 0\
    furosemide | 0\
    hydralazine | 0\
    β-blocker | 0\
    dyslipidemia | 0\
    iron deficiency anemia | 0\
    ferrous sulphate | 0\
    chronic kidney disease | 0\
    dementia | 0\
    reduced oral intake | -168\
    recurrent vomiting | -168\
    decreased level of consciousness | -168\
    severely dehydrated | 0\
    hypotensive (92/58) | 0\
    mildly tachypneic (20) | 0\
    heart rate of 87 | 0\
    Glasgow coma scale of 11 | 0\
    melena | 0\
    leukocytosis (12 × 10^9) | 0\
    low hemoglobin (12.3 g/dL) | 0\
    high C-reactive protein (106 mg/L) | 0\
    high urea (53 mmol/L) | 0\
    acute kidney injury | 0\
    chronic kidney disease | 0\
    elevated lactate (4.6 mmol/L) | 0\
    elevated procalcitonin (4.88 ng/mL) | 0\
    urinary tract infection | 0\
    admitted to intensive care unit | 0\
    severe sepsis | 0\
    secondary to urinary tract infection | 0\
    acute on top of chronic kidney injury | 0\
    upper gastrointestinal bleeding | 0\
    hemoglobin dropped to 9.7 g/dL | 48\
    hiatus hernia | 0\
    Hill's classification grade 4 | 0\
    7-mm sessile polyp | 0\
    Paris classification 0-Is | 0\
    polyp removed by snaring | 0\
    extensive gray to black speckles on gastric corpus | 0\
    duodenal pseudomelanosis | 0\
    gastric pseudomelanosis | 0\
    intact lining epithelium | 0\
    preserved architecture | 0\
    brownish-black pigment-laden macrophages | 0\
    Perl's Prussian blue stain positive | 0\
    iron deposition confirmed | 0\
    pseudomelanosis diagnosis | 0\
    duodenal polyp hyperplastic | 0\
    urosepsis managed with antibiotics | 0\
    kidney injury managed conservatively | 0\
    intravenous fluids | 0\
    supportive measures | 0\
    clinical improvement | 120\
    transferred to wards | 120\
    renal function back to baseline | 288\
    septic markers improved | 288\
    discharged home | 288\
    full recovery | 288\
    melena | 0\
    drop in hemoglobin | 48\
    esophagogastroduodenoscopy | 0\
    pseudomelanosis incidental finding | 0\
    no relation to upper gastrointestinal bleeding | 0\
    no long-term sequelae | 0\
    clinically insignificant | 0\
    charcoal ingestion | 0\
    ferrous sulfide | 0\
    hemosiderin | 0\
    lipofuscin | 0\
    pseudomelanin deposition | 0\
    calcium deposition | 0\
    magnesium deposition | 0\
    differential diagnosis excluded | 0\
    malignant melanoma excluded | 0\
    brown bowel syndrome excluded | 0\
    hemosiderosis excluded | 0\
    hemochromatosis excluded | 0\
    Masson-Fontana stain not done | 0\
    ethical approval obtained | 0\
    no conflict of interest | 0\
    no funding received | 0\
    case report drafted | 0\
    literature review | 0\
    critical revision | 0\
    editing | 0\
    final approval | 0\
    data available | 0\
    histopathology images provided | 0\
    figures included | 0\
    table included | 0\
    informed consent obtained | 0\
    IRB approval | 0\
    references cited | 0\
    authors acknowledged | 0\
    figures descriptions provided | 0\
    differential diagnosis table | 0\
    differential diagnosis characteristics | 0\
    organs involved | 0\
    histopathology findings | 0\
    metastatic melanoma | 0\
    gastric siderosis | 0\
    brown bowel syndrome | 0\
    melanosis coli | 0\
    chronic constipation | 0\
    laxatives use | 0\
    dark mucosal staining | 0\
    malignant melanoma | 0\
    hemosiderosis | 0\
    hemochromatosis | 0\
    iron supplementation | 0\
    vitamin E deficiency | 0\
    malabsorption syndromes | 0\
    celiac disease | 0\
    Crohn's disease | 0\
    post-gastric bypass | 0\
    alcohol abuse | 0\
    lipofuscin-like pigment deposits | 0\
    smooth muscle cells | 0\
    muscularis mucosa | 0\
    muscularis propria | 0\
    cytological atypia | 0\
    increased nuclear cytoplasmic ratio | 0\
    enlarged hyperchromic nuclei | 0\
    prominent nucleoli | 0\
    frequent mitoses | 0\
    immunohistochemical stains | 0\
    Melan-A | 0\
    S100 | 0\
    HMB45 | 0\
    SOX-10 | 0\
    yellow-brown hemosiderin | 0\
    stains positive for iron | 0\
    alcohol-related liver disease | 0\
    repeated blood transfusion | 0\
    primary skin melanoma | 0\
    multiple flat or polypoid lesions | 0\
    GI tract involvement | 0\
    dark-blackish discoloration | 0\
    primary condition identified | 0\
    detailed history taken | 0\
    vitamin E deficiency | 0\
    alcohol abuse | 0\
    chronic constipation | 0\
    long-term laxatives use | 0\
    melanosis coli | 0\
    benign condition | 0\
    histopathological examination | 0\
    confirmation of diagnosis | 0\
    exclusion of metastatic melanoma | 0\
    incidental finding | 0\
    critically ill | 0\
    upper gastrointestinal bleeding | 0\
    melena | 0\
    hemoglobin drop | 48\
    sepsis managed | 0\
    culture-guided antibiotics | 0\
    conservative management | 0\
    intravenous fluids | 0\
    supportive measures | 0\
    clinical improvement | 120\
    transfer to wards | 120\
    renal function recovery | 288\
    septic markers improvement | 288\
    discharge after 12 days | 288\
    full recovery | 288\
    pseudomelanosis linked to chronic kidney disease | 0\
    diabetes mellitus | 0\
    hypertension | 0\
    ferrous sulphate | 0\
    hydralazine | 0\
    furosemide | 0\
    β-blockers | 0\
    rare endoscopic finding | 0\
    speckled dark pigmentations | 0\
    lamina propria macrophages | 0\
    iron deposition | 0\
    Prussian blue stain | 0\
    hyperplastic polyp | 0\
    snaring removal | 0\
    sessile polyp | 0\
    Paris classification | 0\
    Hill's classification | 0\
    hiatus hernia | 0\
    gastric corpus | 0\
    duodenum | 0\
    gastric mucosa | 0\
    preserved architecture | 0\
    brownish-black pigment | 0\
    macrophages | 0\
    Perl's stain | 0\
    positive iron | 0\
    pseudomelanosis confirmed | 0\
    differential diagnosis | 0\
    excluded malignancies | 0\
    benign nature confirmed | 0\
    no specific etiology | 0\
    contributing factors | 0\
    medications | 0\
    comorbidities | 0\
    incidental findings | 0\
    no long-term effects | 0\
    clinically insignificant | 0\
    histopathology confirmation | 0\
    exclusion of melanoma | 0\
    iron supplements | 0\
    propranolol | 0\
    hydrochlorothiazide | 0\
    hemochromatosis | 0\
    gastrointestinal bleeding | 0\
    chronic kidney disease | 0\
    diabetes mellitus | 0\
    hypertension | 0\
    medications list | 0\
    ferrous sulphate | 0\
    hydralazine | 0\
    furosemide | 0\
    β-blockers | 0\
    chronic conditions | 0\
    dementia follow-up | 0\
    acute presentation | 0\
    dehydration | 0\
    hypotension | 0\
    tachypnea | 0\
    heart rate | 0\
    Glasgow coma scale | 0\
    laboratory abnormalities | 0\
    leukocytosis | 0\
    hemoglobin | 0\
    CRP | 0\
    urea | 0\
    AKI | 0\
    CKD | 0\
    lactate | 0\
    procalcitonin | 0\
    urine analysis | 0\
    UTI | 0\
    ICU admission | 0\
    sepsis diagnosis | 0\
    UTI source | 0\
    AKI on CKD | 0\
    upper GI bleeding | 0\
    hemoglobin drop day 2 | 48\
    EGD findings | 0\
    histology results | 0\
    iron deposition confirmed | 0\
    management steps | 0\
    antibiotics | 0\
    fluids | 0\
    supportive care | 0\
    transfer to wards day 5 | 120\
    renal recovery | 288\
    sepsis resolution | 288\
    discharge day 12 | 288\
    recovery achieved | 288\
    pseudomelanosis characteristics | 0\
    endoscopic features | 0\
    pigment deposition | 0\
    iron in macrophages | 0\
    other minerals | 0\
    differential diagnoses | 0\
    exclusion process | 0\
    ethical considerations | 0\
    consent obtained | 0\
    IRB approval | 0\
    no conflicts | 0\
    funding sources | 0\
    author contributions | 0\
    data availability | 0\
    acknowledgments | 0\
    figures included | 0\
    table included | 0\
    references cited | 0\
    case report details | 0\
    patient demographics | 0\
    clinical course | 0\
    management outcomes | 0\
    pseudomelanosis discussion | 0\
    differential diagnosis table | 0\
    histopathology images | 0\
    stain results | 0\
    endoscopic images | 0\
    polyp removal | 0\
    sepsis management | 0\
    kidney injury management | 0\
    discharge outcome | 0\
    full recovery confirmed | 288\
    pseudomelanosis incidental | 0\
    no relation to GI bleeding | 0\
    benign nature | 0\
    histopathology needed | 0\
    melanoma excluded | 0\
    iron confirmed | 0\
    Prussian blue positive | 0\
    hemosiderin excluded | 0\
    lipofuscin excluded | 0\
    pseudomelanin excluded | 0\
    mineral deposits | 0\
    calcium | 0\
    magnesium | 0\
    differentials excluded | 0\
    melanoma features | 0\
    siderosis features | 0\
    brown bowel features | 0\
    hemosiderosis features | 0\
    hemochromatosis features | 0\
    Masson-Fontana not used | 0\
    immunohistochemical markers | 0\
    melanoma stains | 0\
    siderosis stains | 0\
    brown bowel features | 0\
    clinical insignificance | 0\
    no sequelae | 0\
    incidental finding | 0\
    critical illness | 0\
    upper GI bleed | 0\
    melena present | 0\
    hemoglobin drop | 48\
    EGD performed | 0\
    pseudomelanosis found | 0\
    management successful | 0\
    recovery achieved | 288\
    patient demographics | 0\
    comorbidities listed | 0\
    medications listed | 0\
    acute symptoms | 0\
    examination findings | 0\
    lab results | 0\
    diagnosis made | 0\
    ICU admission | 0\
    treatment given | 0\
    procedures done | 0\
    histopathology results | 0\
    management steps | 0\
    outcome described | 0\
    discussion points | 0\
    ethics statement | 0\
    conflicts statement | 0\
    funding statement | 0\
    author contributions | 0\
    data statement | 0\
    acknowledgments | 0\
    figures and tables | 0\
    references | 0\
    patient age | 0\
    patient sex | 0\
    presenting symptoms | 0\
    examination signs | 0\
    lab tests | 0\
    imaging | 0\
    endoscopic findings | 0\
    histology | 0\
    stains used | 0\
    diagnosis confirmation | 0\
    treatment administered | 0\
    response to treatment | 0\
    discharge status | 0\
    follow-up | 0\
    case rarity | 0\
    literature review | 0\
    differentials discussed | 0\
    management approach | 0\
    patient outcome | 0\
    ethical compliance | 0\
    author roles | 0\
    data sharing | 0\
    acknowledgments made | 0\
    figures description | 0\
    table description | 0\
    references cited | 0\
    patient history | 0\
    chronic conditions | 0\
    acute conditions | 0\
    diagnostic process | 0\
    therapeutic interventions | 0\
    clinical course | 0\
    recovery timeline | 0\
    pseudomelanosis features | 0\
    histopathological confirmation | 0\
    differential exclusion | 0\
    management details | 0\
    outcome details | 0\
    ethics details | 0\
    conflict details | 0\
    funding details | 0\
    author details | 0\
    data details | 0\
    acknowledgment details | 0\
    figure details | 0\
    table details | 0\
    reference details | 0\
    pseudomelanosis duodeni | 0\
    gastric pseudomelanosis | 0\
    duodenal pseudomelanosis | 0\
    endoscopic findings | 0\
    histology findings | 0\
    iron deposition | 0\
    pigment-laden macrophages | 0\
    Prussian blue positivity | 0\
    hyperplastic polyp | 0\
    sessile polyp | 0\
    snare removal | 0\
    Hill's classification | 0\
    Paris classification | 0\
    hiatus hernia | 0\
    gastric corpus | 0\
    duodenum | 0\
    ICU stay | 0\
    ward transfer | 0\
    discharge day 12 | 288\
    full recovery | 288\
    pseudomelanosis incidental | 0\
    upper GI bleeding | 0\
    melena | 0\
    hemoglobin drop | 48\
    sepsis management | 0\
    antibiotics | 0\
    fluids | 0\
    supportive care | 0\
    renal recovery | 288\
    septic recovery | 288\
    discharge home | 288\
    pseudomelanosis factors | 0\
    chronic kidney disease | 0\
    diabetes mellitus | 0\
    hypertension | 0\
    medications | 0\
    ferrous sulphate | 0\
    hydralazine | 0\
    furosemide | 0\
    β-blockers | 0\
    rare condition | 0\
    benign nature | 0\
    histopathology needed | 0\
    melanoma excluded | 0\
    iron confirmed | 0\
    management successful | 0\
    patient recovered | 288\
    case reported | 0\
    ethics obtained | 0\
    no conflicts | 0\
    no funding | 0\
    authors involved | 0\
    data available | 0\
    pathologist acknowledged | 0\
    figures provided | 0\
    table included | 0\
    references cited | 0\
    pseudomelanosis duodeni | 0\
    gastric pseudomelanosis | 0\
    endoscopic appearance | 0\
    histology confirmation | 0\
    management approach | 0\
    patient outcome | 0\
    ethical compliance | 0\
    author contributions | 0\
    data sharing | 0\
    acknowledgments | 0\
    figures and tables | 0\
    references | 0