83 years old | 0  
    male | 0  
    osteoarthritis | -624  
    right knee osteoarthritis | -624  
    magnetic resonance imaging | 0  
    lesions in medial femoral condyle cartilage | 0  
    lesions in weight-bearing region | 0  
    TKA operation | 0  
    left primary TKA | -1800  
    severe pain | 0  
    warfarin use | 0  
    paroxysmal atrial fibrillation | 0  
    smoking history | 0  
    cholecystectomy | -17520  
    normal femoral pulses | 0  
    normal popliteal pulses | 0  
    normal ankle pulses | 0  
    ABI right 1.06 | 0  
    ABI left 1.04 | 0  
    echocardiography | 0  
    warfarin hold | -72  
    INR 1.72 | 0  
    enoxaparin sodium administration | 0  
    spinal anesthesia | 0  
    tourniquet inflated to 300 mmHg | 0  
    anterior parapatellar approach | 0  
    blood loss 350 mL | 0  
    tourniquet time 96 minutes | 0  
    compressive dressing applied | 0  
    transfer to recovery room | 0  
    warm lower limb | 0  
    intact dorsalis pedis artery pulsation | 0  
    mental state decline | 0  
    drowsiness | 0  
    decreased respiration | 0  
    blood pressure 80/40 mmHg | 0  
    transfer to ICU | 0  
    CT brain | 0  
    CT lungs | 0  
    supportive therapy | 0  
    vital signs recovery | 24  
    unstable mental status | 24  
    delirium | 24  
    trembling | 24  
    attempted to get out of bed | 24  
    sedative administration | 24  
    restraint band use | 24  
    drain tube removal | 48  
    Hemovac drain 60 mL | 48  
    compressive dressing removal | 48  
    pulse not checked | 48  
    temperature not checked | 48  
    Cnoxane administration | 48  
    warfarin administration | 48  
    INR 1.83 | 48  
    air pressure device use | 48  
    warfarin dosage same | 72  
    necrosis of foot | 60  
    no dorsalis pedis artery pulsation | 60  
    no capillary filling | 60  
    CT angiography | 60  
    femoral artery occlusion | 60  
    cardiovascular consultation | 60  
    angiography | 60  
    embolic occlusion | 60  
    Fogarty thrombectomy | 60  
    unsatisfactory reperfusion | 60  
    no back bleeding | 60  
    open thrombectomy | 60  
    flow maintenance | 60  
    sepsis suspicion | 96  
    rhabdomyolysis suspicion | 96  
    drowsiness | 96  
    blood pressure 70/50 mmHg | 96  
    rapid necrosis deterioration | 96  
    above-knee amputation | 408  
    discharge | 408  
    wheelchair use | 408  
    monitoring for 6 months | 408  

