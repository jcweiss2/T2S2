29 years old | 0
male | 0
admitted to the hospital | 0
muscle pain | -144
joint pain | -144
general weakness | -144
fever | -144
liver dysfunction | -144
total bilirubin 5.7 mg/dl | -144
serum glutamic oxaloacetic transaminase 633 U/L | -144
serum glutamic pyruvate transaminase 412 U/L | -144
gamma-glutamyl transferase 161 U/L | -144
lactate dehydrogenase 1668 U/L | -144
C-reactive protein 519 mg/l | -144
procalcitonin 1.28 ng/ml | -144
increased leukocyte levels | -144
acute respiratory failure | 0
altered state of consciousness | 0
continuous sedation | 0
muscle relaxation | 0
intubation | 0
mechanical ventilation | 0
FiO2 100% | 0
SpO2 88.7% | 0
hemodynamic instability | 0
norepinephrine 0.6 μg/kg/min | 0
vasopressin not available | 0
broad-spectrum empirical antimicrobial therapy | 0
meropenem | 0
azithromycin | 0
oseltamivir | 0
methylprednisolone | 0
stress ulcer prophylaxis | 0
thromboprophylaxis | 0
drug doses adjusted for renal function | 0
prone position | 0
chest CT | 0
massive bilateral pneumonia | 0
minimal pleural effusions | 0
bedside focus ultrasound | 0
acute renal failure | -144
CRRT | -144
CytoSorb adsorber | -168
combined therapy | -168
norepinephrine requirements lowered | -168
norepinephrine discontinued | -144
inflammatory marker levels reduced | -168
CRP decreased | -168
leukocyte levels normalized | -168
ventilation parameters improved | -168
lung function improved | -168
ICU delirium | 0
antipsychotics | 0
percutaneous tracheostomy | 0
hemodynamic status stable | 0
recovery gradual | 0
weaned off ventilator | 0
transferred to general ward | 1152
transferred to rehabilitation clinic | 1152
influenza A (H1N1) | -144
bilateral pneumonia | -144
sepsis | -144
septic shock | -144
cytokine storm | -144
COVID-19 | -144
CRRT and CytoSorb application | -168
patient recovery | 1152
hemodynamic stabilization | -168
inflammation markers decreased | -168
ventilation parameters improved | -168
lung function improved | -168
vasopressors discontinued | -144