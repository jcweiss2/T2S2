57 years old|0
    male|0
    obese|0
    body mass index 39|0
    resident of province with domestic animals|0
    transferred to clinic|0
    treated with bed rest for 2 weeks for spine fracture|-336
    misdiagnosis|-336
    claims dyspnea|0
    severe back pain of 2-month duration|0
    left knee pain|0
    left knee swelling|0
    recent asymptomatic consumption of domestic poultry|-1344
    no pathologic neurological findings|0
    left osteoarthritic knee swollen|0
    chest roentgenogram shows pleural effusion on left side|0
    lateral plain roentgenogram reveals destruction of T12 vertebral body and intervertebral discs T11-T12 and T12-L1|0
    computed tomography scan reveals paravertebral abscess formation|0
    white blood cells 17.5 k/μl|0
    C-reactive protein 23.1 mg/dL|0
    ESR 86 mm/1st h|0
    tuberculosis antibody test normal|0
    virological tests normal|0
    rheumatologic tests normal|0
    Widal-Wright normal|0
    urine cultures normal|0
    stool cultures normal|0
    blood cultures reveal Salmonella enteritis|0
    thoracic drainage tube inserted|0
    seropurulent fluid evacuated|0
    gradual improvement of respiratory function|0
    knee puncture evacuates purulent fluid|0
    percutaneous transpedicular biopsy taken from T12 vertebra|0
    specimen culture taken|0
    cultures isolate Salmonella enteritis|0
    phage typing not available|0
    T12 biopsy discloses chronic osteomyelitis|0
    quinolone given intravenously|0
    3rd generation cephalosporin given intravenously|0
    left thoracotomy with resection of 11th rib|0
    left lung stuck to parietal pleura|0
    residual empyema|0
    meticulous mobilization|0
    purulent material evacuated from paravertebral space|0
    T12 vertebrectomy performed|0
    disc resection|0
    bone debridement to healthy tissue|0
    titanium mesh cage inserted|0
    resected rib bone graft inserted|0
    minimally invasive posterior instrumentation|0
    neurologically intact|0
    severe back pain|0
    obesity|0
    breathing constrained disturbances|0
    pleural effusion|0
    chest tube|0
    breathing unable to cope with needs|0
    paravertebral abscess formation|0
    instability|0
    breathing difficulty|0
    surgery decision|0
    knee fused with Illizarov device 1 month following admission|720
    post-operative course complicated with superficial wound infection|720
    thoracotomy skin infection|720
    knee arthrodesis incision infection|720
    left L2 screw insertion infection|720
    Acinetobacter infection|720
    local debridement|720
    secondary closure|720
    left knee fused completely 3 months following surgery|2160
    antibiotic susceptibility pattern basis for treatment|0
    quinolone given intravenously|0
    ceftriaxone given intravenously|0
    3 months IV antibiotic treatment|0
    discharged with monthly inflammatory marker checks|0
    6-month follow-up CRP normal|4320
    6-month follow-up ESR normal|4320
    radiograms show good fusion|4320
    CT scan shows good fusion|4320
    patient free of pain|4320
    returned to daily routine|4320
    no sign of recurrence|4320
    2 months later became anxious|6240
    family found with altered state of consciousness|6240
    admission to hospital|6240
    lost consciousness|6240
    intubated|6240
    transferred to intensive care unit|6240
    brain CT scan reveals edema|6240
    hydrocephalus|6240
    drainage tube installation|6240
    lumbar puncture cerebrospinal fluid indicative of viral infection|6240
    EEG shows slow waves|6240
    blood cultures reveal Salmonella enteritis|6240
    patient did not recover from meningoencephalitis|6240
    relatives decided to disconnect ventilator|6240
    clinically dead|6240
    SE infection recurrence causes immunosuppression|6240
    central nervous system viral infection|6240

    