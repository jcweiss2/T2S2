65 years old | 0
female | 0
admitted to the hospital | 0
diabetes mellitus | -10080
glimepiride | -10080
vildagliptin | -10080
metformin | -10080
voglibose | -10080
fatigue | -336
appetite loss | -336
cough | -336
dyspnea | -336
elevated white blood cell count | -672
elevated C-reactive protein | -672
no fever | -672
no pain | -672
pitting edema | 0
elevated WBC | 0
elevated CRP | 0
pleural effusion | 0
air in the left pleural cavity | 0
collapse of the left lung | 0
mediastinal shift to the right | 0
tension pyopneumothorax | 0
loss of respiratory variability | 0
elevated lactate level | 0
intensive care unit | 0
thoracostomy tube | 0
drainage | 0
foul odor | 0
yellow viscous pus | 0
Actinomyces sp. | 0
anaerobic bacteria | 0
intravenous sulbactam | 72
intravenous ampicillin | 72
thoracic cavity wash | 72
urokinase | 72
analgesics | 0
no fever | 0
chest CT | 216
pulmonary or bronchopleural fistula | 216
thoracostomy tube removal | 408
antibiotics discontinuation | 432
discharged | 504
recovered from pyopneumothorax | 504
chest CT | 6048
full expansion of the left lung | 6048
slight fibrosis in the lung | 6048