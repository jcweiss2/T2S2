37 years old | 0
    woman | 0
    congenital diagnosis of transposition of the great arteries | 0
    ventricular septal defect | 0
    pulmonary stenosis | 0
    surgical correction during infancy with atrial switch procedure (Mustard operation) | 0
    ventricular septal defect closure | 0
    implant of a valved conduit between the left ventricle and the pulmonary artery | 0
    not under specialized ACHD care | 0
    developed high-grade atrioventricular block | 0
    permanent transvenous PMK implant | 0
    PMK implant performed at local hospital | 0
    drug-resistant pneumonia | -24
    treated with i.v. antibiotics | -24
    full remission | -24
    discharged home | -24
    recurrence of fever spikes | -24
    hospitalization due to recurrent fever spikes | -24
    significantly raised inflammatory markers | -24
    referred to ACHD centre | 0
    admission | 0
    critical conditions due to septic shock | 0
    severe acute respiratory failure | 0
    mechanical ventilation | 0
    transferred to intensive care unit | 0
    stabilization of vital parameters | 0
    transthoracic echocardiography | 0
    transoesophageal echocardiography | 0
    three-dimensional acquisitions | 0
    multiple mobile vegetations in subpulmonary left ventricle | 0
    vegetations attached to PMK lead | 0
    vegetations attached to mitral valve leaflets | 0
    mobile mass in right ventricular outflow tract | 0
    intraventricular abscess in systemic right ventricle | 0
    systemic embolization | 0
    pulmonary septic embolization | 0
    necrosis of the extremities | 0
    total-body CT | 0
    pleural-based peripheral thickenings with triangular morphology | 0
    hypodense ischemic areas in spleen | 0
    hypodense ischemic areas in both kidneys | 0
    cerebral CT | 0
    large haemorrhage involving left fronto-parieto$occipital region | 0
    intraventricular extension into lateral ventricles | 0
    effacement of cortical sulci | 0
    midline shift of 11 mm | 0
    blood cultures positive for MRSA | 0
    diagnosis of infective endocarditis (IE) | 0
    started on antibiotic therapy with daptomycin | 0
    cardiac surgery not deemed feasible | 0
    percutaneous extraction of infected PMK leads | 0
    temporary device implant | 0
    urgent surgical haematoma evacuation | 0
    severe refractory multiorgan failure | 0
    death | 24