48 years old | 0
male | 0
admitted to the hospital | 0
history of hypertension | -672
history of dyslipidemia | -672
sudden onset of chest pain | 0
electrocardiogram revealed ST-segment elevation | 0
ST-segment elevation on leads I, aVL, and V1–V6 | 0
ST-segment depression on leads II, III, and aVF | 0
echocardiography demonstrated severely impaired motion of the anterolateral wall of the left ventricle | 0
white blood cell count of 19100/μL | 0
lactase dehydrogenase level of 213 IU/L | 0
creatinine kinase level of 77 mg/dL | 0
C-reactive protein level of 0.6 mg/dL | 0
D-dimer level of 1.85 μg/mL | 0
AMI on the anterolateral wall of the left ventricle | 0
emergent coronary angiography | 1
severe narrowing of the LMT | 1
PCI with IVUS guidance | 2
intimal flap extending from the aortic wall of the ascending aorta to the ostium of the LMT | 2
pooling of blood in the false channel of the localized aortic dissection | 2
sudden collapse with sustained ventricular tachycardia | 3
resuscitated with tracheal intubation | 3
recovered with normal sinus rhythm | 3
placement of 4.0 mm × 23 mm and 4.0 mm × 28 mm drug-eluting stents | 4
severe hypotension | 4
veno-arterial extracorporeal membrane oxygenation (VA-ECMO) | 5
transferred to the operating room for emergency surgery | 6
exposure of the ascending aorta through a median sternotomy | 7
localized hematoma on the posterior wall of the ascending aorta | 7
trans-esophageal echocardiography showed localized dissection of the posterior wall of the aorta | 7
cardiopulmonary bypass (CPB) with tepid hypothermia | 8
aortic cross clamping with antegrade and retrograde cardioplegia | 9
distal side coronary artery bypass grafting to the LAD and the circumflex branch | 10
additional cardioplegic solution given selectively from the SVGs | 11
dissecting part of the ascending aorta transversely opened | 12
entry found at a 15-mm distal site above the LMT orifice | 12
LMT dissection (Neri’s classification type B) | 12
localized dissection repaired by obliterating the false lumina | 13
proximal side coronary artery bypass grafting | 14
unsuccessful weaning from CPB | 15
support of VA-ECMO and intra-aortic balloon pumping (IABP) | 15
transferred to the intensive care unit | 16
maximum creatine kinase level of 7712 U/L | 20
postoperative contrast-enhanced computed tomography showed successful repair | 24
cardiac dysfunction persisted 5 days after the operation | 120
transferred to a highly specialized hospital for implantation of a left ventricular assist device | 120
died of severe sepsis | 3360