6-day-old | 0
male | 0
3,000-g | 0
born by Cesarean section | -144
38+4 weeks of gestation | -144
Down syndrome | -672
pulmonary atresia with ventricular septal defect (PA-VSD) | -672
icteric | -144
cyanotic | -144
SpO2 of 78% on room air | -144
continuous intravenous prostaglandin | -144
10 μg/kg/min | -144
meconium normally | -144
normal complete blood count | -144
unconjugated hyperbilirubinemia | -144
mildly elevated C-reactive protein of 10.0 mg/L | -144
normal renal function test | -144
mild electrolyte disturbance | -144
abdominal distention | -120
refused to feed | -120
fever of 38.5°C | -120
no tachypnea | -120
oxygen saturation at 60–70% on 3 L of oxygen | -120
lung clear to auscultation | -120
abdomen distended without obvious tenderness or erythema | -120
hypoactive bowel sounds | -120
abdominal X-ray | -120
ultrasound | -120
no pneumoperitoneum or free fluid | -120
no intestinal pneumatosis or portal venous gas | -120
normal leukocyte count of 4,210/µL | -120
diagnosis of NEC, Bell stage IA | -120
empiric intravenous antibiotics with ceftriaxone, amikacin, and metronidazole | -120
nil by mouth | -120
nasogastric tube inserted with intermittent suction | -120
abdominal distention increased | -96
generalized tenderness and erythema of the abdomen | -96
no blood on per rectal examination | -96
repeat abdominal ultrasound | -96
pneumoperitoneum and moderate ascites | -96
bowel loops distended up to 28 mm | -96
no portal venous gas or pneumatosis intestinalis | -96
leukocytosis of 11,780/µL with 68.1% neutrophils | -96
C-reactive protein markedly elevated at 224.3 mg/L | -96
diagnosis of peritonitis due to perforated hollow viscus | -96
exploratory laparotomy | -96
midline incision | -96
entire bowel loops distended | -96
peritoneal cavity filled with turbid and yellowish fluid | -96
fibrinous exudate distributed mainly at the right iliac fossa around the cecum | -96
appendix inflamed and perforated at its middle portion | -96
Vicryl 2.0 suture to secure the base | -96
appendix transected by scalpel | -96
peritoneal cavity irrigated with warm normal saline | -96
peritoneal fluid sent for culture | -96
peritoneal drainage placed at the Douglas pouch | -96
abdomen closed by interrupted suture | -96
pathologic analysis of the appendix | -96
grossly inflamed appendix measuring 4 mm in diameter and 2.5 cm in length | -96
microscopic analysis showed marked infiltration of inflammatory cells | -96
appendiceal mucosa completely necrotic | -96
empiric broad-spectrum antibiotic therapy with meropenem and amikacin | 0
died on postoperative day 5 | 120
worsening sepsis | 120
decompensated hemodynamic instability | 120