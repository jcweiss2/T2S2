36-week gestation | 0
    female | 0
    caucasian | 0
    newborn | 0
    delivered | 0
    26-year-old mother | 0
    primigravida | 0
    spontaneous vaginal delivery | 0
    pregnancy uneventful | 0
    parents not related | 0
    parents healthy | 0
    no family history of gastrointestinal disease | 0
    amniotic fluid stained with thick meconium | 0
    resuscitation | 0
    tracheal suctioning | 0
    positive pressure ventilation | 0
    birth weight 2800 g | 0
    Apgar score 4 at 1 min | 0
    Apgar score 6 at 5 min | 0
    Apgar score 7 at 10 min | 0
    transferred to neonatal intensive care unit | 0
    nasal continuous positive airway pressure | 0
    physical examination unremarkable | 0
    marked pallor | 0
    normocytic normochromic anemia | 0
    hemoglobin 10.6 g/dL | 0
    hematocrit 31.9% | 0
    C-reactive protein normal | 0
    kidney function tests normal | 0
    serum electrolyte levels normal | 0
    no signs of hemolysis | 0
    no fetomaternal hemorrhage | 0
    histopathological examination of placenta revealed chorioamnionitis | 0
    received intravenous antibiotics | 0
    received blood transfusion | 0
    stable after first few hours | 24
    no respiratory distress | 24
    spontaneous breathing | 24
    oral feeding started with breast and formula feeding | 48
    irritable | 72
    lethargic | 72
    severe dehydration | 72
    lost 25% body weight | 72
    adequate urine output | 72
    hyperchloremic metabolic acidosis | 72
    pH 7.18 | 72
    HCO3 12.3 mmol/L | 72
    base excess –14.9 mmol/L | 72
    Cl- 129 mmol/L | 72
    hypernatremic dehydration | 72
    Na+ 155 mmol/L | 72
    glucose levels normal | 72
    lactate levels normal | 72
    sepsis workup negative | 72
    loose watery bloodless stools with mucus | 72
    kept nil per os | 72
    volume expansion with normal saline | 72
    fluid replacement therapy | 72
    sodium bicarbonate replacement therapy | 72
    total parenteral nutrition initiated | 72
    central venous line | 72
    dependent on TPN | 72
    attempts to deliver oral feeding resulted in weight loss | 72
    hyponatremia | 72
    metabolic acidosis | 72
    urinary catheterization performed | 72
    diarrhea profuse | 72
    diarrhea misinterpreted as urine | 72
    diarrhea persisted despite fasting | 72
    stool output up to 120 ml/kg/day | 72
    intravenous fluids replacement | 72
    high sodium requirements up to 10 mmol/kg/day | 72
    stool reducing substance negative | 72
    fecal pH 8 | 72
    stool Na+ concentration 83 mmol/L | 72
    fecal ion gap <50 | 72
    secretory diarrhea pattern confirmed | 72
    initiated octreotide | 456
    no improvement | 456
    developed cholestasis | 456
    catheter-related sepsis | 456
    exhaustive etiological investigation performed | 456
    repeated blood cultures | 456
    repeated stool cultures | 456
    repeated urine cultures | 456
    culture for cytomegalovirus | 456
    metabolic screen | 456
    immunoreactive trypsinogen levels | 456
    renal testing | 456
    hepatic testing | 456
    endocrinological testing | 456
    specific serum cow milk IgE levels | 456
    testing for immunodeficiency | 456
    testing for autoimmune enteropathy | 456
    cerebral ultrasound | 456
    abdominal ultrasound | 456
    cardiac ultrasound | 456
    renal ultrasound | 456
    all test results normal | 456
    congenital enterocyte defect suspected | 456
    MVID suspected | 456
    endoscopy with duodenal biopsy planned | 288
    endoscopy performed on day 12 | 288
    duodenal biopsy performed on day 12 | 288
    duodenal sections revealed unspecific inflammatory enteropathy | 288
    further biopsy performed at three months | 2160
    biopsy showed microvillus atrophy | 2160
    no PAS staining abnormalities | 2160
    EM examination showed no significant changes | 2160
    DNA sequencing revealed MYO5B mutations | 2160
    compound heterozygous mutations of MYO5B gene | 2160
    diagnosis of MVID confirmed | 2160
    parents heterozygous carriers | 2160
    genetic counseling offered | 2160
    discharged home at three months | 2160
    TPN dependence | 2160
    liver function deterioration by five months | 3600
    died at nine months | 6480
    septic shock secondary to catheter-related infection | 6480
