54 years old | 0
male | 0
admitted to the hospital | 0
pre-syncope | 0
syncope | 0
left-sided chest tightness | 0
generalized fatigue | -672
weight loss | -672
diffuse erythematous rash | 0
blood pressure 96/60 mm Hg | 0
unremarkable cardiac examination | 0
unremarkable respiratory examination | 0
normal sinus rhythm | 0
raised troponin concentration | 0
eosinophil count 7.6 × 10^9/l | 0
referred to cardiology | 0
myocarditis | 0
cardiac magnetic resonance imaging | 24
eosinophilic myocarditis | 24
coronary angiography | 24
no coronary artery disease | 24
skin biopsy | 24
cardiac biopsy | 24
edoxaban 30 mg once daily | 48
prednisolone 40 mg once daily | 48
discharged | 48
missed appointment | 1344
presented to cardiology clinic | 1344
neck swelling | 1344
urgently admitted to hospital | 1344
eosinophil count 19.7 × 10^9 cells/l | 1344
increased prednisolone to 100 mg once daily | 1344
computed tomography of neck | 1344
lymphadenopathy | 1344
T-cell lymphoma | 1344
cyclophosphamide therapy | 1344
sepsis | 1368
cholecystitis | 1368
new onset seizures | 1368
reduction in consciousness | 1368
Glasgow Coma Scale 9/15 | 1368
head CT | 1368
multiple bilateral acute infarctions | 1368
transferred to intensive care unit | 1368
hepatitis B | -10000
asthma | -10000
intravenous drug use | -10000
excessive use of alcohol | -10000
diffuse subendocardial late gadolinium enhancement | 1440
mild LV systolic impairment | 1440
eczematous changes | 1440
bone marrow biopsy | 1440
no increase in eosinophils | 1440
axillary lymph node biopsy | 1440
T-cell lymphoma | 1440
infarcts involving frontal, parietal, and left temporo-occipital regions | 1440
apical tear | 1440
intramural myocardial tear | 1440
small apical cavity | 1440
mobile structures attached to dissected myocardium | 1440
diastolic flow in apical cavity | 1440
systolic flow out of apical cavity | 1440
cyclophosphamide therapy | 1440
partial response | 1440
reduction of eosinophil count | 1440
palliation | 1500 
deterioration | 1500 
poor prognosis | 1500