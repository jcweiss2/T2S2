44 years old| 0
    male | 0
    admitted to the hospital | 0
    shortness of breath | -48
    nonproductive cough | -48
    fever | 0
    tachycardia | 0
    hypotension | 0
    hypoxemia | 0
    obesity | 0
    type 2 diabetes | 0
    bilateral hazy opacities | 0
    positive SARS-CoV-2 PCR | 0
    metabolic acidosis (pH 7.09) | 0
    hyperlactatemia (12 mmol/l) | 0
    acute respiratory distress syndrome (ARDS) | 0
    leukocytosis (27.8×10³/μl) | 0
    elevated creatinine (1.88 mg/dl) | 0
    elevated high-sensitivity troponin-T (46 ng/l) | 0
    elevated N-terminal pro-BNP (14,535 pg/ml) | 0
    elevated ferritin (3,495 ng/l) | 0
    elevated D-dimer (>20 μg/ml) | 0
    prolonged prothrombin time (17.0 s) | 0
    left ventricular ejection fraction 45% | 0
    right ventricular dilation | 0
    right ventricular dysfunction | 0
    clot in transit (right ventricle) | 0
    intubation | 0
    admitted to ICU | 0
    hypotension requiring vasopressors | 0
    intravenous methylprednisolone (1 mg/kg/day) | 0
    tissue plasminogen activator (tPA) administration | 0
    unfractionated heparin anticoagulation | 0
    dobutamine infusion | 0
    consideration for ECMO | 0
    resolution of clot in transit | 24
    improved right ventricular function | 24
    negative lower extremity venous Doppler | 24
    oropharyngeal bleeding | 120
    continued systemic anticoagulation | 120
    planned oral anticoagulation post-discharge | 0
    hospitalization ongoing | 0
  