53 years old | 0
Caucasian | 0
male | 0
admitted to the hospital | 0
acute New York Heart Association Class IV dyspnoea | -336
reduced exercise tolerance | -336
intermittent chest pain | -336
multiple hospital attendances in the preceding 8 weeks | -1344
recurrent viral pericarditis | -1344
recent viral illness | -1344
non-steroidal anti-inflammatories | -1344
colchicine | -1344
4 weeks of prednisolone | -1344
asthma | 0
allergic rhinitis | 0
hypertension | 0
hypercholesterolaemia | 0
obesity | 0
treated obstructive sleep apnoea | 0
no history of recent surgery | 0
no history of recent travel | 0
no history of ill contacts | 0
no active dental infection | 0
afebrile | 0
normoxic | 0
normotensive | 0
tachycardic | 0
heart rate 112 beats/min | 0
tachypnoeic | 0
respiratory rate 24 | 0
soft dual heart sounds | 0
decreased breath sounds at bilateral lung bases | 0
no pulsus paradoxus | 0
jugular venous pressure not elevated | 0
multiple previous dental fillings | 0
adequate dental health | 0
no over gingival inflammation | 0
no dental abscesses | 0
no dental decay | 0
sinus tachycardia | 0
no diffuse ECG changes | 0
no electrical alternans | 0
normal white cell count | 0
elevated C-reactive protein | 0
unremarkable chest X-ray | 0
unremarkable NTproBNP | 0
unremarkable autoimmune screens | 0
mild left ventricular dysfunction | 0
large asymmetric pericardial effusion | 0
organized echogenic material adjacent to the right ventricle | 0
diastolic collapse | 0
significant tricuspid and mitral inflow variation | 0
dilated and fixed inferior vena cava | 0
urgent pericardiocentesis | 0
150 mL blood-stained fluid drained | 0
symptom relief | 0
pericardial fluid lactate dehydrogenase 3584 U/L | 0
fluid/serum lactate dehydrogenase ratio 12 | 0
pericardial fluid cholesterol 1.7 mmol/L | 0
pigtail catheter placed | 0
catheter removed | 48
clinical improvement | 48
minimal output | 48
total 240 mL drained | 48
improved inflammatory markers | 48
purulent debris in the catheter | 48
small residual effusion | 48
akinetic and adherent right ventricular free wall | 48
ventricular interdependence | 48
minimally collapsing dilated inferior vena cava | 48
gram-positive bacillus in pericardial fluid culture | 48
intravenous vancomycin commenced | 48
intermittent nocturnal fevers | -720
intermittent nocturnal sweats | -720
attributed to viral upper respiratory tract infection | -720
mild dyspnoea | 72
no chest pain | 72
no fevers | 72
no chills | 72
no rigors | 72
negative septic screening | 72
improved inflammatory markers | 72
unchanged echodense space adjacent to right ventricle | 72
persistent ventricular interdependence | 72
worsening mitral inflow variation | 72
cardiac magnetic resonance imaging | 72
pericardial effusion adjacent to the right ventricle | 72
marked thickening and fibrosis of the pericardium | 72
constrictive effusive pericarditis | 72
increasing pericardial effusion | 120
septal shift | 120
adhered right ventricular free wall | 120
fixed and dilated inferior vena cava | 120
Actinomyces meyeri identified | 120
antibiotics changed to benzylpenicillin | 120
referral to Cardiothoracic Surgery | 120
clinically stable | 168
down-trending C-reactive protein | 168
multidisciplinary meeting | 168
surgical timing discussed | 168
planned 72-hour monitoring | 168
long-term peripheral cannula established | 168
outpatient surgical management planned | 168
worsening exertional dyspnoea | 240
oxygen saturation 93-94% | 240
up-trending C-reactive protein | 240
inpatient surgical intervention planned | 240
surgical pericardiectomy | 312
washout of pericardial collection | 312
transferred to ICU | 312
extubated | 336
no growth on surgical culture aspirate | 312
no bacteria seen on microscopy | 312
organizing fibrous and fibrinous pericarditis | 312
thickened pericardium | 312
reactive stromal cells | 312
reactive endothelial cells | 312
no malignancy | 312
negative acid-fast bacilli culture | 312
negative acid-fast bacilli microscopy | 312
negative blood cultures | 312
negative urine cultures | 312
negative sputum cultures | 312
transferred to Cardiothoracic Surgery ward | 360
clinically stable | 360
down-trending C-reactive protein | 360
febrile episodes | 384
temperature 38.2°C | 384
stable C-reactive protein | 384
reviewed by Infectious Diseases | 384
no septic source | 384
no drug fever | 384
no antibiotic changes | 384
negative blood cultures | 384
negative urine culture | 384
negative chest drain tip culture | 384
repeat transthoracic echocardiogram | 384
small pericardial space | 384
no effusions | 384
no vegetations | 384
normal right ventricle size | 384
preserved left ventricular function | 384
no further febrile episodes | 432
improved C-reactive protein | 432
discharged | 432
plan for intravenous antibiotics | 432
plan for oral antibiotics | 432
no chest discomfort | 432
no dyspnoea | 432
low mood | 432
care from primary care physician | 432
completed 6 weeks of intravenous benzylpenicillin | 432
de-escalation to oral antibiotics | 432
ongoing oral amoxicillin | 432
no recurrent episodes | 432
satisfied with physical recovery | 432
