65 years old | 0
male | 0
admitted to the hospital | 0
4-day history of gradually increasing shortness of breath | -96
fever | -96
dry cough | -96
fatigue | -96
reduced breath sounds in lower lung segments | 0
oxygen saturation (SpO2) 93% | 0
bilateral peripheral ground-glass attenuation | 0
patchy consolidation | 0
lung involvement 60%-70% | 0
SARS-CoV-2 RT-PCR positive | 0
symptoms worsened | 0
increased temperature remained | 0
oxygen saturation decreased to 90% | 0
white cell count 7.93 х 109/L | 0
hemoglobin 159 g/l | 0
platelet count 468 х 109/l | 0
Westergren ESR 41 mm/h | 0
interleukine 6 102 pg/ml | 0
С-reactive protein 142 mg/l | 0
ferritin 939.92 μg/ml | 0
D-dimer 609 ng/ml | 0
procalcitonin 0.11 ng/ml | 0
dexamethasone | 0
heparin | 0
tocilizumab | 0
acetylcysteine | 0
pantoprazole | 0
nadroparin calcium | 0
oxygen supplementation 4 l/min | 0
chest radiography on Day 15 | 360
air in right pleural cavity | 360
pleural effusion in right pleural cavity | 360
collapse of right lung | 360
transferred to ICU | 360
thoracentesis | 360
thoracostomy | 360
evacuated 1400 ml yellowish opaque liquid | 360
follow-up chest radiograph showed lack of air | 360
persistence of fluid remains | 360
lung expansion | 360
linezolid therapy initiated | 360
imipenem/cilastatin therapy initiated | 360
oxygen supplementation increased to 8-10 l/min | 360
daily drainage volume 300-1000 ml | 360
chest CT on day 3 after thoracentesis | 432
pleural effusion with gas bubbles | 432
right lung reduced in volume by half | 432
focal area of subpleural infiltration with central cavity | 432
air layer up to 47 mm anterior chest wall | 432
left side hydropneumothorax | 432
pleural effusion 25 mm anteroposterior depth | 432
air layer 19 mm anterior chest wall | 432
multiple bilateral ground glass infiltrates | 432
exudative lymphocytic-rich effusion | 432
no growth of acid-fast bacteria | 432
gram-negative bacteria Acinetobacter baumannii | 432
gram-negative bacteria Pseudomonas aeruginosa | 432
urine culture positive for Klebsiella pneumoniae | 432
needle thoracocentesis | 432
new pleural drainage established | 432
aspirated air and creamy purulent mass | 432
serofibrinous hemorrhagic fluid drawn daily | 432
chest CT showed air and pleural effusion | 432
pleural empyema confirmed | 504
transferred to Surgical Department | 504
right pleural space irrigated with antiseptic | 504
lung expansion by vacuum aspiration | 504
encapsulated pleural effusion identified | 720
ultrasound-guided puncture | 720
new drainage installed | 720
antibiotic therapy with colistimethatum natrium | 0
antibiotic therapy with imipenem/cilastatin | 0
discharged from hospital | 672
oxygen saturation (SpO2) 97% | 672
small amount of fluid in right pleural cavity | 672
lab tests normal | 672
С-reactive protein 11.7 mg/l | 672
procalcitonin <0.1 ng/ml | 672
plasma D dimer 2424 ng/ml | 504
