69 years old | 0
male | 0
referred to department of family medicine | 0
chronic weakness | -87600
recurrent admissions | -87600
untreated and undiagnosed longstanding pancytopenia | -87600
pancytopenia persisted for 10 years | -87600
severe splenomegaly | -87600
treated for fungal pneumonia | -87600
aspergilloma | -87600
Pneumocystis jirovecii pneumonia | -87600
past medical history of right thyroidectomy | -87600
thyroid cancer | -87600
posterior right coronary artery stenting | -87600
chronic stable angina pectoris | -87600
paroxysmal atrial fibrillation | -87600
repeated admissions | -87600
current admission for exacerbation of fungal pneumonia | 0
initial evaluation | 0
afebrile | 0
body temperature 36.5°C | 0
blood pressure 99/66 mm Hg | 0
heart rate 77 beats per minute | 0
respiratory rate 20 per minute | 0
poor nutritional status | 0
weight 48.7 kg | 0
height 169 cm | 0
BMI 17.05 kg/m² | 0
cachectic | 0
exhausted by prolonged admission | 0
initial laboratory studies | 0
pancytopenia | 0
neutropenia | 0
absolute neutrophil count 150/μL | 0
hyponatremia 131 mmol/L | 0
increased prothrombin time 12.9 seconds | 0
increased partial thromboplastin time 41.1 seconds | 0
elevated C-reactive protein 40.3 mg/L | 0
elevated erythrocyte sedimentation rate 59 mm/h | 0
no evidence of cytomegalovirus infection | 0
negative blood culture | 0
negative sputum culture | 0
urine culture with Gram-positive cocci 1,000 CFU/mL | 0
chest X-ray multiple nodular consolidations | 0
chest CT scan multiple nodular consolidations | 0
small left pleural effusion | 0
pericardial effusion | 0
no enlarged lymph nodes | 0
enlarged spleen 21.4 cm | 0
initial medications: aspirin | 0
nicorandil | 0
trimetazidine | 0
bisoprolol | 0
levothyroxine | 0
total parenteral nutrition initiated | 0
antibiotic therapy commenced with trimethoprim/sulfamethoxazole | 0
meropenem | 0
amphotericin B | 0
chest CT scan minimal possibility of active Pneumocystis pneumonia | 0
negative PCR for Pneumocystis jirovecii | 0
amphotericin B as sole antifungal agent | 0
prophylactic antibacterial agents reduced to cefepime | 0
fever subsided | 0
consultations from hematology | 0
rheumatology | 0
infection | 0
differential diagnosis focused on splenomegaly | 0
peripheral blood smear normochromic, normocytic anemia | 0
reticulocyte percentage 0.65% | 0
iron deficiency anemia screening | 0
anemia of chronic disease | 0
elevated ferritin 3,308.5 ng/mL | 0
low transferrin 98 mg/dL | 0
normal serum iron 79 μg/dL | 0
no deficiency of B12 | 0
no deficiency of folate | 0
bone marrow biopsy average cellularity 60% | 0
no signs of bone marrow failure | 0
prior bone marrow biopsies failed to indicate diagnosis | -87600
primary hematologic disease unlikely | 0
investigations for autoimmune causes | 0
positive ANA titer 320:1 | 0
rheumatoid factor 23 IU/mL | 0
weakly-positive anti-DNA 19 IU/mL | 0
weakly-positive anti-cardiolipin IgM 11 MPL-U/mL | 0
negative anti-beta2-glycoprotein 1 antibodies | 0
negative lupus anticoagulant | 0
low serum C3 36.7 mg/dL | 0
normal C4 11.98 mg/dL | 0
oral ulcer found | 0
no skin rash | 0
no arthritis | 0
no muscular weakness | 0
no uveitis | 0
no Reynaud phenomenon | 0
elevated cystatin C 1.53 mg/L | 0
cystatin C-based eGFR 42.6 mL/min/1.73 m² | 0
normal creatinine 0.82 mg/dL | 0
ongoing infection | 0
renal failure deemed indeterminate | 0
follow-up anti-DNA antibodies 10 IU/mL | 408
elevation of rheumatologic antibodies considered by-product of infection | 408
splenomegaly suspected cause of pancytopenia | 0
pancytopenia progressively worsened | 264
day 11 hospitalization | 264
WBC 540/μL | 264
neutrophil 35.9% | 264
hemoglobin 6.8 g/dL | 264
platelet count 57×10³/μL | 264
suspected sepsis | 264
body temperature 37.0°C | 264
blood pressure 86/52 mm Hg | 264
pulse rate 84 | 264
infusion of 1.5 L fluid | 264
blood pressure not raised | 264
filtered red blood cells transfused | 264
norepinephrine 4 mL/h | 264
indeterminate diagnosis | 264
deteriorating general condition | 264
splenectomy considered | 264
surgical splenectomy deemed hazardous | 264
partial splenic embolization considered | 264
consultations sought | 264
failure to establish definite diagnosis | 264
partial splenic embolization undertaken on day 17 | 408
iodixanol contrast agent | 408
ultrasound guidance for arterial access | 408
right common femoral artery access | 408
celiac angiography | 408
splenic angiography | 408
70% spleen embolized with gelfoam | 408
day after embolization | 432
no serious complications | 432
increased WBC 820/μL | 432
hemoglobin 10.0 g/dL | 432
platelet count 45×10³/μL | 432
2 days after procedure | 456
temperature rose to 38.5°C | 456
temperature drop to 35.7°C | 456
blood pressure 84/56 mm Hg | 456
pulse rate 148 | 456
septic shock suspected | 456
norepinephrine infused | 456
fluids infused | 456
chest CT scan | 456
abdominal CT scan | 456
no pulmonary embolism | 456
no bowel perforation | 456
increased rales in lungs | 456
oxygen saturation 55% | 456
mechanical ventilation initiated | 456
refusal of ICU admission | 456
cardiac arrest | 456
CPR commenced | 456
spontaneous circulation not established | 456
death | 456
