27 years old | 0
female | 0
Mayer Rokitansky Syndrome | -0
Mullerian agenesis | -0
sigmoid neovaginoplasty | -7560
lower abdominal pain | 0
bilateral pelvic pain | 0
denies routinely irrigating or dilating her neovagina | 0
penetrative sexual intercourse | -0
life stressors | -0
no intercourse in a few months | -0
CT imaging of the abdomen | 0
tubular, heterogenous, fluid-filled structure | 0
blind ending | 0
outpatient referral to the gynecologist | 0
abdominal pain acutely worsened | 24
diaphoresis | 24
significant distress due to pain | 24
leukocytosis | 24
absolute neutrophils | 24
repeat abdominal CT | 24
increasing inflammatory process | 24
empiric intravenous piperacillin-tazobactam | 24
transferred emergently to hospital | 24
hypotensive | 24
tachycardic | 24
afebrile | 24
tachypneic | 24
oxygen saturation | 24
IV fluid boluses | 24
antimicrobials changed to IV ceftriaxone, IV vancomycin, and IV metronidazole | 24
exploratory laparotomy | 24
cystoscopy | 24
vaginoscopy | 24
normal bladder | 24
normal urethra | 24
obliterated introitus | 24
diffuse intra-abdominal spillage of the mucus | 24
perforated sigmoid neovagina | 24
purulent fluid drained | 24
intrabdominal drains placed | 24
intubated | 24
mechanical ventilation | 24
septic shock | 24
vasopressor agents | 24
antimicrobials transitioned to IV cefepime, IV vancomycin, and IV metronidazole | 24
peritoneal culture growing gram-negative rods | 24
blood cultures remained negative | 24
peritoneal cultures finalized to Bacterioides thetaioaomicron, Bacteroides caccae, and Actinomyces species | 168
antimicrobials changed to IV piperacillin-tazobactam | 168
weaned off vasopressors | 192
extubated | 192
transferred to the general floor | 288
Infectious Diseases team consulted | 288
discharged home | 360
abdominal wound vacuum | 360
IV piperacillin-tazobactam for four weeks | 360
readmitted with sepsis | 504
generalized malaise | 504
diffuse abdominal pain | 504
white blood count | 504
absolute neutrophil count | 504
d-dimer | 504
lactate | 504
CT of the chest, abdomen and pelvis | 504
bilateral pleural effusions | 504
loculated left pleural effusion | 504
multiple new abdominal abscesses | 504
transcutaneous drainage catheter in pelvis | 504
open anterior midline wound with wound vacuum | 504
hypoxemia | 504
transferred to the intensive care unit | 504
IV piperacillin-tazobactam continued | 504
placement of a right perihepatic drain | 504
aspiration of purulence | 504
unsuccessful drainage of peri-splenic collection | 504
blood cultures remained negative | 504
interventional radiology reconsulted | 504
drained 350 mL of pus from the right perinephric abscess | 504
drained 90 mL of pus from her perisplenic abscess | 504
broad-spectrum PCR sent on the drained fluid | 504
improved clinically | 768
antimicrobials narrowed to IV ampicillin-sulbactam | 768
discharged | 768
broad spectrum PCR from the fluid positive for Gleimia europaea, Alistipes onderdonkil, Varibaculum timonense, and Jonquetella anthropi | 768
followed up at the adult infectious diseases clinic | 1056
continued on ampicillin-sulbactam | 1056
plans to reimage | 1056
improved clinically | 1056
repeat CT abdomen demonstrated decreased in the size of right and left sub-phrenic abscesses | 1056
transitioned from IV ampicillin-sulbactam to oral amoxicillin-clavulanate | 1056
complete resolution of the abscesses | 1056