30-year-old man | 0
admitted to the emergency room | 0
mechanical ileus | 0
enterocutaneous fistula | 0
abdominal pain | 0
difficulty in defecation | 0
sudden changes in mental status | 0
stupor after vomiting | 0
sepsis | 0
blood pressure 60/40 mmHg | 0
heart rate 140 beats/min | 0
MELAS syndrome diagnosis | -61368
partial seizure | -61368
carbamazepine | -61368
valproic acid | -61368
mental retardation | -61368
cerebral infarction left middle cerebral artery | -61368
cerebral infarction right posterior inferior cerebellar artery | -61368
history of lactic acidosis | -61368
white blood cells 2.9 × 103 /μl | 0
lactic acid 142.1 mg/dl | 0
aspartate transaminase 141.1 U/L | 0
alanine transaminase 124.7 U/L | 0
creatine kinase 353.0 U/L | 0
CK-MB 20.79 ng/ml | 0
blood urine nitrogen 36.7 mg/dl | 0
creatinine 1.10 mg/dl | 0
prothrombin time 17.7 s | 0
international normalized ratio 1.57 | 0
activated partial thromboplastin time 56.7 s | 0
metabolic acidosis | 0
pH 7.170 | 0
PaO2 129.5 mmHg | 0
PaCO2 36.8 mmHg | 0
base excess −15.2 mM/L | 0
HCO3- 13.6 mM/L | 0
lactic acidosis | 0
lactate 131.7 mg/dl | 0
ST-elevation anterior lead | 0
Wolff–Parkinson–White syndrome | 0
high sensitivity troponin-T 205 ng/L | 0
pro B-type natriuretic peptide 313.7 pg/ml | 0
hypoglycemia 55.1 mg/dl | 0
dobutamine 10 μg/kg/min | 0
norepinephrine 0.5 μg/kg/min | 0
drowsy-to-stupor mental status | 0
emergency total colectomy | 0
terminal ileostomy | 0
anesthesia induction with propofol | 0
dexmedetomidine infusion | 0
remifentanil infusion | 0
propofol effect-site concentration increased | 0
BIS score 44 | 0
propofol discontinued | 0
rocuronium 0.6 mg/kg | 0
endotracheal intubation | 0
mechanical ventilation | 0
oxygen 60% | 0
tidal volume 600 ml | 0
respiratory rate 12 breaths/min | 0
esophageal temperature monitoring | 0
body cooling with ice bag | 0
fluid management | 0
stroke volume variation | 0
plasma solution | 0
hypotension event | 80
BP 47/18 mmHg | 80
HR 42 beats/min | 80
epinephrine 1 mg | 80
vasopressin 5U | 80
dexmedetomidine infusion stopped | 180
remifentanil target Ce adjusted to 0 | 205
BIS score 97 | 205
opened eyes upon verbal command | 205
sugammadex 200 mg | 205
TOF ratio 13% | 205
extubation | 205
TOF ratio 100% | 205
spontaneous breathing restored | 205
total propofol 50 mg | 205
total dexmedetomidine 225 μg | 205
total remifentanil 2.15 mg | 205
glucose supplement | 205
50% dextrose in water | 205
glucose 8 g/h | 205
blood glucose 101 mg/dl | 205
sodium bicarbonate 120 mEq | 205
pH 7.2 | 205
respiratory rate adjusted | 205
tidal volume adjusted | 205
end-tidal CO2 below 40 mmHg | 205
ice bag application axilla | 205
body temperature 37°C | 205
forced air warmer | 205
temperature above 36°C | 205
surgery duration 210 min | 210
transferred to intensive care unit | 210
ABGA pH 7.278 | 210
PaO2 256.0 mmHg | 210
PaCO2 33.1 mmHg | 210
base excess −11.3 mM/L | 210
HCO3) 15.6 mM/L | 210
lactate 64.1 mg/dl | 210
crystalloids 3,000 ml | 210
urine output 1,100 ml | 210
estimated blood loss 100 ml | 210
critical care for one month | 720
sepsis persisted | 720
condition worsened | 720
cardiac arrest | 720
cardiopulmonary resuscitation not performed | 720
death due to septic shock | 720
