diagnosed with mild COVID-19 illness | -36
sore throat | -36
loss of sense of smell | -36
positive COVID-19 PCR | -36
full recovery by resolution of symptoms | -14
reverting to negative PCR | -14
received the first dose of inactivated SARS-CoV-2 vaccine | 0
remained asymptomatic and well | 0
received the second dose of inactivated SARS-CoV-2 vaccine | 30
started to experience headache | 30
started to experience fatigue | 30
developed fever | 34
developed sore throat | 34
developed abdominal pain | 34
presented to the emergency department | 38
high-grade fever | 38
myalgia | 38
nausea | 38
vomiting | 38
diarrhoea | 38
faint erythematous non-itchy rash over his torso | 38
dry irritant cough | 38
no shortness of breath | 38
no chest discomfort | 38
no urinary symptoms | 38
no pain or swelling of his joints | 38
temperature of 39°C | 38
systolic blood pressure of 110 mm Hg | 38
tachycardia, 140 beats per minute | 38
dry mucous membranes with congested throat | 38
bilateral conjunctival injection | 38
left conjunctival haemorrhage | 38
generalised erythematous maculopapular rash | 38
peripheral lymph nodes were not enlarged | 38
no audible cardiac murmurs | 38
chest was clear to auscultation | 38
abdomen examination was unremarkable | 38
SARS-CoV-2 PCR from nasopharyngeal swab was negative | 38
SARS-CoV-2 IgG from serum was strongly positive | 38
throat swab was negative for group A streptococcus | 38
sputum culture showed mixed flora | 38
bacterial blood cultures were negative | 38
urinalysis showed significant proteinuria | 38
ANA, dsDNA, c-ANCA and p-ANCA titres were all negative | 38
C3 and C4 were reduced | 38
admitted to the intensive care unit | 38
treated empirically with ceftriaxone and levofloxacin | 38
given intravenous hydrocortisone | 38
given intravenous fluids for resuscitation | 38
blood pressure stabilised | 40
fever initially improved | 40
developed facial puffiness | 40
developed generalised body oedema | 40
remained tachycardic | 40
diarrhoea persisted | 40
myalgia persisted | 40
renal impairment with significant proteinuria | 42
ECG showed sinus tachycardia with non-specific T-wave abnormalities | 42
troponin-I was raised | 42
pro-BNP over 8000 pg/mL | 42
transthoracic echocardiogram showed severe tricuspid regurgitation | 42
pulmonary hypertension | 42
right atrium and ventricle were moderately dilated | 42
left ventricle cavity size was normal | 42
mildly reduced ejection fraction | 42
thin rim of pericardial effusion | 42
computed topography scan of the chest showed bilateral moderate pleural effusion | 42
computed topography scan of the chest showed basal atelectasis | 42
discontinued hydrocortisone | 44
shifted to the medical ward | 44
high-level fever began to recur | 46
diagnosed with multisystem inflammatory syndrome in adults | 48
treated with intravenous steroids, dexamethasone | 48
condition improved markedly | 50
generalised oedema subsided | 50
skin rash resolved | 50
conjunctivitis resolved | 50
white blood cell count normalised | 50
renal function improved | 50
inflammatory markers came down to normal levels | 50
repeat transthoracic echocardiography showed trace tricuspid regurgitation | 50
dexamethasone continued for 8 days | 50
switched to oral prednisolone | 58
discharged home with a tapering dose of prednisolone | 60
symptoms resolved | 74
general weakness and fatigue | 74
repeat echocardiogram was completely normal | 74