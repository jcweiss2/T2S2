31-year-old male | 0
motor vehicle accident | -864
severe head injury | -864
cervical spine fracture | -864
spine fixed with plate and screw | -864
intubated | -864
paraplegic | -864
recurrent chest infections | -1440
antibiotics | -1440
widened mediastinum | -1440
Hemoglobin 11.3 g/dL | -1440
hematocrit 35% | -1440
Mean corpuscular volume 67.7 fL | -1440
mean corpuscular hemoglobin 21.8 pg | -1440
albumin 2.7 g/L | -1440
creatinine 0.5 μmol/L | -1440
Na 135 mmol/L | -1440
erythrocyte sedimentation rate 93 mm/h | -1440
superior mediastinal collection | -1440
chronic esophageal perforation | -1440
upper esophageal perforation | -1440
cervical spine plate and screw erosion into esophagus | -1440
neck exploration | -1440
plate removed | -1440
perforation repaired with interposition muscle flap | -1440
limited thoracotomy | -1440
extensive pleural adhesions | -1440
feeding jejunostomy tube | -1440
surgical site infection at cervical wound | -24
exploration and drainage | -24
antimicrobial therapy | -24
admissions to ICU | 0
repeated episodes of sepsis | 0
bronchoscopies | 0
exchanging tracheostomy | 0
acute surgical abdomen | 0
exploration and drainage of intra-abdominal abscess collections | 0
persistent status epilepticus | 0
cardiac arrest | 0
XDR-P. aeruginosa isolated from urinary tract | 0
sepsis | 0
PA179 grown from blood cultures | 0
discharge | 0
death | 0
</|eot_id|>
