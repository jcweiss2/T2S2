45 years old | 0
female | 0
gravidity 5 | 0
parity 2 | 0
body mass index 24 kg/m2 | 0
admitted to the hospital | 0
major placenta previa | -240
antepartum hemorrhage | -240
previous uneventful spontaneous vaginal deliveries | -10000
no remarkable medical history | 0
scheduled for an elective lower segment cesarean delivery | -240
combined spinal-epidural block | 0
electrocardiogram | 0
noninvasive blood pressure | 0
oxygen saturation monitoring | 0
initial blood pressure 120/80 mm Hg | 0
heart rate 105/min | 0
peripheral oxygen saturations 96% | 0
uncomplicated CSE | 0
sensory block to T4 bilaterally | 0
Bromage score of 3 | 0
blood pressure 120/75 mm Hg | 0
phenylephrine infusion of 2 mg/h | 0
heart rate 90-120/min | 0
Spo2 96% | 0
delivery of a live infant | 0
Apgar score 9 at 1 and 5 minutes | 0
nausea | 0
dizziness | 0
bradycardia of 35/min | 0
loss of consciousness | 0
blood pressure 70/35 mm Hg | 0
atropine 600 µg IV | 0
succinylcholine 100 mg | 0
endotracheal intubation | 0
carotid pulse absent | 0
electrocardiogram demonstrating a sinus rhythm of 100/min | 0
pulseless electrical activity | 0
cardiopulmonary resuscitation | 0
epinephrine 1 mg IV | 0
chest compressions | 0
asynchronous ventilation | 0
capnography | 0
endotracheal intubation confirmed | 0
effective chest compressions | 0
lungs ventilated with 100% oxygen | 0
volume-controlled mode | 0
obstetricians delivered the placenta | 0
exteriorized the uterus | 0
monitored effectiveness of thoracic compressions | 0
return of spontaneous circulation | 9
pulseless electrical activity | 19
chest compressions | 19
TEE performed during resuscitation | 19
dilated right ventricle | 19
severely reduced systolic function | 19
left ventricle underfilled | 19
moderate globally reduced systolic function | 19
noradrenaline infusion at 40 µg/min | 30
well-defined mass in the right pulmonary artery | 30
abdominal drains | 30
prophylactic Bakri intrauterine balloon | 30
vaginal packs | 30
abdomen closed | 30
bleeding from the vagina | 40
bleeding from the oropharynx | 40
bleeding from peripheral access sites | 40
massive hemorrhage | 40
institutional massive transfusion protocol activated | 40
lactic acidosis | 40
anemia | 40
ROTEM performed | 40
fibrin formation and polymerization | 40
hypofibrinogenemia | 40
extrinsic coagulation pathway | 40
EXTEM clotting time | 40
hyperfibrinolysis | 40
fibrinogen concentrate | 60
platelets | 60
cryoprecipitate | 60
tranexamic acid | 60
volume resuscitation | 60
balanced electrolyte solution | 60
albumin | 60
calcium gluconate | 60
ROTEM showed improvement | 120
hypofibrinogenemia | 120
fibrinogen concentrate | 120
uterus contracted | 120
core temperature 35.5°C | 120
hemodynamic stability | 120
noradrenaline infusion at 17 µg/min | 120
transferred to the intensive care unit | 120
transthoracic echocardiography | 180
improved LV contractility | 180
ejection fraction 0.55-0.60 | 180
severely dilated RV | 180
impaired systolic function | 180
mild pulmonary hypertension | 180
milrinone | 180
vasopressin | 180
ROTEM results | 180
uterine bleeding | 180
anemia | 180
hysterectomy | 240
packed red blood cells | 240
coagulopathy resolved | 240
formal laboratory tests | 240
hemoglobin concentration stabilized | 240
interhospital transfer | 240
computerized tomography pulmonary angiogram | 360
saddle embolus | 360
ultrasound of the lower limbs | 360
deep venous thrombosis excluded | 360
abdominal ultrasound investigation | 360
right ovarian thrombosis | 360
discharged home | 504
transthoracic echocardiography | 504
normal LV size | 504
low normal systolic function | 504
ejection fraction 0.54 | 504
normal RV | 504
low normal systolic function | 504
anticoagulation treatment | 504
neurophysiological deficits | 504
formal neuropsychology review | 504
intact cognition | 504