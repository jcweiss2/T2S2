64 years old | 0
male | 0
hypertension | -105168
type II diabetes mellitus | -105168
alcohol consumer | -105168
left-sided hemiparesis | 0
right-sided facial deviation | 0
slurring of speech | 0
Broca's aphasia | 0
UMN type VIIth cranial nerve palsy | 0
up-going plantar reflex on the left side | 0
left upper limb power 3/5 | 0
left lower limb power 4/5 | 0
total leukocytes count 15.5 | 0
neutrophil 65% | 0
hemoglobin 14.8 g/dl | 0
platelet count 213 | 0
urea 41 mg/dl | 0
creatinine 1.2 mg/dl | 0
sodium 140 mEq/L | 0
potassium 5.1 mEq/L | 0
bilirubin total 1.1 mg/dl | 0
bilirubin direct 0.4 mg/dl | 0
alkaline phosphatase 85 U/L | 0
ALT 20 U/L | 0
AST 23 U/L | 0
prothrombin time 13.1 sec | 0
INR 1.0 | 0
HbA1C 13.9% | 0
random blood glucose 331 mg/dL | 0
NCCT head showed right temporo-parietal infarction | 0
ischemic stroke | 0
admitted to medical ward | 0
ramipril 5 mg OD | 0
amlodipine 5 mg OD | 0
metformin 500 mg OD | 0
sitagliptin 100 mg OD | 0
empaglifozin 10 mg OD | 0
insulin 10 units OD | 0
aspirin 75 mg OD | 0
statins 10 mg OD | 0
GRBS 186 mg/dL | 0
GRBS 103 mg/dL | 24
GRBS 117 mg/dL | 48
GRBS 145 mg/dL | 72
drowsy | 96
rapid breathing | 96
GCS E3V4M5 | 96
GRBS 218 mg/dL | 96
oxygen saturation 98% | 96
blood pressure 120/80 mmHg | 96
ABG pH 7.124 | 96
HCO3 4.1 | 96
PaCO2 12.7 mmHg | 96
PaO2 90 mmHg | 96
anion gap 25 | 96
lactate 1.86 | 96
urine acetone positive | 96
euglycemic DKA | 96
alcoholic cause ruled out | 96
nasogastric tube feeding | 96
bicarbonate level low | 96
starvation ketosis ruled out | 96
renal function test normal | 96
lactic acid level lower | 96
no salicylates | 96
no antidepressants | 96
empaglifozin therapy | 96
NaHCO3 50 mEq IV | 96
ABG pH 7.214 | 96
HCO3 5.1 | 96
PaCO2 13 mmHg | 96
PaO2 116 mmHg | 96
lactate 1.71 | 96
shifted to HCU | 96
normal saline infusion 100 ml/hour | 96
NaHCO3 50 mEq TID | 96
piperacillin/tazobactam 4.5 gm TDS | 96
insulin infusion 2 units/hour | 96
empaglifozin stopped | 96
shifted to ICU | 96
ABG bicarbonate 13.4 mEq/L | 120
anion gap normal | 120
GCS poor | 168
tachypneic | 168
intubated | 168
mechanically ventilated | 168
sepsis | 168
qSOFA score 2 | 168
blood pressure 110/80 mmHg | 168
respiratory rate 28 | 168
GCS 11/15 | 168
levofloxacin 750 mg OD | 168
vancomycin 15 mg/kg/dose Q8H | 168
linezolid 600 mg Q12H | 168
colistin 300 mg LD | 168
colistin 150 mg BID | 168
spontaneous CPAP | 312
shifted to HCU | 312
insulin glargine 10 units OD | 312
insulin aspart 4 units TDS | 312
stable vital parameters | 312
bedside mobilization | 312
chest physiotherapy | 312
limb physiotherapy | 312
discharged | 432
