46 years old | 0
male | 0
obesity | 0
body mass index 42 kg/m2 | 0
admitted to the hospital | 0
right lower extremity weakness | -24
nausea | -24
generalized weakness | -24
SARS-CoV-2 infection | -1440
mild flu-like symptoms | -1440
diagnosed with SARS-CoV-2 infection | -1440
positive total antibodies | -1440
nasopharyngeal polymerase chain reaction (PCR) for SARS-CoV-2 | -1440
hypotensive | 0
hypoxic | 0
oxygen saturation 89 % | 0
bilateral rhonchi | 0
right lower extremity strength 3/5 | 0
no skin rashes | 0
negative nasopharyngeal PCR | 0
positive total antibody test for SARS-CoV-2 | 0
SARS-CoV-2 total antibodies 238 signal/cut-off (s/co) ratio | 0
IgG 11 s/co ratio | 0
inflammatory markers elevated | 0
ferritin 962 ng/mL | 0
IL-6 121.09 pg/mL | 0
C-reactive protein (CRP) 2.9 mg/dL | 0
lactate dehydrogenase (LDH) 802 units/L | 0
procalcitonin 0.678 ng/mL | 0
acute kidney injury | 0
elevated creatinine 4.10 mg/dL | 0
high anion gap metabolic acidosis | 0
lactic acidosis | 0
left retrocardiac opacity | 0
non-ST elevation myocardial infarction (NSTEMI) | 0
elevated troponin 0.282 ng/mL | 0
brain natriuretic peptide (BNP) 3590 pg/mL | 0
grossly normal ejection fraction | 0
borderline elevated right ventricular systolic pressure (RVSP) | 0
dependent ground glass opacities | 0
hepatic steatosis | 0
right ataxia | 0
mild right hemiparesis | 0
left hemianesthesia | 0
hypoxia | 0
oxygen support with 6 L of nasal cannula | 0
diffuse bilateral mixed interstitial and airspace opacities | 24
tachypneic | 24
worsening hypoxemia | 24
high-flow nasal cannula | 24
transferred to the Intensive Care Unit (ICU) | 24
invasive mechanical ventilation | 24
norepinephrine | 24
ceftriaxone 2 gm daily | 24
azithromycin 500 mg daily | 24
dexamethasone 6 mg daily | 24
unfractionated heparin | 24
negative nasopharyngeal SARS-CoV-2 PCR | 24
negative SARS-CoV-2 PCR from bronchoalveolar lavage (BAL) sample | 72
tocilizumab 8 mg/kg | 72
steroids | 72
elevated troponins | 72
elevated BNP | 72
RVSP 39.4 mmHg | 72
normal left ventricle | 72
normal left ventricular wall thickness | 72
normal left ventricular wall motion | 72
normal right ventricle | 72
continuous veno-venous hemodialysis (CVVH) | 96
no documented clinical improvement | 96
inflammatory markers continued to uptrend | 96
ferritin 1993 ng/mL | 96
IL-6 1412.44 pg/mL | 96
LDH 4773 units/L | 96
d-dimer 0.62 mcg/mL | 96
CRP 8.3 mg/dL | 96
liver and kidney function continued to worsen | 96
troponins were persistently elevated | 96
multiorgan failure | 96
clinical improvement | 144
less ventilator support | 144
no longer needing pressors | 144
hypotensive | 192
febrile | 192
thick foul-smelling respiratory secretions | 192
respiratory cultures only grew Candida albicans | 192
empiric broad spectrum antibiotics | 192
vancomycin | 192
cefepime | 192
norepinephrine restarted | 192
ferritin >100,000 ng/mL | 192
LDH > 12,000 units/L | 192
SARS-CoV-2 RT PCR (plasma) repeated | 192
below limit of detection | 192
whole genome sequencing of Spike (S) gene from BAL | 192
no SARS-CoV-2 RNA detected | 192
hydrocortisone 50 mg q6h | 216
severe refractory acidosis | 216
hyperkalemia | 216
arrhythmia | 240
death | 240