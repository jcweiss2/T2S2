78 years old | 0
male | 0
admitted to the hospital | 0
benign prostatic hyperplasia | 0
coronary artery disease | 0
atrial fibrillation | 0
leukocytosis | 0
worsening renal function | 0
hyperkalemia | 0
Pseudomonas aeruginosa urinary tract infection | 0
hemodynamic instability | 0
septic shock | 0
cefepime | 0
vasopressor support | 0
fever | -168
pustular rash | -168
erythematous base | -168
upper extremities | -168
trunk | -168
mucosal involvement | 0
neutrophilia | -168
elevated C-reactive protein | -168
chest X-ray | -168
bilateral interstitial opacities | -24
consolidation | -24
COVID-19 | -168
SARS-CoV-2 RNA nasopharyngeal swab | -168
real-time reverse transcription polymerase chain reaction | -168
skin biopsy | -24
papillary dermal edema | -24
subcorneal/intracorneal pustules | -24
mixed inflammatory infiltrate | -24
lymphocytes | -24
neutrophils | -24
eosinophils | -24
EuroSCAR study group criteria | -24
definite diagnosis of AGEP | -24
discontinuation of cefepime | 24
topical emollients | 24
resolution of exanthem | 48
post-pustular desquamation | 48
discharged | 168