36 years old | 0
female | 0
admitted to the hospital | 0
dyspnea | 0
severe vomiting | -48
poor oral intake | -48
bronchial asthma | -252 months
near-fatal asthma | -252 months
asthma medication | -252 months
increased asthma attack frequency | -168
rescue medication | -168
agitated | 0
tachypnea | 0
inspiratory and expiratory wheezing | 0
Kussmaul breathing | 0
mixed respiratory alkalosis | 0
metabolic acidosis | 0
no hypoxia | 0
supplemental oxygen | 0
high-dose short-acting beta-agonist | 0
ipratropium | 0
intravenous steroids | 0
intubated | 2
pressure-control ventilation | 2
hydration with 0.9% saline | 2
fetal viability monitored | 2
cardiotocography | 2
elevated C-reactive protein | 2
leucocyte count | 2
normal renal function | 2
normal liver function | 2
normal creatinine kinase | 2
random capillary blood glucose | 2
normal glycosylated hemoglobin | 2
urinalysis | 2
acetone | 2
no glycosuria | 2
no proteinuria | 2
admitted to ICU | 8
adjusted ventilator settings | 8
inhaled short-acting beta-agonist | 8
inhaled corticosteroid | 8
intravenous magnesium sulfate | 8
breathless | 8
deep and labored breathing | 8
dynamic hyperinflation | 8
intrinsic end-expiratory pressure | 8
sedated with propofol | 8
subcutaneous emphysema | 10
suspected pneumomediastum | 10
rapid decrease in bicarbonate levels | 10
increased anion gap | 10
lactic acidosis | 10
sepsis work-up | 10
no evidence of infection | 10
serum ketone levels | 29
pH | 29
bicarbonate levels | 29
diagnosed with starvation ketoacidosis | 29
emergency caesarean section | 29
betamethasone | 27
delivered a 2.3-kg girl | 29
umbilical cord arterial pH | 29
5-min Apgar score | 29
intensive care for 2 days | 31
grade II respiratory distress syndrome | 31
successfully extubated | 49
rapid resolution of metabolic derangement | 49
superficial gastritis | 49
discharged | 72
note: some events have been condensed or rephrased for clarity and brevity.