74 years old | 0
    male | 0
    admitted to the emergency department | 0
    lower abdominal pain | -96
    signs of infection | -96
    deterioration in overall well-being | -96
    uncontrolled diabetes mellitus | 0
    metformin | 0
    right femur fracture | -175200
    sequela of stroke | 0
    motor aphasia | 0
    facial paralysis | 0
    urethral stenosis | 0
    recurrent urinary tract infections | 0
    most recent urinary tract infection episode | -1296
    intravenous antibiotics (previous) | -1296
    dysuria | 0
    fever | 0
    pneumaturia | 0
    lower abdominal tenderness | 0
    hyperglycemia (3.18 g/L) | 0
    elevated C-reactive protein (143 mg/L) | 0
    elevated lactate (4.07 mmol/L) | 0
    normal renal function | 0
    normal hepatic function | 0
    urine dipstick positive for leukocytes | 0
    urine dipstick positive for nitrites |: 0
    abdominal and pelvic CT | 0
    diffuse thickening of the bladder wall | 0
    multiple circumferentially arranged air bubbles in bladder wall | 0
    urinary analysis white blood cells (3500/mm³) | 0
    urinary analysis red blood cells (28000/mm³) | 0
    emphysematous cystitis diagnosis | 0
    ceftriaxone | 0
    metronidazole | 0
    gentamicin | 0
    urinary catheter insertion | 0
    drainage of 500 ml cloudy urine with gas | 0
    urine culture positive bacteriological growth | 0
    transfer to intensive care unit | 0
    close clinical monitoring | 0
    biochemical monitoring | 0
    surveillance for complications | 0
    intravenous antibiotics (current) | 0
    insulin therapy | 0
    improvement in overall condition | 288
    discharged | 480
    <|eot_id|>
    74 years old|0
    male|0
    admitted to the emergency department|0
    lower abdominal pain|-96
    signs of infection|-96
    deterioration in overall well-being|-96
    uncontrolled diabetes mellitus|0
    metformin|0
    right femur fracture|-175200
    sequela of stroke|0
    motor aphasia|0
    facial paralysis|0
    urethral stenosis|0
    recurrent urinary tract infections|0
    most recent urinary tract infection episode|-1296
    intravenous antibiotics (previous)|-1296
    dysuria|0
    fever|0
    pneumaturia|0
    lower abdominal tenderness|0
    hyperglycemia (3.18 g/L)|0
    elevated C-reactive protein (143 mg/L)|0
    elevated lactate (4.07 mmol/L)|0
    normal renal function|0
    normal hepatic function|0
    urine dipstick positive for leukocytes|0
    urine dipstick positive for nitrites|0
    abdominal and pelvic CT|0
    diffuse thickening of the bladder wall|0
    multiple circumferentially arranged air bubbles in bladder wall|0
    urinary analysis white blood cells (3500/mm³)|0
    urinary analysis red blood cells (28000/mm³)|0
    emphysematous cystitis diagnosis|0
    ceftriaxone|0
    metronidazole|0
    gentamicin|0
    urinary catheter insertion|0
    drainage of 500 ml cloudy urine with gas|0
    urine culture positive bacteriological growth|0
    transfer to intensive care unit|0
    close clinical monitoring|0
    biochemical monitoring|0
    surveillance for complications|0
    intravenous antibiotics (current)|0
    insulin therapy|0
    improvement in overall condition|288
    discharged|480