history of SLE | -8760
history of stage IV lupus nephritis | -8760
history of prior stroke | -8760
history of intravenous drug use | -8760
history of three prior mitral valve replacements | -168
cardiogenic shock | 0
mental status changes | 0
elevated jugular venous pressure | 0
prominent v wave | 0
body temperature 36.3°C | 0
blood pressure 95/66 mm Hg | 0
heart rate 94 beats/min | 0
hemoglobin of 10.3 g/dL | 0
white blood cell count of 18.9 × 10^9/L | 0
platelet count of 64 × 10^9/L | 0
international normalized ratio of 3.6 | 0
creatinine level of 1.7 mg/dL | 0
drug studies positive for narcotics | 0
drug studies positive for cannabis | 0
antiphospholipid serology performed | 0
antiphospholipid serology reported as normal | 0
blood cultures collected | 0
blood cultures remained negative | 0
intravenous antibiotics initiated | 0
broad-spectrum intravenous antibiotics advised | 0
serologic studies assessing for Coxiella | 0
serologic studies assessing for Legionella | 0
serologic studies assessing for Chlamydia | 0
serologic studies assessing for Bartonella | 0
serologic studies assessing for Brucella | 0
serologic studies assessing for Tropheryma whipplei | 0
serologic studies assessing for human immunodeficiency virus | 0
serologic studies assessing for hepatitis | 0
operative cultures sent for Gram staining | 0
operative cultures sent for anaerobic and aerobic cultures | 0
operative cultures sent for fungal smear and culture | 0
operative cultures sent for acid-fast smear | 0
operative cultures sent for mycobacterial culture | 0
operative cultures sent for pathologic examination | 0
operative cultures sent for 16s recombinant ribonucleic acid testing | 0
transthoracic echocardiography (TTE) showed dehisced mitral valve prosthesis | 0
transthoracic echocardiography (TTE) showed severe mitral regurgitation | 0
transesophageal echocardiography (TEE) | 0
transesophageal echocardiography (TEE) showed posterior annulus dehiscence | 0
transesophageal echocardiography (TEE) showed loculated cavity | 0
transesophageal echocardiography (TEE) showed perivalvular regurgitation | 0
patient and family counseled regarding high-risk nature of planned procedure | 0
patient decided to proceed with procedure | 0
fourth sternotomy | 12
mitral valve prosthesis dehisced along majority of posterior annulus | 12
mitral valve prosthesis sitting high in left atrium | 12
true mitral annulus displaced apically | 12
large cavity at intervalvular fibrosa with multiloculations debrided | 12
surgical pathology showed bland fibrin thrombus and fibrous tissue with mild chronic inflammation | 12
surgical pathology negative for microorganisms | 12
extensive reconstruction of fibrous skeleton of heart and atria | 12
mitral valve annulus reconstructed integrating 33-mm bioprosthesis | 12
large patch of bovine pericardium used to reconstruct left atrial dome and interatrial septal incision | 12
postbypass TEE showed well-seated mitral valve bioprosthesis | 24
postbypass TEE showed mean gradient of 3 mm Hg | 24
postbypass TEE showed no regurgitation | 24
patient required extracorporeal membrane oxygenation | 24
patient required multiple blood product transfusions | 24
TEE in intensive care unit showed layered thrombus in left atrium adjacent to mitral valve | 120
surgical clot removal | 120
thrombus reaccumulated | 120
extracorporeal membrane oxygenation support withdrawn | 120
patient died | 120
autopsy declined | 120