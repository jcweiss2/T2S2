35 years old | 0
female | 0
Caucasian | 0
admitted to the emergency department | 0
low-grade fever | 0
chills | 0
nonspecific abdominal pain | 0
nonbilious emesis | 0
no associated cough | 0
no dysuria | 0
no skin rashes | 0
history of CD | -2640
status postright hemicolectomy | -2640
adhesion-related small bowel obstruction | -720
status postadhesiolysis | -720
off disease-modifying therapy | -120
generalized anxiety disorders | 0
bipolar disorders | 0
not on any regular medications | 0
tachycardiac | 0
hypotensive | 0
febrile | 0
diffuse tenderness | 0
no focal guarding | 0
no rigidity | 0
low hemoglobin | 0
leucopenic count | 0
low platelets count | 0
elevated serum lactate | 0
raised C-reactive protein | 0
acute kidney injury | 0
elevated serum creatinine | 0
high serum calcium | 0
normal total bilirubin | 0
slightly raised alanine transaminase | 0
abnormal alkaline phosphatase | 0
negative urinalysis | 0
unremarkable Chest X-rays | 0
admitted to the intensive care unit | 0
presumed intra-abdominal sepsis | 0
treated with aggressive fluid resuscitation | 0
treated with empiric broad-spectrum antibiotics | 0
mild gallbladder wall thickening | 24
pericholecystic fluids | 24
no calcified gallstones | 24
no evidence of active Crohn’s flare-up | 24
mild cholecystitis | 48
normal appearance of biliary ducts | 48
continued to spike fevers | 48
underwent an uneventful cholecystectomy | 72
acalculous cholecystitis | 72
liver biochemistry worsened | 96
ALT up trended | 96
ALP rose | 96
total bilirubin increased | 96
predominantly direct component | 96
normal postoperative changes | 96
no collections | 96
normal biliary ducts | 96
nonreactive viral serologies | 120
negative autoimmune screening | 120
normal total IgG | 120
normal IgM | 120
normal IgA | 120
normal transferrin saturation | 120
normal ferritin | 120
normal ceruloplasmin | 120
no known hepatotoxic medication | 120
hepatology consultation | 120
liver biopsy advised | 120
marked acute hepatitis | 144
focal necrosis | 144
noncaseating granulomas | 144
giant cells | 144
no primary biliary cirrhosis | 144
no primary sclerosing cholangitis | 144
no autoimmune hepatitis | 144
infectious workup | 144
negative acid-alcohol fast bacilli | 144
negative Giemsa fungal staining | 144
negative QuantiFERON gold assay | 144
negative Coccidiosis | 144
negative Brucella | 144
negative Bartonella | 144
negative Coxiella | 144
negative urine screening for Histoplasma antigens | 144
hypercalcemia responsive to fluid therapy | 144
renal function normalized | 144
slightly below normal parathyroid hormones | 144
normal PTH-related peptide | 144
normal Vitamin D3 1,25-OH | 144
normal angiotensin-/ (ACE) levels | 144
no pulmonary sarcoidosis | 144
small nonspecific ground-glass pulmonary nodules | 144
discontinuation of antibiotics | 168
plan of re-institution | 168
interdisciplinary discussions | 168
hepatic granulomas possibly represent extraintestinal manifestation of CD | 168
hepatic granulomas possibly represent extrapulmonary sarcoidosis | 168
oral steroids instituted | 168
discharged on prednisone taper | 192
completed 8-week course of steroids | 336
clinically well | 336
normalization of ALT | 336
normalization of ALP | 336