29 years old | 0
female | 0
admitted to the hospital | 0
complex regional pain syndrome | -1096
sports-related injury | -1096
shoulder surgery | -1096
recurrent shoulder infections | -1096
Pseudomonas aeruginosa | -1096
Sphingomonas paucimobilis | -1096
Candida colliculosa | -1096
Staphylococcus aureus | -1096
left shoulder tendon release and revision | -240
development of CRPS | -240
severe pain | -240
allodynia | -240
edema | -240
muscle spasms | -240
temperature changes | -240
electromyography evaluation | -240
brachial plexus injury | -240
asthma | -720
selective IgG3 deficiency | -720
oral medical management | -240
opioids | -240
antidepressants | -240
antispasmodics | -240
left stellate ganglion blockade | -240
continuous cervical epidural infusions | -240
placement of a left C6–C7 interlaminar epidural catheter | 0
fluoroscopic guidance | 0
preprocedure labs | 0
antibiotic prophylaxis | -1
vancomycin | -1
epidural infusion | 0
0.25% bupivacaine | 0
hydromorphone | 0
clonidine | 0
oral home medications | 0
methadone | 0
diazepam | 0
baclofen | 0
amitriptyline | 0
decrease in pain | 24
improved sleep | 24
decrease in LUE spasms and edema | 24
febrile | 120
increase in temperature | 120
wean the infusion | 120
remove the epidural catheter | 120
progressive headache | 126
neck pain | 126
increase in temperature | 126
neurological examination | 126
nontender to palpation | 126
no signs of active infection | 126
blood and urine cultures | 126
chest x-ray | 126
increase in white count | 126
cephalosporin | 126
cefepime | 126
abatement of fever | 132
decrease in white count | 132
MRI of the cervical spine | 132
epidural collection | 132
compression of the left C5 and C6 nerve roots | 132
effacement of the thecal sac | 132
interstitial edema | 132
transfer to the neurosciences intensive care unit | 132
hourly neurological examination | 132
intractable nausea and vomiting | 156
left arm weakness | 156
emergent decompression and evacuation | 156
C3 to C7 cervical laminectomies | 156
C4–C5 and C5–C6 left foraminotomies | 156
intraoperative cultures | 156
P aeruginosa | 156
susceptible to cefepime | 156
vancomycin stopped | 156
cefepime continued | 156
resolution of arm weakness | 180
uneventful postoperative course | 180
discharged home | 180
intravenous cefepime | 180