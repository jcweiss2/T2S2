40 years old | 0
female | 0
admitted to the intensive burn care unit | 0
assault chemical burn | -1.5
conjugal violence | -1.5
burned surface area 35% | 0
third degree burn | 0
severe bilateral eyes and ears lesions | 0
injury due to sulfuric acid | -1.5
irrigation with water started | 0
fluid resuscitation | 0
orotracheal intubation | 0
sedated for hospital transfer | 0
arterial blood pressure 70/30 mmHg | 0
pulse 110 bpm | 0
SpO2 >90% | 0
normal lung auscultation | 0
admission electrocardiogram | 0
chest X-ray examination | 0
metabolic acidosis | 0
pH 6.92 | 0
PaCO2 42 mmHg | 0
total bicarbonate 8.6 mEq/l | 0
base deficit 23.4 mEq/l | 0
sodium 148 mEq/l | 0
potassium 4.1 mEq/l | 0
chloride 117 mEq/l | 0
calcium 6.1 mg/dl | 0
phosphorus 15.1 mg/dl | 0
lactate level 1.7 mmol/L | 0
renal function preserved | 0
serum creatinine 0.83 mg/dl | 0
no evidence for rhabdomyolysis | 0
blood coagulation tests disturbed | 0
fibrinogen 117 mg/dl | 0
activated partial thromboplastin time (APTT) 69 s | 0
International Normalized Ratio (INR) 2.23 | 0
platelets count 169 000/mm3 | 0
administration of sodium bicarbonate | 0
administration of lactate from Hartmann's solution | 0
progressive development of thoracic rigidity | 12
mechanical ventilation | 0
percutaneous tracheostomy | 720
mild inotropic support | 0
dobutamine 5 μg/kg/min | 0
echocardiography | 0
moderate alteration of the left ventricular function | 0
urine output maintained | 0
continuous venovenous hemofiltration | 168
multiple episodes of wound-related sepsis | 0
antimicrobial therapy | 0
iterative surgery | 0
excision and grafting | 0
left the intensive care unit for rehabilitation | 120 
discharged from hospital | 5040