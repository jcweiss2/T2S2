22 years old | 0
male | 0
admission to the hospital | 0
somnolent patient | 0
unclear aetiology | 0
intubation | 0
insertion of an arterial catheter | 0
insertion of a central venous line | 0
entry intensive care unit | 5
septic shock | 11
measurement of SvO2 from blood of the central venous line | 15
SvO2 100% | 15
pO2 198 mmHg | 15
control of the result from 14:15 | 15.25
SvO2 100% | 15.25
pO2 200 mmHg | 15.25
measurement of arterial blood gas values | 15.5
SaO2 98% | 15.5
pO2 90-111 mmHg | 15.5
chest X-ray | 16
central venous catheter tip appeared on the left side of the heart | 16
echocardiography | 16.75
aortic positioning of the central venous line was not evident | 16.75
electrocardiogram (ECG) | 17
venous pressure-like curve was seen | 17
computed tomography image showed placement of the catheter in the upper left pulmonary vein | 17.5
aspiration pneumonia | -72
insertion of the central venous line into the left jugular vein | 0
blood saturation was determined | 0
saturation 100% | 0
pO2 198 mmHg | 0
pCO2 46 mmHg | 0
arterial blood gas analysis | 0
saturation 98% | 0
pO2 111 mmHg | 0
pCO2 48 mmHg | 0
cervical ultrasound showed that the catheter was inserted correctly in the left jugular vein | 17.5
persistent left superior vena cava | -672
persistent foramen ovale | -672
atrial septal defect | -672
partial anomalous pulmonary venous return (PAPVR) | 17.5
discharge from the hospital | 720
follow-up | 8760
conservative treatment | 720