preterm baby | 0 | 0 | Factual
male | 0 | 0 | Factual
born by emergency cesarean section | 0 | 0 | Factual
severe preeclampsia in the mother | -672 | 0 | Factual
gestational week 25 6/7 | 0 | 0 | Factual
birthweight 665 g | 0 | 0 | Factual
intubated | 0 | 0 | Factual
mechanical ventilation | 0 | 0 | Factual
total parenteral nutrition | 24 | 0 | Factual
minimal enteral nutrition with breast milk | 24 | 0 | Factual
delayed meconium passage | 48 | 72 | Factual
abdominal distension | 48 | 72 | Factual
increased gastric residuals | 48 | 72 | Factual
necrotizing enterocolitis | 72 | 120 | Factual
gastric free drainage | 120 | 0 | Factual
broad-spectrum antibiotic therapy | 120 | 0 | Factual
perforated NEC | 144 | 144 | Factual
surgery | 144 | 144 | Factual
short bowel syndrome | 168 | 0 | Factual
thyroid screening tests | 336 | 336 | Factual
low fT4 | 336 | 336 | Factual
low TSH | 336 | 336 | Factual
cortisol 5.75 µg/dL | 336 | 336 | Factual
serum total bilirubin level 12.12 mg/dL | 336 | 336 | Factual
direct reacting bilirubin 11.48 mg/dL | 336 | 336 | Factual
enteral levothyroxine 5 µg/kg/day | 336 | 432 | Factual
no response to treatment | 432 | 432 | Factual
enteral levothyroxine 10 µg/kg/day | 432 | 504 | Factual
still no response to treatment | 504 | 504 | Factual
rectal levothyroxine 10 µg/kg/day | 504 | 0 | Factual
increasing fT4 levels | 576 | 576 | Factual
decreasing direct bilirubin levels | 576 | 576 | Factual
death | 1848 | 1848 | Factual
severe bronchopulmonary dysplasia | 1848 | 1848 | Factual
surgical NEC | 1848 | 1848 | Factual
short bowel syndrome | 1848 | 1848 | Factual
sepsis | 1848 | 1848 | Factual