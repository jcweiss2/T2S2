30 years old | 0
woman | 0
African American | 0
presented to the emergency department | 0
shortness of breath on exertion | 0
chest pain with deep inspiration | 0
no indication of recent infections | 0
physical examination did not yield any abnormalities or concerns | 0
VQ scan indicated high probability for pulmonary emboli in right lobe | 0
chest x ray showed possible small bilateral pleural effusions |EOL
chest x ray showed multiple nodular opacities scattered throughout the lungs | 0
chest x ray showed nodular opacities more prominent than before | 0
CT scan of the abdomen showed moderate alveolar consolidation in right lower lobe | 0
CT scan consistent with pulmonary infarct or pneumonia | 0
EKG normal | 0
2D echocardiograms normal | 0
no indication of endocarditis | 0
admitted for treatment of acute pulmonary embolism | 0
Heparin drip initiated | 0
developed high fevers | 0
developed tachycardia | 0
blood cultures positive (four out of four bottles) | 0
Gram positive cocci in pairs and clusters indicative of Staphylococcus species | 0
identified as S. caprae | 0
initially started on vancomycin | 0
S. aureus ruled out | 0
antibiotics changed to Kefzol 2 gm IV every 8 hours | 0
fever resolved | 0
significant clinical improvement | 0
urinalysis indicated presence of E. coli | 0
E. coli sensitive to all 17 antimicrobial agents | 0
three days of Ciprofloxacin administered | 0
echocardiogram no evidence of endocarditis | 0
unclear cause of infection | 0
no recent visit to farm | 0
no contact with goats | 0
no risk factors such as transplants, internal fixation, or foreign subject implants | 0
contracted S. caprae during hospital stay | 0
S. caprae misidentified in past | 0
identity established by Vitek 2 GP system | 0
isolate produced acid from mannitol | 0
isolate urease positive | 0
S. caprae strains with methicillin resistance | 0
slime production | 0
biofilm formation | 0
discharged | 0
