57 years old | 0
male | 0
hypertension | -2160
admitted to the hospital | 0
fever | -216
chills | -216
shortness of breath | -216
malaise | -216
poor appetite | -216
oxygen saturation 64% on room air | 0
bilateral crackles | 0
leukocyte count 8.17 K/μL | 0
procalcitonin 0.41 ng/mL | 0
nasopharyngeal swab positive for SARS-CoV-2 | 0
sputum Gram stain 10–25 WBCs/LPF | 0
sputum culture positive for methicillin susceptible Staphylococcus aureus | 0
sputum culture positive for oropharyngeal microbiota | 0
chest radiograph bilateral patchy airspace disease | 0
chest radiograph increased interstitial opacities | 0
dexamethasone 6 mg daily | 0
remdesivir | 0
oxygen support via non-rebreather mask | 0
azithromycin 500 mg daily | 0
ceftriaxone 1 g daily | 0
persistent hypoxia | 120
inability to wean from non-rebreather mask | 120
steroids continued beyond day 10 | 120
cyanotic | 168
dyspneic | 168
endotracheal intubation | 168
chest radiograph progression of infiltrates | 168
vancomycin | 168
meropenem | 168
methylprednisolone 40 mg three times per day | 168
worsening renal function | 216
continuous renal replacement therapy | 216
hypotension | 216
diarrhea | 396
Candida colitis | 396
nystatin 1 million units 6 times a day | 396
hypoxic | 432
hypotensive | 432
methylprednisolone changed to hydrocortisone 100 mg three times a day | 432
midodrine 10 mg three times a day | 432
blood cultures revealed yeast | 432
micafungin 100 mg every 24 hours | 432
antibiotics discontinued | 432
yeast identified as Cryptococcus neoformans | 456
lumbar puncture | 456
opening pressure 28 cm H2O | 456
cerebrospinal fluid 185 WBCs/μL | 456
cerebrospinal fluid 65,000 RBCs/μL | 456
positive India ink | 456
cerebrospinal fluid culture confirmed Cryptococcus neoformans | 456
cerebrospinal fluid cryptococcal antigen positive | 456
HIV 1/2/P24 combination screen negative | 456
HIV-1 Real Time PCR test negative | 456
micafungin discontinued | 456
liposomal amphotericin B 400 mg daily | 456
flucytosine 2000 mg via gastrostomy tube every other day | 456
lumbar puncture repeated | 480
new skin nodules | 480
disseminated cryptococcal infection | 480
died during hypotensive episode | 504
adrenal gland heterogeneity | 504
CT scan | 504