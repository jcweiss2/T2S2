28 years old | 0
male | 0
sickle cell trait | 0
history of intravenous drug use | 0
admitted to the hospital | 0
fever | -216
right-sided chest pain | -216
abdomen pain | -216
flank pain | -216
dysuria | -216
intermittent hematuria | -216
blood pressure 129/68 mmHg | 0
heart rate 129 beats per minute | 0
respiratory rate 19 breaths per minute | 0
temperature 39.4°C | 0
oxygen saturation 99% | 0
elevated white blood cells | 0
c-reactive protein | 0
abnormal liver function tests | 0
urine dipstick analysis 3+ urobilinogen | 0
urine dipstick analysis 3+ erythrocytes | 0
diffuse bilateral nodular densities on chest radiograph | 0
electrocardiography normal sinus rhythm | 0
referred to surgeons | 0
acute abdominal pain | 0
ultrasound possible acalculous cholecystitis | 0
ultrasound ill-defined mass near liver | 0
abdominal/pelvic computed tomography | 0
bowel perforation or infection | 0
cryptogenic organizing pneumonia | 0
admitted pending repeat CT | 0
drowsy | 2
ill-looking | 2
tachypneic | 2
profusely sweating | 2
tachycardia | 2
hypotension | 2
suspected IE | 2
pulmonary septic emboli | 2
CT with oral contrast | 2
pyelonephritis | 2
diagnosed with possible acute chest syndrome | 2
echocardiography confirmed vegetation | 4
tricuspid valve vegetation | 4
treated with intravenous vancomycin | 4
treated with cefepime | 4
antibiotics switched to flucloxacillin | 8
blood cultures confirmed methicillin-sensitive Staphylococcus aureus | 8
blood cultures confirmed viridans group streptococci | 8
urine culture no growth | 8
radiologist re-evaluated CT | 12
renal infarction | 12
multiple cortical wedge-shaped areas of delayed striated contrast enhancement | 12
condition improved | 60
discharged | 61
follow up with cardiology clinic | 61
tests for human immunodeficiency virus negative | 61
tests for hepatitis negative | 61
tests for thrombophilia negative | 61