85 years old | 0
male | 0
farmer | 0
active lifestyle | 0
admitted to the hospital | 0
transferred to rehabilitation unit | 0
past medical history of atrial fibrillation | -672
past medical history of benign prostatic hypertrophy | -672
injured leg | -1344
trismus | -1344
hypertonia | -1344
C. tetani infection | -1344
treatment with immunoglobulins | -1344
tetanus vaccination | -1344
metronidazole | -1344
transferred to ICU | -672
tracheostomy | -672
mechanical ventilation | -672
vasoactive support | -672
respiratory failure | -672
seizures | -672
treated with baclofen | -672
treated with midazolam | -672
treated with diazepam | -672
electroencephalography | -672
severely slow cerebral activity | -672
opacity on chest radiography | -672
peripheral leukocytosis | -672
possible ventilator-associated pneumonia | -672
blood cultures | -672
tracheal secretion samples | -672
Klebsiella pneumoniae | -672
methicillin-sensitive Staphylococcus aureus | -672
antibiotic therapy with piperacillin-tazobactam | -672
transferred to geriatric unit | -336
coma | -336
breathed spontaneously | -336
supplemental oxygen | -336
tracheal cannula | -336
antibiotic therapy switched to linezolid | -336
treated with meropenem | -336
septic shock | -336
gradually awoke | -168
feeding tube removed | -168
cholestasis | -168
acute edematous pancreatitis | -168
endoscopic treatment postponed | -168
urinary tract infection | -168
treated with colistin | -168
treated with amoxicillin-clavulanate | -168
multidrug-resistant organisms | -168
K. pneumoniae | -168
Acinetobacter baumannii | -168
Enterococcus faecalis | -168
clinical condition improved | 0
considered eligible for rehabilitation | 0
MDRO isolation | 0
tracheal supplemental oxygen | 0
bladder catheter | 0
pressure ulcers | 0
sarcopenic | 0
low handgrip strength | 0
appendicular skeletal mass | 0
rehabilitative evaluations | 0
rehabilitation with good compliance | 24
Clostridioides difficile infection | 24
treated with oral vancomycin | 24
atrial fibrillation | 72
third-degree atrioventricular block | 72
heart rate 30 beats/min | 72
transferred to cardiac ICU | 72
single-chamber pacemaker implantation | 72
hyperkinetic delirium | 96
Pseudomonas aeruginosa bloodstream infection | 120
treated with ceftazidime-avibactam | 120
treated with amikacin | 120
SARS-CoV-2 | 120
treated with remdesivir | 120
droplet isolation | 120
second recurrence of C. difficile | 144
treated with fidaxomicin | 144
bloodstream infection | 168
Candida parapsilosis | 168
MSSA | 168
Candida tropicalis | 168
treated with caspofungin | 168
treated with cefazolin | 168
intravenous catheter replaced | 168
bloodstream infection | 216
P. aeruginosa | 216
treated with piperacillin-tazobactam | 216
treated with aztreonam | 216
treated with ceftazidime-avibactam | 216
antibiotic resistance | 216
treated with cefepime | 240
tracheostomy closure | 240
nutritional supplementation | 240
malnutrition | 240
sarcopenia | 240
motor reconditioning | 240
respiratory reconditioning | 240
postural transition training | 240
aided transfers | 240
axial stability | 240
balance improvement exercises | 240
breath-movement coordination exercises | 240
thoracic expansion exercises | 240
girdle opening exercises | 240
inhalation-exhalation exercises | 240
wheelchairs | 240
walkers | 240
rehabilitation follow-up | 240
ENT follow-up | 240
geriatric follow-up | 240
discharged | 720