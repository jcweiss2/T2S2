72 years old | 0
male | 0
current smoker | 0
dysuria | 0
subjective fever | 0
mild confusion | 0
dizziness | 0
denied shortness of breath | 0
denied loss of consciousness | 0
foley catheter removal | -48
obstructive uropathy | -48
benign prostatic hyperplasia | -48
stage II chronic kidney disease | 0
multiple kidney stones | 0
status post lithotripsy | 0
road traffic accident 15 years ago | -131400
surgery | -131400
right hip osteoarthritis | 0
avascular necrosis | 0
status post replacement | 0
nonalcoholic | 0
denied illicit substance use | 0
mild fever | 0
tachycardia | 0
hypotension | 0
tachypnea | 0
cardiopulmonary examination unremarkable | 0
abdominal examination unremarkable | 0
bilateral edematous swelling | 0
right leg swelling | 0
arterial blood gases normal | 0
leukocyte count elevated | 0
hemoglobin 10.9 mg/dl | 0
serum bicarbonate 22 mEq/L | 0
creatinine 3.4 mg/dl | 0
blood urea nitrogen 39 mg/dl | 0
lactic acid 3.2 mg/dl | 0
urinalysis positive leukocyte esterase | 0
urinalysis high white cell count | 0
electrocardiogram normal | 0
serum troponin levels normal | 0
septic shock suspected | 0
blood cultures ordered | 0
broad spectrum intravenous antibiotics started | 0
hypotension persistent | 0
central venous catheter placed | 0
high doses intravenous norepinephrine required | 0
bedside ultrasonography performed | 0
ultrasound revealed good cardiac contractility | 0
ultrasound showed no intra-abdominal bleeding | 0
ultrasound bilateral noncompressible femoral veins | 0
deep vein thrombosis | 0
pulmonary embolism suspected | 0
echocardiogram performed | 0
ejection fraction 60% | 0
normal right ventricular ejection fraction | 0
normal right ventricular dimensions | 0
computed tomography pulmonary embolism protocol negative | 0
CT abdomen showed bilateral nonobstructive renal stones | 0
CT abdomen stranding suspicious for small retroperitoneal hematoma | 0
reevaluation of patient history with family | 0
road traffic accident complicated with DVT right leg 15 years ago | -131400
inferior vena cava filter placement 15 years ago | -131400
obstructive shock secondary to IVC obstruction suspected | 0
venography performed | 0
complete occlusion of IVC at filter level | 0
filling defects in distal IVC | 0
filling defects in bilateral common iliac veins | 0
filling defects in bilateral external iliac veins | 0
filling defects in common femoral veins | 0
thrombus present | 0
collateral arising from left common iliac vein hypertrophy | 0
mechanical thrombectomy performed | 0
