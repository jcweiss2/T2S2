75 years old | 0
male | 0
admitted to the hospital | 0
congestive heart failure | -672
non-ST elevated myocardial infarction | -672
hypertension | -672
diabetes | -672
bronchial asthma | -672
hyperuricemia | -672
intubated | 0
percutaneous coronary angioplasty | 0
refractory respiratory failure | 0
pulmonary edema | 0
pneumonia | 0
intravenous methylprednisolone | 0
oral prednisone | 0
ceftriaxone | 96
intubated three times | 0
extubated | 432
pneumomediastinum | 432
subcutaneous emphysema | 432
subdiaphragmatic free air | 432
afebrile | 432
mild tachycardia | 432
abdominal bloating | 432
abdominal pain denied | 432
crepitation all over his body | 432
abdomen distended and soft | 432
white cell count 1.21x10∧9/L | 432
blood urea nitrogen 89.6 mg/dL | 432
creatinine 4.35 mg/dL | 432
non-contrast CT | 432
extensive subcutaneous emphysema | 432
pneumomediastinum | 432
massive pneumoperitoneum | 432
pneumoretroperitoneum | 432
diffuse mesenteric emphysema | 432
acute care surgery service consulted | 432
upper gastrointestinal study | 432
no contrast leakage | 432
lower gastrointestinal contrast study refused | 432
diagnostic laparoscopy discussed | 432
exploratory laparotomy | 432
gush of air evacuated | 432
no free fluid in the peritoneum | 432
diffuse emphysema in the small and large intestinal mesenteries | 432
mild emphysema and edema from the descending colon to the sigmoid colon | 432
diverticula not observed | 432
no perforation or discoloration | 432
abdomen closed | 432
transferred to the surgical intensive care unit | 432
extubated on postoperative day 1 | 480
transferred to the ward on postoperative day 2 | 528
fever spiked | 936
left lower quadrant pain | 936
septic shock | 936
blood, sputum, and urine specimens sent to the laboratory | 936
CT of the chest and abdomen with intravenous and oral contrast | 936
fat stranding and extraluminal air | 936
free fluid around the descending colon | 936
re-exploration | 936
small abscess cavity identified | 936
Hartmann’s procedure | 936
resected specimen revealed a tiny diverticulum | 936
pathological analysis results compatible with perforated diverticulitis | 936
prolonged mechanical ventilation | 936
tracheostomy | 936
discharged to a rehabilitation hospital | 3528