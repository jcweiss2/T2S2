44 years old | 0
female | 0
admitted to the emergency department | 0
left groin and inner thigh redness | -72
left groin and inner thigh pain | -72
left groin and inner thigh swelling | -72
fever | -72
chills | -72
vomiting | -72
treated with intravenous vancomycin | -24
discharged on oral antibiotics | -24
afebrile | 0
normotensive | 0
tachycardia | 0
mild tachypnea | 0
left inner thigh and groin induration | 0
morbidly obese | 0
BMI>45 kg/m2 | 0
lactate 3.5 mmol/L | 0
WBC 18.2 × 103 per mm3 | 0
hemoglobin 12.3 g/dL | 0
sodium 136 mmol/dL | 0
glucose 225 mg/dL | 0
creatinine 1.8 mg/dL | 0
LRINEC score of 6 | 0
bedside ultrasound | 0
positive subcutaneous thickening | 0
positive air | 0
positive fascial fluid | 0
started on intravenous vancomycin | 0
started on piperacillin/tazobactam | 0
surgery consulted | 0
operative debridement of the left groin and perineum | 2
excision of 15 cm × 23 cm of tissue | 2
extensive washout | 2
admitted to the surgical intensive care unit | 2
septic shock | 2
requiring vasopressors | 2
ventilator dependence | 2
repeat washouts with minor debridements | 26
lactate normalization | 74
down-trending WBC to 13.5 × 103 per mm3 | 74
extubated | 122
transferred to a step-down unit | 122
plastic surgery consulted | 122
evaluate for possible skin graft | 122
deemed to be a poor graft candidate | 218
wound vacuum-assisted closure (V.A.C.) device placed | 218
transferred to the plastic surgery service | 218
discharged home with a wound V.A.C. | 672
received a skin graft | 672