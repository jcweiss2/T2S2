55 years old | 0
female | 0
admitted to the hospital | 0
abdominal pain | -240
diabetes mellitus | -18000
coronary by-pass operation | -8760
left infrapatellar amputation | -2880
chronic renal failure | -1752
hemodialysis treatment | -876
no history of abdominal trauma | 0
White Blood Cell: 15 100/mm3 | 0
Hemoglobin: 8.5 g/dL | 0
C-reactive protein: 40 mg/dL | 0
Urea: 37.9 mg/dL | 0
Creatinine: 2.25 mg/dL | 0
Albumin: 2.4 g/dL | 0
Sodium: 134 mmol/L | 0
Potassium: 3.1 mmol/L | 0
Calcium: 7.9 mg/dL | 0
Glucose: 329 mg/dL | 0
diffusely tender abdomen | 0
guarding | 0
rebound tenderness | 0
blood temperature: 38.7°C | 0
abdominal ultrasonography | 0
diffuse intraabdominal free fluid collection | 0
abdominal computed tomography | 0
free fluid collections in all abdominal quadrants | 0
intraabdominal minimal free air images | 0
air-fluid images in the splenic parenchyma | 0
radiology department reported gastrointestinal perforation | 0
urgently operated | 0
intraabdominal seropurulent fluid aspirated | 0
diffuse fibrin matrixes in the entire peritoneum | 0
no intestinal perforation | 0
perforated abscess pouch | 0
splenectomy | 0
drainage | 0
abdominal cavity irrigated | 0
postoperatively monitored in intubated state | 0
no proliferation in blood culture | 0
Escherichia coli isolated from abscess culture | 0
Meropenem treatment | 0
Metronidazole treatment | 0
dialysis program maintained | 0
died on postoperative Day 25 | 600
septic shock | 600
multiple organ failure | 600
histopathologic examination | 600
suppurative inflammation | 600
abscess formation of the splenic tissue | 600