59 years old | 0
male | 0
unhealthy | 0
admitted to the emergency department | 0
generalized weakness | -12
chest pain | -12
dyspnea | -12
back pain | -12
chronic obstructive pulmonary disease | -8760
coronary artery disease | -8760
bypass surgery | -8760
insulin dependent diabetes mellitus | -8760
obstructive sleep apnea | -8760
morbid obesity | -8760
urinary retention | -8760
indwelling urinary catheter | -8760
Do Not Resuscitate order | 0
tachycardia | 0
hypertensive | 0
increasing oxygen requirements | 0
leukocytosis | 0
acute renal insufficiency | 0
scrotal cystocele | -8760
mild hydronephrosis | -8760
ureters inserting into the bladder cephalad to the symphysis pubis | -8760
distended bladder within the right hemiscrotum | 0
bladder trigone migrated outside of the pelvis | 0
ureters coursing anterior and distal to the pubic symphysis | 0
catheter removed | 0
hypotensive | 12
transferred to the intensive care unit | 12
bedside ultrasound | 12
holding sutures into the anterior scrotum | 12
14fr catheter placed | 12
stabilized in the ICU | 24
discharged | 120
follow up cystoscopy | 720
catheter exchanges | 720
no symptomatic infections | 720
neocystotomy tube | 12