3 years 2 months | 0
female | 0
admitted to the hospital | 0
personality changes | -336
behavioral regression | -288
unsteady gait | -288
headache | -288
irritable crying | -288
catatonia-like response | -288
generalized choreoathetoid movements | -288
orofacial dyskinesia | -288
collapsed lung | -288
transferred to the pediatric intensive care unit | -288
cerebrospinal fluid analysis | -288
pleocytosis with predominance of lymphocytes | -288
brain magnetic resonance imaging | -288
leptomeningeal enhancement at bilateral frontoparietal area | -288
nodular enhancement along the tentorium | -288
tiny white-matter lesions over bilateral frontal lobes | -288
global cortical dysfunction | -288
electroencephalogram | -288
no epileptiform discharge | -288
empirically treated with acyclovir | -288
empirically treated with azithromycin | -288
cerebrospinal fluid NMDA receptor antibody study | -288
reported positive results | -288
treated with intravenous immunoglobulin | 0
treated with pulse methylprednisolone therapy | 0
treated with maintenance oral prednisolone | 0
aripiprazole | 0
midazolam sedation | 0
choreoathetosis recovered partially | 168
orofacial dyskinesia recovered partially | 168
discontinued prednisolone | 504
episodic sepsis | 504
autonomic instability | 504
poorly-controlled gastrointestinal bleeding | 504
plasmaphoresis | 744
anaphylactic reactions | 744
bilateral pneumonia | 744
collapsed lung | 744
rituximab | 1008
cyclophosphamide pulse therapy | 1008
azathioprine | 1344
passive range-of-motion exercise | 1008
intensive facilitation | 1344
postural training | 1344
temporary percutaneous endoscopic gastrostomy | 1344
discharged | 1680
outpatient rehabilitation | 1680
physical therapy | 1680
occupational therapy | 1680
speech therapy | 1680
cognitive deficits | 1680
cognitive–behavioral therapy | 2160
intelligence quotient | 2160
mild mental retardation | 2160
full IQ = 62 | 2160
performance IQ | 2160
verbal IQ | 2160
reached full development in gross-motor milestones | 3024
regained control of continence sphincters | 3024
communicate in complete sentences | 3024
improved reasoning | 3024
IQ test | 4320
no significant change | 4320
performance IQ improvement | 4320
mild mental retardation | 4320
mildly impulsive personality | 4320
easily distracted | 4320