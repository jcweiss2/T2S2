68 years old | 0
male | 0
type II diabetes mellitus | -672
peripheral neuropathy | -672
hypertension | -672
chronic obstructive pulmonary disease | -672
bipolar depression | -672
gastroesophageal reflux | -672
shortness of breath | -336
cough | -336
decrease in exercise tolerance | -336
intermittent diarrhea | -336
admitted to the hospital | 0
treated with vancomycin | 0
treated with piperacillin/tazobactam | 0
transferred to the medical intensive care unit | 0
dopamine started for hypotension | 0
presumed sepsis | 0
condition stabilized | 24
transferred to a medical floor | 24
pulmonary embolus | 48
colonic distension | 48
profuse watery diarrhea | 48
diagnosed with colonic pseudo-obstruction | 48
nasogastric tube placed | 48
rectal tube placed | 48
renal service consulted for hypokalemia | 48
aspirin 81 mg daily | 0
atorvastatin 80 mg daily | 0
budesonide/formoterol | 0
levalbuterol | 0
tiotroprium | 0
insulin | 0
pantoprazole 40 mg daily | 0
piperacillin/tazobactam | 0
potassium chloride 100 mEq daily | 48
blood pressure 103/50 mm Hg | 48
pulse 102 beats per minute | 48
respiratory rate 24 breaths per minute | 48
tachypneic | 48
using accessory muscles | 48
rhonchi in the anterior lung fields | 48
abdomen distended | 48
hypoactive bowel sounds | 48
tenderness to palpation in the right upper quadrant | 48
tenderness to palpation in the midepigastric area | 48
trace lower extremity edema | 48
Foley catheter in place | 48
rectal tube in place | 48
serum sodium concentration 146 mmol/l | 48
serum chloride 118 mmol/l | 48
serum potassium 2.7 mmol/l | 48
serum bicarbonate 19.9 mmol/l | 48
blood urea nitrogen 6.1 mmol/l | 48
serum creatinine 110 μmol/l | 48
arterial blood gases pH 7.27 | 48
arterial blood gases pCO2 36.9 mm Hg | 48
arterial blood gases bicarbonate 17.1 mEq/l | 48
urine sodium 49 mmol/l | 48
urine potassium 20 mmol/l | 48
urine chloride 90 mmol/l | 48
urine anion gap -21 | 48
24-hour urine collection 9.1 mmol potassium excreted | 72
stool sodium concentration <10 mmol/l | 72
stool potassium concentration 139.7 mmol/l | 72
marked colonic distension | 72
radiographic examination of the abdomen | 72
diagnosis of severe gastrointestinal potassium wasting | 72
large doses of potassium chloride | 72
serum potassium concentrations maintained in the 3.5–4.0 mmol/l range | 96
respiratory status deteriorated | 120
family decided to withdraw care | 120
patient expired | 144