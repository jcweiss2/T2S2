51 years old | 0
indigenous woman | 0
back pain | -120
radiating to the left flank | -120
dehydration | -120
insulin dependent type two diabetes mellitus | 0
medically managed ischaemic heart disease | 0
hypertension | 0
chronic lower back pain | 0
intra-muscular anti-inflammatories | -120
discharged | -120
vomiting | -96
flank pain | -96
confusion | -96
transferred to a regional health service | -96
blood pressure 76/53 mmHg | -96
tachypnoeic at 55bpm | -96
impaired consciousness | -96
oliguria | -96
sepsis | -96
non-ketotic high anion gap metabolic acidosis | -96
pH 7.15 | -96
lactate 10.1mmol/L | -96
hyperglycaemia | -96
blood glucose 23.5mmol/L | -96
acute kidney injury | -96
serum creatinine 348μmol/L | -96
urinalysis demonstrated leukocytes | -96
haemolysed blood | -96
protein | -96
no nitrites | -96
inflammatory markers elevated | -96
white cell count 14x10^9 | -96
CRP 156mg/L | -96
hyponatraemic | -96
thrombocytopaenic | -96
septic shock | -96
broad-spectrum antibiotics | -96
piperacillin-tazobactam | -96
gentamicin | -96
resuscitation | -96
non-contrast computed tomography scan | -96
marked oedema of the left kidney | -96
hydronephrosis | -96
extensive loculated and mottled areas of gas | -96
emphysematous pyelonephritis | -96
trace perinephric gas | -96
no fluid levels | -96
no drainable collection | -96
simple cyst of the superior pole | -96
admitted to the intensive care unit | -96
vasopressor support | -96
antibiotics | -96
strict fluid balance | -96
indwelling catheter | -96
continuous veno-venous haemodialysis | -96
insulin infusion | -96
urine and blood cultures | -96
Klebsiella Pneumoniae | -96
antibiotic therapy narrowed | -48
ceftriaxone | -48
metronidazole | -48
8Fr nephrostomy tube | 0
CT guidance | 0
nephrostomy drainage | 0
organ support | 0
ability to cease CVVHD | 72
failed to show significant improvement | 72
persisting confusion | 72
high grade fevers | 72
tachycardia | 72
dependence on vasopressors | 72
parenteral analgesia infusion | 72
new anaemia | 72
Hb 82g/L | 72
persisting inflammatory rise | 72
WCC 13.6x10^9 | 72
thrombocytopaenia | 72
114x10^9 | 72
recurring deterioration in renal function | 72
Cr 142μmol/L | 72
post CVVHD nadir | 72
71μmol/L | 72
repeat imaging | 72
no parenchymal improvement | 72
open nephrectomy | 144
subcapsular approach | 144
fibrous adhesions | 144
intraoperatively | 144
post-operatively | 168
recovered well | 168
intravenous antibiotics transitioned to oral | 168
discharged | 192
creatinine 106 μmol/L | 192