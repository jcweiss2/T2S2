49 years old | 0
leucodermal | 0
male | 0
admitted to the hospital | 0
non-specific malaise | 0
feeling of postprandial infarction | 0
colic-like abdominal pain | -1440
bloodless diarrhoea | -1440
asthenia | -720
oedema of the lower limbs | -720
oedema of the face | -720
polydipsia | -720
polyuria | -720
cutaneous trunk hyperpigmentation | -720
cutaneous face hyperpigmentation | -720
non-productive cough | 0
no recent weight changes | 0
hypertension | -6720
treated with lisinopril | -6720
treated with furosemide | -6720
tobacco history | -25200
alcohol habit | -25200
dyslipidaemia | -25200
hyperuricaemia | -25200
treated with statin | -25200
treated with colchicine | -25200
lived in Brazil | -8760
lived in Angola | -8760
lived in Guinea | -8760
mild melanoderma | 0
apyrexia | 0
conscious | 0
temporally and spatially oriented | 0
weighed 96.6 kg | 0
height of 192 cm | 0
body mass index of 26.2 kg/m2 | 0
cardiac auscultation revealed no changes | 0
pulmonary auscultation revealed bilateral wheezing | 0
pulmonary auscultation revealed snoring | 0
blood pressure was 196/76 mmHg | 0
symmetrical soft oedema of the lower limbs | 0
no palpable adenopathies | 0
severe metabolic alkalosis | 0
hypokalaemia | 0
moderate hypoxaemia | 0
elevated serum adrenocorticotropic hormone | 0
elevated urinary cortisol levels | 0
bilateral pulmonary opacity | 0
renal and suprarenal ultrasonographic examination was normal | 0
admitted to the Endocrinology Department | 0
diagnostic hypotheses of Cushing’s syndrome | 0
diagnostic hypotheses of ectopic ACTH production | 0
admitted to the Intensive Care Unit | 48
diagnosis of community-acquired pneumonia | 48
invasive mechanical ventilation | 48
empirically medicated with ceftriaxone | 48
empirically medicated with azithromycin | 48
urinary screening for urinary antigens from Legionella pneumophila was negative | 48
urinary screening for urinary antigens from Streptococcus pneumoniae was negative | 48
multiple polymerase chain reaction tests for gastroenteritis were negative | 48
upper digestive endoscopy | 72
swollen duodenal folds | 72
biopsied | 72
inflammatory lamina propria infiltrate with eosinophils | 72
presence of larvae and eggs of parasitic structures compatible with Strongyloides stercoralis | 72
ultrasound-guided liver biopsy | 96
metastasis of small cell neuroendocrine carcinoma | 96
immunohistochemical profile suggesting pulmonary origin | 96
treated with ivermectin | 120
haemodynamic support | 120
ventilatory support | 120
etomidate therapy | 120
metyrapone therapy | 120
tracheostomy | 1056
transferred to the Pulmonology Department | 1680
died | 1950
eosinophilia of 8.4% | -720
eosinophilia of 7.2% | -8760
eosinophils 0.4% | 0
self-infection phenomenon | -8760
cerebral intraparenchymal haemorrhage | 1008
diffuse metastasis of carcinoma | 1008
primary lesion in the head of the pancreas | 1008
Strongyloides stercoralis infection | -8760
hyperinfection syndrome | 0
disseminated disease | 0
immunosuppressive condition | 0
spread of Strongyloides stercoralis infection | 0