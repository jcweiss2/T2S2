Here is the table of events and timestamps:

18 years old | 0
male | 0
cactus plant prick | -72
progressive left leg swelling | -72
worsening of erythema | -72
pain | -72
felt generally unwell | -72
Primary Sclerosing Cholangitis | -672
mild Ulcerative Colitis | -672
long-standing deranged liver function tests | -672
admitted to the intensive care unit (ICU) | 0
Blood Pressure (BP): 71/41mmHg | 0
Mean Arterial Pressure (MAP): 48mmHg | 0
Respiratory Rate: 36 breaths per minute | 0
Heart Rate (HR): 125 beats per minute | 0
sinus tachycardia | 0
Temperature: 39°C | 0
Oxygen Saturation: 86% with 0.21 FiO2 | 0
pH 7.15 | 0
PO2 84 | 0
HCO3 15 | 0
Lactate 7.6 | 0
Sodium (Na) 134 | 0
Urea 7.6 | 0
Creatinine (sCr) 173 | 0
eGFR 27 | 0
White Cell Count (WCC) 13.8 | 0
C-reactive protein (CRP) 22 | 0
Hemoglobin (Hb) 114 | 0
Platelet (Plt) 81 | 0
Liver Function Test (LFT)- Total Bilirubin (Bili) 99 | 0
Alanine transaminase (ALT) 61 | 0
Aspartate aminotransferase (AST) 83 | 0
Alkaline Phosphatase (ALP) 96 | 0
Piperacillin-Tazobactam IV 4.5g stat | 0
Meropenem IV 2g | 0
Lincomycin IV 600mg | 0
Vancomycin IV 2g | 0
Emergency left lower limb fasciotomy, debridement and below knee amputation | 0
extensive left foot and below knee tissue necrosis | 0
“dishwasher fluid” in appearance along with liquefied fat | 0
large areas of unviable skin and muscle | 0
Histopathology was undertaken to confirm diagnosis | 0
oliguria 10-14ml/hour | 24
severe acidosis | 24
severe acidosis requiring left internal jugular vascath insertion | 24
Continuous Renal Replacement Therapy (CRRT) | 24
pH 7.28 | 24
Lactate 4.7 | 24
Na 130 | 24
sCr 206 | 24
Hb 89 | 24
Plt 105 | 24
WCC 17 | 24
CRP 78 | 24
International normalized ratio (INR) 2.2 | 24
Activated Partial Thromboplastin Time (APTT) 150 | 24
Initial blood cultures (BCs) isolated Group B Streptococcus pneumoniae (GBSPn) | 24
Ventilation sedation: Propofol 170mg/hr | 24
Fentanyl 40mcg/hr | 24
CRRT (Day 1) on heparin circuit commenced | 24
Renal dose - 30ml/kg/hr | 24
Triple vasopressor support continued: Noradrenaline 23mcg/min | 24
Adrenaline 18mcg/min | 24
Vasopressin 0.04units/min | 24
Antibiotics (MLV): Meropenem IV 2g TDS | 24
Lincomycin IV 600mg TDS | 24
Vancomycin IV 2g BD | 24
Intravenous Immunoglobin G (IVIgG) therapy 100g was initiated | 24
taken back to theatre to confirm source control and the viability of the left stump | 48
no evidence of necrotic tissue | 48
Remained intubated but developed new onset of Rapid Atrial Fibrillation (RAF) with HR 110bpm | 48
patient remained oliguric 7-25ml/hour | 48
pH 7.40 | 48
Lactate 3.9 | 48
Na 131 | 48
sCr 116 | 48
WCC 26 | 48
CRP 105 | 48
Procalcitonin (PCT) 21.18 μg/L | 48
Hb 83 | 48
Plt 63 | 48
INR 3.1 | 48
Fibrinogen 2.4 | 48
Echocardiography: Moderate segmental left ventricular dysfunction | 48
Ejection Fraction 40-45% | 48
Dilated atria bilaterally | 48
Raised Right Atrial Pressure | 48
Amiodarone loading dose 300mg over 1 hour | 48
Amiodarone infusion | 48
Antibiotics remained unchanged (MLV) | 48
CRRT (Day 2) – AN69 anti-inflammatory heparin laden adsorbing filter applied | 48
Oxiris Filter | 48
Citrate based anticoagulation circuit applied | 48
developed features consistent with Sepsis Induced Coagulopathy (ISTH -SIC criteria) | 72
bedside surgical debridement was performed by surgical team | 72
pH 7.31 | 72
Lactate 2.4 | 72
Na 135 | 72
sCr 79 | 72
WCC 27 | 72
CRP 127 | 72
Hb 78 | 72
Plt 50 | 72
INR 2.0 | 72
Histopathology consistent with NF | 72
Wound culture for microscopy culture and sensitivity (MCS) had medium growth of GBSPn | 72
Tissue culture (intraoperatively) had medium growth of GBSPn | 72
Vasopressor support - weaning: Noradrenaline 20mcg/min | 72
Adrenaline weaned off | 72
Vasopressin 2.4units/min | 72
Antibiotics remained unchanged (MLV) | 72
CRRT (Day 3) - ongoing | 72
patient remained oliguric (6-20ml/hr) | 96
despite being challenged with a single dose Furosemide IV 250mg stat | 96
Citrated based CRRT was continued | 96
new onset purpura over the right forearm | 96
multiple weeping skin tears on right upper thigh | 96
Ongoing RAF HR 130 | 96
pH 7.36 | 96
Lactate 1.5 | 96
Na 130 | 96
sCr 116 | 96
WCC 33 | 96
CRP 103 | 96
PCT 15.37 | 96
Hb 91 | 96
Plt 53 | 96
INR 1.7 | 96
LFT - Bili 131 | 96
AST 127 | 96
ALP 121 | 96
Double inotropic support: Noradrenaline 20mcg/min | 96
Vasopressin 2.4units/min | 96
Antibiotics remained unchanged (MLV) | 96
CRRT (Day 4) | 96
Amiodarone infusion | 96
patient developed fulminant hepatic failure/ encephalopathy | 120
refractory oliguria 0-5ml/hr | 120
pH 7.39 | 120
Lactate 1.2 | 120
Na 134 | 120
sCr 124 | 120
WCC 39.5 | 120
CRP 74 | 120
Hb 116 | 120
Plt 49 | 120
INR 1.5 | 120
LFT- Bili 139 | 120
AST 69 | 120
ALT 97 | 120
ALP 140 | 120
Dual inotropic support: Noradrenaline 20mcg/min | 120
Vasopressin weaned off | 120
Antibiotics remained unchanged (MLV) | 120
CRRT (Day 5) | 120
patient was severely deconditioned | 144
developed ICU acquired weakness | 144
unarousable and had no response to noxious stimuli | 144
Remained intubated and ventilated on Pressure Support Ventilation | 144
Refractory oliguria at 5ml/hr | 144
pH 7.44 | 144
Lactate 1.1 | 144
WCC 43.5 | 144
CRP 109 | 144
Hb 90 | 144
Plt 57 | 144
INR 1.5 | 144
LFT - Bili 150 | 144
AST 95 | 144
ALP 154 | 144
Sedation weaned off | 144
Off vasopressor | 144
Noradrenaline weaned off | 144
Antibiotic de-escalation: Lincomycin and Vancomycin ceased | 144
Meropenem IV 2g TDS continued | 144
CRRT (Day 6) | 144
Hyper-Ammonium Therapy initiated - Rifaximin NGT 550mg BD | 144
Lactulose NGT 20ml TDS | 144
2 units of PRBCs transfusion | 144
patient developed jaundice | 168
hypoactive delirium | 168
remained deeply sedated despite being off sedation with a RASS -5 | 168
new onset lateralizing signs to the left upon painful stimuli compared to the right side | 168
Refractory oliguria | 168
CT Brain: No acute intracranial pathology | 168
Ultrasound abdomen: Acute Calculous Cholecystitis noted | 168
pH 7.44 | 168
Lactate 1.1 | 168
WCC 44.3 | 168
CRP 109 | 168
Hb 129 | 168
Plt 66 | 168
INR 1.3 | 168
LFT - Bili 235 | 168
AST 75 | 168
ALP 175 | 168
Conjugated Bilirubin 142 | 168
Meropenem IV 2g TDS | 168
CRRT (Day 7) on a Heparin circuit | 168
anuria was established by this stage | 192
hypotensive BP 71/33 | 192
MAP 51mmHg | 192
Febrile 39°C | 192
RAF HR 160 | 192
Significant deterioration despite ongoing medical therapy | 192
patient was commenced on palliative care pathway | 192
deceased shortly post treatment withdrawal | 192
Troponin 616 | 192
Ammonia 158 | 192
LFT - Bili 352 | 192
AST 100 | 192
ALP 299 | 192
CRRT (Day 8) Renal recovery assessment | 192
challenged with combination of Furosemide IV 250mg and Acetazolamide IV 500mg | 192
Recommenced Vasopressor support; Noradrenaline 2.5mcg/min | 192
Antibiotic regimen: Lincomycin IV 600mg TDS – recommenced as antitoxin | 192
Meropenem IV 2g TDS – continued | 192
Digoxin IV 500mcg | 192
Metoprolol IV 15mg | 192