83 years old | 0
    female | 0
    atrial fibrillation | 0
    hypertension | 0
    hyperlipidemia | 0
    type 2 diabetes mellitus | 0
    small bowel obstruction | 0
    exploratory laparotomy | 0
    ventral hernia repair | 0
    abdominal wound infections | 0
    multiple debridements | 0
    discharge | 0
    fever | 0
    chills | 0
    purulent drainage from abdominal wounds | 0
    sepsis | 0
    7.5 Fr triple lumen right internal jugular vein CVC placement | 0
    post-procedure chest X-ray demonstrating possible arterial cannulation | 0
    contrasted computed tomography scan | 0
    CVC penetration of right internal jugular vein | 0
    CVC penetration into right subclavian artery | 0
    CVC termination in aortic arch | 0
    right-sided aortic arch anatomical variant | 0
    separate origins of RSCA and RCCA | 0
    tortuous course of arch vessels | 0
    LCCA arising from aorta most proximally | 0
    RCCA | 0
    RSCA | 0
    LSCA with Kommerel’s diverticulum | 0
    transfer to intervention facility | 0
    endovascular intervention of central arterial stent graft placement via open brachial access | 0
    right brachial artery cutdown | 0
    systemic heparinization with 5000 units of unfractionated heparin | 0
    modified Seldinger technique access | 0
    intravascular ultrasound | 0
    angiography | 0
    vertebral artery origin identified | 0
    proximity of vertebral artery to CVC entry site | 0
    imaging suggested suitable landing zone for stent graft | 0
    deployment of 11 × 29 mm Gore VBX stent graft | 0
    stent graft deployment in proximal subclavian artery | 0
    proximal portion overhang into aortic arch | 0
    CVC removal from between stent graft and arterial wall | 0
    balloon angioplasty with 14 × 40 mm balloon | 0
    completion angiogram revealing no contrast extravasation | 0
    extubation | 0
    observation in surgical intensive care unit | 0
    500 unit/hr flat-rate heparin infusion | 0
    transition to home anticoagulant (apixaban) on postoperative day 2 | 48
    transfer to floor on postoperative day 1 | 24
    discharge on postoperative day 7 | 168
    apixaban therapy | 168
    aspirin therapy | 168
    oral doxycycline | 168
    cefpodoxime | 168
    arterial duplex at 1-month follow-up | 720
    normal arterial duplex | 720
    medication regimen transition to apixaban monotherapy | 720
