65 years old | 0
male | 0
diabetes | -4800
admitted to the hospital | 0
fever | -120
headache | -120
dizziness | -120
cough | -120
poorly managed diabetes mellitus | -4800
cranial MRI | 0
multiple abnormal signals | 0
encephalitis | 0
chest CT scan | 0
multiple lung inflammations | 0
pleural adhesions | 0
pleural effusion | 0
C-reactive protein (CRP) level | 0
severe infection | 0
neck stiffness | 0
deep coma | 0
Glasgow Coma Scale score of 5 | 0
weakness | 0
nausea | 0
repeated vomiting | 0
intensive care unit (ICU) admission | 0
lumbar puncture | 24
cerebrospinal fluid (CSF) analysis | 24
cloudiness | 24
white blood cell count | 24
glucose level | 24
microprotein level | 24
Pan's test | 24
HvKP infection | 48
metagenomic next-generation sequencing (mNGS) | 48
virulence factors | 48
rmpA | 48
iutA | 48
iucA | 48
iucB | 48
iucC | 48
iucD | 48
iroB | 48
iroC | 48
iroD | 48
fimH | 48
drug sensitivity analysis | 48
resistance to piperacillin | 48
resistance to levofloxacin | 48
sensitivity to amikacin | 48
severe intracranial infection | 0
community-acquired HvKP pathogen | 0
meropenem | 0
amikacin | 0
fever subsided | 72
vital signs stabilized | 72
blood sugar levels monitoring | 72
repeat CSF analysis | 216
clarity | 216
colorlessness | 216
no presence of microorganisms | 216
regained consciousness | 264
endotracheal tube extubated | 264
antimicrobial treatment | 504
discharged | 504