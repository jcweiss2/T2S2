57 years old | 0
male | 0
Chinese | 0
admitted to the hospital | 0
fever | -72
lumbago | -72
right flank pain | -72
fatigue | -72
poorly controlled diabetes | -8760
smoking | -10950
drinking | -10950
stopped smoking | -72
stopped drinking | -72
POCUS | 0
hyperechoic spotted or patchy foci | 0
dirty shadowing | 0
comet-tail artifacts | 0
falls sign | 0
septic shock | 0
transferred to ICU | 0
abdominal CT scan | 0
gas in the right perirenal space | 0
enlarged right kidney | 0
perinephric fat stranding | 0
mild right hydronephrosis | 0
no urinary stones | 0
leukocytosis | 0
neutrophils | 0
hemoglobin | 0
thrombocytopenia | 0
elevated serum creatinine | 0
inflammation markers | 0
elevated glycosylated hemoglobin | 0
heavy pyuria | 0
white blood cell count | 0
arterial blood gas analysis | 0
pH | 0
partial pressure of carbon dioxide | 0
partial pressure of oxygen | 0
bicarbonate | 0
elevated lactate | 0
blood culture | 0
urine culture | 0
Escherichia coli bacteremia | 0
broad-spectrum antibiotic therapy | 0
meropenem | 0
tigecycline | 0
fluid resuscitation | 0
insulin infusion | 0
vasopressor support | 0
CT-guided PCD | 72
percutaneous catheter drainage | 72
abscess in the right perirenal space | 72
pig-tail catheter | 108
discharged | 336
oral levofloxacin | 336
follow-up | 504
repeat urinary CT scan | 504
normal kidney imaging | 504
stable blood glucose control | 504
normal renal function | 504