79 years old | 0
female | 0
admitted to the intensive care unit | 0
thoracoabdominal aortic aneurysm | 0
surgical interposition graft | 0
hypertension | 0
chronic obstructive pulmonary disease | 0
chronic kidney disease | 0
creatinine 105 μmol/l | 0
MDRD 44 ml/min | 0
transcatheter aortic valve implantation | 0
percutaneous coronary intervention of the right coronary artery | 0
vascular graft of the abdominal aorta below the renal arteries | 0
acute-on-chronic kidney failure | 0
continuous veno-venous haemofiltration | 0
persistent chylous leakage | 0
re-thoracotomy | 0
third-degree atrioventricular block | 0
pacemaker implanted | 0
surgical tracheostomy | 0
mechanical ventilator | 0
Staphylococcus aureus bacteraemia | -840
infected thoracotomy wound | -840
pleural fluid cultures positive for Staphylococcus aureus | -840
continuous intravenous flucloxacillin 12 g/24 hours | -840
high flucloxacillin blood concentrations | -816
flucloxacillin dosage decreased to 3 g/24 hours | -816
flucloxacillin dosage changed to 6 g/24 hours | -720
acetaminophen 3 g per day | -840
appendicitis | -576
surgery postponed | -576
antibiotics (piperacillin-tazobactam) | -576
supportive care | -576
reduced consciousness | -432
controlled mechanical ventilation | -432
severe respiratory acidosis | -432
high anion gap metabolic acidosis | -432
pH 7.16 | -432
pCO2 7.1 kPa | -432
pO2 14.9 kPa | -432
bicarbonate 18.5 mmol/l | -432
base excess −9.6 mmol/l | -432
lactate 1.1 mmol/l | -432
sodium 143 mmol/l | -432
potassium 3.7 mmol/l | -432
chloride 107 mmol/l | -432
albumin 13 g/l | -432
creatinine 158 μmol/l | -432
MDRD-GFR 27 ml/min | -432
5-oxoprolinaemia | -432
acetaminophen prescription stopped | -432
progression of abdominal pain | -408
CT scan of the abdomen | -408
intra-abdominal abscesses | -408
ICU treatment stopped | -408
patient died | -408
urinary 5-oxoproline 1,721 μmol/mmol/creatinine | -408
creatinine 1.69 mmol/l | -408
