65 years old | 0
female | 0
nausea | -8760
vomiting | -8760
loss of appetite | -8760
weight loss | -8760
open cholecystectomy | -10440
cure for eventration | -10320
admitted to the hospital | 0
afebrile | 0
normal respiratory rate | 0
normal resting heart rate | 0
midline vertical scar | 0
no palpable masses | 0
digital rectal exam normal | 0
digital examination of the vagina normal | 0
Eso-gastro-duodenal fibroscopy | 0
extrinsic compression of the lesser curvature | 0
erythematous mucosa | 0
biopsy | 0
mixed dense lymphoid infiltrate | 0
abdominal CT scan | 0
heterogeneous formation | 0
duodenal mass | 0
multiple parietal and central calcifications | 0
thoracic CT scan | 0
no secondary lesions | 0
CA 19-9 slightly raised | 0
ACE normal | 0
preanesthesic assessment | 0
surgery | 0
tumor ablation | 0
laparotomy | 0
irregular contour mass | 0
release of the mass from the duodenum | 0
biopsies of the duodenal edges | 0
atypical segmental hepatectomy | 0
kellyclasia | 0
abdomen closed | 0
counts of surgical items | 0
surgical sponge found | 0
histological report confirmed necrotic textiloma | 0
extubated | 6
respiratory distress | 72
thoraco-abdominal CT | 72
lesion related to infection lung | 72
treated by ATB | 72
transferred to intensive care unit | 72
intubated | 72
ventilated | 72
hypotension | 72
tachycardia | 72
cardio-respiratory arrest | 240
died | 240