71 years old | 0
    woman | 0
    admitted to the emergency department | 0
    dyspnea | 0
    thyroid excision | -2400
    spinal fusion | -2400
    follicular thyroid cancer | -2400
    lung metastasis | -2400
    cranial bone metastasis | -2400
    vertebrae metastasis | -2400
    spinal metastasis recurrence | -2400
    acetaminophen | -2400
    loxoprofen | -2400
    morphine | -2400
    pulse 118 beats per minute | 0
    blood pressure 121/86 mmHg | 0
    respiratory rate 28 breaths per minute | 0
    oxygen saturation 96% | 0
    no significant heart murmurs | 0
    ST-segment elevation in leads I, aVL, V2-5 | 0
    cardiothoracic ratio 71% | 0
    pulmonary congestion | 0
    infiltrative shadow | 0
    apical akinesis | 0
    basal hyperkinesis |