84 years old | 0
female | 0
diabetes mellitus | 0
hypertension | 0
paroxysmal atrial fibrillation | 0
old cerebrovascular event | 0
left middle cerebral artery infarction | 0
no residual weakness | 0
ambulatory | 0
acceptable cardiorespiratory status | 0
admitted to hospital | 0
left intertrochanteric femur fracture | 0
Gama nailing of femur | 24
postoperative course uneventful | 24
right-sided hemiparesis | 168
altered mental status | 168
Glasgow coma scale 10/15 | 168
noncontrast computed tomography of brain | 168
bilateral cerebrospinal fluid hygroma | 168
left parietal Burr hole | 168
evacuation of CSF hygroma | 168
general anesthesia | 168
extubated | 168
intensive care unit | 168
Glasgow coma scale 15/15 | 168
persistent right-sided hemiparesis | 168
generalized tonic-clonic seizures | 174
Glasgow coma scale 5/15 | 174
intubation | 174
sedation | 174
fentanyl | 174
midazolam | 174
mechanical ventilation | 174
levetiracetam | 174
computed tomography of brain | 174
near-complete evacuation of bilateral CSF hygroma | 174
development of classic “Mount Fuji” sign | 174
tension pneumocephalus | 174
maintenance in flat position | 174
100% oxygen | 174
sedation | 174
antiepileptic | 174
brain-protective measures | 174
left frontoparietal decompressive craniectomy | 174
general anesthesia | 174
intensive care unit | 174
sedation | 216
computed tomography of brain | 216
near-complete resolution of pneumocephalus | 216
sedation stopped | 216
Glasgow coma scale 9/15 | 216
tracheotomy | 474
low GCS | 474
ventilator-associated pneumonia | 474
sepsis | 474
acute kidney injury | 474
multi-organ failure | 474
death | 600
consent for publication | 600
case report approved | 600