83 years old | 0
female | 0
admitted to hospital | 0
chest pain | 0
abdominal pain | 0
severe hypotension | 0
normal ECG | 0
no change in cardiac enzymes levels | 0
ileus | 0
hypovolemic shock | 0
septic shock | 0
admitted to intensive care unit | 0
feculent vomiting | 1
cardiorespiratory arrest | 1
resuscitation | 1
unsuccessful resuscitation | 1
autopsy | 60
pallor of the entire body skin | 60
fibrosis of myocardial muscle | 60
hypertrophy of myocardial muscle | 60
pulmonary oedema | 60
cerebral oedema | 60
hematoma in left hypochondrium | 60
liver cyanosis | 60
fatty changes in liver | 60
splenic cyanosis | 60
right kidney with single cyst | 60
left kidney surrounded by hematoma | 60
chronic gastric ulcer | 60
no signs of acute hemorrhage | 60
arteries severely atherosclerotically changed | 60
abdominal aortic rupture | 60
pulmonary cyanosis | 60
pulmonary myelolipoma | 60
well-circumscribed yellow-brown nodule | 60
calcified nodule | 60
mature adipose tissue | 60
hematopoietic cells | 60
myeloid cells | 60
megakaryocytes | 60
erythroid cells | 60
mature bony tissue | 60
no foci of extramedullary hematopoiesis | 60
death | -1 
abdominal aortic rupture diagnosis | 60 
myelolipoma diagnosis | 60 
no symptoms related to myelolipoma | 0 
no treatment of myelolipoma | 60 
monitoring of myelolipoma | 60 
no malignant transformation of myelolipoma | 60 
distinguishing myelolipoma from malignant lesions | 60 
surgical removal of myelolipoma | 60 
myelolipoma rupture | 60 
life threatening hemorrhage | 60 
compression of adjacent structures | 60