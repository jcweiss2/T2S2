55 years old | 0
female | 0
admitted to the oncology centre | 0
abdominal distension | -168
ovarian cancer | -8760
hysterectomy | -8760
bilateral salpingo-oophorectomy | -8760
chemotherapy | -8760
normochromic normocytic anaemia | 0
healthy liver function | 0
healthy kidney function | 0
normal clotting limits | 0
ascites | 0
pleural effusion | 0
pelvic mass | 0
diffuse large B cell lymphoma (DLBCL) | 0
pleuritic tap | 0
cytology | 0
biopsy | 0
pleural effusion drained | 0
ascites drained | 0
persistent tachycardia | 168
respiratory failure | 168
intubation | 168
ventilation | 168
metabolic acidosis | 168
respiratory compensation | 168
pH 7.29 | 168
CO2 29mmHg | 168
pO2 77mmHg | 168
FiO2 0.5 | 168
BE -11.7 | 168
HCO3- 13mmol/L | 168
lactate 5.7mmol/L | 168
anion gap 18 | 168
pneumoperitoneum | 168
left lower zone lung consolidation | 168
emergency exploratory laparotomy | 168
septic shock | 168
hypoperfusion | 168
tissue hypoxia | 168
noradrenaline infusion | 168
fluid boluses | 168
blood pressure 82/50 mmHg | 168
blood pressure 90/60 mmHg | 168
Vancomycin | 168
Caspofungin | 168
Meropenem | 168
broad-spectrum empirical antibiotics | 168
feculent peritonitis | 168
hospital-acquired pneumonia | 168
Fentanyl infusion | 168
postoperative analgesia | 168
Noradrenaline infusion weaned off | 192
tachycardia | 192
lactic acidosis | 192
urine output 0.5-1ml/kg/hr | 192
PlasmaLyte infusion | 192
20% human albumin solution | 192
positive fluid balance | 192
left shift neutrophilia | 192
liver function tests normal | 192
renal function tests normal | 192
respiratory failure resolved | 336
hyperlactatemia plateaued | 336
Type A LA | 336
Type B LA | 336
intra-abdominal sepsis | 336
Klebsiella pneumoniae | 336
Candida tropicalis | 336
blood cultures | 336
Meropenem-resistant | 336
Ceftazidime-Avibactam | 336
respiratory wean | 336
severe tachypnoea | 336
spontaneous respiratory rate 35-45 breaths/min | 336
pressure support ventilation | 336
respiratory compensation | 336
lactic acidosis | 336
LDH elevated | 432
DLBCL activity | 432
CRRT | 432
lactate clearance | 432
chemotherapy | 432
cyclophosphamide | 432
rituximab | 432
etoposide | 432
Type B LA resolved | 504
extubated | 672
transferred out of ICU | 672
succumbed to DLBCL | 10080