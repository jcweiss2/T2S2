48 years old | 0
male | 0
admitted to the hospital | 0
pain | 0
distension of abdomen | 0
low-grade fever | -720
cough | -720
scanty expectoration | -720
weight loss | -720
bilateral upper zone opacities | 0
anti-tubercular therapy | -720
Directly Observed Treatment Shortcourse-Category I | -720
sputum negative for acid fast bacilli | -720
pulse rate 112/min | 0
blood pressure 134/86 mm Hg | 0
respiratory rate 36/min | 0
temperature 100°F | 0
abdomen distended | 0
abdomen tender | 0
rigidity | 0
guarding | 0
tenderness aggravated by movement | 0
tenderness aggravated by cough | 0
tympanitic percussion note | 0
vesicular breath sounds diminished intensity | 0
coarse crackles bilaterally over infraclavicular areas | 0
perforated hollow viscous abdomen | 0
hemoglobin 110 g/L | 0
total leukocyte count 11.2 × 10^9/L | 0
neutrophil 68% | 0
lymphocytes 27% | 0
polymorphonuclear leukocytosis | 0
no parasite | 0
no premature cell | 0
aspartate transaminase 64 U/L | 0
alanine transaminase 78 U/L | 0
alkaline phosphatase 156 U/L | 0
random plasma glucose 98 mg/dL | 0
blood urea nitrogen 12 mmol/L | 0
creatinine 1.1 μmol/L | 0
sodium 134 mEq/L | 0
potassium 3.4 mEq/L | 0
serum amylase normal | 0
serum lipase normal | 0
routine urine examination normal | 0
HbSAg negative | 0
anti-hepatitis C virus negative | 0
HIV test negative | 0
chest radiograph infiltrations in bilateral upper zones | 0
increased broncho vascular markings | 0
X-ray abdomen erect posture free gas under diaphragm | 0
ultrasonography abdomen intraperitoneal gaseous distension | 0
intraperitoneal free fluids with internal echogenicity | 0
exploratory laparotomy | 0
midline incision | 0
purulent fluid 500 ml | 0
two small perforations 1cm apart | 0
ileocaecal junction 20 cm proximal | 0
pus sample collected for microbiological study | 0
peritoneal lavage | 0
perforations sealed with omental fat | 0
pelvic drain | 0
incision closed in single layer | 0
postoperative tidal volume low | 24
postoperative respiratory distress | 24
shifted to intensive care unit | 24
mechanical ventilation | 24
intravenous piperacillin-tazobactam | 24
intravenous amikacin | 24
Gram-negative bacilli with bipolar staining | 24
pus culture lactose fermenting pink colonies MacConkey's agar | 24
dry and wrinkled colonies on day 4 | 96
B. pseudomallei suspected | 96
ceftazidime 2g 8h | 144
amikacin continued | 144
organism confirmed B. pseudomallei | 144
oxidase positive | 144
nitrate reduction test positive | 144
arginine dihydrolase activity | 144
glucose oxidation | 144
lactose oxidation | 144
imipenem sensitive | 144
doxycyclin sensitive | 144
cotrimoxazole sensitive | 144
imipenem 1g 8h | 216
doxycyclin 100mg twice daily | 216
ventilator weaned off | 216
T-piece ventilation with oxygen | 216
T-piece removed | 288
oxygen saturation maintained in room air | 288
imipenem continued | 336
doxycyclin continued | 336
cotrimoxazole 160+800mg | 336
discharged | 576
cotrimoxazole continued for 4 months | 576
follow-up after 6 months | 4320
no relapse | 4320
abdomen tender |(Output exceeds around 1000 words. Complete the answer. Then explain why you think so)
