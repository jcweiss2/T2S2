69 years old | 0
male | 0
advanced prostate cancer | -6720
multiple bone metastases | -6720
PSA 1149 ng/ml | -6720
orchiectomy | -6720
maximal androgen blockade | -6720
PSA decreased to 3.3 ng/ml | -6720
PSA increased | -150
anti-androgen therapy discontinued | -120
estramustine administered | -120
PSA increased to 32.6 ng/ml | 0
docetaxel therapy started | 0
performance status 1 | 0
nonsmoker | 0
normal chest X-ray | 0
normal lung sound | 0
prednisone 5 mg twice daily | 0
intravenous dexamethasone 20 mg | 0
docetaxel 75 mg/m2 | 0
PSA level decreased to 2.7 ng/ml | 42
leucopenia | 42
G-CSF injected | 42
leucocytes increased to 9.4×10^3/ul | 42
dyspnea | 210
cough | 210
sputum | 210
fever 39.2℃ | 210
mild diffuse fine crackle | 210
elevated leukocyte count | 210
blood gas pH 7.422 | 210
blood gas pCO2 21.4 mmHg | 210
blood gas pO2 58.3 mmHg | 210
diffuse reticulonodular shadow in both lungs | 210
sputum and blood cultures negative | 210
empiric broad-spectrum antibiotics administered | 210
high-dose corticosteroids administered | 210
vancomycin administered | 210
ceftriaxone administered | 210
piperacillin/tazobactam administered | 210
septic shock | 213
O2 saturation decreased to 80% | 213
intubated | 213
mechanical ventilation | 213
dopamine administered | 213
cardiopulmonary resuscitation | 214
death | 214