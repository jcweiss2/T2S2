32 years old | 0
female | 0
family history of polycystic kidney disease | 0
admitted to the hospital | 0
hemorrhagic left renal cyst | - hours unknown, assume -24 
stable vital signs | 0
abdomen distended | 0
left kidney palpable | 0
hemoglobin level of 9.6 g/dl | 0
creatinine level: 64 μmol/l | 0
enhanced Computed Tomography (CT) of the abdomen | 0
polycystic kidneys | 0
enlarged left kidney with a hemorrhagic component | 0
no signs of active bleeding | 0
discharged home | 24
followed as an outpatient | 24
seen in the clinic 10 days later | 240
abdominal pain | 240
abdomen distended more | 240
admit her electively for angioembolization | 240
repeated enhanced CT | 240
left complex renal cyst with thick septation | 240
enhancement with contrast extravasation | 240
suggesting active bleeding | 240
angiogram | 240
no evidence of extravasation | 240
tortuous arteries in the lower pole | 240
embolized | 240
increasing in the abdominal distention | 240
dropping of hemoglobin | 240
symptomatic | 240
surgical intervention | 240
evacuate the hematoma | 240
capsulated mass around 30 cm | 240
bleeding around it | 240
radical nephrectomy | 240
bowel injury | 240
repaired primarily intraoperative | 240
post operatively | 240
chyle leak | 240
managed conservatively | 240
histopathology revealed the diagnosis of embryonal rhabdomyosarcoma | 240
tumor board | 240
planned for chemotherapy | 240
multiple peritoneal metastatic deposit | 240
liver and bone metastasis | 240
received first cycle of Dactinomycin, Vincristine, Cyclophosphamide | 240
complicated by sepsis | 240
pulmonary embolism | 240
profound neutropenia | 240
intensive care unit admission | 240
passed away 88 days post-operatively | 2088
disease progression | 2088