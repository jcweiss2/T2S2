78 years old | 0
    woman | 0
    presented to the emergency room | 0
    progressively worsening non-bloody diarrhea | -336
    approximately 5 bowel movements per day | -336
    left lower-quadrant dull abdominal pain | -72
    nausea | -72
    non-bloody vomiting | -72
    no fever | 0
    no headache | 0
    no cough | 0
    no shortness of breath | 0
    no jaw claudication | 0
    no joint pain | 0
    no visual disturbances | 0
    lived in Wisconsin | 0
    not travelled outside of the state recently | 0
    reported no sick contacts | 0
    immunized against COVID-19 with the Moderna mRNA vaccine | -2880
    past medical history: poorly controlled type 2 diabetes mellitus (A1C 8.4%) | 0
    hypertension | 0
    CKD 3b A2 | 0
    depression | 0
    hypertriglyceridemia | 0
    anemia with CKD | 0
    surgical history: bilateral cataract surgery | -87600
    compliant with her medications | 0
    could not take medications due to nausea and vomiting | -24
    aspirin 81 mg daily | -24
    atorvastatin 40 mg daily | -24
    famotidine 20 mg twice daily as needed | -24
    glargine insulin 18 units subcutaneous at bedtime | -24
    aspart insulin 20 units subcutaneous 3 times daily | -24
    metformin 1000 mg twice daily | -24
    metoprolol tartrate 25 mg twice daily | -24
    losartan 100 mg daily | -24
    torsemide 20 mg daily | -24
    sertraline 150 mg daily | -24
    denied recent medication changes | 0
    taken metformin since 2005 | -175200
    former smoker | 0
    denied history of alcohol use | 0
    denied illicit drug use |9 0
    family history negative for cerebrovascular disease | 0
    family history negative for vasculitides | 0
    temperature of 36.3°C | 0
    blood pressure 165/67 mmHg | 0
    heart rate 104 beats per minute | 0
    respiratory rate 16 breaths per minute | 0
    oxygen saturation normal on ambient air | 0
    alert | 0
    pale | 0
    no distress | 0
    pupils round | 0
    pupils equal 2–3 mm | 0
    reactive to light | 0
    reactive to accommodation | 0
    dry mucous membranes | 0
    heart sounds regular | 0
    tachycardia | 0
    no murmurs | 0
    no rubs | 0
    lungs clear to auscultation | 0
    mild tenderness to palpation of the left lower quadrant | 0
    no guarding | 0
    no rebound tenderness | 0
    normal neurological exam | 0
    leukocytosis 10.2×109/L | 0
    neutrophilia | 0
    lymphopenia | 0
    hemoglobin 10.6 g/dL | 0
    mild thrombocytosis 438×109/L | 0
    lactate 6.4 mmol/L | 0
    sodium 135 mmol/L | 0
    hypochloremia 86 mmol/L | 0
    hyperkalemia 6.2 mmol/L | 0
    anion gap elevated metabolic acidosis | 0
    bicarbonate 6 mmol/L | 0
    anion gap 43 | 0
    no osmolar gap | 0
    glucose 269 mg/dL | 0
    blood urea nitrogen 83 mg/dL | 0
    creatinine 8.47 mg/dL | 0
    baseline creatinine 1.2–1.4 mg/dL | 0
    normal liver transaminases | 0
    normal total bilirubin | 0
    creatine kinase 110 U/L | 0
    venous blood gas pH <6.80 | 0
    pCO2 17 mmHg | 0
    beta-hydroxybutyrate 1.8 mmol/L | 0
    SARS CoV-2 PCR test negative | 0
    urinalysis: no signs of infection | 0
    glucose 500 mg/dL | 0
    ketones 80 mg/dL | 0
    CT scan of the abdomen and pelvis without IV contrast | 0
    extensive colonic diverticula | 0
    inflammatory change in the fat around the descending colon | 0
    mild diverticulitis | 0
    no free air | 0
    no abscess collection | 0
    administered IV ceftriaxone | 0
    administered Flagyl | 0
    2 L NaCl 0.9% fluid bolus | 0
    300 mEq bicarbonate bolus | 0
    bicarbonate drip | 0
    repeat lactate increase to 9.6 mmol/L | 0
    imaging of the abdomen and pelvis with IV contrast | 0
    ruled out acute mesenteric ischemia | 0
    admitted to the Intensive Care Unit | 0
    insulin drip initiated | 0
    2-L NaCl 0.9% fluid bolus | 0
    confusion | 3
    lethargy | 3
    hypothermia 32.2°C | 3
    sudden painless bilateral vision loss | 3
    blood pressure stable | 3
    heart rate stable | 3
    pupils equal at 3–4 mm | 3
    no light pupillary reaction | 3
    absent blink to threat | 3
    normal remaining neurological exam | 3
    no change in abdominal exam | 3
    CT head negative for acute abnormalities | 3
    ophthalmology evaluation: preserved extraocular motility | 3
    no retinopathy | 3
    no macular edema | 3
    no acute glaucoma | 3
    no embolic phenomena | 3
    confirmed no pupillary reaction to light | 3
    confirmed absent blink to threat | 3
    cortical blindness considered | 3
    MRI of the brain revealed no acute abnormalities | 3
    ruled out acute stroke | 3
    repeated blood work 7 hours after initial presentation | 7
    worsening lactic acid of 14.2 mmol/L | 7
    sodium 138 mmol/L | 7
    hypochloremia 92 mmol/L | 7
    hyperkalemia 6.0 | 7
    bicarbonate <5 | 7
    anion gap unable to calculate | 7
    glucose 264 | 7
    venous blood gas pH 6.87 | 9
    pCO2 29 mmHg | 9
    worsening lactic acid of 16.1 | 9
    persistent metabolic disturbances | 9
    development of new neurologic deficit | 9
    suspected MALA with vision loss | 9
    initiated on emergent CRRT | 9
    hypotension | 9
    norepinephrine infusion initiated | 9
    TTE revealed preserved left ventricular ejection fraction | 9
    no segmental wall motion abnormalities | 9
    no intracardiac mass | 9
    no thrombus | 9
    ruled out cardiogenic etiology of shock | 9
    volatile serum screen: high acetone at 18 mg/dL | 9
    negative for methanol | 9
    negative for ethanol | 9
    negative for isopropanol | 9
    metabolic acidosis improved | 11
    vision started to improve | 11
    vision returned to baseline | 11
    mental status returned to baseline | 11
    hypothermia resolved | 11
    bicarbonate infusion discontinued | 11
    lactic acid normalized | 11
    insulin drip transitioned to subcutaneous insulin | 11
    weaned off norepinephrine within 7 hours | 11
    infectious diseases work-up: negative blood cultures | 11
    infectious diseases work-up: negative urine cultures | 11
    abdominal exam remained benign | 11
    no recurrence of diarrhea | 11
    empiric antibiotics discontinued | 48
    sepsis deemed unlikely | 48
    dialysis discontinued after 18 hours | 18
    creatinine improved to 2.93 mg/dL | 18
    hyperkalemia resolved | 18
    discharged home | 48
    adjusted insulin regimen | 48
    indefinite discontinuation of metformin | 48
    