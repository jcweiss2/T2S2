48 years old | 0
female | 0
non-alcoholic | 0
non-smoker | 0
cough | -168
generalized myalgia | -168
arthralgia | -168
fever | -168
temperature 36.9°C | 0
pulse 76/m | 0
blood pressure 132/78 mmHg | 0
oxygen saturation 96% | 0
body mass index 26 | 0
diffuse arthralgia | 0
myalgia | 0
no previous medical history | 0
no chronic diseases | 0
no previous treatment with any medication | 0
no previous medical family history | 0
elevated erythrocyte sedimentation rate | 0
elevated C-reactive protein level | 0
elevated creatine kinase levels | 0
nasopharyngeal swab confirmed COVID-19 | 0
mild disease | 0
mild pulmonary infiltrations | 0
hospitalized in COVID-19 isolation department | 0
confusion | 72
high fever 39.8°C | 72
tachycardia 125/m | 72
hypotension 75/40 mmHg | 72
Glasgow score 10/15 | 72
elevated White blood cells | 72
elevated erythrocyte sedimentation rate | 72
elevated C-reactive protein level | 72
elevated Creatine phosphokinase | 72
elevated myoglobin | 72
elevated Aspartate aminotransferase | 72
elevated Alanine aminotransferase | 72
elevated urea | 72
elevated creatinine | 72
treated with oxygen | 72
treated with intravenous normal saline | 72
treated with bicarbonate | 72
treated with epinephrine | 72
treated with azithromycin | 72
treated with methyl prednisone | 72
treated with enoxaparine | 72
intubated and mechanically ventilated | 72
dialysis therapy | 72
cardiac arrest | 96
death | 96