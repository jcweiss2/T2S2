57 years old | 0
male | 0
admitted to the hospital | 0
fever | -48
cough | -48
sputum | -48
dyspnea | -24
hypothermia (35.5°C) | 0
tachypnea (29 bpm) | 0
hypoxemia (SpO2 78%) | 0
tachycardia (118 bpm) | 0
blood pressure 115/50 mmHg | 0
bilateral lung moist rale | 0
arterial blood gas analysis hypoxygen (PaO2 68.8 mmHg) | 0
metabolic acidosis | 0
hyperlactatemia (7.09 mmol/L) | 0
white cell count 4.31 ×10^9/L | 0
neutrophil 88.2% | 0
platelet count 48 ×10^9/L | 0
hemoglobin 150 g/L | 0
C-reactive protein 295.92 g/L | 0
procalcitonin >200.00 ng/ml | 0
NT-proBNP >35000 pg/mL | 0
troponin T 40.76 pg/mL | 0
CK 2639.00 U/L | 0
CK-MB 63.00 U/L | 0
blood urea nitrogen 18.16 mmol/L | 0
creatinine 513.00 μmol/L | 0
total bilirubin 72.5 μmol/L | 0
alanine aminotransferase 41.00 U/L | 0
aspartate aminotransferase 88.00 U/L | 0
cholinesterase 3.97 U/mL | 0
septic shock | 0
multiple organ dysfunction syndrome (MODS) | 0
fluid resuscitation | 0
continuous renal replacement therapy | 0
organ protective therapy | 0
blood culture | 0
sputum culture | 0
empiric antibiotic therapy (piperacillin tazobactam and moxifloxacin) | 0
nasal intubation | 0
mechanical ventilation | 0
prone position ventilation | 0
Klebsiella pneumoniae culture positive | 72
antimicrobial susceptibility sensitive to piperacillin tazobactam | 72
hvKP confirmed (string test and wax moth larvae test) | 72
hypoxemia improved slightly | 72
airway secretion requiring bronchoscope suction | 72
hemodynamic instability | 72
norepinephrine 0.5-0.8 μg/kg/min | 72
second thoracic CT on day 10 | 240
lung consolidation in right upper lobe | 240
abscess formation | 240
CEUS performed on day 12 | 288
sulfur hexafluoride microbubble contrast agent | 288
CEUS-guided drainage with pigtail tube | 288
hypoxemia improvement | 336
hemodynamic improvement | 336
ventilator weaning on day 16 | 384
third thoracic CT on day 21 | 504
lung lesion improvement | 504
