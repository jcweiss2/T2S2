72 years old | 0
female | 0
cirrhosis caused by autoimmune hepatitis | 0
hepatic encephalopathy | 0
ascites | 0
admitted to the hospital | 0
bilious vomiting | -48
diffuse abdominal pain | -48
oliguria | -48
headache | -48
esophagogastroduodenoscopy showing gastritis | 0
grade IV esophageal varices | 0
nadolol | 0
spironolactone | 0
furosemide | 0
azathioprine | 0
esomeprazole | 0
lactulose | 0
temperature 36.06°C | 0
blood pressure 82/32 mm Hg | 0
pulse 92 beats/min | 0
lethargy | 0
bibasilar rales | 0
tender abdomen | 0
tense ascites | 0
no jaundice | 0
no lower extremity edema | 0
no focal neurological deficits | 0
white blood count 9,400 cells/mm3 | 0
bandemia | 0
macrocytic anemia | 0
thrombocytopenia | 0
hemoglobin 9.6 g/dl | 0
hematocrit 28.5% | 0
platelets 116,0000/μl | 0
MCV 115.9 fl | 0
INR 1.98 | 0
prothrombin time 16 s | 0
renal failure | 0
creatinine 5 mg/dl | 0
metabolic acidosis | 0
lactic acid 6.7 mmol/l | 0
serum ammonia 16 μmol/l | 0
sodium 128 meq/l | 0
potassium 5 meq/l | 0
chloride 101 meq/l | 0
bicarbonate 13 meq/l | 0
BUN 70 mg/dl |3c72
cirrhotic liver | 0
splenomegaly | 0
no ruptured viscus | 0
no obstruction | 0
large volume paracentesis | 0
serosanguinous ascitic fluid drained | 0
albumin concentration in fluid <1 mg/dl | 0
serum albumin 2.6 mg/dl | 0
