30 years old | 0
first pregnancy | 0
persistent nausea | -72
vomiting | -72
generalized abdominal pain | 0
abdominal distension | 0
moderate tenderness | 0
increased depth of palpation | 0
intravenous ceftriaxone | 0
limited ultrasound | 0
abdominal magnetic resonance imaging | 24
dilated loops of the colon | 24
sigmoid colon dilation | 24
fluid-gas levels | 24
tarry stools | 24
upper gastrointestinal bleeding | 24
gastroscopy | 24
rapid deterioration | 24
significant increase in inflammatory parameters | 24
symptoms of septic shock | 24
exacerbation of abdominal pain | 24
intravenous Meropenem | 24
intravenous Vancomycin | 24
intravenous Fluconazole | 24
midline laparotomy | 72
serous fluid | 72
large intestine dilation | 72
serosal membrane damage | 72
ruptures sutured | 72
appendectomy | 72
cecostomy | 72
safety drains | 72
acute intestinal pseudo-obstruction diagnosis | 72
respiratory insufficiency | 72
intubation | 72
mechanical ventilation | 72
enteral nutrition | 72
parenteral nutrition | 72
antibiotic therapy continued | 72
elevated inflammatory markers | 72
transferred to Intensive Care Unit | 72
transfer to Department of Surgery | 264
transfer to obstetrics ward | 312
delivered a healthy baby | 312
restore gastrointestinal continuity | 456
adhesions released | 456
completed treatment | 456
no further surgical interventions | 456
family doctor care | 456
