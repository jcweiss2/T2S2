24 years old | 0
female | 0
gravida 2 | 0
para 1 | 0
admitted to the hospital | 0
fever | -72
right low abdominal pains | -72
ovarian cyst | -672
dichorionic-diamniotic twin pregnancy | -672
increased fetal heart rate | -72
intrauterine hypoxia | -72
ascites | -72
WBC count 19.85×10^9/L | -72
neutrophils 84.9% | -72
C-reactive protein 20.22mg/L | -72
oral cephalosporin | -72
TORCH tests | -672
intrauterine death of one fetus | -24
transferred to our hospital | -24
temperature 36.6°C | -24
WBC count 22.14×10^9/L | -24
neutrophils 81.6% | -24
CRP 195.76mg/L | -24
intravenous injection of cefuroxime sodium | -24
intramuscular injection of dexamethasone sodium phosphate | -24
chest distress | -48
nasal cannula oxygen therapy | -48
supplement with calcium and potassium | -48
temperature 39.5°C | -24
blood pressure 105/59 mmHg | -24
WBC count 12.6×10^9/L | -24
RBC count 3.71×10^12/L | -24
hemoglobin 80g/L | -24
neutrophils 86.5% | -24
lymphocyte 6.8% | -24
Ca2+ 2.00mmol/L | -24
K+ 3.4mmol/L | -24
Na+ 134mmol/L | -24
albumin 29g/L | -24
BNP 175.0pg/mL | -24
blood culture | -24
chest Computed Tomography (CT) | -24
cardiac insufficiency | -24
pulmonary edema | -24
anti-infection with ampicillin-sulbactam | -24
caesarean section | 0
septic shock | 0
one alive fetus delivered | 0
Apgar score 8, 10, 10 | 0
one dead fetus | 0
amniotic fluid aeruginous | 0
uterus limp and feeble | 0
bilateral uterine artery ligation | 24
B-Lynch suture | 24
postpartum hemorrhage | 24
blood transfusion | 24
exploratory laparotomy | 24
Listeria monocytogenes infection identified | 96
blood culture result positive | 96
placenta tissue culture positive | 144
ampicillin-sulbactam continued | 0
patient discharged | 432
readmitted with fever | 1008
blood culture result negative | 1008
CT scan of the chest | 1008
brain MRI | 1008
newborn admitted to NICU | 24
neonatal dehydration | 24
premature and low birth weight infant | 24
suspected neonatal sepsis | 24
intracranial infection | 24
lumbar puncture | 24
cerebrospinal fluid examination | 24
aerobic cultures of whole blood and CSF | 24
brain MRI | 24
coagulation function disordered | 24
anti-infection and nutrition support | 24
condition deteriorated | 696
neonatal sepsis | 696
meropenem and immune globulin | 696
feeding refusal | 696
abdominal distension | 696
abdominal plain radiography | 696
potential neonatal necrotizing enterocolitis | 696
transferred to Department of Pediatric Surgery | 696