21 years old | 0
male | 0
presented to the hospital | 0
high-velocity motorcycle accident | -168
comminuted pelvic fractures | -168
multiple extremity fractures | -168
catastrophic degloving injury of the buttocks and perineum | -168
gross wound soilage | -168
vascular injuries | -168
bilateral iliac arteries angioembolization | -168
rapidly progressing necrotizing soft tissue infection | -168
polymicrobial infection | -168
Acinetobacter spp. | -168
Pseudomonas spp. | -168
Stenotrophomonas maltophila | -168
Trichosporon asahii | -168
Saksenaea spp. | -168
Fusarium spp. | -168
daily or alternating-day operative debridement | -168
broad-spectrum parenteral and topical antibacterial therapy | -168
broad-spectrum parenteral and topical antifungal therapy | -168
ceftazidime | -168
metronidazole | -168
trimethoprim-sulfamethoxazole | -168
micafungin | -168
amphotericin B | -168
posaconazole | -168
VERAFLO vac instillation | -168
multisystem organ failure | -168
shock | -168
debridement of >3000 cm2 of skin, subcutaneous tissue, and muscle | -168
perineum involvement | -168
bilateral thighs involvement | -168
buttocks involvement | -168
circumferential abdominal wall involvement | -168
persistently positive cultures for Trichosporon asahii | -168
persistently positive cultures for Saksenaea spp. | -168
invasive fungal elements on histopathological exam | -168
increased lymphocyte count | -168
persistent lymphopenia | -168
neutrophilia | -168
recombinant human IL-7 therapy initiation | 0
IL-7 administered (3 µg/kg) | 0
IL-7 dosage increased to 10 µg/kg | 24
significant clinical improvement | 96
slowed progression of invasive soft tissue necrosis | 96
improved wound healing | 96
healthier-appearing tissue margins | 96
improvement of fever curve | 96
improvement of tachycardia | 96
improvement of tachypnea | 96
progressive decreases in total white blood cell count | 96
increasing absolute lymphocyte counts | 96
absolute lymphocyte count increased to >4000 lymphocytes/µL | 96
persistently negative fungal cultures | 120
negative fungal tissue histology | 120
healthy granulation tissue development | 120
skin grafting | 120
negative blood cultures | 720
negative wound cultures | 720
negative bone cultures | 720
definitive closure of >90% of open wounds | 720
exposed pelvic bone | 720
persistent perineal wound | 720
urine drainage | 720
recent biopsy positive for Trichosporon asahii | 720
extended course of isavuconazonium | 720
increased number of activated IFN-γ-producing T cells | 96
increased proportion of activated T cells | 96
increased CD3+ T cells in wound margins | 96
increased pSTAT5 expression in CD4-T cells | 96
increased pSTAT5 expression in CD8-T cells | 96
informed consent obtained | 0
test dose of IL-7 well tolerated | 0
small region of exposed pelvic bone | 720
persistent perineal wound remains open | 720
pending reconstruction | 720
no recurrence of necrotizing fasciitis | 720
