86 years old | 0
female | 0
right hip replacement | -2880
altered mental status | 0
not feeling well | -48
respiratory distress | 0
tachycardia | 0
tachypnea | 0
dehydration | 0
no evidence of trauma | 0
rapid shallow respiration | 0
wheezing | 0
mild pedal edema | 0
WBC count 6.5 × 10^3 per µL | 0
normal differential count | 0
Hemoglobin 3.2 gm/dL | 0
hematocrit 9.6% | 0
MCV 127 fL | 0
platelets 59 × 10^3 per µL | 0
retic count 7.5% | 0
corrected retic 1.6% | 0
LDH 7077 IU/L | 0
haptoglobin very low | 0
severe metabolic acidosis | 0
high anion gap | 0
renal functions impaired | 0
BUN 34 mg/dL | 0
creatinine 1.9 mg/dL | 0
serum glucose 93 mg/dL | 0
osmolality 308 mOsm/L | 0
lactic acid 20.3 mmol/L | 0
hyperbilirubinemia | 0
total bilirubin 3.7 mg/dL | 0
direct bilirubin 1 mg/dL | 0
aspartate transaminase 51 IU/L | 0
alanine transaminase 22 IU/L | 0
alkaline phosphatase 41 IU/L | 0
BNP 670 pg/mL | 0
troponin negative | 0
INR elevated | 0
PT 29 s | 0
aPTT 24 s | 0
toxicology screen negative | 0
mild cardiomegaly | 0
CT head negative | 0
CT abdomen negative | 0
CT PE protocol negative | 0
intubated | 0
intravenous antibiotics | 0
blood transfusion | 0
received 3 units of blood | 0
improved significantly after blood transfusion | 10
lactic acid normalized | 10
antibiotics discontinued | 10
acute kidney injury resolved | 10
mentation improved | 10
weaned off ventilator | 48
fecal occult blood tests negative | 48
ferritin 588 ng/mL | 48
TIBC 194 µg/dL | 48
transferrin 155 mg/dL | 48
iron saturation 91% | 48
peripheral smear showed large RBCs | 48
hypersegmented neutrophils | 48
schistocytes | 48
poikilocytes | 48
anisocytosis | 48
mixed picture of megaloblastic anemia and hemolytic anemia | 48
vitamin B12 38 pg/mL | 48
methylmalonic acid 753 nmol/L | 48
homocysteine 99.3 µmol/L | 48
anti-parietal antibodies 21.7 units | 48
anti-intrinsic factor antibodies 4.7 AU/mL | 48
direct Coombs test negative | 48
indirect Coombs test negative | 48
fibrinogen 185 mg/dL | 48
D-dimer 5170 ng/mL | 48
serology negative for HIV and hepatitis virus | 48
diagnosed with pernicious anemia | 48
diagnosed with pseudo-TTP | 48
started on parenteral vitamin B12 | 48
hematological parameters improved | 120
clinical condition improved | 120
discharged | 120