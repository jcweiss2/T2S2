61 years old | 0
male | 0
presented to the emergency department | 0
pleuritic chest pain | 0
pulmonary vein isolation (PVI) by cryothermal ablation | -240
paroxysmal atrial fibrillation | -240
diabetes mellitus | 0
hypertension | 0
atrial fibrillation | 0
treated with empagliflozin | 0
treated with dabigatran | 0
treated with bisoprolol | 0
pericardial friction rub | 0
diffuse ST-elevation | 0
PR depression | 0
troponin levels within normal limits | 0
preserved ventricular function | 0
small to medium circumferential pericardial effusion | 0
hospitalized | 0
presumptive diagnosis of pericarditis | 0
treated with prednisone | 0
treated with colchicine | 0
clinical improvement | 0
discharged | 96
presented to the emergency department again | 144
severe weakness | 144
fatigue | 144
syncopal episode | 144
blood-tinted vomitus | 144
pleuritic chest pain | 144
blood pressure 80/50 mmHg | 144
temperature 38.5°C | 144
oxygen saturation 96% | 144
haemoglobin 11.2 gr/dL | 144
mild neutrophilia 9.23 103/uL | 144
creatinine 1.72 mg/dL | 144
urea 114.1 mg/dL | 144
troponin levels normal | 144
nasogastric tube inserted | 144
coffee-ground matter drainage | 144
no active bleeding | 144
TTE showed no differences from previous study | 144
presumptive diagnosis of mediastinitis due to AOF | 144
received intravenous fluids | 144
received norepinephrine | 144
received amoxicillin clavulanate | 144
received fluconazole | 144
non-gated CT angiography | 144
multiple mediastinal lymph nodes | 144
small amount of fluid in mediastinum | 144
small amount of fluid in pericardium | 144
no extravasation of contrast medium | 144
no pneumomediastinum | 144
no pneumopericardium | 144
brain CT showed no focal lesion | 144
developed multiorgan failure | 168
haemoglobin declined to 9.7 mg/dL | 168
creatinine rose to 1.83 mg/dL | 168
intubated | 168
mechanically ventilated | 168
no definitive proof of AOF | 168
third TTE | 168
same amount of pericardial effusion | 168
preserved biventricular function | 168
no air in cardiac cavities | 168
injection of agitated saline through nasogastric tube | 168
bubbles appeared in left atrium | 168
bubbles appeared in left ventricle | 168
diagnosis of atrial–oesophageal fistula (AOF) | 168
transferred to operating room | 168
surgical repair of left atrium necrotic rupture | 168
gastroscopy performed | 168
12 mm tear in low oesophagus | 168
closed with endoclips | 168
postoperative high-grade fever | 168
postoperative haemodynamic instability | 168
treated with meropenem | 168
treated with micafungin | 168
positive polymicrobial pleural fluid cultures | 168
discharged after 30 days | 720
deceased | N/A
