24 years old | 0
female | 0
severe headache | -72
projectile vomiting | -72
no fever | -72
no convulsions | -72
no focal neurological deficit | -72
symptomatic treatment | -72
admission to hospital | 0
provisional diagnosis of metabolic encephalopathy | 0
symptomatic treatment | 0
altered sensorium | 12
Glasgow Coma Scale-9 | 12
high-grade fever | 12
chills | 12
dyselectrolytemia | 12
low serum phosphate | 12
neutrophilic leukocytosis | 12
empirical treatment with ceftriaxone | 12
Gram stain of CSF | 12
polymorphs and lymphocytes in CSF | 12
Gram-positive bacilli in CSF | 12
culture of CSF | 24
L. monocytogenes in CSF | 24
blood culture | 0
Gram-positive bacilli in blood culture | 0
L. monocytogenes in blood culture | 24
switch to meropenem | 24
clinical improvement | 48
microbiological improvement | 48
discharge | 120