15 years old | 0
female | 0
acute myelogenous leukemia | -1008
standard induction treatment | -1008
2 cycles of chemotherapy | -1008
pancytopenia | -504
broad anti-infective treatment | -504
ciprofloxacin | -504
linezolid | -504
meropenem | -504
tobramycin | -504
liposomal amphotericin | -504
admitted to the pediatric intensive care unit | 0
tachycardia | -24
hypotension | -24
lactic acidosis | -24
transthoracic echocardiography | 0
severely impaired left ventricular ejection fraction | 0
electrocardiogram | 0
sinus tachycardia | 0
incomplete right bundle branch block | 0
N-terminal prohormone of brain natriuretic peptide | 0
high-sensitive troponin T | 0
fluid therapy | 0
noradrenaline | 0
dobutamine | 0
milrinone | 0
deep sedation | 0
mechanical ventilation | 0
respiratory insufficiency | 0
va-ECMO | 0
cannulation of the left femoral artery and vein | 0
va-ECMO blood flow | 0
extracorporeal blood flow | 0
mean arterial pressure | 0
noradrenaline | 0
vasopressin | 0
levosimendan | 0
hydrocortisone | 0
continuous venovenous hemodiafiltration | 0
anti-infective therapy | 0
meropenem | 0
ciprofloxacin | 0
metronidazole | 0
cotrimoxazole | 0
liposomal amphotericin B | 0
acyclovir | 0
linezolid | 0
vancomycin | 0
procalcitonin | 0
C-reactive protein | 0
leukocytes | 0
high-sensitive troponin T | 0
creatine kinase MB | 0
total creatine kinase | 0
microbial specimens | 0
viral myocarditis | 0
myocardial biopsy | 0
second day with va-ECMO | 24
mean arterial blood pressure | 24
LVEF | 24
levosimendan infusion | 24
acute ischemic injury | 24
right femoral artery | 24
Dacron conduit | 24
second arterial cannula | 24
ECMO circuit | 24
Y-connector | 24
ECBF | 24
venous drainage pressures | 24
inspiratory oxygen fraction | 24
harlequin syndrome | 24
arterial oxygen partial pressure | 24
broad-complex tachycardia | 48
esmolol | 48
metoprolol | 48
left ventricular function | 48
aortic valve | 48
pulmonary edema | 48
intracardiac clot formation | 48
second venous cannula | 48
left atrium | 48
percutaneous atrioseptostomy | 48
catheter lab | 48
ECBF | 48
lactate levels | 48
mean arterial pressure | 48
cerebral oximetry | 48
near infrared spectroscopy | 48
regional oxygen saturation | 48
unfractionated heparin | 48
partial thrombin time | 48
PCT | 72
CRP | 72
leukocytes | 72
high-sensitive troponin T | 72
creatine kinase MB | 72
total creatine kinase | 72
day 5 | 120
ECMO cannulas | 120
left femoral vessels | 120
day 7 | 168
ECMO | 168
operating theater | 168
LVEF | 168
mean arterial pressures | 168
transseptal cannula | 168
CVVHDF | 168
renal function | 168
leucocyte count | 168
day 13 | 312
day 30 | 720
respirator weaning | 792
day 33 | 792
allogenic stem cell transplantation | 1008
6 weeks later | 1008
rehabilitation facility | 1008
critical illness | 1008
polyneuropathy | 1008
LVEF | 1008
ventricular dilatation | 1008