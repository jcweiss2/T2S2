11 years old | 0
girl | 0
presented to her primary care physician with concern for pallor of the lips | 0
variable duration episodes (minutes to days) | 0
episodes not associated with obvious trigger | 0
no fever | 0
no illness | 0
no dizziness | 0
no fatigue | 0
low free T4 | 0
normal TSH | 0
referral to endocrinology | 0
uncomplicated full-term gestation | -105120
delivery by emergency cesarean section | -105120
fetal distress | -105120
maternal fever of 104°F | -105120
2-week neonatal intensive care unit stay | -105120
rule out sepsis | -105120
received phototherapy for hyperbilirubinemia | -105120
family history negative for sudden death | -105120
unremarkable developmental history | -105120
past medical history notable for several urinary tract infections prior to 1 year of age | -105120
prolonged hospitalization at age 5 for septic shock and multi-organ dysfunction | -105120
presented to emergency department at age 5 with nausea | -52560
vomiting | -52560
diarrhea | -52560
fever | -52560
abdominal pain | -52560
hypotension | -52560
tachycardia | -52560
tachypnea | -52560
admitted for presumed gastroenteritis | -52560
intravenous fluid resuscitation | -52560
rule out sepsis | -52560
cultures drawn | -52560
empiric ceftriaxone provided | -52560
became unresponsive | -52560
intubated | -52560
hypoglycemia | -52560
received multiple dextrose 25% boluses without significant improvement | -52560
transferred to another facility for higher level of care | -52560
5-week PICU stay | -52560
received broad-spectrum antibiotics | -52560
intravenous fluids | -52560
pressor support | -52560
hypotension persisted | -52560
developed acute renal failure requiring dialysis | -52560
high-dose intravenous glucocorticoids initiated | -52560
clinical findings improved | -52560
hospitalized at age 6 for observation | -52560
febrile illness | -52560
sore throat | -52560
dry cough | -52560
temperature 102.5°F | -52560
blood pressure 114/69 mm Hg | -52560
temperature spiked to 105°F | -52560
blood, urine, throat, and stool cultures obtained | -52560
started on empiric antibiotic therapy | -52560
no hospitalizations or health concerns for next 5 years | -52560
onset of episodic lip pallor | -52560
initial endocrinology evaluation | 0
reports dry skin | 0
denies cold intolerance | 0
denies constipation | 0
denies fatigue | 0
denies weakness | 0
denies recent change in weight | 0
well appearing | 0
weight at 70th percentile | 0
height at 60th percentile | 0
growth records showing plateau over previous 6 months | 0
mid-parental height at 10th percentile | 0
mildly delayed deep tendon reflexes | 0
Tanner stage B3PH1 | 0
thyroid gland not enlarged | 0
no proximal muscle weakness | 0
mildly elevated TSH | 0
low IGF-binding protein-3 | 0
low IGF-1 ECL | 0
low estradiol | 0
undetectable early morning cortisol | 0
low peak cortisol post ACTH | 0
elevated prolactin serum | 0
non-elevated titers of thyroid peroxidase antibodies | 0
non-elevated titers of thyroglobulin antibodies | 0
bone age not skeletally mature | 0
predicted adult height 62.8 inches | 0
ectopic posterior pituitary gland | 0
severely hypoplastic and anteriorly displaced pituitary stalk | 0
diagnosis of central hypothyroidism | 0
panhypopituitarism due to PSIS | 0
hydrocortisone started | 0
thyroid hormone replacement initiated | 24
estrogen provided via oral contraceptive | 0
growth hormone treatment | 0
no significant illnesses or emergency visits | 0
responded well to growth hormone treatment | 0
initial annualized growth velocity 7.2 cm/year | 0
first-year height gain 6.8 cm | 0
final height 5’7” | 0
developed hypertension | 0
acute tubular injury | 0
history of hypotensive crisis | 0
well-managed with low-dose lisinopril | 0
