42 years old | 0
male | 0
Brazilian | 0
alcohol withdrawal | 0
altered mental status | 0
chronic alcohol abuse | -672
chronic cocaine abuse | -672
admitted to the medical floors | 0
elevated heart rate | 0
elevated blood pressure | 0
hypoxic | 0
agitation | 0
expiratory wheezes | 0
elevated WBC count | 0
elevated serum creatinine | 0
positive urine drug screen for cocaine | 0
elevated blood alcohol level | 0
CT scan of the head without contrast | 0
normal CT scan of the head | 0
possible right small pleural effusion | 0
Chest X-ray | 0
CT pulmonary angiogram | 0
moderate hiatal hernia | 0
mild debris in the left main stem bronchus | 0
aspiration pneumonia | 0
started on CIWA protocol | 0
started on antibiotics | 0
started on oxygen supplementation | 0
COVID-19 test | 0
negative COVID-19 test | 0
coffee ground vomitus | 0
started on IV Protonix | 0
gastroenterology department consultation | 0
no active bleeding | 0
normal hemoglobin value | 0
worsening mental status | 24
transferred to the intensive care unit | 24
worsening delirium tremens | 24
respiratory distress | 24
increasingly hypoxic | 24
decreased breath sounds on the right side of the chest | 24
repeat CXR | 24
large right-sided pleural effusion | 24
thoracic surgery consultation | 24
insertion of the right inferior chest thoracostomy tube | 24
draining of dark fluid | 24
exudative effusion | 24
likely empyema | 24
fluid cultures positive for Candida Albicans | 48
infectious diseases department consultation | 48
switched to meropenem and vancomycin | 48
added antifungal agent micafungin | 48
transferred to the medical floor | 48
worsening agitation | 72
admitted to the ICU | 72
treated with lorazepam infusion | 72
persistently febrile | 72
leukocytosis | 72
repeat CT scan of the chest | 72
multiple right-sided loculated pleural effusions | 72
air-fluid levels | 72
no growth in blood cultures | 72
thoracic surgery department consultation | 72
poor surgical candidate | 72
high risk of operative complications | 72
insertion of two chest tubes | 96
removal of initially inserted chest tube | 96
draining of pus | 96
draining of purulent fluid and air | 96
pleural fluid cultures showed candida and staphylococcus epidermidis | 96
fluid analysis suggestive of empyema | 96
changed antibiotic regimen to meropenem, vancomycin, and fluconazole | 96
insertion of 3rd chest tube | 120
increased effusion size in basilar portion of right lung | 120
removal of two upper chest tubes | 120
switched meropenem to ampicillin-sulbactam | 120
improved mental status | 360
started oral feeding | 360
repeat CT chest showed empyema on the right side | 360
moderate left pleural effusion | 360
food contents in chest tube | 360
high chest tube output | 360
contrast esophagogram showed leak from right side of distal esophagus | 360
preferential passage of contrast into right pleural space | 360
gastroenterology and thoracic surgery departments consultation | 360
decision to proceed with feeding tube placement and esophageal stent insertion | 360
percutaneous endoscopic gastrostomy (PEG) | 672
endoscopic findings confirmed esophageal defect | 672
endoscopic esophageal stent placement | 672
stopped vancomycin | 672
switched to ampicillin-sulbactam | 672
completed fluconazole treatment after discharge | 720