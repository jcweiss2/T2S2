80 years old | 0
    male | 0
    consulted to the urology department | 0
    scrotal mass suspected to be an abscess | 0
    history of urethral catheter replacement every 2 weeks for 4 months | -4320
    urinary retention | -4320
    purulent discharge from left scrotal wall | -120
    fever | -120
    urethral catheter replaced one day before admission | -24
    pain | -24
    lump on the left scrotum | -24
    referred to Hasan Sadikin Hospital | -24
    blood pressure 90/60 mmHg | 0
    heart rate 120 beats per minute | 0
    respiratory rate 24 times per minute |7 0
    body temperature 37.5 °C | 0
    lump in the left scrotum | 0
    cystic on palpation | 0
    pus coming out from the left scrotum | 0
    purulent fluid inside the urethral catheter tube | 0
    scrotal ultrasound examination revealed balloon catheter in the left scrotum | 0
    hyperechoic lesion with acoustic shadow in the posterior urethra | 0
    KUB x-ray showed two radio opaque shadows in the pelvic area | 0
    white blood cell count 19.790 WBC/mL | 0
    hemoglobin 7.8 g/dL | 0
    serum BUN 103.14 mg/dL | 0
    serum creatinine 5.29 mg/dL | 0
    serum lactate 2.1 | 0
    blood glucose level 114 mg/dL | 0
    urinalysis >50/hpf red blood cells | 0
    urinalysis >50/hpf white blood cells | 0
    Fournier Gangrene Scoring Index 18 points | 0
    correction of fluid and electrolyte imbalance | 0
    third generation cephalosporin | 0
    emergency necrotomy debridement | 0
    retrograde urethrography showed contrast extravasation at the pendulare area | 0
    open vesicolithotomy performed | 0
    two stones extracted from bladder and urethra | 0
    bladder stone size 45x20x15 mm | 0
    urethral stone size 20x18x12 mm | 0
    cystostomy tube inserted | 0
    incision drainage | 0
    necrotomy debridement of the scrotum | 0
    5 cm defect on the urethra | 0
    level of consciousness E3M6V4 | 0
    white cell count 16000 WBC/mL | 0
    hemoglobin 9.5 g/dL | 0
    serum BUN 67.2 mg/dL | 0
    serum creatinine 2.4 mg/dL | 0
    shortness of breath | 48
    consulted to the internal medicine department | 48
    diagnosed with hospital-acquired pneumonia | 48
    respiratory problem worsened | 72
    intubated | 72
    moved to the ICU | 72
    patient's condition not improved | 72
    died due to respiratory failure | 72
    