22 years old | 0
male | 0
MADD | -0
born | -7920
parents healthy | -7920
parents first cousins | -7920
three older siblings died | -7920
suffered from MADD | -7920
one younger sibling suffered from MADD | -7920
two younger siblings did not suffer from MADD | -7920
genetic counseling | -7920
prenatal diagnostic testing | -7920
DNA sequencing | -7920
homozygous c.1074G > C variant | -7920
ETF dehydrogenase | -7920
arginine substitution | -7920
myristate oxidation reduction | -7920
standard treatment | 0
diet | 0
riboflavin supplements | 0
L-carnitine supplements | 0
numerous crises of hypoglycemia | -0
metabolic decompensation | -0
trivial infections | -0
intravenous glucose | -0
acute kidney failure | -0
acute respiratory distress syndrome | -0
hemodialysis | -0
assisted ventilation | -0
full recovery | -0
routine exams | 0
moderate liver steatosis | 0
lipid storage myopathy | 0
mild exercise intolerance | 0
muscle weakness | 0
muscle pain | 0
elevated plasma-creatine kinase | 0
acyl-carnitine profile | 0
normal free carnitine | 0
increased acyl-carnitines | 0
hospitalized with acute hypoglycemia | -720
metabolic acidosis | -720
intestinal Clostridium difficile infection | -720
intravenous glucose | -720
antibiotics | -720
recovered | -720
hospitalized again | -576
acute hypoglycemia | -576
metabolic acidosis | -576
recurrent CDI | -576
treated with glucose | -576
antibiotics | -576
recovered | -576
hospitalized again | -432
abdominal pain | -432
CT scan | -432
enlarged spleen | -432
normal liver | -432
fecal microbiota transplantation | -432
septicemia | -288
staphylococcal bacteria | -288
treated with glucose | -288
antibiotics | -288
recovered | -288
hospitalized again | -168
progressive abdominal pain | -168
bloating | -168
mushy stools | -168
jaundiced | -168
febrile | -168
abdomen distended | -168
prolonged coagulation | -168
elevated transaminases | -168
elevated bilirubin | -168
impaired synthesis function | -168
acute necrosis of liver cells | -168
CT scan | -168
cirrhotic-looking liver | -168
parenchymal micro-abscesses | -168
liver decompensation | -168
ascites | -168
rectal portosystemic shunt | -168
splenomegaly | -168
severe colitis | -168
no stigmata of chronic liver disease | -168
negative hepatitis tests | -168
unchanged amino acids | -168
unchanged acylcarnitines | -168
ultrasound images | -168
CT angiography | -168
patent vessels | -168
no biliary dilatation | -168
severe portal hypertension | -168
hepato-fugal portal venous flow | -168
liver biopsy | -168
parenchymal damage | -168
macro-vesicular steatosis | -168
micro-vesicular steatosis | -168
glycogen accumulation | -168
copper accumulation | -168
Mallory bodies | -168
cirrhotic liver | -168
no malignancy | -168
no infection | -168
rapidly deteriorating liver function | -168
died | 0
intensive care unit | 0
acute liver failure | 0
no liver transplant surgery | 0
no trans-jugular intrahepatic portosystemic shunt | 0
family declined autopsy | 0