21 years old | 0
male | 0
blunt abdominal trauma | -72
major liver laceration | -72
liver packing | -72
received 20 units of packed red blood cells | -72
received fresh frozen plasma | -72
transferred to the Armed Forces Hospital | -24
required more blood | -24
required more fresh frozen plasma | -24
continued to bleed from the site of the liver laceration | -24
underwent emergency right hepatectomy | -24
intubated with mechanical ventilation | 0
in intensive care unit | 0
pneumothorax | 24
sepsis | 24
bed sores | 24
renal failure | 24
coagulopathy | 24
cardiac arrest | 360
deranged liver enzymes | 0
abnormal liver function | 0
abdominal distension | 0
drain of bile from the abdominal drainage | 0
endoscopic retrograde cholangiopancreatography | 72
major bile leak from one of the main branches of the left main bile duct | 72
10 Fr 5 cm plastic stent inserted | 72
sphincterotomy not performed | 72
improvement in abdominal distension | 168
improvement in bile drainage | 168
improvement in liver function | 168
abdominal distension | 504
deranged liver chemistry | 504
high bilirubin | 504
high alkaline phosphate | 504
second ERCP | 504
stent replacement | 504
major leak from the right hepatic duct stump | 504
plastic stent removed | 504
leaking bile branch selectively cannulated | 504
metallic endovascular coil deployed | 504
injection of NBCA and lipidol | 504
improvement in liver enzymes | 528
improvement in bile drainage | 528
discharged home | 720
endovascular coil remained in place | 2160
abdominal pain | 4320
low grade fever | 4320
mild elevation in liver enzymes | 4320
preserved liver function | 4320
CT abdomen revealed mildly dilated CBD | 4320
radio-opaque object most likely migrated endovascular coil | 4320
treated with antibiotics | 4320
ERCP performed | 4332
CBD found to be patent | 4332
most likely passed the endovascular coil | 4332