53 years old | 0
male | 0
rheumatoid arthritis | -8760
methotrexate | -8760
prednisolone | -8760
dog bite | -96
fever | -72
dyspnea | -72
admitted to primary care physician | -72
diagnosed as viral infection | -72
discharged home | -72
symptoms worsened | -48
transferred to emergency department | -48
admitted to hospital | 0
bite wound | 0
no signs of cellulitis | 0
no signs of erythema | 0
blood pressure 63/52 mmHg | 0
heart rate 129 beats/min | 0
respiratory rate 40/min | 0
body temperature 38.0 ° Celsius | 0
oxygen saturation 100% | 0
pancytopenia | 0
high-grade inflammatory status | 0
renal impairment | 0
coagulation studies showed prolonged prothrombin time-international normalized ratio | 0
coagulation studies showed increased fibrin/fibrinogen degradation products | 0
septic shock | 0
disseminated intravascular coagulation | 0
ground-glass opacity with consolidation in bilateral lower lobes | 0
blood samples collected for culture analysis | 0
transferred to intensive care unit | 0
massive fluid replacement | 0
administered meropenem | 0
platelet transfusion | 0
nafamostat mesilate | 0
noradrenaline | 0
hydrocortisone | 0
hypotension | 24
respiratory condition worsened | 24
repeat CT showed progression of consolidations | 24
acute respiratory distress syndrome | 24
mechanical ventilation | 24
GNR isolated from blood cultures | 24
pupillary dilation | 72
no light reflex | 72
cerebral hemorrhage | 72
cerebral herniation | 72
died | 120
slow-growing GNR subcultured | 120
grew well on sheep blood agar plates | 120
positive for catalase and oxidase | 120
multiple rods within cytoplasm of neutrophils | 120
identified as C. canimorsus | 120
sensitive to carbapenems | 120
sensitive to macrolides | 120
sensitive to β-lactam drugs | 120
sensitive to penicillin G | 120