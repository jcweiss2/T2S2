24 years old | 0
    male | 0
    admitted to the hospital | 0
    fever | -72
    cough | -72
    fatigue | -72
    blood in nasopharynx | 0
    no oral injury | 0
    no urinary incontinence | 0
    no bowel incontinence | 0
    no neck stiffness | 0
    vomited coffee ground emesis | 0
    hematemesis | 0
    oxygen saturation 99% | 0
    blood pressure 126/84 mmHg | 0
    temperature 39.4°C | 0
    deteriorated consciousness | 0
    intubated | 0
    normal chest X-ray | 0
    severe deranged liver function | 0
    SARS-CoV-2 positive | 0
    started on chloroquine | 0
    started on azithromycin | 0
    started on oseltamivir | 0
    started on tocilizumab | 0
    received acetylcysteine infusion | 0
    received lactulose | 0
    received vitamin K | 0
    received rifaximin | 0
    received pantoprazole | 0
    received 4F-PCC | 0
    received fresh frozen plasma | 0
    received fibrinogen | 0
    started on sustained low-efficiency dialysis | 0
    no intracranial hemorrhage | 0
    normal brain parenchyma | 0
    no hydrocephalus | 0
    no midline shift | 0
    no mass effect | 0
    liver normal size | 0
    coarse liver parenchyma | 0
    no liver foci | 0
    patent common bile duct | 0
    spleen normal size | 0
    kidneys normal size | 0
    fluctuating temperature | 0
    disseminated intravascular coagulation | 0
    bleeding from IV site | 0
    bleeding from endotracheal tube | 0
    multiorgan failure | 240
    acute liver failure | 240
    acute renal failure | 240
    death | 240
    