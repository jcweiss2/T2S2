68 years old | 0
    male | 0
    admitted to the hospital | 0
    abdominal pain | -168
    chronic inflammation of the lungs | 0
    thickening of the lower esophageal wall | 0
    enlarged mediastinal lymph nodes | 0
    esophageal malignancy | 0
    radical surgery for esophageal carcinoma | 264
    pathological mitosis in the tumor cells | 264
    tumor infiltration to the deep muscular layer | 264
    cancer metastasis in periesophageal lymph nodes (4/6) | 264
    no nerve invasion | 264
    positive expression of p40 | 264
    positive expression of CK5/6 | 264
    positive expression of EGFR | 264
    positive expression of p53 | 264
    negative expression of CK7 | 264
    negative expression of p16 | 264
    negative expression of CD34 | 264
    negative expression of S-100 | 264
    stage IIIa moderately differentiated ulcerative esophageal squamous cell carcinoma (T2N1M0) | 264
    high fever (38.3°C) | 300
    dyspnea | 300
    blood pressure 80/50 mmHg | 300
    clean and dry neck wound | 300
    white blood cells 34.38 × 10^9/L | 300
    neutrophils 95.7% | 300
    C-reactive protein 207.26 mg/L | 300
    procalcitonin >100 ng/mL | 300
    urinary leukocytes 62.20/µL | 300
    leukocytes per high-power field 11.20 | 300
    increased exudative lesions in both lungs | 300
    postoperative changes in the esophagus | 300
    sepsis | 300
    severe septic shock | 300
    meropenem administration | 300
    E. fergusonii bacteremia | 300
    sensitive to cefuroxime | 300
    sensitive to cefuroxime axetil | 300
    sensitive to ceftazidime | 300
    sensitive to ceftriaxone | 300
    sensitive to cefepime | 300
    sensitive to cefoxitin | 300
    sensitive to amoxicillin–clavulanic acid | 300
    sensitive to piperacillin–tazobactam | 300
    sensitive to cefoperazone–sulbactam | 300
    sensitive to imipenem | 300
    sensitive to ertapenem | 300
    sensitive to amikacin | 300
    sensitive to tigecycline | 300
    sensitive to cotrimoxazole | 300
    fever subsided | 312
    clinical indicators improved | 312
    negative blood culture | 552
    recovered | 336
    discharged | 336
    postoperative adjuvant radiation therapy | 1440
    