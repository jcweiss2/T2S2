43 years old | 0
male | 0
diabetes mellitus | 0
hypertension | 0
COVID-19 infection | -120
recovered from COVID-19 | -120
blurred vision | -120
impaired vision | -120
retro-orbital pain | -90
denies diplopia | 0
denies scalp tenderness | 0
denies weight loss | 0
denies jaw claudication | 0
treated with IV methylprednisolone | -60
treated with oral corticosteroid therapy | -60
transient relief of symptoms | -30
recurrence of symptoms | 0
visual acuity 6/36 | 0
visual acuity 6/6 | 0
impaired abduction | 0
impaired upward movement | 0
Humphrey Visual Field testing | 0
RAPD | 0
brisk reflex | 0
blurred disc margin | 0
flat retina | 0
hematocrit 42% | 0
white blood cell count 14,500/uL | 0
erythrocytes sedimentation rate 31 mm/h | 0
MRI of brain and orbits | -120
optic neuritis | -120
T2W hyper-intense signal foci | -120
mild post-contrast enhancement | -120
inflammatory changes | -120
treated with IV methylprednisolone | 0
improvement in visual acuity | 30
recurrence of pain and vision impairment | 60
no light perception | 60
initiation of prednisolone | 60
orbital MRI | 62
heterogeneously enhancing lesion | 62
encasing and compressing optic nerve | 62
focal asymmetric enhancement | 62
paranasal CT scan | 64
heterogeneously enhancing soft tissue | 64
widening of canal | 64
extension into sphenoid sinus | 64
excision biopsy | 66
histopathological examination | 66
PAS stain | 66
aspergillosis | 66
yellowish-white tissue | 66
purulent discharge | 66