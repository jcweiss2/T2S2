60 years old | 0
male | 0
injured in a motor-vehicle accident | -96
4th to 9th right side rib fractures | -96
bilateral pneumothorax | -96
left hip dislocation | -96
fractures of spinous processes of 5th to 8th thoracic vertebrae | -96
obese | 0
BMI = 39 kg/m2 | 0
quit smoking | -8760
left lower lobectomy for carcinoid | -8760
admitted to regional hospital | -96
thoracic cavity drained | -96
hip dislocation reduced | -96
general anaesthesia | -96
mechanical ventilation dependence | -96
transferred to ICU | 0
respiratory insufficiency | 0
haemodynamic instability | 0
acute renal failure | 0
haemodialysis | 0
massive SE of face, neck, thoracic and abdominal wall | 0
CT scans | 0
persistent bilateral pneumothorax | 0
pneumomediastinum | 0
pneumoperitoneum | 0
subcutaneous emphysema extending to the pelvis | 0
thoracic drains replaced | 0
continuous venovenous haemodiafiltration | 0
septic | 0
multi-resistant Acinetobacter baumanii isolated | 0
Bilevel positive airway pressure mode of mechanical ventilation | 0
high inspiratory airway pressure | 0
high positive end-expiratory pressure | 0
low dynamic compliance | 0
respiratory status deteriorated | 120
high inspired oxygen fraction | 120
control CT | 120
surgical decompression | 120
subclavicular blowhole incisions | 120
NPWT dressing applied | 120
swift regression of SE | 132
improvement in ventilatory parameters | 132
transition to pressure support mode of mechanical ventilation | 132
NPWT dressing removed | 192
wounds sutured | 192
surgical tracheostomy | 192
weaned off ventilator | 240
renal function improved | 240