69 years old| 0
male| 0
admitted to the intensive care unit| 0
septic shock| 0
bloody diarrhea| -504
hypertension| 0
cardiomyopathy| 0
chronic obstructive pulmonary disease| 0
laryngeal carcinoma (T3N0)| 0
amoxicillin/clavulanic acid| -1344
laryngitis| -1344
confused mental state| 0
hypotension (77/28 mmHg)| 0
temperature (35.6°C)| 0
diffuse abdominal tenderness| 0
increased leucocytes (38.9 × 10^9/l)| 0
increased C-reactive protein (318 mg/l)| 0
renal insufficiency (creatinine 534 umol/l)| 0
low albumin (23 g/l)| 0
normal lactate (1.6 mmol/l)| 0
broad-spectrum antibiotics| 0
abdominal CT-scan (diffuse colonic wall thickening)| 0
C. difficile isolated (PCR-ribotype 001)| 0
severe CDI diagnosis| 0
oral vancomycin| 0
metronidazole intravenously| 0
vasopressor support dependence| 216
progressive abdominal distension| 216
delirium| 216
metabolic acidosis| 216
surgical consultation for colectomy| 216
FMT consideration| 216
FMT delivered via nasoduodenal tube| 288
vancomycin stopped| 276
metronidazole stopped| 276
fidaxomicin started| 276
fidaxomicin continued| 288
abdominal distension decrease| 360
C. difficile negative on PCR| 360
fidaxomicin continued until nine days post-FMT| 432
discharged from ICU| 432
no recurrent CDI| 432
