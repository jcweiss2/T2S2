19 years old | 0
male | 0
gunshot wound to the right temporal region | 0
recreational drug use | 0
alcohol use | 0
unconscious | 0
intubated | 0
Glasgow coma score 3E | 0
skin incision in right temporal region | 0
soft tissue defects in right temporal region | 0
negative light reflexes | 0
negative corneal reflexes | 0
absent spontaneous breathing | 0
heart rate 56 beats/min | 0
blood pressure 80/40 mmHg | 0
body temperature below 36°C | 0
central venous pressure 1 cm H2O | 0
bone fragments in right temporal region | 0
hemorrhagic contusion area in right frontotemporal area | 0
edema in right frontotemporal area | 0
temporal lobe inferomedially | 0
midline structures | 0
minimal left shift | 0
mechanical ventilation | 0
crystalloid fluid administration | 0
dopamine infusion | 0
mannitol therapy | 0
furosemide | 0
metoclopramide HCl | 0
famotidine | 0
acetylcysteine | 0
noradrenaline infusion | 0
enteral feeding | -24
eye opening | -72
eye closing | -72
blinking | -72
positive light reflexes | -72
positive corneal reflexes | -72
absent spontaneous limb movement | -72
absent response to pain stimuli | -72
percutaneous tracheotomy | -144
locked-in syndrome diagnosis | -168
vertical eye movements | -168
meaningful blinking | -168
quadriplegia | -168
minimal pressure in pons and mesencephalon | -168
partial compression in fourth ventricle | -168
hyperdense area in left cerebellar hemisphere | -168
hemodynamic problems | -168
fever | -168
infection | -168
antibiotic treatment | -168
pulmonary edema | -168
acute respiratory distress syndrome | -168
adjusted ventilation modes | -168
melena | -408
decreased hemoglobin | -408
decreased hematocrit | -408
blood product replacement | -408
omeprazole | -408
multiorgan failure | -864
death | -864
cerebellar ischemia | -864
normal vertebrobasilar artery system | -864
pneumonia | -864
respiratory arrest | -864
respiratory failure | -864
pulmonary embolism | -864
sepsis | -864
gastrointestinal hemorrhage | -864
disseminated intravascular coagulation | -864
pontine abscess | -864
