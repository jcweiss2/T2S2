63 years old | 0
male | 0
admitted to the hospital | 0
ingestion of wild mushrooms | -36
weakness | 0
nausea | 0
vomiting | 0
diarrhea | 0
hypertension | -6720
colon carcinoma | -6720
surgery | -1344
chemotherapy | -1344
no metastasis in the liver | 0
no alcohol consumption | 0
no medication use | 0
awake and fully oriented | 0
normal vital signs | 0
dehydration | 0
normal arterial blood gas analysis | 0
nonreactive hepatitis B surface antigen | 0
nonreactive hepatitis B core antibody | 0
nonreactive immunoglobulin M | 0
nonreactive antihepatitis C antibody | 0
negative hepatitis B virus DNA analysis | 0
gastric lavage | 0
activated charcoal | 0
rehydration | 0
silibinin | 0
acetylcysteine | 0
penicillin G | 0
multivitamin | 0
alpha lipoic acid | 0
vitamin K | 6
severe nausea | -29
severe vomiting | -29
severe diarrhea | -29
increased AST | 6
increased ALT | 6
increased LDH | 6
increased total bilirubin | 6
increased direct bilirubin | 6
prolonged PT | 6
elevated INR | 6
metabolic acidosis | 12
respiratory alkalosis | 12
fresh frozen plasma | 12
hemodialysis | 12
somnolent | 30
mildly tachypneic | 30
flapping tremor | 48
hepatic encephalopathy | 48
hepatorenal syndrome | 84
sedated and intubated | 84
cardiac arrest | 90
resuscitation | 90
second cardiac arrest | 98
death | 98