45 years old | 0
male | 0
cardiac transplantation | -2016
ischaemic cardiomyopathy | -2016
atrial fibrillation/flutter | 0
hypertension | 0
dyslipidaemia | 0
depression | 0
cardiac biopsy | -336
mild rejection | -336
tacrolimus | -336
mycophenolate mofetil | -336
prednisolone | -336
worsening rejection | -350
first-degree heart block | -350
second-degree heart block | -350
isoprenaline | -350
methylprednisolone | -350
sepsis | -720
dialysis-dependent acute kidney injury (AKI) | -720
haemopericardium | -720
peripheral limb ischaemia | -720
below-knee amputation | -720
severe upper abdominal pain | -240
investigated for severe upper abdominal pain | -240
haemoglobin reduced | -240
elevated white cell count | -240
reduced platelets | -240
elevated bilirubin | -240
elevated gamma-GT | -240
elevated alkaline phosphatase | -240
elevated transaminases | -240
non-contrast CT abdomen | -240
hyperdense haemobilia | -240
haemoperitoneum | -240
abdominal ultrasound | -240
contiguous haematoma | -240
gallbladder wall defect | -240
emergency laparoscopic cholecystectomy | 0
abdominal washout | 0
necrotic and perforated gallbladder | 0
moderate-volume haemoperitoneum | 0
bradycardic | 2
loss of cardiac output | 2
resuscitation | 2
epinephrine infusion | 2
follow-up ultrasound | 216
no collection or biliary obstruction | 216
protracted recovery | 216
cardiac arrest | 360
automated implantable cardioverter-defibrillator (AICD) insertion | 360
fungal infective endocarditis | 360
post-transplant lymphoproliferative disorder | 360
pulmonary embolism | 360
discharged from ICU | 1800
readmission to ICU | 1800
sepsis | 1800
hypotension | 1800
AKI resolved | 1800
discharged home | 5760
physical rehabilitation | 5760
ongoing antirejection regimen | 5760
everolimus | 5760
tacrolimus | 5760
prednisolone | 5760
physiotherapy | 5760
occupational therapy | 5760
consideration of lower limb prostheses | 5760