42 years old | 0 | 0 
male | 0 | 0 
admitted to the hospital | 0 | 0 
generalized weakness | -2160 | 0 
fever | -2160 | 0 
cough | -2160 | 0 
weight loss | -2160 | 0 
lived in Guatemala | -8760 | -720 
HIV-antibody test positive | -720 | -720 
sputum AFB smear positive | -720 | -720 
AIDS diagnosis | -720 | -720 
HIV-1 Western blot test positive | -720 | -720 
CD4 cell count 10/µL | -720 | -720 
HIV RNA titer 18,000 copies/mL | -720 | -720 
anti-tuberculosis medications started | -720 | -480 
fluconazole started | -720 | -480 
trimethoprim/sulfamethoxazole started | -720 | -480 
generalized weakness persisted | -480 | 0 
fever persisted | -480 | 0 
oral thrush | 0 | 0 
hepatosplenomegaly | 0 | 0 
ascites | 0 | 0 
hemoglobin 10.6g/dL | 0 | 0 
white blood cell 2,700/µL | 0 | 0 
platelet 58,000/µL | 0 | 0 
total bilirubin 2.4mg/dL | 0 | 0 
AST/ALT 131/48IU/L | 0 | 0 
ALP 114IU/L | 0 | 0 
GGT 133 IU/L | 0 | 0 
costophrenic angle blunting | 0 | 0 
fluid shifting in the right hemithorax | 0 | 0 
mild pneumonic infiltration in left lung | 0 | 0 
disseminated tuberculosis suspected | 0 | 0 
anti-retroviral agents started | 0 | 0 
pancytopenia progressed | 24 | 120 
hemoglobin 7.4g/dL | 24 | 24 
white blood cell 1,070/µL | 24 | 24 
platelet 13,000/µL | 24 | 24 
rifampin discontinued | 24 | 24 
zidovudine discontinued | 24 | 24 
trimethoprim/sulfamethoxazole discontinued | 24 | 24 
new pulmonary infiltrates | 120 | 120 
septic shock | 120 | 120 
piperacillin/tazobactam started | 120 | 120 
mechanical ventilator support started | 144 | 144 
bone marrow aspiration and biopsy performed | 216 | 216 
Histoplasma capsulatum identified | 216 | 216 
disseminated histoplasmosis diagnosed | 216 | 216 
death | 240 | 240 
refractory septic shock | 240 | 240 
hypoxia | 240 | 240