70 years old | 0
female | 0
chronic obstructive pulmonary disease | 0
smoking | 0
hypertension | 0
dyslipidemia | 0
osteoporosis | 0
appendectomy | -122640
left partial mastectomy | -113880
right femoral hernia repair | -8760
ruptured abdominal aortic aneurysm | 0
retroperitoneal hematoma | 0
infra-renal aortic prosthesis | 0
ligated inferior mesenteric artery |0
bilateral iliac thrombosis | 0
aorto-bifemoral bypass | 24
non ST-elevating myocardial infarction | 24
occluded circumflex artery | 24
right brachial artery thrombosis | 48
brachial embolectomy | 48
post-operative ileus | 168
diffuse abdominal pain | 576
leukocytosis | 576
no fever | 576
hemodynamically stable | 576
no peritonitis | 576
air in left retroperitoneum | 576
possible free air above bladder | 576
descending colon wall thickening | 576
contrast extravasation | 576
left colic perforation | 576
ischemic colitis | 576
exploratory laparotomy | 576
ischemia of small bowel | 576
ischemia of descending colon | 576
ischemia of sigmoid colon | 576
ischemia of rectum | 576
small bowel resection | 576
primary anastomosis | 576
left colectomy | 576
sigmoidectomy | 576
proctectomy | 576
terminal colostomy | 576
JP drains placement | 576
failed extubations | 912
exacerbated COPD | 912
volume overload | 912
splenic infarction | 912
left renal artery thrombosis | 912
non-enhancing left kidney | 912
peri-renal air bubbles | 912
intra-abdominal fluid collections | 912
JP drains well positioned | 912
dilated small bowel | 912
non-viable small bowel resection | 912
primary anastomosis | 912
colostomy takedown | 912
splenic necrosis | 912
left kidney necrosis | 912
splenectomy | 912
left nephrectomy | 912
terminal colostomy | 912
jejunal feeding tube | 912
abdominal fluid culture | 912
Gram stain | 912
Pseudomonas aeruginosa | 912
piperacillin-tazobactam | 912
fungal culture positive | 1032
voriconazole | 1032
sepsis | 1032
respiratory failure | 1032
acute kidney injury | 1032
diffuse abdominal pain | 1032
JP drain enteric formula | 1032
enteral feeds stopped | 1032
CT abdomen perforated small bowel | 1032
anastomotic leak | 1032
Mucor sp. culture | 1032
liposomal amphotericin B | 1032
comfort measures | 1032
death | 1032
