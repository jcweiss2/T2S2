48 years old | 0
female | 0
weight loss | -720
fever | -720
general weakness | -720
hyperparathyroidism | -720
febrile shock | -720
admitted to another hospital | -720
transferred to our hospital | 0
blood pressure 86/54 mmHg | 0
pulse rate 136/min | 0
body temperature 38.5℃ | 0
respiratory rate 28/min | 0
coarse breathing sounds | 0
crackles in both lower lung zones | 0
severe dyspnea | 0
serum urea 37 mg/dL | 0
creatinine 2.3 mg/dL | 0
calcium 14.1 mg/dL | 0
ionized calcium 7.8 mg/dL | 0
phosphorus 2.3 mg/dL | 0
intact PTH 635.30 pg/mL | 0
WBC 24,460/mm3 | 0
pH 7.235 | 0
PaCO2 61.8 mmHg | 0
PaO2 75.9 mmHg | 0
HCO3 25.6 mmol/L | 0
O2 saturation 94% | 0
patchy bilateral airspace consolidation | 0
airspace consolidation in bilateral lower lobes | 0
multifocal patchy ground-glass opacities | 0
parathyroid adenoma | 0
hyperparathyroidism-associated hypercalcemia | 0
pneumonia-complicated septic shock | 0
mechanical ventilator care | 0
ACMV | 0
CRRT | 0
bronchoscopy | 0
bronchoalveolar lavage | 0
MRSA | 0
parathyroidectomy | 24
improved from sepsis | 24
weaned from mechanical ventilation | 24
bilateral pulmonary airspace consolidations remained | 24
HRCT | 48
geographic high-attenuation consolidation | 48
ground-glass opacities | 48
metastatic calcifications | 48
bone scintigraphy | 48
Tc-99m MDP | 48
dense accumulation of radioactive tracer | 48
exertional dyspnea | 48
severely restrictive physiology | 48
low diffusion capacity | 48
percutaneous lung biopsy | 72
metastatic pulmonary calcification | 72
surgical resection of parathyroid | -2160
serum calcium level maintained within normal range | 2160
pulmonary function test showed nearly complete recovery | 2160
recovered health without symptoms | 2160