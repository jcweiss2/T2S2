32 years old | 0
male | 0
admitted to the hospital | 0
abdominal pain | -432
recurrent ascites | -432
nausea | -24
dizziness | -24
sodium level of 120 mEq/L | -24
paracentesis | -24
ceftriaxone | -24
dyspnea | -24
increased oxygen requirements | -24
pleural fluid analysis | -24
Cryptococcal antigen positive | -24
titer 1:256 | -24
IV fluconazole | -24
transferred to hospital | 0
cryptogenic cirrhosis | 0
right hypothalamic juvenile pilocytic astrocytoma | 0
status-post resection | 0
radiation | 0
bilateral occipital ventriculoperitoneal shunt placement | 0
panhypopituitarism | 0
oral hydrocortisone | 0
desmopressin | 0
hypernatremic | 0
afebrile | 0
normal white blood cell count | 0
blood cultures negative | 0
HIV test negative | 0
ALT 28 units/L | 0
AST 35 units/L | 0
viral hepatitis panel negative | 0
stress-dose steroids | 0
IV hydrocortisone | 0
symptomatic relief of dyspnea | 24
thoracentesis | 24
transudative fluid | 24
paracentesis | 48
ceftriaxone discontinued | 48
CT thorax | 48
massive left-sided pleural effusion | 48
atypical pneumonia | 48
reactive lymphadenopathy | 48
serum Cryptococcal Ag positive | 72
liposomal amphotericin B | 72
flucytosine | 72
flucytosine toxicities monitored | 72
transudative pleural fluid Cryptococcal Ag positive | 96
blood cultures grew C. neoformans | 96
pleural and abdominal fluid cultures grew C. neoformans | 120
fungemia | 120
transthoracic echo | 120
no vegetation | 120
CT of the head | 120
no ventriculitis | 120
lumbar puncture | 120
CSF positive for Cryptococcal Ag | 120
CSF culture positive | 144
neurologic intensive care unit | 144
removal of VP shunt | 144
placement of external ventricular drain | 144
lethargic | 264
altered mental status | 264
EEG consistent with non-convulsive status epilepticus | 264
levetiracetam | 264
lacosamide | 264
intubated | 264
midazolam drip | 264
ketamine | 264
pressor support | 264
nephrology consulted | 264
anuric AKI | 264
acute tubular necrosis | 264
furosemide diuresis stopped | 264
continuous veno-venous hemofiltration | 264
flucytosine renally adjusted | 264
septic shock | 312
negative repeat blood cultures | 312
piperacillin/tazobactam | 312
vancomycin | 312
meropenem | 312
daptomycin | 312
five pressors | 312
sodium bicarbonate infusion | 312
increase in stress steroids | 312
shock liver | 312
disseminated intravascular coagulopathy | 312
bleeding from nasogastric tube | 336
transfusions of blood | 336
transfusions of platelets | 336
transfusions of fresh frozen plasma | 336
transfusions of cryoprecipitate | 336
comfort care measures | 360
died | 360