10 years old | 0 | 0 
male | 0 | 0 
pre-term | 0 | 0 
gestational age of 33 weeks and 2 days | 0 | 0 
developmental delays in growth | 0 | 0 
developmental delays in motor function | 0 | 0 
short stature | -1440 | -1440 
Russell–Silver syndrome | -1440 | -1440 
proteinuria | -1440 | -1440 
hypoalbuminemia | -1440 | -1440 
nephrotic syndrome | -1440 | -1440 
high-dose steroid | -1440 | -720 
calcineurin inhibitor | -1440 | -720 
renal function deterioration | -720 | 0 
right renal vein thrombosis | -720 | -720 
pulmonary embolism | -720 | -720 
anticoagulants | -720 | -720 
persistent pulmonary hypertension | -720 | 0 
sildenafil | -720 | 0 
living donor kidney transplantation | 0 | 0 
immunosuppression | 0 | 215 
prednisolone | 0 | 215 
mycophenolate mofetil (MMF) | 0 | 70 
tacrolimus | 0 | 215 
discontinued MMF | 70 | 70 
steroid tapered | 70 | 215 
pneumocystis pneumonia | 90 | 104 
mechanical ventilation | 90 | 104 
intravenous sulfamethoxazole/trimethoprim | 90 | 104 
steroid increased | 90 | 215 
dysuria | 135 | 215 
gross hematuria | 135 | 215 
blood urea nitrogen (BUN) 24 mg/dL | 135 | 135 
creatinine (Cr) 0.56 mg/dL | 135 | 135 
C-reactive protein (CRP) 0.42 mg/dL | 135 | 135 
urinalysis revealed a red blood cell (RBC) count > 100/high power fields (HPF) | 135 | 135 
urinalysis revealed a white blood cell (WBC) count > 100/HPF | 135 | 135 
urine culture for bacteria negative | 135 | 135 
urine BK virus negative | 135 | 135 
urine John Cunningham (JC) virus polymerase chain reaction (PCR) positive | 135 | 135 
urine adenovirus culture positive | 135 | 135 
hemorrhagic cystitis | 135 | 215 
hydration | 135 | 215 
pain control | 135 | 215 
fever | 159 | 215 
general weakness | 159 | 215 
chest tightness | 159 | 215 
mild cough | 159 | 215 
persistent dysuria | 159 | 215 
persistent hematuria | 159 | 215 
BUN at 175 mg/dL | 159 | 159 
Cr at 8.29 mg/dL | 159 | 159 
CRP at 30.23 mg/dL | 159 | 159 
emergent hemodialysis | 159 | 215 
piperacillin/tazobactam | 159 | 215 
sputum culture negative | 159 | 159 
blood culture negative | 159 | 159 
urine culture negative | 159 | 159 
adenovirus real-time PCR of sputum positive | 159 | 159 
blood cytomegalovirus (CMV) antigen positive | 159 | 159 
disseminated adenovirus infection | 159 | 215 
immunosuppression reduction | 159 | 215 
ganciclovir | 159 | 215 
renal allograft biopsy | 159 | 159 
diffuse necrotizing granulomatous tubulointerstitial nephritis | 159 | 159 
infectious tubulointerstitial nephritis | 159 | 159 
staining for CD3 negative | 159 | 159 
staining for C4d negative | 159 | 159 
JC virus PCR positive | 159 | 159 
serum CMV PCR positive | 159 | 159 
coinfection | 159 | 215 
ganciclovir targeting CMV | 159 | 215 
antibiotic therapy | 159 | 215 
granulocyte colony-stimulating factor | 159 | 215 
immunoglobulin | 159 | 215 
transfusion | 159 | 215 
hemodialysis | 159 | 215 
cidofovir | 167 | 215 
nephrotoxicity | 167 | 215 
serum adenovirus PCR positive | 167 | 215 
cerebrospinal fluid adenovirus PCR positive | 167 | 215 
renal function not recovered | 167 | 215 
generalized tonic-clonic seizure | 167 | 215 
vancomycin | 167 | 215 
meropenem | 167 | 215 
acyclovir | 167 | 215 
anemia | 167 | 215 
leukopenia | 167 | 215 
thrombocytopenia | 167 | 215 
bone marrow suppression | 167 | 215 
mechanical ventilation | 167 | 215 
continuous renal replacement therapy | 167 | 215 
death | 215 | 215