42 years old | 0
male | 0
Hispanic | 0
admitted to the hospital | 0
bilateral lower extremity pain | -504
bilateral lower extremity pain located at the upper thighs with radiation down the legs | -504
severe and constant bilateral lower extremity pain | -504
non-radiating severe frontal throbbing headache | -168
diplopia | -168
nausea | -96
vomiting | -96
low-grade fever | -96
20 pack year history of smoking | -33600
chronic alcohol intake | -33600
construction worker | 0
somnolent but arousable patient | 0
hypereflexia of the right brachioradialis | 0
hypereflexia of the right biceps | 0
decrease of muscle strength of bilateral lower extremities | 0
mild hyponatremia | 0
mild transaminase elevation | 0
hyperbilirubinemia | 0
ammonia level in the upper normal range | 0
urinalysis negative | 0
urine toxicology screen negative | 0
alcohol level negative | 0
hepatitis serology panel negative | 0
HIV negative | 0
chest x-ray unremarkable | 0
CT of the brain with multiple intraaxial hyperdense lesions | 0
CT of the brain with surrounding vasogenic edema | 0
hematogenous spread suggested | 0
Chest-CT with bilateral cavitary nodules | 0
Chest-CT with right hilar lymphadenopathy | 0
empiric antibiotics started | 0
vancomycin 1 gram every 12 hours | 0
ceftriaxone 2 grams every 12 hours | 0
dexamethasone 6mg IV every 8 hours | 0
MRI of the brain | 24
MRI of the brain with multiple bilateral supratentorial and infratentorial rim enhancing lesions | 24
pulmonary service consulted | 48
bronchoscopy | 48
bronchoalveloar lavage (BAL) | 48
BAL cultures negative | 48
AFB stain negative | 48
infectious disease service consulted | 48
PPD recommended | 48
Quaniferon Gold recommended | 48
coccidiodies serology recommended | 48
aspergillus antigen recommended | 48
toxoplasma IgG antibody recommended | 48
serum crytococcal antigen recommended | 48
lumbar puncture recommended | 48
cerebrospinal fluid (CSF) analysis | 48
CSF analysis with elevated WBC count | 48
no evidence of vegetations on echocardiogram | 48
neurosurgery consulted | 96
brain biopsy suggested | 96
brain biopsy not possible | 96
mental status deteriorated | 240
disoriented to time and place | 240
oriented to person | 240
weakness of the left upper extremity | 288
unsteady antalgic gait | 288
weakness of the right upper extremity | 312
ptosis | 312
right lower facial weakness | 312
cardiothoracic surgery consulted | 312
video-assisted thoracoscopic surgery with biopsy of cavitary lung lesions recommended | 312
location of the lesion unsuitable for surgical access | 312
GCS decreased to 7 | 336
bradycardic | 336
complete right sided paralysis | 336
positive right side babinski | 336
transferred to the medical intensive care unit (MICU) | 336
repeat head-CT with contrast | 336
multiple ring enhancing lesions | 336
no evidence for acute intracranial hemorrhage | 336
no evidence for herniation | 336
no evidence for mass effect | 336
no evidence for midline shift | 336
amphotericin B started | 336
albendazole started | 432
pyrimethamine started | 432
sulfadiazine started | 432
leukovorin started | 432
tachycardic | 456
desaturated to <80% | 456
intubated | 456
mechanical ventilation support started | 456
expired | 480
autopsy performed | 480
macroscopic findings of respiratory system with bilateral serosanguineous pleural effusions | 480
lung abscess at the right hilum | 480
microscopic examination of the right hilum abscess with foci of necrosis | 480
microscopic examination of the right hilum abscess with acute inflammation | 480
microscopic examination of the right hilum abscess with microabscess formation | 480
macroscopic findings of the brain with multiple bilateral cavities | 480
microscopic examination findings with foci of acute inflammation | 480
microscopic examination findings with microabscess formation | 480
Grocott methena mine silver (GMS) stain positive | 480
grain stain positive | 480
Fite’s stain positive | 480
tissue samples from the brain abscess lesions and lung cavitary lesions sent for cultures | 480
cultures grew nocardia species | 480
PCR analysis revealed nocardia wallacei species | 480
resistance to ceftriaxone | 480
resistance to levofloxacin | 480
resistance to aminoglycosides (amikacin) | 480
resistance to sulfonamides (trimethoprim-sulfamethoxazole – TMP-SMX) | 480
sensitive to imipenem | 480
final autopsy diagnosis with nocardia pneumonitis | 480
final autopsy diagnosis with nocardia encephalitis | 480
cause of death stated as systemic nocardiosis | 480