57 years old | 0
male | 0
admitted to the hospital | 0
hepatitis B virus | -1200
alcoholic liver cirrhosis | -1200
hepatic failure | -1200
esophageal varix bleeding | -36
hepatic encephalopathy | -36
Child-Pugh grade C | -36
intensive medical care | -36
left bipolar hemiarthroplasty | -12
left femoral neck fracture | -12
decompensated liver cirrhosis | -12
liver transplant candidate | -12
MELD score of 28 points | -12
painful anal swelling | -24
dysuria | -24
icteric sclera | -24
abdominal distension | -24
hepato-renal syndrome | -24
ICU admission | -24
Fournier’s gangrene | -24
wide debridement of the wound | -24
T-colostomy | -24
bleeding control surgery | -24
norepinephrine administration | -24
vasopressin administration | -24
bleeding control | -12
DDLT | 0
Enterococcus faecium detection | -12
Candida albicans detection | -12
vancomycin-resistant Enterococcus | -12
Achromobacter xylosoxidans detection | -12
Pseudomonas aeruginosa detection | -12
varix bleeding | -12
wound bleeding | -12
coagulopathy | -12
blood transfusions | -12
hemoglobin level dropped | -12
tazocin administration | -24
meropenem administration | -24
vancomycin administration | 0
teicoplanin administration | 0
amphotericin B administration | 0
micafungin administration | 0
C-reactive protein levels decreased | 12
immunosuppressant treatment | 0
FK-506 trough level adjustment | 0
mycomofetil administration | 0
steroids administration | 0
recovered | 24
discharged | 168