72 years old | 0
male | 0
admitted to the hospital | 0
weakness | -336
fatigue | -336
dyspnoea on exertion | -96
no chest pain | -96
no palpitations | -96
no ankle oedema | -96
increased urinary frequency | -96
dark urine | -96
no dysuria | -96
no dysphagia | -96
no bleeding per rectum | -96
no abdominal pain | -96
no weight loss | -96
no fever | -96
no rigours | -96
no recent travel | -96
benign prostatic hyperplasia | 0
Dutasteride/tamsulosin 0.5/0.4 mg | 0
tachycardia | 0
fever | 0
temperature 39.1°C | 0
C-reactive protein 101 mg/L | 0
high-sensitivity troponin T 500 ng/L | 0
N-terminal pro-B-type natriuretic peptide 4337 pg/mL | 0
ferritin 1498 ng/mL | 0
sinus tachycardia | 0
diffuse non-territorial ischaemic changes | 0
pulmonary oedema | 0
bilateral pleural effusions | 0
ground glass change | 0
interlobular septal thickening | 0
pericardial fluid | 0
pericardial thickening | 0
systemic inflammatory response syndrome | 0
investigated for COVID-19 | 0
nasal-pharyngeal swabs negative | 0
first presentation of heart failure | 48
ischaemic aetiology | 48
audible murmur | 48
abnormal electrocardiogram | 48
elevated NT-proBNP | 48
pulmonary embolism | 48
cardiology team consulted | 96
coronary angiogram | 144
occlusion of right coronary artery | 144
collateralization from left coronary system | 144
left coronary system free of significant coronary disease | 144
intravenous diuretic therapy | 144
disease-modifying HF therapies | 144
discharged home | 216
ischaemic HF with LV involvement | 216
RCA occlusion | 216
pantoprazole 40 mg | 216
aspirin 75 mg | 216
clopidogrel 75 mg | 216
furosemide 40 mg | 216
atorvastatin 80 mg | 216
ramipril 2.5 mg | 216
bisoprolol 1.25 mg | 216
re-presentation to hospital | 600
acute decompensation | 600
New York Heart Association class III symptoms | 600
fatigue | 600
night sweats | 600
palpitations | 600
intravenous diuresis | 600
severe MR | 600
restricted motion of posterior mitral valve leaflet | 600
large LV saccular outpouching | 600
basal inferior wall | 600
CMR viability study | 624
dilated LV | 624
focal posterior saccular outpouching | 624
basal to mid-inferior wall | 624
transmural late gadolinium enhancement | 624
thrombus | 624
intact pericardium | 624
organizing thrombus | 624
inferior free wall rupture | 624
saccular outpouching | 624
narrow neck | 624
attenuated layer | 624
LV pseudoaneurysm | 624
severe secondary MR | 624
tethered chordae | 624
restricted motion of posterior mitral leaflet | 624
bed rest | 624
close monitoring | 624
coronary care unit | 624
surgical replacement of mitral valve | 744
repair of LVP | 744
Perimount Magna Ease mitral valve | 744
cuff of pericardium | 744
direct closure | 744
no immediate complications | 744
postoperative course | 744
arrhythmia | 744
cardiogenic shock | 744
ischaemic sigmoid colitis | 744
bowel perforation | 744
sepsis | 744
intensive rehabilitation | 1032
discharged home | 1032
fully independent | 1032
atorvastatin 80 mg | 1032
bisoprolol 7.5 mg | 1032
furosemide 40 mg | 1032
aspirin 75 mg | 1032
apixaban 5 mg | 1032
pantoprazole 40 mg | 1032
ramipril 7.5 mg | 1032
severely depressed LV systolic function | 1032
ejection fraction 26% | 1032
inferior and infero-lateral walls akinetic | 1032
mitral valve prosthesis functioning well | 1032
no significant transvalvular or paravalvular regurgitation | 1032