born | -72 
breech presentation | -72 
cord prolapse | -72 
mechanical ventilation initiated | 0 
central umbilical catheters inserted | 0 
total parenteral nutrition initiated | 0 
empiric antibiotics initiated | 0 
skin sensors for monitoring applied | 0 
late-onset sepsis secondary to Escherichia coli bacteremia | -216 
antimicrobial therapy with cefepime initiated | -216 
antimicrobial therapy with cefepime discontinued | -156 
adhesive patch removed | -144 
skin abrasion | -144 
erythema | -120 
induration | -120 
plaque with necrotic center | -120 
ulcer with extension to subcutaneous cell tissue | -96 
necrotic area progression | -96 
intensive treatment by wound care team initiated | -96 
thermic instability | -48 
metabolic acidosis | -48 
hyperglycemia | -48 
hypotension | -48 
cutaneous mucormicosis suspected | -48 
skin biopsy | -48 
empiric antifungal treatment with liposomal amphotericin B initiated | -48 
fungal biomarkers not performed | -48 
general condition deterioration | -24 
refractory shock | -12 
renal failure | -12 
death | 0 
fungal cultures obtained | -24 
Rhizopus spp. identified | -24 
histopathology report | -24 
broad aseptate hyphae with right angle branching identified | -24 
mass spectroscopy performed | -24 
polymerase chain reaction performed | -24 
Rhizopus arrhizus identified | -24 
fungal blood cultures collected | -72 
fungal blood cultures negative | -72 
autopsy not performed | 0 
skin abscesses not found | 0 
necrotizing fasciitis not found | 0 
clostridial gas gangrene not found | 0 
sepsis-associated purpura fulminans not found | 0 
bacterial cellulitis not found | 0 
pyoderma gangrenosum not found | 0 
surgical debridement not performed | 0 
antifungal treatment with L-AmB continued | 0 
antifungal treatment with L-AmB discontinued | 0 
infection control not achieved | 0 
case report approved by Institutional Ethics Committee | 0 
case report published | 0