39 year old|0
male|0
admitted for septic shock|0
malaise|-168
encephalopathy|-168
blood cultures grew MSSA|0
fluid cultures obtained from left elbow olecranon bursa grew MSSA|0
fluid cultures obtained from right foot abscess grew MSSA|0
concern for endocarditis|0
systemic emboli|0
chest radiograph notable for retained foreign objects|0
abdominal radiograph notable for retained foreign objects|0
transesophageal echocardiography negative for vegetation|0
CT chest showed multiple bilateral peripheral nodular opacities|0
developing central cavitation|0
MSSA pulmonary septic emboli|0
retained foreign body in right upper pulmonary artery sub-segmental branch|0
CT abdomen and pelvis showed retained guide wire|0
retained guide wire extending from IVC to left iliac and left common femoral vein|0
motor vehicle accident|-140160
trauma intensive care stay|-140160
femoral central venous access placement|-140160
sixteen years prior to current presentation|-140160
aware of guide wire presence|0
initial plan for re-imaging and retrieval|0
lost to follow up|0
interventional radiology removed IVC portion of wire|0
unable to retrieve right pulmonary artery portion|0
completely epithelialized|0
started on appropriate antibiotic regimen|0
clearance of bacteremia|0
source control|0
resolution of bacteremia|0
resolution of symptoms|0
lack of exposed hardware|0
did not require chronic lifelong suppression therapy|0
retained pulmonary artery fragment of guide wire|0
