37 years old | 0
    female | 0
    diagnosed with late-onset OTCD | -288576
    seizures at age 7 | -288576
    hyperammonemia after valproic acid administration | -288576
    liver biopsy examination | -288576
    liver OTC enzyme activity 30% of control | -288576
    visited emergency room for hyperammonemia | -21600
    hemodialysis for impaired consciousness at age 18 | -21600
    hemodialysis for impaired consciousness at age 21 | -21600
    self-restricted protein diet | -21600
    L-carnitine treatment | -21600
    natural pregnancy at age 37 | 0
    delivered male baby at 41 weeks and 1 day gestation | 0
    blood ammonia 68 μmol/L at delivery | 0
    blood ammonia 59 μmol/L at 10 hours after delivery | 10
    blood ammonia 54 μmol/L at 24 hours after delivery | 24
    hyperammonemia 194 μmol/L 4 days after delivery | 96
    discharged 6 days after delivery | 144
    consumed hamburger and 250g beef after discharge | 144
    hospitalized on emergency basis at midnight | 168
    hyperammonemia 180 μmol/L | 168
    impaired consciousness | 168
    blood ammonia decreased to 82 μmol/L with arginine | 168
    hemodialysis and continuous hemodiafiltration | 168
    blood ammonia increased to 339 μmol/L | 168
    grade III hepatic coma | 168
    high-calorie infusion 2500 kcal/d | 168
    arginine 80 mg/kg per day | 168
    citrulline 150 mg/kg per day | 168
    sodium benzoate 150 mg/kg per day | 168
    sodium phenylbutyrate 140 mg/kg per day | 168
    hyperammonemia improved | 168
    attempted extubation | 168
    reintubated due to respiratory failure | 168
    blood ammonia increased to 210 μmol/L after extubation stress | 168
    ammonia levels decreased to 60 μmol/L | 168
    sepsis | 168
    managed in ICU for 43 days | 168
    atrophy of bilateral frontal and temporal lobes | 168
    decreased blood flow on SPECT | 168
    discharge from hospital | 168
    brain MRI and SPECT 7 months after delivery | 168
    able to raise child | 168
    developed hepatic coma requiring respirator | 168
    resumed breathing without assistance after 40 days | 168
    improved consciousness | 168
    maternal milk production continued for a month | 168
    hyperammonemia persisted after stopping maternal milk | 168
    candidate for liver transplantation | 168
    <|eot_id|>
    