85 years old | 0
woman | 0
hypertension | 0
dyslipidemia |6
chest pain | -72
presented to emergency room | 0
dyspnea | 0
elevated troponin T level | 0
ST depression in V2–5 | 0
pulmonary congestion | 0
severe mitral regurgitation | 0
P2 prolapse | 0
99% stenosis of mid-portion of left circumflex artery | 0
intra-aortic balloon pumping initiated | 0
intubated in intensive care unit | 0
papillary muscle rupture | 0
diagnosed acute mitral regurgitation with papillary muscle rupture as complication of acute myocardial infarction | 0
cardiogenic shock | 0
hemodynamics managed with intra-aortic balloon pumping and inotrope support | 0
emergency percutaneous coronary intervention performed | 0
mitral valve replacement via minithoracotomy performed | 0
cardiopulmonary bypass established | 0
right femoral arterial cannulation | 0
right femoral and jugular venous drainage | 0
cardiac arrest achieved with antegrade cardioplegia | 0
approached mitral valve through left atriotomy | 0
partial anterolateral papillary muscle rupture observed | 0
mitral valve replacement performed with 29-mm Epic mitral stented tissue valve | 0
weaned from cardiopulmonary bypass | 0
minimal inotrope support | 0
hemodynamic status stabilized | 0
intra-aortic balloon pumping discontinued | 24
extubated | 48
sepsis | 96
rectal ulcer | 96
antibacterial treatment | 96
discharged from intensive care unit | 144
normal cardiac function | 144
normal bioprosthetic valve function | 144
walking 200 m independently | 0
transferred to another hospital | 0
