87 years old | 0
male | 0
admitted to the hospital | 0
diabetic ketoacidosis | 0
uncontrolled diabetes mellitus | -672
chronic renal failure | -672
left below knee amputation | -672
penetrating keratoplasty | -240
generalized weakness | 0
afebrile | 0
confused | 0
generally weak | 0
incoherent | 0
complete ophthalmoplegia | 0
non-reactive pupils | 0
no view of the posterior fundus | 0
reduction in right visual acuity | 0
infiltration of the right globe | 0
cavernous sinus thrombosis | 0
orbital cellulitis | 0
intravenous meropenem | 0
vancomycin | 0
heparin | 0
deteriorated level of consciousness | 24
seizures | 24
worsened orbital involvement | 24
poor enhancement of the right cavernous sinus | 24
lumbar puncture | 24
negative for microorganisms | 24
provisional diagnosis of mucormycosis | 24
micronasal abscesses | 24
right alar blackish discoloration | 24
intravenous amphotericin B | 24
caspofungin | 24
partial opacification of the maxillary and sphenoid sinuses | 48
fluid levels denoting acute insult | 48
increased right pre-septal thickening | 48
abnormal infiltration of the right eye | 48
rapid progression to the orbit | 48
gangrenous area on the tip of the nose | 48
suspicion of mucormycosis confirmed | 48
surgical debridement discussed | 48
written informed consent obtained | 48
right orbital exenteration | 72
widespread deep excision of the necrotic area | 72
peri-operative intravenous antibiotics | 72
peri-operative antifungals | 72
post-operative support | 72
Glasgow Coma Score of three | 96
clinically septic | 96
extension of necrotic tissue | 96
involvement of the right ear and left eye | 96
refused further surgical intervention | 96
negative blood cultures | 96
microscopic examination of tissue samples | 96
invasive broad fungal hyphae yeast cells | 96
acute and chronic inflammatory cells | 96
necrotic tissue | 96
suppurative microabscesses | 96
death | 96