29 years old | 0
    man | 0
    admitted to the hospital | 0
    intermittent fevers | -48
    fever | -48
    forehead headache | -48
    nausea absence | -48
    consumed unpasteurized cooked beef | -48
    type 2 diabetes mellitus | 0
    fatty liver | 0
    smoking | 0
    drinking | 0
    denied family history of hypertension | 0
    denied family history of stroke | 0
    nuchal rigidity | 0
    high glucose | 0
    high C-reactive protein | 0
    high erythrocyte sedimentation rate | 0
    normal white blood cells | 0
    normal red blood cells | 0
    normal hemoglobin | 0
    normal urea | 0
    normal creatinine | 0
    normal serum minerals | 0
    normal autoimmune antibodies | 0
    turbid cerebrospinal fluid | 0
    leukocytes 2090/mm3 | 0
    CSF protein 233.85 mg/dL | 0
    CSF glucose 1.4 mmol/L | 0
    serum glucose 9 mmol/L | 0
    CSF pressure > 33 cmH2O | 0
    CSF Gram-positive rods | 0
    negative CSF fungi | 0
    negative CSF acid-fast bacilli | 0
    blood cultures yielded L. monocytogenes | 192
    L. monocytogenes susceptible to ampicillin | 192
    susceptible to erythrocin | 192
    susceptible to meropenem | 192
    susceptible to penicillin | 192
    resistant to sulfamethoxazole | 192
    CSF cultures negative | 192
    urine cultures negative | 192
    CSF WBCs decreased | 336
    CSF protein decreased | 672
    unremarkable brain CT | 0
    bilateral bronchopneumonia | 0
    brain MRI T2-FLAIR hyperintense right pons | 96
    prominent temporal horns | 96
    ventricular enlargement | 96
    brain CT hemorrhage right pons | 336
    hydrocephalus | 336
    bilateral lateral ventricular hydrocephalus | 336
    third ventricle hydrocephalus | 336
    cerebral CT significant dilatation fourth ventricle | 528
    no remission lateral ventricles | 528
    brain CT rehaemorrhagia lateral ventricle | 696
    larger ventricular system | 696
    diagnosed Listeria rhombencephalitis | 0
    diagnosed hydrocephalus | 0
    diagnosed intracranial hemorrhage | 0
    empiric antibiotic therapy | 0
    ceftriaxone 2g every 12h | 0
    meropenem 1g every 8h | 48
    new symptoms | 120
    fever | 120
    sinus tachycardia | 120
    tachypnea | 120
    confusion | 120
    Glasgow Coma Scale score 12/15 | 120
    bilateral horizontal nystagmus | 120
    bilateral abducens nerve palsy | 120
    dysarthria | 120
    weakness of all four limbs | 120
    transferred to ICU | 120
    coma | 192
    Glasgow Coma Scale score 5/15 | 192
    intubated | 192
    ventilated | 192
    ampicillin | 192
    etimicin | 192
    meropenem | 192
    etimicin discontinued | 288
    afebrile | 288
    extraventricular drainage | 528
    rehaemorrhagia lateral ventricle | 696
    condition deteriorated | 696
    Glasgow Coma Scale score 3/15 | 696
    anisocoria | 696
    died | 744

<|eot_id|>
