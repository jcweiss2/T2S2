64 years old | 0
male | 0
Caucasian | 0
admitted to the hospital | 0
type 2 diabetes | -672
hypertension | -672
kidney transplant recipient | -672
immunosuppressive drugs | -672
tacrolimus | -672
mycophenolic acid | -672
prednisone | -672
shortness of breath | -96
fever | -96
cough | -96
emergency department visit | 0
serum creatinine 0.7 mg/dL | 0
glomerular filtration rate >60 ml/min/1.73 m2 | 0
chest radiography | 0
diffuse interstitial and airspace opacities | 0
multifocal pneumonia | 0
gram stain negative | 0
rapid influenza test negative | 0
pneumococcal and legionella urinary antigen test negative | 0
SARS-CoV-2 infection | 0
nasopharyngeal swab positive | 0
intensive care unit admission | 0
elective intubation | 0
hydroxychloroquine | 0
azithromycin | 0
cefepime | 0
mycophenolic acid suspension | 0
tacrolimus reduction | 0
prednisone continuation | 0
mechanical ventilation | 0
low tidal volume lung-protective strategy | 0
prone positioning | 0
neuromuscular blockade | 0
sedation | 0
high positive end-expiratory pressure therapy | 0
sputum sample redrawn | 72
increased endotracheal secretions | 72
worsening chest radiography results | 72
hypoxemia | 72
high dose corticosteroids | 72
methylprednisolone | 72
sputum examination positive for gram-negative bacilli | 96
S. maltophilia identification | 120
TMP/SMX initiation | 120
cefepime discontinuation | 120
AKI development | 168
worsening serum creatinine | 168
oliguria | 168
fluid administration | 168
immunosuppressive drugs continuation | 168
TMP/SMX discontinuation | 192
levofloxacin initiation | 192
kidney function deterioration | 192
serum creatinine increase | 192
GFR decrease | 192
hyperkalemia | 192
hemodialysis initiation | 192
urinalysis | 192
eosinophiluria absence | 192
white cell casts absence | 192
steroids continuation | 192
tacrolimus therapeutic levels | 192
kidney biopsy consideration | 192
comfort care measures | 264
death | 288