11 years old | 0
    female | 0
    systemic methicillin-resistant staphylococcus aureus (MRSA) infection | 0
    transferred to our hospital for rehabilitation | 0
    right knee pain | -1008
    back pain | -1008
    fevers | -1008
    purulent spider bite | -1008
    COVID-19 infection | -1008
    dehydration | -1008
    presented to an emergency department | -1008
    altered mental status | -1008
    incontinence | -1008
    febrile | -1008
    tachypneic | -1008
    tachycardic | -1008
    hypoxic | -1008
    admitted to the pediatric intensive care unit (PICU) | -1008
    blood culture positive for MRSA | -1008
    intravenous antibiotic therapy | -1008
    persistent symptoms | -1008
    magnetic resonance imaging (MRI) of the spine | -1008
    computed tomography (CT) of chest, abdomen, and pelvis | -1008
    multifocal fluid collections | -1008
    inflammation | -1008
    right psoas muscle involvement | -1008
    right thoracolumbar paraspinal soft tissues involvement | -1008
    cervical and thoracic prevertebral soft tissues involvement | -1008
    multifocal septic arthritis | -1008
    bilateral pleural effusions | -1008
    multifocal opacities | -1008
    multiple pulmonary nodules | -1008
    septic emboli | -1008
    MRI of the brain | -1008
    meningitis | -1008
    ventriculitis | -1008
    lumbar puncture | -1008
    cerebrospinal fluid positive for MRSA | -1008
    multiarticular surgical washouts | -1008
    washout of paraspinal abscesses | -1008
    bilateral chest tubes placed for empyema | -1008
    antibiotics continued | -1008
    clearing of blood cultures | -936
    clinical improvement | -936
    transfer to our facility for rehabilitation | -0
    clinically well appearing | 0
    afebrile | 0
    normal vital signs | 0
    CT imaging of chest, abdomen, and pelvis | 192
    decrease in most fluid collections | 192
    increased size of right psoas collection | 192
    MRI showing increased T1 signal intensity | 192
    blood products in right psoas collection | 192
    CT angiography | 192
    enhancing lesions in left medial lower lobe | 192
    enhancing lesions in right posterior mediastinum | 192
    enhancing lesions in right psoas | 192
    pseudoaneurysms | 192
    retrospective review of prior imaging | 192
    lesions present 2 weeks prior | -432
    hematocrit level stable | 0
    no need for blood transfusion | 0
    consultation with interventional radiology (IR) service | 192
    embolization of pulmonary lesion | 192
    right common femoral vein access | 192
    left pulmonary artery catheterization | 192
    diagnostic angiogram | 192
    pseudoaneurysm in left lower lobe artery | 192
    embolization with detachable coils | 192
    no antegrade flow postembolization | 192
    left common femoral artery access | 192
    diagnostic angiography of right L2-L3 lumbar artery | 192
    pseudoaneurysm in right psoas | 192
    embolization of lumbar artery pseudoaneurysm | 192
    angiography of right T9 intercostal artery | 192
    active hemorrhage | 192
    embolization of intercostal artery pseudoaneurysm | 192
    return to PICU | 192
    clinical stability | 192
    transfer to rehabilitation medicine service | 216
    CT angiogram postprocedure | 288
    stable embolization coils | 288
    no recurrent pseudoaneurysms | 288
    decrease in right psoas collection | 288
    uneventful clinical course | 336
    discharge | 336
    follow-up CT angiogram | 432
    further decrease in fluid collections | 432
    no new or recurrent pseudoaneurysms | 432