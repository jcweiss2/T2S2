66 years old | 0
female | 0
admitted to the hospital | 0
unconscious | 0
coma | 0
blood pressure 115/70 mm Hg | 0
heart rate 85/min | 0
oxygen saturation 97% | 0
temperature 36.0°C | 0
tachypnoeic | 0
bilateral miosis | 0
fingers in ulnar deviation | 0
absent reflexes | 0
discrete pretibial oedema bilateral | 0
no clonus | 0
no extrapyramidal signs | 0
hypotension 70/50 mm Hg | 2
decrease in SaO 85% | 2
pulmonary oedema | 2
miosis | 2
no pupillary reflexes on light | 2
no nuchal rigidity | 2
absent limb’s reflexes | 2
GCS 3 | 2
pulmonary crackles bilaterally | 2
respiration rate 25–30/min | 2
non-invasively monitored | 2
WBC 7.9 | 0
Plt 339 | 0
Hb 148 | 0
RBC 4.7 | 0
Htc 0.42 | 0
CRP 2.5 | 0
Glycemia 12.2 | 0
BUN 4.3 | 0
Creatinine 59.6 | 0
Na 136 | 0
K 3.76 | 0
Ca 2.3 | 0
AST 17.9 | 0
ALT 12.1 | 0
GGT 15.3 | 0
AF 85.5 | 0
Myoglobin 49.6 | 0
Troponin 11.1 | 0
D-dimer 3254.36 | 0
Ketones + | 0
Proteins 30 | 0
Ethanol 526 | 0
PT 10.67 | 0
aTPP 26.37 | 0
TT 20 | 0
pH 7.26 | 0
pCO2 3.5 | 0
SaO 94% | 0
HCO3 14 | 0
BE -15.4 | 0
Anion gap 21.7 | 0
Lactates >2 | 0
symptomatic treatment | 2
pulmonary aspiration | 2
intravenous colloids 500 mL | 2
NaCl 0.9% 500 mL | 2
oxygen support with nasal cannula 4–5 L/min | 2
amp furosemide 10 mg i.v. | 2
stable hemodynamic condition | 4
increase in blood pressure 110/70 mm Hg | 4
HR 110–120/min | 4
urine output 3.5 mL/min | 4
persistence of coma | 4
absence of reflexes | 4
toxicological screening | 4
low benzodiazepine levels 477 ng/mL | 4
excluded opiates | 4
excluded tramadol | 4
excluded methadone | 4
excluded cannabis | 4
hypotensive reaction 80/60 mm Hg | 6
drop of SaO 85% | 6
tachypnoea 35–40/min | 6
shallow respirations | 6
family indicated missing 250 mL of 70% ethanol-disinfectants | 6
BAC 526 mg/dL | 6
metabolic acidosis | 6
calculated osmolality 403–421 | 6
DD 3254 ng/mL | 6
anaesthesiology consultant recommended mask-oxygen | 6
no mechanical ventilation | 6
treatment with standard protocol | 8
D5 NS 100 mL/h | 8
potassium 10 mmoL/h | 8
thiamine 100 mg i.v. | 8
oxygen 4–5 L/min | 8
persistent areflex coma | 8
oscillation of BP 90/60 mm Hg | 8
PCR test for SARS-COV-2 negative | 8
hemodynamic instability | 10
age with reduced biotransformation activity | 10
risk of fluids overload | 10
immunocompromised condition | 10
high susceptibility to infections | 10
haemodialysis | 12
femoral catheter | 12
discontinued after 2.5 hours | 14.5
increased blood coagulation | 14.5
nadroparin 0.6 mL | 14.5
stuporous | 14.5
restoration of reflexes | 14.5
post-dialysis alcoholaemia 250 mg/dL | 14.5
ABGA corrected | 14.5
DD increased | 14.5
glycemia controlled | 16
lowest recorded values 5.0 mmol/L | 16
further treatment | 16
D5NS 100 mL/h | 16
amp ceftriaxone 2.0 g | 16
amp famotidine 20 mg i.v. tid | 16
nadroparin 0.6 mL tid | 16
LOC improved to mild somnolence | 24
pronounced depressed mood | 24
alcoholaemia 104 mg/dL | 24
no gastric discomfort | 24
no haematemesis | 24
no reduction in haemogram | 24
denied taking more than regular 5-HTP tablets | 24
specific therapy for RA discontinued | 24
transferred to psychiatric clinic | 48
stable hemodynamic and mental status | 48
recommended to use LMWH | 48
control haemostatic parameters | 48
continue regular therapy | 48