87 years old | 0
male | 0
admitted to the oncologic center | 0
abnormal prostate-specific antigen | -672
prostate cancer | -672
hypertension | -672
chronic kidney disease | -672
amlodipine | -672
hydrochlorothiazide | -672
no personal or familial history of abnormal bleeding | -672
no altered blood clotting test | -672
surgical castration | -1344
decrease of the PSA determinations | -1344
castration-resistant disease | -728
PSA levels rose | -728
peripheral anti-androgen blockade with bicalutamide | -728
decline in transient PSA determinations | -728
rising PSA | -480
second-line therapy with prednisone | -480
stabilization of the PSA levels | -480
gross hematuria | 0
back pain | 0
spontaneous skin hematomas | 0
severe anemia | 0
hemoglobin determination of 4.8 g/dL | 0
red-blood-cell transfusion | 0
prothrombin time of 14.7 seconds | 0
active partial thromboplastin time of 97.7 seconds | 0
fibrinogen level of 406 mg/dL | 0
liver function tests were normal | 0
abnormal bleeding | 0
inhibitor of the coagulation factor | 0
diagnosis of AHA | 0
FVIII < 1% | 0
FVIII inhibitor | 0
PSA level was stable | 0
computerized tomography scan | 0
no signs of new metastasis | 0
no evidence of cancer progression | 0
iliopsoas hematoma | 0
treatment with prednisone | 0
no improvement | 48
azathioprine | 48
hematuria ceased | 72
hemoglobin level remained stable | 72
no signs of new skin hematomas | 72
homeostatic agents were not necessary | 72
new CT study | 120
no further enlargement of the iliopsoas hematoma | 120
hematoma-associated back pain improved | 120
patient became asymptomatic | 408
discharged | 408
progressive fall of the inhibitor titles | 936
increase of the coagulation FVIII levels | 936
no other hemorrhage phenomenon | 936
admitted to the Intensive Care Unit | 1116
diagnosis of pneumonia | 1116
died due to septic shock | 1116