69 years old | 0
man | 0
Child–Pugh class C cirrhosis | 0
presented to the Emergency department | 0
slipped on wet grass | -unknown
fell on his left side | -unknown
glasgow coma score 15/15 | 0
pulse rate 78/min | 0
respiratory rate 13/min | 0
blood pressure 113/54 mm Hg | 0
SpO2 100% in air | 0
left hip tenderness | 0
no ecchymosis to the abdomen | 0
no ecchymosis to the flank | 0
no ecchymosis to the thigh | 0
radiograph of pelvis | 0
undisplaced fracture of left acetabulum | 0
fracture of anterior column | 0
fracture of posterior column | 0
blood tests confirmed liver dysfunction | 0
pH 7.271 | 0
base excess minus 7.3 | 0
PT 18.2 | 0
INR 1.5 | 0
APTT ratio 1.42 | 0
platelets 73 | 0
bilirubin 63 mmol/l | 0
Hb 124 g/l | 0
18 g intravenous cannula insertion | 0
warmed Hartmanns one litre infusion commenced | 0
referred to Orthopaedic on call team | 0
initial delay due to pressure in Emergency department | 0
blood pressure dropped to 75/51 mm Hg | -unknown
tachycardic | -unknown
serum lactate 9 mmol/l | -unknown
FAST examination | -unknown
intraabdominal fluid | -unknown
decompensated liver disease | -unknown
low energy fall | -unknown
haemorrhagic shock not considered | -unknown
treated for sepsis in Emergency department | -unknown
intensive care attendance | -unknown
orthopaedic attendance | -unknown
general registrar attendance | -unknown
pH 7.227 | -unknown
base excess −17.9 | -unknown
serum lactate 16.3 mmol/l | -unknown
Hb 75 g/l | -unknown
arterial blood pressure 90/60 mm Hg | -unknown
pulse rate 90/min | -unknown
left lower abdominal quadrant swelling | -unknown
upper thigh swelling | -unknown
ecchymosis | -unknown
diagnosis of haemorrhagic shock | -unknown
massive transfusion pathway activation | -unknown
transfusion of 4 units of Blood | -unknown
transfusion of 4 units of FFP | -unknown
transfusion of 2 adult therapeutic doses of platelets | -unknown
transfusion of 10 units of cryoprecipitate | -unknown
noradrenaline infusion | -unknown
pelvic binder in place | -unknown
pelvic binder not tightened | -unknown
lateral compression injury | -unknown
CT scan deemed necessary | -unknown
on call radiology team attendance | -unknown
vascular surgeons attendance | -unknown
CT abdomen confirmed fracture of left acetabulum | -unknown
significant haematoma on left pelvic sidewall | -unknown
8 mm enhancing nodule suggestive of internal iliac artery pseudoaneurysm | -unknown
ill-defined blush of contrast within haematoma | -unknown
extra-peritoneal haematoma inseparable from bladder | -unknown
cirrhotic liver | -unknown
incidental 6.7 cm infra-renal aortic aneurysm | -unknown
transfer to intensive care unit | -unknown
further stabilization | -unknown
invasive cardiovascular monitoring | -unknown
CT Angiogram next morning | 24
no arterial bleed | 24
discussion with vascular team | 24
further review of images | 24
recommended for prophylactic embolization | 24
gelfoam embolization of anterior division segmental branches of left internal iliac artery | 48
gelfoam embolization of posterior division segmental branches of left internal iliac artery | 48
consultation with regional pelvic surgeon | 48
10 lb skeletal traction application | 48
discharged to orthopaedic ward after 5 days in ICU | 120
uncontrollable bleeding from pin site | -unknown
skeletal traction removal | -unknown
continuous pressure applied to wound | -unknown
died | 1224
chronic liver disease | 1224
print(f"{event[0]} | {event[1]}")
