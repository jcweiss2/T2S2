23 years old | 0\
male | 0\
history of methicillin-resistant Staphylococcus aureus (MRSA) impetigo at the forearm | -8760\
right tibia fracture | -8760\
treated with intramedullary fixation (IMN) | -8760\
interlocking screws removed | -8760\
skin irritation | -8760\
pain | -8760\
redness and swelling at the surgical site | -336\
diagnosed with stitch abscess | -336\
cultures from the surgical site were positive for MRSA | -336\
oral antibiotic treatment | -336\
fever | -168\
right groin pain | -168\
viral infection | -168\
systemic fever | -168\
myalgia | -168\
difficult and painful ambulation | -168\
right forearm cellulitis | -168\
right sudden onset uveitis | -168\
systemic rash | -168\
right hip lymphadenopathy | -168\
increased CRP | -168\
increased WBC count | -168\
elevated hepatic enzymes | -168\
elevated lactic dehydrogenase (LDH) | -168\
elevated creatine phosphokinase (CPK) levels | -168\
radiograph of both hips in anterior-posterior view was unremarkable | -168\
intravenous (IV) antibiotics | -168\
deterioration | -168\
positron emission tomography-computed tomography (PET-CT) scan | -168\
OIM abscess with systemic manifestations | -168\
blood cultures were positive for MRSA bacteria | -168\
hemodynamic deterioration | -168\
fulminant MRSA sepsis | -168\
admitted to the intensive care unit (ICU) | -168\
ultrasound-guided drainage | -168\
full-body CT scan | -120\
enlargement of the abscesses diameter | -120\
persistent fever | -120\
elevated CRP level | -120\
elevated WBC count | -120\
consulting the orthopaedic team | -120\
surgical intervention | -120\
surgical plan | -120\
combined approach of Smith-Peterson and modified Stoppa | -120\
surgery | 0\
improving general condition | 24\
less frequent fever spikes | 24\
decrease in CRP and WBC levels | 24\
additional antibiotic treatment | 24\
almost complete recovery | 336\
able to ambulate normally | 336\
no pain | 336\
no functional limitations | 336\
returned to daily activities | 336