21 years old | 0
lady | 0
presented to emergency department | 0
shock | 0
respiratory distress | 0
vague abdominal discomfort | -336
abdominal distension | -336
suspicion of abdominal sepsis | 0
fever | 0
cough | 0
breathing difficulty | 0
loose stools | -672
reported from red zone area | -672
IgM/IgG rapid test | 0
negative IgM/IgG rapid test | 0
abdominal examination revealed peritonism | 0
bowel sounds normal | 0
intubated | 0
mechanical ventilation | 0
ionotropic support | 0
coronavirus disease ICU | 0
RT-PCR test | 0
positive RT-PCR | 0
haemoglobin 7.2 g/dl | 0
total leucocyte count 16 ×109/L | 0
platelet count 99 ×109/L | 0
ultrasound abdomen showed large thick-walled collection | 0
percutaneous pigtail drainage | 0
purulent output | 0
chest X-ray showed bilateral lower lobe atelectasis | 0
prominent bronchovascular markings | 0
stabilisation of blood pressure | 0
CECT thorax | 0
bilateral basal atelectasis | 0
ground-glass opacities | 0
CO-RADS score 4 | 0
CECT abdomen reported sealed off perforation | 0
localized large pelvic collection | 0
diagnosis of sealed off enteric perforation | 0
suspicion of severe acute SARS-CoV-2 | 0
exploratory laparotomy | 0
faecopurulent peritoneal collection | 0
dense interbowel adhesions | 0
greater omentum smeared to clumped bowel loops | 0
adhesiolysis | 0
five perforations in distal ileum | 0
jejunal perforation near duodenojejunal junction | 0
perforations repaired | 0
loop ileostomy created | 0
loop ileostomy technically challenging | 0
short broad mesentery | 0
friable inflamed bowel | 0
small bowel mesentery mobilised | 0
oversized abdominal wall defect | 0
flush to skin loop ileostomy fashioned | 0
nasojejunal tube inserted | 0
tip negotiated beyond repaired jejunal perforation | 0
repeat second COVID-19 RT-PCR test | 120
negative RT-PCR | 120
stomal viability assessed by pinprick test | 120
fresh blood | 120
lubricated transparent tube inserted | 120
pink mucosa on torch illumination | 120
nasojejunal tube feeding started | 48
HPE report showed granulomatous inflammation | 120
Ziehl-Neelsen staining demonstrated acid-fast bacilli | 120
possibility of pulmonary tuberculosis | 120
sputum examination | 120
no acid-fast bacilli | 120
GenXpert-Mtb/Rif test | 120
detected Mycobacterium tuberculosis | 120
diagnosis of disseminated tuberculosis | 120
anti-tubercular regime started | 120
low output enterocutaneous fistula | 168
midline wound | 168
managed conservatively | 168
sepsis subsided | 336
accepted oral feeds | 336
nasojejunal tube removed | 336
