3 years old | 0
female | 0
no significant past medical problems | 0
unknown immunization history | 0
dry cough | -336
dyspnea | -336
no fever | -336
no upper respiratory tract infection | -336
weight loss | -168
progressive fatigue | -168
admitted to local hospital | -48
weakness of both lower limbs | -48
inability to walk | -24
flaccid weakness of lower limbs | -24
dyspnea worsened | -24
central cyanosis | -24
referred to tertiary center | 0
severely dyspneic | 0
central cyanosis | 0
respiratory rate of 50 cycles/minute | 0
SpO2 of 85% on room air | 0
loss of sphincter control | 0
bladder palpable | 0
catheterization | 0
supraclavicular lymph nodes | 0
poor air entry in right lung | 0
flaccid paraparesis | 0
loss of tone and reflexes | 0
equivocal Babinski reflex | 0
opsoclonus-myoclonus movement | 0
normal pupils | 0
ventilated with SMV | 0
normal serum electrolyte levels | 0
respiratory acidosis | 0
MRI showed large right posterio-superior mediastinal mass | 0
heterogeneous enhancement | 0
pleural effusion | 0
direct invasion of dorsal spine | 0
canal stenosis | 0
liver normal | 0
no metastasis | 0
whole-spine MRI showed extension of tumor | 0
high levels of urine VMA | 0
bone marrow biopsy confirmed neuroblastoma | 0
thoracotomy | 24
total resection of mass | 24
spinal decompression | 24
relief of canal stenosis | 24
pedicle screw instrumentation | 24
histopathological examination detected poorly differentiated neuroblastoma | 48
supraclavicular lymph node biopsy detected neuroblastoma | 48
high-risk neuroblastoma | 48
postoperative period passed smoothly | 72
improvement of dyspnea | 72
weaning from ventilator | 72
residual lower limb weakness | 72
opsoclonus myoclonus eye movement | 72
loss of bladder control | 72
induction chemotherapy | 96
cyclophosphamide | 96
etoposide | 96
vincristine | 96
died during induction phase | 168
severe pancytopenia | 168
overwhelming septicemia | 168
renal impairment | 168