26 years old | 0
male | 0
inflammatory bowel disease | -672
ulcerative colitis | -672
admitted to the acute surgical unit | 0
folliculitis | 0
multiple carbuncles | 0
debridement | 0
wound management | 0
tachycardic | 24
hypotensive | 24
vasopressor support | 24
ICU admission | 24
broad-spectrum antibiotics | 24
steroid therapy | 48
multi-organ dysfunction | 48
creatinine of 125 µmol/L | 48
mild ALT rise | 48
INR of 1.8 | 48
pancytopenia | 48
increasing oxygen requirements | 48
negative growth on blood cultures | 48
negative growth on wound swabs | 48
negative QuantiFERON assay | 48
negative treponemal serology | 48
negative HIV | 48
negative hepatitis serology | 48
negative acid-fast bacilli | 48
negative fungal elements | 48
central chest histology showed severe active inflammation | 48
large numbers of neutrophils | 48
leucocytes | 48
necrosis | 48
microabscess formation | 48
no organisms identified | 48
lesions continued to heal well with steroid therapy | 96
almost complete resolution at ∼2 months of follow-up | 1440
discharged | 1440