42 years old | 0
gravida 7 | 0
para 4 | 0
mechanical mitral valve replacement | 0
reduced fetal movement | 0
no history of trauma | 0
enoxaparin 80 mg twice daily | -560
switched to warfarin 10 mg/day | -280
warfarin | -280
INR 4.7 | 0
prothrombin time 49 s | 0
activated partial thromboplastin time 44 s | 0
fibrinogen 3.4 g/L | 0
platelets 309,000/mL | 0
hemoglobin 9 g/dL | 0
cardiotocography demonstrated instability of fetal heart rate | 0
ultrasound revealed crescent hyperechoic collection | 0
SDH | 0
emergency cesarean section | 0
warfarin stopped 36 h prior to the surgery | -36
baby born non-vigorous | 0
no respiratory effort | 0
pale | 0
heart rate 40 BPM | 0
resuscitation | 0
bagging for 30 s | 0
heart rate increased to >100 BPM | 0
no breathing | 0
intubated at 1 min of age | 0
oxygen saturation 72-82% | 0
poor perfusion | 0
pale color | 0
umbilical venous catheter inserted | 0
bolus of normal saline administered | 0
blood transfusion | 0
Apgar score 2, 5, 6, and 8 | 0
surfactant given | 0
oxygen saturation improved | 0
fraction of inspired oxygen 21% | 0
transferred to the neonatal intensive care unit | 0
stable condition | 0
birthweight 2,010 g | 0
length 43 cm | 0
head circumference 31 cm | 0
bulged anterior fontanelle | 0
swelling in the right scrotum | 0
capillary blood gas revealed pH 7.11 | 0
PCO2 58 mm Hg | 0
base excess −11.6 mmol/L | 0
bicarbonate 18.4 mmol/L | 0
complete blood count with hematological profile | 0
hemoglobin 10.4 g/dL | 0
platelets 119,000/mL | 0
INR 3.7 | 0
prothrombin time 38.8 s | 0
activated partial thromboplastin time 71.9 s | 0
vitamin K prophylaxis | 0
brain ultrasound on day 1 of life | 24
crescent shape hypoechoic collection | 24
SDH | 24
layering of the hematoma | 24
clotted blood | 24
no midline shift or ventricular dilatation | 24
ultrasound for testes on day 1 of life | 24
large turbid fluid collection | 24
hemorrhagic fluid | 24
normal appearance and perfusion of both testes | 24
computed tomography scan of the head on day 2 of life | 48
bilateral SDH | 48
subarachnoid hemorrhage | 48
diffuse brain edema | 48
midline structures shifted at least 6 mm to the right | 48
brain ultrasound at 20 days of life | 480
large subacute/chronic SDH | 480
midline shift to the right side | 480
cystic changes involving both cerebral hemispheres | 480
PVL | 480
cephalomalacia | 480
dilated lateral ventricles | 480
MRI at 24 days of life | 576
large bilateral acute on subacute SDH | 576
encephalomalacic changes | 576
cerebral hemispheres | 576
basal ganglionic region | 576
frontotemporal area | 576
posterior fossa structures | 576
conservative management | 0
no seizure activity | 0
no evidence of hydrocephalus | 0
right scrotal hemorrhage self-resolved | 336
late onset sepsis | 336
urine culture positive for Klebsiella pneumoniae | 336
antibiotics for 2 weeks | 336
discharged at 4 weeks of age | 672
spastic quadriplegic cerebral palsy | 8760
gross motor function classification system level 5 | 8760
kyphotic posture | 8760
severe global delays | 8760
no grasp | 8760
blindness | 8760
non-recognized speech | 8760