47 years old | 0
    nulliparous woman | 0
    two-week history of increasing abdominal girth | -336
    two-day history of fever | -48
    brought to the Accident and Emergency department | 0
    no previous significant medical or surgical history | 0
    nonsmoker | 0
    in a stable relationship | 0
    no history of sexually transmitted disease | 0
    never used an intra-uterine copper device | 0
    no previous gynecological problems | 0
    temperature 38.5 C | 0
    pulse 113 beats per minute | 0
    blood pressure 76/46 mm Hg | 0
    pale | 0
    clammy | 0
    cachectic | 0
    abdomen grossly distended | 0
    abdomen tense | 0
    large mass felt on the right side | 0
    whole abdomen generally tender | 0
    bowel sound not audible | 0
    large umbilical hernia noted | 0
    hemoglobin 7.8 g/dl | 0
    WBC 21.7 | 0
    CRP 205 | 0
    chest X-ray showed clear lung fields | 0
    abdominal X-ray raised possibility of extensive intra-abdominal fluid | 0
    CT showed large ovarian mass 33x23 cm | 0
    CT showed large ascites | 0
    left ureter obstructed | 0
    malignant ovarian mass | 0
    super imposed infection | 0
    started on cefuroxime | 0
    started on Metronidazole | 0
    laparotomy performed | 0
    total abdominal hysterectomy (TAH) | 0
    bilateral salpingo-oophorectomy (BSO) | 0
    repair of umbilical hernia | 0
    midline laparotomy performed | 0
    six liters of pus aspirated from abdominal cavity | 0
    large cystic mass originating from right adnexa | 0
    extending to the right hemi diaphragm | 0
    both tubes edematous | 0
    five liters of thick pus drained from ovarian cyst | 0
    necrosis inside the cavity wall | 0
    uterus large with multiple fibroids | 0
    fibroids measuring approximately 20 weeks of gestation | 0
    subtotal (supra cervical) hysterectomy | 0
    left ovary adherent to posterior pelvic wall | 0
    endometriotic cysts | 0
    left ovary removed as much as possible | 0
    hernial sac excised | 0
    hernia repaired | 0
    no apparent bowel perforation | 0
    appendix normal | 0
    abdominal wash out with saline performed | 0
    two drains inserted | 0
    mass closure of the abdomen performed | 0
    estimated blood loss one liter | 0
    admitted to intensive care | 0
    maximum ventilatory support | 0
    inotropic cardiac support | 0
    received six units of blood transfusion | 72
    decision of early tracheostomy | 48
    pus culture grew Bacteroides fragilis | 0
    no other bacteria grew from blood or pus culture | 0
    Mycobacterium species not grew from blood or pus culture | 0
    antibiotics changed to Tazocine 4.5g TDS | 72
    inflammatory markers rising | 72
    apyrexial after laparotomy | 0
    remained on antibiotics for 10 days | 0
    histology confirmed multiple fibroids | 0
    right ovarian cyst wall showed marked inflammation | 0
    glandular foci in cyst wall representing endometriosis origin | 0
    endometriosis identified on ovary surface | 0
    endometriotic cyst confirmed in left ovary | 0
    CRP 33 on fourth postoperative day | 96
    good recovery | 336
    discharged home on 14th postoperative day | 336
    primary infertility | 0
    acute abdomen | 0
    peritonitis | 0
    sepsis | 0
    symptoms that brought patient to emergency department | 0
    