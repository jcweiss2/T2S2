66 years old | 0
male | 0
presented to the emergency department | 0
dyspnea | -168
chest pain | -168
body temperature 38.6°C | 0
heart rate 140 beats/min | 0
blood pressure 75/36 mm Hg | 0
respiratory rate 26 breaths/min | 0
oxygen saturation 92% | 0
respiratory distress | 0
accessory muscle use | 0
erythema over the sternum | 0
pitting edema in both lower extremities | 0
feet cool to touch | 0
rapid heart rate | 0
regular rhythm | 0
soft systolic murmur | 0
jugular venous distension | 0
pulsus paradoxus | 0
tachypnea | 0
clear lung auscultation | 0
aortic stenosis | 0
surgical mechanical aortic valve replacement | -504
chronic obstructive pulmonary disease | 0
cirrhosis | 0
hypertension | 0
hyperlipidemia |# | 0
septic shock | 0
sternal wound infection | 0
endocarditis | 0
cardiogenic shock | 0
tamponade | 0
postpericardiotomy syndrome | 0
postsurgical bleed | 0
warfarin anticoagulation | -504
bacterial pneumonia | 0
viral pneumonia | 0
acute coronary syndrome | 0
pneumothorax | 0
pulmonary embolism | 0
acute heart failure exacerbation | 0
chronic obstructive pulmonary disease exacerbation | 0
pericardial effusion | 0
tamponade physiology | 0
pericardiocentesis | 0
hemopericardium | 0
hemodynamic improvement | 0
pericardial effusion decreased | 0
pericardial effusion reaccumulated | 24
pericardial drain | 0
suspected ongoing bleeding | 0
elevated international normalized ratio | 0
fresh frozen plasma | 0
vitamin K | 0
admitted to cardiac intensive care unit | 0
vasopressor support | 0
sternal erythema | 0
fever | 0
blood cultures | 0
pericardial cultures | 0
broad-spectrum antibiotics | 0
chest CT | 48
mid to lower sternotomy wound dehiscence | 0
broken sternal wires | 0
fractured wire penetrated pericardium | 0
RV free wall injury | 0
intubated | 48
surgical exploration | 48
RV free wall laceration | 48
hypotension | 0
shock | 0
blood cultures positive for Staphylococcus aureus | 48
pericardial cultures positive for Staphylococcus aureus | 48
sternal osteomyelitis | 48
ongoing shock | 48
acute kidney injury | 48
acute liver injury | 48
purulent exudate from sternal wound | 48
repeat sternal debridement | 72
nonhealing sternal wound | 336
blood cultures positive | 336
TEE | 336
vegetation on mitral valve | 336
endocarditis | 336
comfort care | 336
passed away | 336
RV free wall injury confirmed | 336
infective endocarditis | 336
