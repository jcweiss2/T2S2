18 years old | 0
female | 0
severe headache | -72
projectile vomiting | -72
no history of fever | -72
no history of convulsions | -72
no history of focal neurological deficit | -72
treated symptomatically | -72
metabolic encephalopathy | 0
symptomatic treatment | 0
deteriorated | 12
altered sensorium | 12
Glasgow Coma Scale-9 | 12
high-grade fever | 12
chills | 12
dyselectrolytemia | 12
serum potassium 3.7 mEq/L | 12
low serum phosphate | 12
serum phosphate 1.57 mg/dL | 12
neutrophilic leukocytosis | 12
total leukocyte count 24,170/μl | 12
neutrophils 91% | 12
cerebrospinal fluid sent for evaluation | 12
ceftriaxone | 12
Gram stain of the centrifuged deposit of CSF | 12
polymorphs and lymphocytes with Gram-positive bacilli | 12
Listeria monocytogenes | 12
culture of CSF | 12
Gram-positive bacilli | 12
diphtheroids | 12
Listeria monocytogenes | 24
meropenem | 24
corrective measures | 24
clinical improvement | 48
microbiological improvement | 48
Listeria monocytogenes identified by conventional methods | 48
Listeria monocytogenes identified by automated methods | 48
VITEK-2, Biomerieux | 48
healthy young female | 48
preexisting illness | 48
prolonged medication | 48
meningitis by Listeria monocytogenes | 48
lower incidence of meningeal signs | 48
dyselectrolytemia | 48
meningeal signs | 48
Gram stain occurs singly or in pairs | 48
diphtheroids or diplococci | 48
proper diagnosis and treatment | 48