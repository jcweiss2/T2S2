57 years old | 0
female | 0
visited the trauma and emergency department | 0
history of falling | -24
sudden onset of weakness | -72
nausea | -72
vomiting | -72
diarrhea | -72
known smoker | 0
obese | 0
uncontrolled hypothyroidism | 0
leukocytosis | 0
lymphopenia | 0
thrombocytopenia | 0
deteriorated renal function | 0
hyperglycemic hyperosmolar nonketotic state | 0
blood urea 78 mg/dl | 0
serum creatinine 3.1 mg/dl | 0
glycosuria | 0
pyuria | 0
negative results for ketones | 0
blood glucose concentration 1680 mg/dl | 0
glycated hemoglobin 16.3% | 0
diagnosed with hyperglycemic hyperosmolar non-ketotic state | 0
arterial blood gases revealed normal pH | 0
serum osmolarity 335 mosm/lt | 0
C reactive protein 43.2 mg/dl | 0
procalcitonin 56.34 ng/ml | 0
afebrile | 0
vital signs were stable | 0
vigorous intravenous hydration | 0
insulin infusion pump | 0
sedated and intubated | 12
injection ceftriaxone 2 g qDay intravenously | 12
clindamycin 1.8 g/day IV divided q8hr | 12
abdominal and pelvic CT scan | 12
gas within the left kidney | 12
infiltration of septa in the perirenal space | 12
moderate intraosseous gas within the L3 and L4 lumbar vertebral bodies | 12
emphysema in the epidural space | 12
diagnosed with emphysematous pyelonephritis | 12
diagnosed with emphysematous osteomyelitis of the spine | 12
Klebsiella pneumoniae identified in urine culture | 12
antibiotic therapy changed to meropenem 1 g iv q8hr | 12
septic shock | 24
multiple organ dysfunction | 24
died | 48
emphysematous pyelonephritis | 12
emphysematous osteomyelitis of spine | 12