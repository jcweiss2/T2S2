62 years old | 0
male | 0
admitted to the hospital | 0
high fever | 0
dark urine | 0
lumbar vertebral injury | -8760
paralyzed | -8760
sacrococcygeal bedsores | -8760
debridement | -8760
muscle flap application | -8760
repeated dehiscence | -216
exudation of wounds | -216
infected wound | 0
amyotrophy of both lower limbs | 0
disappearance of cutaneous expression of sensation | 0
elevated CK level | 0
debridement | 24
intraoperative exploration | 24
necrotic tissue removal | 24
frequent dressing changes | 24
antimicrobial therapy | 24
correction of electrolyte imbalances | 24
correction of acidosis | 24
nutritional support | 24
suture area dry and clean | 72
dark urine lightened | 24
fever resolved | 72
CK level peaked | 24
CK level decreased | 120
CK level returned to normal | 216
white blood cell count decreased | 168
white blood cell count returned to normal | 168
C-reactive protein concentration decreased | 264
C-reactive protein concentration returned to normal | 264
wound healed | 720
discharged | 720