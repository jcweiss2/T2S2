51 years old | 0
    female | 0
    visited to receive total hip arthroplasty | 0
    osteoarthritis | 0
    acetabular dysplasia | 0
    left hip joint | 0
    no special findings in personal medical history | 0
    no recent physical examination findings | 0
    no chest X-ray findings | 0
    no electrocardiogram findings | 0
    no blood test findings before surgery | 0
    famotidine administered | 0
    glycopyrrolate administered | 0
    intramuscular administration | 0
    spinal block | 0
    bupivacaine injected into subarachnoid space | 0
    lack of sensation in 9th thoracic vertebrae | 0
    midazolam injected | 0
    oxygen administered through face mask | 0
    anesthesia duration approximately two hours | 0
    blood loss 400 ml | 0
    fluid administered 2,100 ml | 0
    urine output 950 ml | 0
    arterial blood gas analysis | 0
    pH 7.386 | 0
    PaCO2 42.5 mmHg | 0
    PaO2 164.7 mmHg | 0
    HCO3 24.6 mM/L | 0
    SaO2 99.8% | 0
    Hb 10.1 g/dl | 0
    blood pressure 110/60 mmHg | 0
    heart rate 65 beats/min | 0
    pulse oximetry 99% | 0
    cold complaint | 0
    shivering | 0
    warm blanket applied | 0
    approximately three hours after arrival in recovery room | 72
    dizziness complaint | 72
    slight cyanosis in lips | 72
    blood test performed | 72
    chemical test performed | 72
    coagulation test performed | 72
    blood pressure 90/50 mmHg | 72
    heart rate 70-95 beats/min | 72
    pulse oximetry 98% | 72
    hemoglobin 7.9 g/dl | 72
    hematocrit 24.3% | 72
    suspected hypovolemia | 72
    central venous catheter insertion decision | 72
    left subclavian catheter insertion | 72
    Trendelenburg position | 72
    left arm internal rotation | 72
    neck turned to the right | 72
    lidocaine administered | 72
    skin punctured with 18 G needle | 72
    J-inducing wire inserted | 72
    expander used | 72
    central venous catheter inserted | 72
    blood aspiration confirmed | 72
    catheter fixed at 15 cm length | 72
    blood pressure 110/60 mmHg | 72
    heart rate 78-100 beats/min | 72
    pulse oximetry 99% | 72
    packed red blood cells injected | 72
    emergency blood test | 72
    50 ml blood drained into Hemovac | 72
    CT decision next morning | 72
    iopromide injected | 96
    contrast medium injection rate 2 ml/s | 96
    total contrast dose 120 ml | 96
    CT abdomen and pelvis | 96
    chest heaviness complaint | 96
    oxygen administered through face mask | 96
    blood pressure 110/66 mmHg | 96
    heart rate 70 beats/min | 96
    arterial blood gas analysis | 96
    pH 7.406 | 96
    PaCO2 36.8 mmHg | 96
    PaO2 109.6 mmHg | 96
    HCO3-11.5 mM/L | 96
    SaO2 99.3% | 96
    no electrocardiogram findings | 96
    no echo cardiogram findings | 96
    no cardiac enzyme test findings | 96
    no allergic reaction signs | 96
    chest X-ray | 96
    central venous catheter tip at brachiocephalic vein | 96
    hydrothorax observed on CT | 96
    hydrothorax detection at radiology department | 96
    Chiba needle inserted | 96
    100 ml pleural effusion drained | 96
    8.5 F pig tail catheter inserted | 96
    transparent fluid aspirated | 96
    contrast medium confirmed | 96
    contrast medium injected through catheter | 96
    vein flow confirmed | 96
    blood suction without resistance | 96
    central venous catheter replacement | 96
    catheter fixed at 20 cm length | 96
    blood aspiration confirmed | 96
    chest X-ray confirmation | 96
    no dyspnea complaint | 96
    no other symptoms | 96
    extracoporeal drainage 20 ml | 96
    chest cavity pig tail catheter insertion | 96
    postoperative observation | 96
    chest X-ray monitoring | 96
    vital signs monitoring | 96
    hydrothorax disappearance | 168
    no side effects | 168
    no cardiopulmonary symptoms | 168
    catheter removed after seven days | 168
    general ward transfer | 168
    discharged after 14 days | 336
