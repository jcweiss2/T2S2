23 years old | 0
    male | 0
    spontaneously delivered at full term | 0
    poor feeding | -72
    decreased tone | -72
    decreased reflexes | -72
    admitted to the neonatal intensive care unit | -72
    sepsis workup | -72
    cranial ultrasonography | -72
    small right-sided choroid plexus cyst | -72
    partial agenesis of corpus collosum | -72
    myoclonic jerks | -72
    hiccups | -72
    lethargy | -72
    unresponsiveness | -72
    central hypotonia | -72
    amino acid analysis of CSF | -72
    amino acid analysis of plasma | -72
    normal liver studies | -72
    normal ammonia level | -72
    negative blood culture | -72
    negative CSF bacterial culture | -72
    negative CSF viral culture | -72
    abnormal electroencephalographic monitoring | -72
    diffuse cortical dysfunction | -72
    partial seizures | -72
    progressive encephalopathy | -72
    respiratory insufficiency | -72
    mechanical ventilation | -144
    MR imaging of the brain | -144
    intraventricular hemorrhage | -144
    partial agenesis of the corpus callosum | -144
    1H-MR spectroscopy | -144
    elevated brain glycine | -144
    elevated glycine peak at 3.55 ppm | -144
    CSF glycine level elevated | -144
    plasma glycine level elevated | -144
    CS-to-plasma glycine ratio elevated | -144
    negative urine organic acid analysis | -144
    treatment with dextromethorphan | -144
    treatment with phenobarbital | -144
    treatment with sodium benzoate | -144
    improved consciousness | -144
    extubation from mechanical ventilation | -360
    decreased plasma glycine concentrations | -360
    periodic plasma glycine elevations | -360
    homozygous GLDC gene mutation | -360
    feeding problems | -360
    poor growth | -360
    recurrent vomiting | -360
    seizures | -360
    