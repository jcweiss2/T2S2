66 years old | 0
male | 0
polycystic kidney disease | 0
polycystic liver disease | 0
kidney dialysis | -8760
admitted to the emergency department | 0
complaining of acute abdominal pain | 0
left flank pain | -168
fever | -168
vomiting | -168
severe diffuse pain | -48
obstipation | -48
temperature of 38, 5°C | 0
enlarged and painful left kidney | 0
diffuse tenderness | 0
purulent urine | 0
white blood count was 10300/mm3 | 0
serum creatinine concentration was 624 μmol/ml | 0
urine culture isolated Escherichia coli | 0
X-ray abdominal exam showed small bowel dilation | 0
enhanced CT scan revealed multiple hepatic cysts | 0
enhanced CT scan revealed bilaterally enlarged polycystic kidneys | 0
communication between heterogenous cyst in left kidney and pericolic space | 0
soft tissue thickening in the left mesocolon | 0
increased amount of peritoneal fluid | 0
diagnosis of peritonitis | 0
laparotomy exploration | 0
generalized peritonitis | 0
purulent collection from a ruptured cyst of a giant polycystic left kidney | 0
peritoneal lavage | 0
drainage after debridement | 0
bacteriol analysis of the collection isolated Escherichia coli | 0
intensive medical support | 0
parenteral antibiotic | 0
septic shock | 72
hemodynamic instability | 72
died on the 3rd post-operative day | 72