8 years old | 0
male | 0
admitted to the hospital | 0
viral prodrome | -168
high fever | -168
malaise | -168
fatigue | -168
anorexia | -168
myalgias | -168
reddish maculopapular skin rashes | -168
pitting edema | -168
pure motor symmetrical progressive weakness | -168
pelvifemoral region muscle pain | -168
flaccid weakness | -120
bedbound | -120
generalized pitting anasarca | -120
normal renal functions | -120
no family history of autoimmune disorders | 0
no Raynaud's phenomenon | 0
no polyarthralgias | 0
no polyarthritis | 0
no bulbar symptomatology | 0
no soft-tissue calcifications | 0
no oral ulceration | 0
flaccid quadriparesis | 0
Grade 1 deep tendon reflexes | 0
diffuse Grade 1/5 Medical Research Council muscular weakness | 0
exquisite pain | 0
symmetric proximal and axial weakness | 0
grotesque pitting swelling | 0
erythematous maculopapular rashes | 0
hypoalbuminemia | 0
hypotension | 0
tachycardia | 0
normal echocardiogram | 0
normal renal functions | 0
normal serum procalcitonin | 0
negative sepsis work up | 0
negative viral serologies | 0
normal complete blood counts | 0
normal serologic tests | 0
normal ANA | 0
normal rheumatoid factor | 0
normal ANA profile | 0
normal perinuclear antineutrophil cytoplasmic antibody | 0
normal cytoplasmic-ANCA | 0
normal antistreptolysin-O titers | 0
normal thyroid functions | 0
normal hepatitis serologies | 0
normal electrocardiography | 0
normal cardiac injury enzymes | 0
normal chest radiography | 0
normal abdominal ultrasonography | 0
elevated creatine phosphokinase | 0
elevated lactate dehydrogenase | 0
rhabdomyolysis | 0
nerve conduction studies normal | 0
electromyography abnormal | 0
increased muscle membrane irritability | 0
low amplitude short duration polyphasic myopathic MUPs | 0
muscle biopsy | 0
Jo-1 IgG antibody positive | 0
anti-Mi2 antibody positive | 0
reduced C3 and C4 complement levels | 0
fulminant SCLS | 0
hemoconcentration | 0
high hematocrit | 0
“shock”-like syndrome | 0
parenteral Tramadol | 0
paracetamol | 0
hemodynamic instability | 0
cardiovascular monitoring | 0
central venous pressure monitoring | 0
aggressive fluid resuscitation | 0
high-dose catecholamine therapy | 0
norepinephrine infusion | 0
pulse methylprednisolone | 24
high-dose intravenous immunoglobulin | 24
theophylline | 24
salbutamol | 24
leukotriene inhibitors | 24
fresh frozen plasma | 24
20% albumin | 24
improvement after 72 hours | 72
immunomodulatory therapy | 72
prednisolone | 72
azathioprine | 72
motoric recovery | 336
amelioration of edema | 336
ambulating | 720
discharged | 720
normal motoric power | 1440
switched to alternate-day glucocorticoid schedule | 1440
reduction of maintenance dose | 1440
taper of prednisolone and azathioprine | 1440
clinical remission | 2880
immunomodulatory therapy tapered off | 2880