65 years old | 0
male | 0
admitted to the hospital | 0
weight loss | -2160
lack of appetite | -2160
generalized fatigue | -2160
dehydrated | 0
cachexic | 0
fluid-responsive hemodynamics | 0
heart rate 109 beats per minute | 0
blood pressure 78/54 mm Hg | 0
respiratory rate 17 per min | 0
oxygen saturation 97% on room air | 0
received 3 L of crystalloids | 0
blood pressure rose to 93/69 mm Hg | 0
no stigmata of chronic liver disease | 0
numerous ecchymoses on his extremities | 0
coarse crepitations bilaterally in his lower lung zones | 0
nontender splenomegaly | 0
palpable nonpulsatile firm periumbilical mass | 0
no lymphadenopathy | 0
no scrotal or pedal swelling | 0
anemia | 0
thrombocytopenia | 0
hypoglycemia | 0
severely elevated anion gap metabolic acidosis | 0
hyperlactatemia | 0
aggressive fluid-resuscitation with crystalloids | 0
blood transfusion | 0
broad-spectrum antibiotics | 0
workup for infection was negative | 0
D-lactate level was normal | 0
diffuse cervical-mediastinal lymphadenopathy | 0
nodular consolidative changes in the left upper lobe | 0
mesenteric mass | 0
persistent hypoglycemia | 0
required continuous dextrose infusion | 0
bronchoscopy | 0
gastrointestinal endoscopies | 0
bone marrow aspiration and biopsy | 432
CD20-positive non-Hodgkin's lymphoma | 432
diffuse large B-cell lymphoma | 432
CD10 and cyclin D1 overexpression | 432
lactate levels climbed steadily | 432
encephalopathy | 648
nosocomial pneumonia from aspiration | 648
sepsis | 648
tumor lysis syndrome | 648
multiorgan failure | 648
mechanical intubation | 648
initiation of vasopressors | 648
continuous renal replacement therapy | 648
withdrew care | 648
died | 648