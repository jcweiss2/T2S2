27 years old | 0
woman | 0
acute myeloblastic leukemia | 0
FAB 6 | 0
secondary to myelodysplastic syndrome | 0
normal karyotype | 0
WT1+ | 0
single mutation of CEBPa | 0
mutation TAD1 from CEBPa | 0
no mutation of NMP1 | 0
complete response after induction chemotherapy | 0
received two cycles of high-dose Ara-C | 0
associated with pegfilgrastim | 0
relapsed | -1080
received Ara-C | -1080
received idarubicine | -1080
second complete response | -1080
no HLA-identical unrelated donor identified | -1080
after 12 weeks of research | -1080
haplo-identical allogeneic HSCT from her mother scheduled | -1080
conditioning regimen with fludarabine | 0
conditioning regimen with cyclophosphamide | 0
conditioning regimen with busulfan | 0
conditioning regimen with antithymocyte globulin | 0
conditioning regimen with cyclophosphamide post graft infusion | 0
GvHD prophylaxis with tacrolimus | 0
GvHD prophylaxis with mycophenolate mofetil | 0
stem cell source PBSC with 4.32×10e6 CD34+/kg | 0
recipient CMV+ | 0
recipient HSV+ | 0
recipient HHV6+ | 0
recipient TOXO+ | 0
recipient EBV+ | 0
recipient VZV+ | 0
transplantation not complicated except SOS | 0
SOS treated with diuretics | 0
SOS treated with ursodeoxycholic acid | 0
tacrolimus stopped at day 21 | 504
developed schizocytes | 504
MMF continued alone | 504
MMF progressive tapering | 504
aim to stop MMF at 6 months after transplantation | 504
hematological recuperation on day 18 | 432
chimerism 100% donor on PB | 432
chimerism 100% donor on BM | 432
discharged on day 27 after transplantation | 648
during first three months of follow-up | 2160
EBV PCR examined | 2160
HHV6 PCR examined | 2160
Toxoplasmosis PCR examined | 2160
CMV PCR examined | 2160
ADV PCR examined | 2160
received monthly serum immunoglobulin | 2160
CMV reactivation at day 56 | 1344
treated with valgancyclovir | 1344
during 6 weeks | 1344
routine follow-up at 3 months after transplantation | 2160
no evidence of relapse | 2160
chimerism 100% donor on PB | 2160
chimerism 100% donor on BM | 2160
blood tests showed CD3 count:16×10e3/mm3 | 2160
CD4 count: 4×10e3/mm3 | 2160
CD8 count: 12×10e3/mm3 | 2160
CD4:CD8 ratio of 0.33 | 2160
IgG:9.07 g/L | 2160
IgA 0.59 g/L | 2160
IgM 0.08 g/L | 2160
Hg 8.1 g/dL | 2160
WC count:2.0×10e3/mm3 | 2160
neutro 1.61×10e3/mm3 | 2160
Platelets count:89×10e3/mm3 | 2160
collect donor lymphocytes | 2160
second CMV reactivation occurred on day 121 | 2904
treated with valgancyclovir | 2904
dose reduced after 1 week | 2904
developed severe toxic pancytopenia | 2904
Hg:7.0 g/dL | 2904
neutro:0.5 G/L | 2904
Plat 30×10e3/mm3 | 2904
started G-CSF three times a week | 2904
received serum immunoglobulin weekly | 2904
DLI of 1×10e5 CD3+/kg administrated on day 134 | 3216
admitted with fever | 3384
fever 38.5° | 3384
nausea | 3384
vomiting | 3384
loss of weight | 3384
loss of appetite | 3384
severe oral candidiasis | 3384
blood tests showed Hg:9.1 g/dL | 3384
WC:2.7×10e3/mm3 | 3384
Plat:56×10e3/mm3 | 3384
CRP:86 mg/L | 3384
Na:135 mmol/L | 3384
K:3.0 mmol/L | 3384
Protein:67 g/L | 3384
creatinine:1.06 mg/dL | 3384
T Bili:0.2 mg/dL | 3384
D Bili <0.1 mg/dL | 3384
AST:228 U/L | 3384
ALT:136 U/L | 3384
ALP:105 U/L | 3384
gamma GT 75 U/L | 3384
posaconazole stopped | 3384
toxic cause suspected | 3384
ursodeoxycholic acid reintroduced | 3384
improvement in hepatic test | 3384
started Ceftazidim | 3384
started Caspofungin | 3384
gastric fibroscopy with biopsies performed | 3384
developed diarrhea within 48h of admission | 3456
bacteriological stool analyses performed | 3456
viral stool analyses performed | 3456
fungal stool analyses performed | 3456
Ceftazidim replaced by Tazocillin | 3456
Ceftazidim replaced by Metronidazole | 3456
tests for fecal biomarkers performed | 3456
MMF discontinued | 3456
short course of steroids started | 3456
Foscavir started | 3456
CMV PCR two times a week | 3456
number of copies decreased progressively | 3456
no evidence of GvHD on gastric biopsies | 3456
oral candidiasis secondary to Candida albicans confirmed | 3456
chest CT showed hypodense lesions in right liver | 3456
abdominal CT showed hypodense lesions in right liver | 3456
pelvic CT showed hypodense lesions in right liver | 3456
liver biopsy scheduled | 3456
postponed due to sepsis | 3456
sepsis with Staphylococcus hominis | 3552
Vancomycin started | 3552
port pulled | 3552
diarrhea stopped | 3552
no evidence of GvHD | 3552
steroids dose rapidly decreased | 3552
presented rash on 20–25% of corporeal surface | 3696
profuse diarrhea | 3696
biopsies of gut | 3696
biopsies of skin | 3696
steroids reached to 2 mg/kg/day for 4 days | 3696
developed hepatomegaly | 3696
pain | 3696
ascitis | 3696
edema | 3696
fever 40°C | 3696
blood test showed pancytopenia | 3792
severe neutropenia | 3792
severe hepatic cytolysis | 3792
cholestasis | 3792
CMV PCR realized | 3792
EBV PCR realized | 3792
HHV6 PCR realized | 3792
toxoplasmosis PCR realized | 3792
adenovirus PCR realized | 3792
HBV PCR realized | 3792
HCV PCR realized | 3792
BM aspiration realized | 3792
no evidence of haemophagocytosis | 3792
no evidence of viral infection on BM | 3792
signs of myelotoxicity due to drug toxicity | 3792
liver biopsy obtained by transjugular approach | 3816
developed disseminated intravascular coagulation | 3816
continued bleeding in jugular vein | 3816
died from hepatic failure | 3840
death occurred in Intensive Care Department | 3840
PCR for ADV positive | 4320
all other results normal | 4320
chimerism on BM 100% donor | 4320
positive adenovirus immunohistochemistry | 4320
patchy necrosis in perivenular areas | 4320
patchy necrosis in parenchyma | 4320
patchy necrosis in periportal areas | 4320
hepatocytes with nuclear inclusion bodies | 4320
confluent hepatic necrosis due to adenovirus infection | 4320
limited macrophages showing hemophagocytosis | 4320
haplo-identical allogeneic HSCT scheduled | -1080
conditioning regimen | 0
GvHD prophylaxis | 0
stem cell source PBSC | 0
tacrolimus stopped | 504
MMF continued | 504
MMF tapering | 504
hematological recuperation | 432
discharged | 648
EBV PCR | 2160
HHV6 PCR | 2160
Toxoplasmosis PCR | 2160
CMV PCR | 2160
ADV PCR | 2160
monthly serum immunoglobulin | 2160
CMV reactivation | 1344
valgancyclovir treatment | 1344
routine follow-up | 2160
no relapse | 2160
chimerism 100% donor | 2160
blood test results | 2160
donor lymphocytes collection | 2160
second CMV reactivation | 2904
valgancyclovir treatment | 2904
dose reduction | 2904
pancytopenia | 2904
G-CSF started | 2904
weekly immunoglobulin | 2904
DLI administered | 3216
admission with fever | 3384
weight loss | 3384
appetite loss | 3384
oral candidiasis | 3384
blood test results | 3384
hepatic test improvement | 3384
antibiotics started | 3384
gastric fibroscopy | 3384
diarrhea developed | 3456
stool analyses | 3456
antibiotic change | 3456
steroids started | 3456
CMV PCR monitoring | 3456
CMV copies decreased | 3456
no GvHD on biopsies | 3456
Candida albicans confirmed | 3456
CT findings | 3456
sepsis | 3552
Vancomycin | 3552
port removal | 3552
diarrhea resolved | 3552
steroids reduced | 3552
rash | 3696
gut biopsy | 3696
skin biopsy | 3696
steroid increase | 3696
hepatomegaly | 3696
ascites | 3696
high fever | 3696
pancytopenia | 3792
neutropenia | 3792
hepatic cytolysis | 3792
viral PCR tests | 3792
BM aspiration | 3792
no haemophagocytosis | 3792
no viral infection | 3792
drug toxicity signs | 3792
liver biopsy | 3816
DIC | 3816
jugular bleeding | 3816
death | 3840
ADV PCR positive | 4320
other tests normal | 4320
chimerism confirmed | 4320
adenovirus confirmed | 4320
hepatic necrosis | 4320
limited haemophagocytosis | 4320
