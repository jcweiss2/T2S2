59 years old | 0
female | 0
admitted to peripheral hospital | -264
peritonitis | -264
perforation of sigmoid diverticulum | -264
sigmoid resection | -264
L-T anastomosis | -264
new widespread peritonitis | -253
emergency re-laparotomy | -253
dehiscence of posterior wall of anastomosis | -253
fecal contamination of abdomen | -253
ileostomy | -253
toilet of peritoneal cavity | -253
wound margins not juxtaposed | -253
transfer to ICU | -231
sedated | -231
intubated | -231
mechanically ventilated | -231
hemodynamically unstable | -231
invasive blood pressure 80/50 mmHg | -231
body temperature 38°C | -231
dehiscence of cutaneous and subcutaneous abdominal layers | -231
chronic obstructive pulmonary disease | 0
gastro-esophageal reflux disease | 0
paroxysmal atrial fibrillation | 0
culture tests collected | -231
surgical wound swab positive for E. coli | -231
surgical wound swab positive for E. faecius | -231
surgical wound swab positive for Bacteroides Ovatum | -231
blood cultures negative | -231
CT scan of abdomen | -231
free air in peritoneal cavity | -231
multiple confluent abscesses | -231
nodules in chest | -231
ipodense areas within spleen | -231
debridement rejected | -231
conservative treatment proposed | -231
broad-spectrum antibiotic therapy | -231
Negative Pressure Therapy (NTP) | -231
VAC therapy | -231
V.A.C. VeraFlo Cleanse | -231
intermittent cleaning cycles | -231
saline infusion | -231
suction phases | -231
formation of granulation tissue | -28
resolution of septic state | -28
hemodynamic stability | -28
conventional GranuFoam Dressings | -28
tissue repair accelerated | -28
progressive juxtaposition of flaps | -28
discharged from ICU | 35
afebrile | 35
clinically stable | 35
hemodynamically stable | 35
spontaneous breathing | 35
oxygen therapy | 35
normal urine output | 35
VAC therapy continued | 35
complete closure of abdominal wall | 77
alive | 156
no complications | 156