female | 0
3.28 kg | 0
40 weeks gestation | 0
caesarean section | 0
scoliosis | -672
right hydronephrosis | -672
active stagnation | -672
suspected intrauterine infection | -672
fever | -2
amniotomy | -2
IV oxytocin | -2
IV cefuroxime sodium | -2
Apgar score 8/9 | 0
amniotic fluid clear | 0
no meconium staining | 0
severe acute chorioamnionitis | 0
moderate umbilical vasculitis | 0
extensive neutrophilic infiltration | 0
cellulose attachment in villi | 0
groaning | 0
spitting | 0
generalized erythematous papular eruption | 0
transient respiratory distress | 0
low-flow oxygen | 0
decreased transmittance chest X-ray | 0
pustules | 72
desquamation | 72
palms and soles affected | 72
skin scrapings negative for Candida spp | 72
no oral or perianal thrush | 72
increased C-reactive protein | 18
leucocytosis with left shift | 18
lumbar puncture | 18
cerebrospinal fluid culture negative | 18
cerebrospinal fluid white blood cell count 15 cells/mm3 | 18
cerebrospinal fluid protein 63.4 mg/dl | 18
cerebrospinal fluid glucose 2.5 mmol/l | 18
empiric antimicrobial therapy | 18
cefoperazone/sulbactam | 18
penicillin | 18
differential diagnosis | 18
congenital herpes simplex virus | 18
congenital syphilis | 18
streptococcal infection | 18
Listeria monocytogenes infection | 18
candidiasis | 18
skin rash desquamated | 168
excoriated lesions persisted | 168
WBC count normal | 168
CRP levels normal | 168
antibiotics stopped | 168
blood culture positive for C. albicans | 168
urine culture positive for C. albicans | 168
skin culture positive for C. albicans | 168
serum (1–3)-β-D-glucan assay negative | 168
IV fluconazole | 168
topical skin antifungal therapy | 168
miconazole nitrate | 168
high-throughput DNA sequencing | 312
no evidence of fungi, bacteria, or viruses | 312
urine cultures negative | 312
cutaneous lesions resolved | 528
recurrent bacterial UTIs | 528
immune deficiency suspected | 528
blood immunity-related genetic analysis | 528
immune function tests | 528
normal immune function | 528
chronic granulomatous disease/galactosemia excluded | 528
vesicoureteral reflux suspected | 528
voiding cystourethrography not performed | 528
IV vancomycin | 720
urine cultures sterile | 720
urine routine examinations normal | 720
audiometry normal | 720
ophthalmologic examination normal | 720
brain magnetic resonance imaging normal | 384
chest computed tomography normal | 312
liver, renal, and bladder ultrasonography normal | 72
99mTc-DMSA static renal scan normal | 1176
echocardiogram | 72
small atrial septal defect | 72
patent foramen ovale | 72
no endocarditis | 72
discharged | 1488
good development | 1488