43 years old | 0
woman | 0
sought medical attention | 0
abdominal pain | -720
lumbar pain | -720
nausea | -720
nonproductive retching | -720
denied fever | 0
symptoms over the past month | -720
progressively worsened | -720
over-the-counter painkillers | -720
cesarean sections | 0
cholecystectomy | 0
hiatoplasty | -52560
hiatal hernia | -52560
ill-looking appearance | 0
pained expression | 0
pale | 0
anicteric | 0
afebrile | 0
normal respiratory pattern | 0
blood pressure 124/82 mmHg | 0
pulse 84 bpm | 0
respiratory rate 20 rpm | 0
room air oximetry 98% | 0
thoracic kyphosis | 0
painful abdominal palpation | 0
negative rebound tenderness | 0
normal bowel sounds | 0
hemoglobin 15.8 g% | 0
creatinine 1.09 mg/dL | 0
hematocrit 48.9% | 0
potassium 3.8 mEq/L | 0
leucocytes 18.4 ×10³/mm³ | 0
sodium 140 mEq/L | 0
bands 0% | 0
ALT 20 U/L | 0
segmented 84% | 0
AST 35 U/L | 0
eosinophil 0% | 0
total bilirubin 0.5 mg/dL | 0
basophil 0% | 0
glucose 178 mg/dL | 0
lymphocyte 9% | 0
amylase 859 U/L | 0
monocyte 7% | 0
lipase 1038 U/L | 0
platelets 265×10³/mm³ | 0
Cai+ 1.06 mmol/L | 0
CRP 180 mg/L | 0
PT INR 1.59 | 0
urea 51 mg/dL | 0
abdominal computed tomography | 0
gastric volvulus | 0
intrathoracic stomach | 0
organoaxial rotation | 0
mesenteroaxial rotation | 0
splenic arteriovenous vascular pedicle displacement | 0
pancreatic tail displacement | 0
tachypnea | 24
decreased oxygen saturation | 24
hypotension | 24
exploratory laparotomy | 24
stomach herniation into chest | 24
gastric volvulus with necrosis | 24
gastric perforation | 24
gastro enteric contents in left pleural cavity | 24
stomach reduction | 24
vertical gastrectomy | 24
thoracic drainage | 24
mediastinal drainage | 24
intensive care unit admission | 24
sedation | 24
mechanical ventilatory support | 24
norepinephrine infusion | 24
hemodynamic stabilization | 24
multiple organ failure | 48
death | 48
foul-smelling enteric liquid in pleural cavity | 48
thick brownish fibrinous material | 48
right lung 403 g | 48
left lung 518 g | 48
wine-colored lung surfaces | 48
congestion | 48
edema | 48
alveolar hemorrhage | 48
pneumonia | 48
diffuse alveolar damage | 48
focal thrombosis | 48
infarction of subpleural parenchyma | 48
acute pleurisy | 48
food debris in pleura | 48
petechiae on pericardial surface | 48
chronic myocarditis | 48
diaphragm laceration | 48
gastric serositis | 48
acute pancreatitis | 48
steatonecrosis | 48
liver congestion | 48
lobular necrosis | 48
microvesicular steatosis | 48
acute tubular necrosis | 48
mucosal hemorrhage | 48
submucosal hemorrhage | 48
potassium 3.8 mEq/L |(Note: This is the correct thinking process.)
