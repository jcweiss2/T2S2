14 years old | 0
girl | 0
diagnosed with ALL | -672
started on induction chemotherapy | -672
Vincristine | -672
Daunorubicin | -672
Prednisone | -672
PEG-Asparaginase | -672
routine outpatient laboratory studies | -24
pancytopenia | -24
absolute neutrophil count of 210/mm3 | -24
developed acute-onset left-lower-extremity pain | -18
presented to the emergency department | -18
worsening bilateral leg pain | -14
worsening hip pain | -14
worsening back pain | -14
progressive weakness of both lower extremities | -14
inability to bear weight | -14
tachycardic | -14
febrile | -14
hypotensive | -14
systolic pressures in the low 80s | -14
physical exam demonstrated nonspecific swelling | -14
significant tenderness of the left thigh | -14
initial laboratory studies confirmed pancytopenia | -14
decreased platelet count (37,000/mm3) | -14
low fibrinogen (78 mg/dL) | -14
elevated thrombin time (19 seconds) | -14
IV fluid bolus | -14
started on gentamycin | -14
started on ceftazadime | -14
left-lower-extremity Doppler ultrasound examination | -14
deep venous thrombosis excluded | -14
acute onset of thigh pain | -14
rapidly developing sepsis | -14
neutropenia | -14
laboratory studies suggestive of disseminated intravascular coagulation | -14
necrotizing deep3soft-tissue infection considered | -14
General Surgery service consulted | -14
inability to localize area of involvement | -14
patient unable to localize specific muscle compartment | -14
altered mental status | -14
cross-sectional imaging performed | -14
CT revealed intramuscular gas | -14
intramuscular gas within multiple muscle compartments | -14
involved muscle compartments identified | -14
blood cultures demonstrated Clostridium perfringens | -14
brought emergently to the operating room | -14
exploration and debridement of necrotizing soft-tissue infection | -14
extensive longitudinal incisions made | -14
access to medial and lateral thigh compartments | -14
access to posterior compartment of the calf and hemipelvis | -14
skin intact | -14
subcutaneous tissue intact | -14
superficial fascia intact | -14
good blood supply | -14
entrance into deep muscle compartments | -14
sweet foul-smelling liquefactive necrosis encountered | -14
myonecrosis confirmed | -14
adductor magnus involved | -14
adductor brevis involved | -14
gracilis involved | -14
gastrocnemius involved | -14
posterior hamstrings involved | -14
muscle bellies debrided | -14
large defects in muscle groups | -14
brought to the Intensive Care Unit | -14
serial washouts performed | 0
further debridement performed | 0
postoperative day 4 | 96
wound bed adequately debrided | 96
Vacuum-Assisted Closure device applied | 96
nonviable skin and subcutaneous tissue excised | 96
no sensory function below either knee | 96
no voluntary motor function below either knee | 96
bilateral above-knee amputations | 96
pedicled myocutaneous flaps based on popliteal artery | 96
transferred to surgical floor | 96
wounds healed well | 96
began physical therapy | 96
rehabilitation initiated | 96
short-interval followup of two months | 1344
