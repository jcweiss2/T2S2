76 years old | 0
    Caucasian | 0
    man | 0
    hypertension | 0
    type two diabetes mellitus | 0
    stage four chronic kidney disease | 0
    obstructive sleep apnoea | 0
    previous pacemaker insertion | 0
    symptomatic bradycardia | 0
    previous bilateral total knee joint replacement | 0
    chest pain | 0
    shortness of breath on exertion | 0
    electrocardiogram showed old left bundle branch block | 0
    serial high-sensitivity troponin levels | 0
    hs-TnT 55 ng/L | 0
    hs-TnT 71 ng/L | 0
    temperature 35.8°C | 0
    TTE showed normal biventricular size and function | 0
    angiography | 0
    99% stenosis in dominant RCA | 0
    stents placed in RCA | 0
    balloon rupture | 0
    discharged home | 72
    progressive shortness of breath | 840
    mild bilateral pedal oedema | 840
    normal heart and lung sounds | 840
    white cell count 14.3 × 10^9/L | 840
    C-reactive protein 110 mg/L | 840
    non-dynamic hs-TnT 85 ng/L | 840
    hs-TnT 82 ng/L | 840
    TTE showed normal biventricular function | 840
    normal valve function | 840
    no endocarditis | 840
    no pericardial effusion | 840
    blood cultures positive | 24
    MSSA | 24
    IV flucloxacillin | 24
    mild trauma to left knee | -120
    knee mildly swollen | 24
    knee tender | 24
    no erythema | 24
    aspirate performed | 24
    white cell count 100 800 × 10^6/L | 24
    no organisms | 24
    arthroscopic washout | 24
    serous fluid | 24
    Staphylococcus epidermidis | 24
    TOE showed no endocarditis | 24
    no pacemaker wire infection | 24
    no pericardial effusion | 24
    worsening shortness of breath | 24
    pleuritic chest pain | 24
    worsening kidney injury | 24
    oliguria | 24
    attempted dialysis | 24
    hypotension | 24
    angina | 24
    admitted to ICU | 24
    dialysis with inotropic support | 24
    focused cardiac ultrasound showed moderate pericardial effusion | 24
    no tamponade | 24
    TTE confirmed moderate circumferential pericardial effusion | 24
    no haemodynamic compromise | 24
    hypoechoic collection around RCA and stent | 24
    TOE confirmed tamponade | 24
    pericardiocentesis | 24
    purulent fluid drained | 24
    white cell count 2540 × 10^6/L | 24
    MSSA | 24
    severe cardiogenic shock | 24
    vasoplegic shock | 24
    hypoxia | 24
    intubated | 24
    escalating vasoactive support | 24
    CT coronary angiography showed RCA aneurysm | 24
    contrast extravasation | 24
    TTE showed severe biventricular failure | 24
    large pericardial effusion | 24
    pericardial drain blocked | 24
    conservative management | 24
    antibiotics escalated to vancomycin | 24
    clindamycin | 24
    cefazolin | 24
    extubated | 168
    percutaneous balloon pericardial window | 168
    discharged from ICU | 168
    discharged from hospital | 168
    lifelong suppression antibiotics with flucloxacillin | 168
    full time work 3 months post discharge | 2160
    no functional limitations | 2160
    repeat TTE showed moderate to severely reduced LV function | 8760
    moderately reduced RV function | 8760
    no significant pericardial effusion | 8760
    