59 years old | 0
female | 0
blood type O | 0
Rh positive | 0
admitted to the hospital | 0
segment-V space-occupying lesion in the liver | -365
transarterial embolization | -348
sorafenib | -304
dizziness | -273
skin ulcers | -273
computed tomography scan | -273
radiation therapy | -14
Piggyback LT | 0
hepatitis B | 0
entecavir | 0
HBV serology test | 0
acute renal failure | 0
hematoma around the liver | 0
intravenous administration of hepatitis B immunoglobulin | 24
immunosuppressive drugs | 24
steroids | 24
tacrolimus | 24
continuous hemodialysis | 24
intermittent infusion of fresh frozen plasma | 24
leukocyte-depleted red blood cells | 24
active bleeding in the abdominal cavity ceased | 48
renal function gradually recovered | 48
pathological analyses | 48
HCC | 48
massive tumor necrosis | 48
liver function began to improve | 240
AST | 240
ALT | 240
GGT | 240
ALP | 240
fevers | 240
procalcitonin levels | 240
rash | 312
obscure red spots | 312
no symptoms such as itching | 312
Nikolsky sign was negative | 312
tacrolimus administration changed to sirolimus | 408
mycophenolate mofetil | 408
sputum culture | 432
Acinetobacter baumannii | 432
methicillin-resistant Staphylococcus aureus | 432
rash advanced into erythematous macules and papules | 456
severe bone marrow suppression | 456
WBC count | 456
PLT count | 456
HGB level | 456
oral examination | 456
white ulcers on both sides of the buccal mucosa and lips | 456
severe bone marrow suppression | 456
bone marrow aspiration | 768
bone marrow pathology report | 768
FISH analysis of the peripheral blood | 792
donor lymphocytes | 792
skin biopsy | 816
epidermal dyskeratosis | 816
basic vacuolization | 816
lymphocytic infiltrates | 816
grade-1 acute lt-GVHD | 816
multidisciplinary team | 816
steroids | 816
tacrolimus | 816
G-CSF | 816
meropenem | 816
voriconazole | 816
rash was significantly reduced | 1104
general condition continued to deteriorate | 1104
serum ferritin levels | 1104
esophageal and oral ulcers | 1104
temperature rose to 39.4°C | 1128
hallucinations | 1128
septic shock | 1320
multiple organ dysfunction syndrome | 1320
death | 1320