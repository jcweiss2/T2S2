70 years old | 0
man | 0
presented to the emergency room | 0
chronic diarrhea | -240
confusion worsening | -240
gout | -1440
colchicine | -1440
allopurinol | -1440
prednisone taper | -1440
diarrhea began | -1440
denied recent surgeries | 0
denied abdominal pain | 0
denied hematochezia | 0
denied melena | 0
denied nausea | 0
denied vomiting | 0
denied fevers | 0
denied chills | 0
denied night sweats | 0
tremulous | 0
weak | 0
worsening fatigue | 0
falls | -168
required 2 L of oxygen | 0
sleep apnea | 0
continuous positive airway pressure | 0
heart failure | 0
furosemide | 0
non-alcoholic steatohepatitis | 0
liver transplant in 2013 | 0
hypertension | 0
coronary artery disease | 0
drug eluting stent placement | 0
60-pack-year smoking history | 0
quit smoking 29 years prior | 0
denied alcohol use | 0
denied drug use | 0
thyroid disease in sister | 0
pulse 117-135 | 0
temperature 36.6°C | 0
respirations 24 | 0
oxygen saturation 96% on 2 L NC | 0
blood pressure 96/72 mmHg | 0
morbidly obese | 0
tachycardia | 0
lethargic | 0
arousable | 0
oriented only to person | 0
intact cranial nerves | 0
normal motor examination | 0
normal sensory examination | 0
no enlargement of thyroid | 0
no nodule of thyroid | 0
no ophthalmopathy | 0
tenderness of thyroid undetermined | 0
white blood cells 4.76 K/cumm | 0
hemoglobin 10.0 g/dL | 0
platelets 106 K/cumm |:0
sodium 134.0 mmol/L | 0
potassium 5.20 mmol/L | 0
BUN 74.0 mg/dL | 0
creatinine 3.3 mg/dL | 0
magnesium 1.7 mg/dL | 0
phosphorus 7.2 mg/dL | 0
INR 1.54 | 0
blood cultures negative | 0
respiratory bacterial culture negative | 0
gastrointestinal PCR negative | 0
herpes simplex virus PCR negative | 0
cytomegalovirus PCR negative | 0
chest x-ray negative | 0
urinalysis negative | 0
VRE culture negative | 0
MRSA culture negative | 0
CT head negative | 0
urine drug screen negative | 0
tacrolimus levels within range | 0
hemoglobin A1c 4.7 | 0
glucose level 286 mg/dL | 0
lithium level <0.1 mmol/L | 0
procalcitonin level 0.09 ng/mL | 0
TSH 0.01 mIU/L | 0
Free T4 5.91 ng/dL | 0
Free T3 14.5 pg/mL | 0
ultrasound of head and neck negative | 0
diffusely mildly hypervascular thyroid | 0
diarrhea | 0
delirium | 0
thyroid storm | 0
denied exogenous thyroid hormone | 0
excluded infection | 0
excluded myocardial infarction | 0
excluded diabetic ketoacidosis | 0
head and neck ultrasound | 0
right thyroid lobe 5.2 × 2.8 × 2.2 cm³ | 0
left thyroid lobe 5.0 × 2.4 × 1.9 cm³ | 0
anti-thyroglobulin antibody 2555.0 IU/mL | 0
Burch-Wartofsky score 50 | 0
confirmed thyroid storm | 0
transferred to ICU | 0
propanol 40 mg every six hours | 0
methimazole 20 mg TID | 0
prednisone 60 mg daily | 0
non-ST-elevation myocardial infarction | 0
demand ischemia | 0
right lower lobe pneumonia | 0
piperacillin-tazobactam for 7 days | 0
thrombocytopenia | 0
liver disease | 0
sepsis | 0
returned to baseline | 504
Free T4 normalized after 9 days | 216
Free T4 rise on hospital day 21 | 504
Free T4 1.64 ng/dL | 504
Free T4 2.01 ng/dL | 504
Free T4 2.23 ng/dL | 504
methimazole washout 6 days | 504
thyroid uptake scan | 504
globally decreased uptake 1.2% | 504
no active nodules | 504
restarted prednisone 40 mg daily | 504
Free T3 2.1 pg/mL | 2160
T4 0.82 ng/dL | 2160
TSH 16.23 mIU/L | 2160
denied hypothyroidism symptoms | 2160
denied hyperthyroidism symptoms | 2160
levothyroxine 50 mcg daily | 2160
euthyroid | 8760
Free T3 2.5 pg/mL | 8760
T4 1.17 ng/dL | 8760
TSH 1.38 mIU/L | 8760
