72 years old | 0 | 0 
male | 0 | 0 
admitted to the hospital | 0 | 0 
high-grade fever | -96 | 0 
influenza B virus infection | -96 | 0 
wife diagnosed with influenza B virus infection | -168 | -168 
daughters diagnosed with influenza B virus infection | -168 | -168 
rapid test positive for influenza B antigens | -96 | -96 
oseltamivir administered | -96 | -96 
persistent fever | -96 | 0 
dyspnea at rest | -96 | 0 
temperature 38.7°C | 0 | 0 
blood pressure 117/80 mmHg | 0 | 0 
heart rate 76 beats/min | 0 | 0 
oxygen saturation level 88% | 0 | 0 
fine crackles in lung fields | 0 | 0 
white blood cell count 7400/mm3 | 0 | 0 
C-reactive protein 18.1 mg/dL | 0 | 0 
aspartate transaminase 91 IU/L | 0 | 0 
L-lactate dehydrogenase 362 IU/L | 0 | 0 
creatine kinase 793 IU/L | 0 | 0 
Krebs von den Lungen-6 1772 U/mL | 0 | 0 
hypoxemia | 0 | 0 
arterial blood gas analysis | 0 | 0 
ground-glass opacity in lung fields | 0 | 0 
chest computed tomography | 0 | 0 
diffuse ground-glass opacity in lung fields | 0 | 0 
high-flow nasal oxygen support | 0 | 129 
intravenous peramivir | 0 | 129 
antibiotics | 0 | 129 
piperacillin/tazobactam | 0 | 129 
levofloxacin | 0 | 129 
reticular shadow on chest CT worsened | 72 | 72 
PaO2/FiO2 ratio deteriorated | 72 | 72 
severe ARDS | 72 | 129 
mechanical ventilation proposed | 72 | 72 
high levels of positive end-expiratory pressure proposed | 72 | 72 
intubation refused | 72 | 72 
polymyxin B-immobilized fiber column hemoperfusion | 72 | 72 
intravenous methylprednisolone | 144 | 144 
noninvasive positive pressure ventilation support | 144 | 129 
immunosuppressant therapy | 144 | 129 
intravenous cyclophosphamide | 144 | 129 
respiratory status did not improve | 144 | 129 
reticular infiltrates on chest CT worsened | 144 | 129 
death | 129 | 129 
autopsy performed | 129 | 129 
diffuse alveolar damage | 129 | 129 
prominent hyaline membranes | 129 | 129 
no specific abnormality in other organs | 129 | 129