40 years old | 0
    female | 0
    liver transplantation | -4320
    cirrhosis | -4320
    nonalcoholic steatohepatitis | -4320
    hypertrophic cardiomyopathy | -4320
    myomectomy | -4320
    hypothyroidism | -4320
    Type II diabetes mellitus | -4320
    chronic kidney disease | -4320
    tacrolimus | -4320
    mycophenolic acid | -4320
    prednisone | -4320
    tacrolimus-related posterior reversible encephalopathy syndrome | -1512
    everolimus-based therapy | -1512
    liver biopsy | -1344
    severe acute cellular rejection | -1344
    high-dose steroids | -1344
    thymoglobulin | -1344
    cyclosporine | -1344
    admitted to ICU | 0
    adult respiratory distress syndrome | 0
    septic shock | 0
    Legionella pneumophila pneumonia | 0
    respiratory failure | 0
    failed extubation | 0
    ventilatory support | 0
    acute on chronic renal failure | 0
    CRRT | 0
    worsening graft dysfunction | 0
    propofol | 0
    opioids | 0
    cyclosporine | 0
    aggressive up-titration | 0
    subtherapeutic levels | 0
    CRRT filter clotting multiple times | 312
    heparin infusion | 312
    activated partial thromboplastin time goal | 312
    right radial artery thrombus | 312
    aPTT stable between 48 s and 64 s | 312
    propofol infusion | 312
    TG level of 3745 mg/dl | 312
    TG level of 156 mg/dl | -4320
    filter and circuits changed | 312
    propofol discontinued | 312
    clotting | 312
    line color change | 312
    filter color change | 312
    TG level of 3865 mg/dl | 312
    normal lipase level | 312
    rising serum potassium of 5.8 mmol/L | 312
    serum bicarbonate of 20 mmol/L | 312
    pH of 7.2 | 312
    intravenous insulin | 312
    heparin | 312
    emergent therapeutic plasma exchange | 312
    TPE initiated | 318
    5% albumin | 318
    citrate anticoagulant | 318
    CRRT resumed | 318
    acid–base balance normalized | 318
    electrolytes normalized | 318
    heparin infusion | 318
    elevated TG levels up to 708 mg/dl | 384
    increasing serum lipase levels peaking at 240 mg/dl | 384
    abdominal pain | 384
    pancreatitis | 384
    two additional TPE sessions | 384
    TG decreased from 708 to 186 mg/dl | 384
    TG decreased from 499 to 212 mg/dl | 504
    cyclosporine with escalating doses | 504
    persistent subtherapeutic serum levels | 504
    liver graft dysfunction | 504
    recurrent hypertriglyceridemia | 504
    persistent hypertriglyceridemia | 504
    oral fibrate | 504
    fish oil | 504
    preventive measures | 504
    combined liver–kidney transplant | 1344
    propofol for sedation intraoperatively | 1344
    cyclosporine postoperatively | 1344
    TGs level of 154 mg/dl | 1344
    lowest TGs level since baseline | 1344
    TGs level remained well-controlled | 1344

