65 years old | 0
female | 0
liver cirrhosis | -8760
chronic hepatitis B | -8760
hepatocellular carcinoma | 0
admitted to the hospital | 0
premedication with glycopyrrolate | 0
general anesthesia induced | 0
intubated and ventilated mechanically | 0
monitored by electrocardiography | 0
monitored by arterial blood pressure | 0
monitored by central venous pressure | 0
monitored by SpO2 | 0
hepatectomy started | 0
CUSA used | 0
sudden decrease in arterial blood pressure | 1
tachycardia | 1
ST elevation on EKG | 1
resuscitation with colloid and catecholamines | 1
intraoperative ultrasonography revealed massive air emboli | 1
diagnosed with VAE and PAE | 1
arterial blood gas analysis | 1
catecholamine administration | 1
systolic blood pressure maintained | 1.17
heart rate maintained | 1.17
central venous pressure maintained | 1.17
end-tidal carbon dioxide restored | 1.17
ABGA at 30 minutes after the occurrence | 1.5
norepinephrine infusion continued | 1.5
fluid resuscitation continued | 1.5
air emboli in left heart disappeared | 2.17
hepatectomy restarted | 2.17
hepatectomy completed | 5
intubated and ventilated mechanically in ICU | 5
responded only to intense pain | 5
systolic pressure maintained | 5
norepinephrine infusion | 5
postoperative laboratory findings | 5
postoperative EKG showed ST elevation | 5
EKG findings recovered normally at POD 1 | 24
trans-thoracic echocardiogram showed unremarkable findings | 24
vital signs stable | 24
norepinephrine infusion tapered out | 24
mental status unchanged at POD 5 | 120
brain CT and MRI revealed multiple acute cerebral infarctions | 120
weaned to spontaneous ventilation with CPAP mode | 264
extubated | 264
vital signs became unstable | 360
intravenous administration of catecholamines started | 360
panperitonitis confirmed | 744
expired due to cardiac arrest caused by septic shock | 744