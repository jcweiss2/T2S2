89 years old | 0
male | 0
admitted to the ICU | 0
COPD | -336
nocturnal oxygen therapy | -336
COPD exacerbation | -336
hospitalized | -336
fever | -168
hypoxemia | -168
bilateral lung infiltrates | -168
RT-PCR positive for SARS-CoV-2 | -168
hydroxychloroquine | -168
azithromycin | -168
intubated | 0
sedated | 0
mechanically ventilated | 0
tidal volume of 6.5 ml/kg | 0
rate of 20 breaths per minute | 0
PEEP of 8cmH2O | 0
physical examination unremarkable | 0
hemodynamically stable | 0
PaO2/FiO2 of 110 | 0
respiratory system compliance 35 ml/cmH2O | 0
airway resistance 18cmH2O/L/sec | 0
intrinsic PEEP of 2cmH2O | 0
CVP of 12 mmHg | 0
ScvO2 of 76 % | 0
ECG showed incomplete RBBB | 0
chest X-ray revealed signs of emphysema and bilateral infiltrates | 0
mild leukocytosis | 0
low lymphocyte count | 0
elevated C-reactive protein | 0
elevated ferritin | 0
elevated interleukin-6 | 0
elevated d-dimer levels | 0
acute circulatory collapse | 24
non-responding to fluid resuscitation | 24
non-responding to high dose of vasopressors | 24
CVP of 18 mmHg | 24
ScvO2 of 58 % | 24
ECG showed new onset infero-lateral ST elevation | 24
high sensitive cardiac troponin I | 24
bedside transthoracic echocardiography | 24
anterior pericardial effusion | 24
right ventricular diastolic collapse | 24
mitral valve inflow variation of 30 % | 24
left ventricular systolic function normal | 24
LVEF of 60 % | 24
echo-guided pericardiocentesis | 24
aspiration of 200 mL of serous fluid | 24
hemodynamic improvement | 24
pericardial drainage maintained in situ | 24
yielded a total of 240 mL of fluid | 48
pericardial fluid tested negative for Gram stain | 24
pericardial fluid tested negative for acid-fast bacilli smear | 24
no growth on bacterial and fungal cultures | 24
molecular testing for Mycobacterium tuberculosis negative | 24
RT-PCR for SARS-CoV-2 negative | 24
fluid cytology yielded no malignant cells | 24
thyroid function tests normal | 24
serologic tests for Coxsackievirus negative | 24
serologic tests for Echovirus negative | 24
serologic tests for hepatitis viruses negative | 24
serologic tests for cytomegalovirus negative | 24
serologic tests for human immunodeficiency virus negative | 24
serologic tests for autoantibodies negative | 24
treatment with colchicine started | 24
rapidly weaned off vasopressors | 48
repeat echocardiograms showed no recurrence of pericardial effusion | 48
septic shock | 144
multi-organ failure | 144
multi-drug resistant Acinetobacter baumanii | 144
died | 144