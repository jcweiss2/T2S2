3-year-old | 0
    female | 0
    Noonan syndrome | 0
    heterozygous RIT1 mutation | 0
    heart murmur | -8760
    hypertrophic cardiomyopathy | -8760
    mid cavity left ventricular outflow tract obstruction | -8760
    severe right ventricular outflow tract obstruction | -8760
    dysplastic stenotic pulmonary valve | -8760
    surgical relief of LVOT obstruction with myectomy | -6864
    surgical relief of RVOT obstruction with muscular resection | -6864
    transannular patch | -6864
    epicardial pacemaker | -6864
    post-operative complete heart block | -6864
    recovered well following the procedure | -6864
    no progression of HCM | -6864
    admitted to intensive care unit | -2184
    respiratory failure | -2184
    parainfluenza 3 infection | -2184
    bilateral pleural effusions | -2184
    pleural effusions requiring drainage | -2184
    chylothorax | -2184
    fluid triglycerides 1.9 mmol/L | -2184
    fluid protein 30 g/L | -2184
    gram stain negative | -2184
    mononuclear white blood cells | -2184
    low fat diet | -2184
    high medium chain triglycerides diet | -2184
    octreotide infusion | -2184
    significant chyle loss | -2184
    low immunoglobulin levels | -2184
    acute deterioration | -2184
    spontaneous bowel perforation | -2184
    terminal ileum resection | -2184
    stoma formation | -2184
    bacterial sepsis | -2184
    candida sepsis | -2184
    antibiotics | -2184
    antifungals | -2184
    immunoglobulin replacements | -2184
    parenteral nutrition | -2184
    refractory pleural effusions | -2184
    high stoma losses | -2184
    MCT diet | -2184
    discharged home | -2184
    reaccumulation of pleural effusions | 0
    multiple chest drains | 0
    respiratory compromise | 0
    pulmonary lymphangiectasia | 0
    residual cardiac anomalies | 0
    surgical damage to thoracic duct | 0
    no residual left ventricular outflow tract obstruction | 0
    no residual right ventricular outflow tract obstruction | 0
    small atrial septal defect | 0
    bidirectional shunt | 0
    restrictive right ventricular physiology | 0
    elevated bi-atrial pressures | 0
    mean pulmonary artery pressure of 20 mmHg | 0
    mildly increased pulmonary vascular resistance | 0
    calculated cardiac index of 3.8 L/min/m2 | 0
    innominate vein wedge angiogram | 0
    thoracic duct entry point not demonstrated | 0
    IV unobstructed | 0
    lymphatic dysplasia | 0
    elevated right-sided filling pressures | 0
    parenteral nutrition | 0
    intense diuresis | 0
    no improvement | 0
    trametinib treatment | 0
    severe eczema | 0
    stoma output increased | 0
    parenteral nutrition | 0
    fat-free oral feeds | 0
    reduction in left ventricular mass | 0
    3-month course of trametinib | 0
    enteral feeds | 0
    MCT diet | 0
    normal fat content diet | 0
    discharged home | 0
    free of chylothorax recurrence | 0
    chest X-ray | 0
    ultrasound | 0
    last pleural drainage | 0
    chylothorax resolution | 2160
    trametinib completion | 2160
    stoma reversal | 2160
    
