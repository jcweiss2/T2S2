61 years old | 0
female | 0
severe community-acquired pneumonia | 0
acute renal failure | 0
type 2 diabetes mellitus | 0
chronic obstructive airway disease | 0
acute tubular necrosis | 0
sepsis | 0
hypotension | 0
urine without red cells or casts | 0
initial stable renal function | 0
rapid worsening renal function | 24
significant fluid overload | 24
4 sessions of haemodialysis | 24
improved renal function | 24
became dialysis independent | 24
discharged home after 45 days | 1080
acute pulmonary oedema | 1080
skin rash | 1080
readmission to ICU within 48h of discharge | 1128
pulmonary hypertension | 1128
splenomegaly | 1128
hepatomegaly | 1128
bilateral pleural effusion | 1128
skin lesions typical of vasculitis | 1128
dysmorphic red cells in urine | 1128
proteinuria | 1128
hypoalbuminaemia | 1128
low complement levels | 1128
positive serology for mixed cryoglobulinaemia | 1128
normal renal ultrasound | 1128
weakly positive rheumatoid factor | 1128
negative HCV RNA | 1128
negative autoimmune screens | 1128
renal biopsy findings | 1128
5 sessions of plasma exchange | 1128
2 sessions of haemodialysis | 1128
prednisolone | 1128
cyclophosphamide | 1128
decrease in cryoglobulin levels within 3 weeks | 168
symptomatic improvement | 168
discontinued cyclophosphamide due to thrombocytopenia | 168
discharged on prednisolone 50 mg | 168
normal renal function on discharge | 168
symptomatic again after 2 weeks | 384
reappearance of rash | 384
positive/high serum cryoglobulins | 384
low complements | 384
worsening proteinuria | 384
significant weight gain | 384
high urea level | 384
5 sessions of plasmapheresis | 384
recommenced cyclophosphamide 50 mg/100 alternate days | 384
discharged again with normal renal function | 384
negative serum cryoglobulin | 384
represented with fluid overload and pneumonia after 12 days | 624
cyclophosphamide ceased due to thrombocytopenia | 624
sepsis | 624
herpes zoster | 624
intermittent haemodialysis | 624
plasmapheresis on alternate days for 1 month | 624
new-onset paraproteinaemia | 624
monoclonal IgM kappa | 624
negative Bence Jones protein | 624
normal skeletal survey | 624
no light chains in serum | 624
bone marrow biopsy showing low-grade lymphoma | 624
CD20 expression on B cells | 624
no clinical improvement | 624
regular dialysis/ultrafiltration | 624
given 600 mg rituximab/week for 3 weeks | 624
responded within 1 week | 744
dramatic improvement in symptoms | 744
