38 years old|0
female|0
presented to the otolaryngology outpatient clinic|0
bleeding from an ulcerating left fungating parotid tumour|0
first noted a pea-sized mass|-43200
fine-needle aspiration cytology of the mass|-43200
ACC|-43200
refused surgery|-43200
lost to follow-up|-43200
tumour slowly increased in size|-43200
rapid growth within the last year|-8760
malnourished|0
14 by 12 cm fungating parotid mass|0
areas of necrosis|0
haemorrhage|0
motor function of the facial nerve could not be assessed properly|0
hemoglobin 9.3 g/L|0
albumin level <10 g/L|0
other blood tests including electrolytes, liver function tests, and coagulation profile were normal|0
admitted for nutritional support|0
hemostasis|0
further management of her parotid malignancy|0
developed acute confusion|48
became agitated|48
computed tomography of the brain showed thrombosis of the contralateral transverse sinus extending into the proximal part of the internal jugular vein|48
Doppler ultrasound scan of the lower limbs revealed thrombosis of the distal part of the right common femoral vein|48
started on warfarin|48
inferior vena caval filter inserted|48
INR value went up to 8.0|288
bled from the tumour site|288
warfarin stopped|288
given Vitamin K|288
fresh-frozen plasma|288
INR came down to 2.0|312
warfarin switched to low-molecular-weight heparin (LMWH)|312
platelet count dropped from 500 to 15 × 109/L|672
serum positive for platelet factor-4 antibodies|672
diagnosis of Type II heparin-induced thrombocytopenia (HIT)|672
heparin switched to lepirudin|672
platelets returned to the normal level after 5 days of stopping heparin|768
condition deteriorated rapidly due to septicemia|792
transferred to the intensive care unit|792
started on broad-spectrum antibiotics|792
nutritional status got worse|792
not having adequate per oral intake|792
refused nasogastric feeding|792
multidisciplinary team recommended the surgery|792
underwent radical left-sided parotidectomy|792
type-1 modified radical neck dissection|792
carcinoma staged as T4|792
neck dissection necessary for facilitation of the latissimus dorsi pedicled muscle flap reconstruction|792
facial nerve sacrificed|792
tumour engulfed all branches of the nerve|792
accessory nerve preserved|792
internal jugular vein preserved|792
part of the zygomatic arch removed|792
tumour found herniating into the oral cavity through the parotid duct opening (Stensen's duct)|792
oral mucosa around the tumour excised and closed primarily|792
latissimus dorsi pedicled muscle flap raised|792
split skin graft used to cover the muscle flap|792
histology confirmed moderately differentiated ACC of the parotid with clear margins|792
noted vascular invasion|792
none of the 61 lymph nodes harvested were positive for malignancy|792
disease staged as pT4pN0M0|792
hematoma formation at the latissimus dorsi flap donor site|792
drained|792
episode of septicemia due to an infected central venous catheter|792
treated with antibiotics|792
part of the split skin graft had to be re-grafted|792
local wound infection|792
discharged from the hospital after 65 days|1560
normalized serum albumin level|1560
underwent adjuvant postoperative radiotherapy|1560
died 19 months after the surgery due to lung metastasis|14160
