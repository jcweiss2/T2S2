59 years old | 0
female | 0
blood type O | 0
Rh positive | 0
segment-V space8occupying lesion in liver | -14400
suspected liver cancer | -14400
transarterial embolization | -14400
sorafenib | -1464
stopped sorafenib | -480
dizziness | -480
skin ulcers | -480
CT scan | -1440
liver segment V lesions enlarged | -1440
radiation therapy | -1440
PTV5400cGy/18f | -1440
dose rate 0.6-1 Gy/min | -1440
Piggyback liver transplantation | 0
hepatitis B | 0
entecavir | 0
HBsAg 113.23 IU/mL | 0
anti-HBs 0 mIU/mL | 0
HBeAg 0.08 PEI µ/mL | 0
anti-HBe >4.4 PEI µ/mL | 0
anti-HBc 8.26 PEI µ/mL | 0
serological tests negative for HIV, hepatitis A, hepatitis C | 0
donor age 21 | 0
male | 0
HLA class-I A11, A30 | 0
HLA-B B13 | 0
HLA-DR 11,15 | 0
HLA-DQ 6,7 | 0
recipient HLA-A 2,11 | 0
HLA-B 13,46 | 0
HLA-DR 14,15 | 0
HLA-DQ 5,6 | 0
acute renal failure | 24
hematoma around liver | 24
hepatitis B immunoglobulin | 24
steroids | 24
tacrolimus | 24
tacrolimus blood level ~10 ng/mL | 24
continuous hemodialysis | 24
fresh frozen plasma | 24
leukocyte8depleted red blood cells | 24
active bleeding ceased | 24
renal function recovery | 24
HCC diagnosis | 24
tumor necrosis ~90% | 24
surviving tumor ~10% | 24
liver function improvement | 240
AST normal | 240
ALT normal | 240
GGT normal | 240
ALP normal | 240
fever 37-39°C | 312
fever peaks at 23:00 daily | 312
PCT 10.3 ng/mL | 312
PCT dropped to 3 ng/mL | 360
blood cultures negative | 360
cytomegalovirus negative | 360
EBV negative | 360
fever persisted | 360
red spots on chest | 360
no itching | 360
Nikolsky sign negative | 360
tacrolimus changed to sirolimus | 408
mycophenolate mofetil added | 408
Acinetobacter baumannii | 432
MRSA | 432
rash advanced to erythematous macules/papules | 456
spread to limbs, palms, neck, face | 456
oral white ulcers | 456
WBC 0.86×109/L | 456
PLT 35×109/L | 456
HGB 70 g/L | 456
transferred to ICU | 456
rash hypothesized as drug reaction | 456
gamma globulin 2500 mg | 456
skin biopsy | 456
FISH peripheral blood | 456
abdominal incision split | 696
sutured again | 696
bone marrow aspiration | 768
bone marrow pathology no special lesions | 768
megakaryocyte production reduced | 768
PLT decreased | 768
FISH detected 3% donor lymphocytes | 792
skin biopsy epidermal dyskeratosis | 792
basic vacuolization | 792
lymphocytic infiltrates | 792
grade-1 acute lt-GVHD | 792
CD4:CD8 ratio reversed 1:13.3 | 792
IgM reduced to 0.3 g/L | 792
PLT 3.2×109/L | 792
steroids continued | 792
tacrolimus continued | 792
G-CSF | 792
meropenem | 792
voriconazole | 792
rash reduced | 792
serum ferritin 11,276.55 ng/mL | 792
esophageal ulcers worsened | 792
oral ulcers worsened | 792
difficulty eating | 792
fever 39.4°C | 1128
hallucinations | 1128
MRSA infection | 1128
Acinetobacter baumannii infection | 1128
Enterococcus faecalis infection | 1128
IgM 0 g/L | 1128
septic shock | 1320
MODS | 1320
death | 1320
