39 years old | 0 | 0 
female | 0 | 0 
palpable mass on her right breast | -168 | 0 
Hodgkin lymphoma | -6336 | -6336 
chemotherapy | -6336 | -6336 
mantle field radiation | -6336 | -6336 
inflammatory colitis | -6336 | -168 
mesalazine | -168 | -168 
family history of myxoid liposarcoma | 0 | 0 
radiological examination of the breast | -168 | 0 
invasive ductal carcinoma | -168 | 0 
triple-negative phenotype | -168 | 0 
MIB1 85% | -168 | 0 
staging CT scan of the thorax and abdomen | -168 | 0 
no distant metastasis | -168 | 0 
neoadjuvant chemotherapy | -168 | 0 
paclitaxel | -168 | 0 
carboplatin | -168 | 0 
first cycle of chemotherapy | -24 | 0 
port-à-cath insertion | 0 | 0 
subcutaneous cellulitis | 12 | 12 
colliquative necrosis | 12 | 12 
elevated white blood cell count | 12 | 12 
neutrophilia | 12 | 12 
elevated C-reactive protein | 12 | 12 
broad-spectrum i.v. antibiotic therapy | 12 | 12 
piperacillin/tazobactam | 12 | 12 
daptomycin | 12 | 12 
PORT rimotion and necrosectomy | 12 | 12 
defervescence | 12 | 12 
improvement in subcutaneous cellulitis | 12 | 12 
improvement in blood works | 12 | 12 
febrile seizure | 14 | 14 
WBC rise | 14 | 14 
worsening of skin lesion | 14 | 14 
second necrosectomy | 14 | 14 
peripheral blood cultures | 14 | 14 
skin plug | 14 | 14 
i.v. catheter tip showed positivity for Klebsiella pneumoniae | 14 | 14 
antibiotic therapy modification | 14 | 14 
meropenem | 14 | 14 
levofloxacin | 14 | 14 
chest/abdomen CT scan | 14 | 14 
mediastinitis | 14 | 14 
bilateral pleural effusion | 14 | 14 
left pulmonary atelectasis | 14 | 14 
thoracoscopy with pleural and mediastinal drainage | 14 | 14 
sepsis | 14 | 24 
broad-spectrum antibiotic and antifungal therapy | 14 | 24 
hemodynamic support | 14 | 24 
non-invasive ventilation | 14 | 24 
specimens of skin and subcutaneous and muscular tissue | 14 | 14 
intensive inflammatory infiltrate | 14 | 14 
neutrophils | 14 | 14 
differential diagnosis of PG | 14 | 14 
systemic methylprednisolone | 24 | 168 
topical cyclosporine | 24 | 168 
seriate chest X-ray | 24 | 168 
CT scan | 24 | 168 
progressive resolution of mediastinitis | 24 | 168 
progressive resolution of pleural effusion | 24 | 168 
wound improvement with scar | 24 | 168 
progressive normalization of blood count | 24 | 168 
progressive normalization of flogosis index | 24 | 168 
breast ultrasound | 168 | 168 
no change in the dimension of the lump | 168 | 168 
multidisciplinary meeting | 168 | 168 
right mastectomy | 168 | 168 
axillary dissection | 168 | 168 
breast surgical wound healing | 168 | 168 
pathology assessment | 168 | 168 
fibroelastosis | 168 | 168 
chronic inflammation | 168 | 168 
isolated neoplastic cells | 168 | 168 
negative axillary nodes | 168 | 168 
restaging brain/chest/abdomen CT | 168 | 168 
no distant metastasis | 168 | 168 
BRCA and p53 mutation tests | 168 | 168 
negative BRCA and p53 mutation tests | 168 | 168 
autologous skin graft | 336 | 336 
no further complications | 336 | 336 
PICC implant | 336 | 336 
resumed chemotherapy | 336 | 336 
carboplatin | 336 | 336 
paclitaxel | 336 | 336 
dose reduction | 336 | 336 
good tolerance | 336 | 504 
follow-up | 504 | 504 
postsurgical PG | 12 | 168 
pathergy | 12 | 168 
immune deregulation | 0 | 504 
tumor and PG diagnoses | 0 | 504 
tumor-related surgery | 168 | 168 
PG improvement | 168 | 504 
anti-tumor therapy | 168 | 504 
aberrant immune surveillance mechanisms | 0 | 504 
paraneoplastic conditions | 0 | 504 
lymphocytic infiltration | 168 | 168 
moderate infiltrate | 168 | 168 
cross-reactive antigens | 0 | 504 
anti-tumor immune response | 0 | 504 
tumor samples | 0 | 504 
pre-treatment sample | -168 | -168 
surgical sample | 168 | 168 
TILs | 168 | 168 
pathological assessment | 168 | 168 
written informed consent | 0 | 0 
conflict of interest statement | 0 | 0 
funding sources | 0 | 0 
author contributions | 0 | 0