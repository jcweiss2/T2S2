62 years old | 0
male | 0
COPD Gold II | 0
Hashimoto's disease | 0
presented to emergency department with shortness of breath | 0
presented to emergency department with coughing | 0
presented to emergency department with fever | 0
presented to emergency department with myalgia | 0
experienced symptoms for ten days | -240
tested positive for SARS-CoV-2 | -168
admitted to intensive care | 0
started treatment with remdesivir | 0
started treatment with dexamethasone | 0
started treatment with high-dose prophylactic LMWH | 0
LMWH dose adjusted to therapeutic range | 0
CTPA showed no pulmonary embolisms | 0
paroxysmal hypoxia | 192
chest pain | 192
macrocirculation stable | 192
SOFA score of 2 | 192
electrocardiogram showed no abnormalities | 192
cardiac markers showed no abnormalities | 192
echocardiography showed no abnormalities | 192
D-dimer increased from 1.73 mg/L to 8.44 mg/L | 192
new CTPA showed large vessel thrombosis of pulmonary arteries | 192
new CTPA showed large vessel thrombosis of thoracic aorta | 192
partial abdominal imaging showed renal infarction | 192
partial abdominal imaging showed spleen infarction | 192
sublingual microcirculation showed hyperdynamic circulation | 192
sublingual microcirculation showed increased total vessel density | 192
sublingual microcirculation showed no thrombosis | 192
isolated respiratory failure | 192
started continuous high molecular weight heparin infusion | 192
APTT adjusted every 6 hours | 192
respiratory status deteriorated | 216
mechanical ventilation needed | 216
Staphylococcus Aureus pneumosepsis | 408
progressive multi-organ failure | 408
patient died | 408
