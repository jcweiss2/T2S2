36 years old | 0
    female | 0
    admitted to the hospital | 0
    diabetes mellitus type II | 0
    obstructive sleep apnea | 0
    hypertension | 0
    hypothyroidism | 0
    morbid obesity | 0
    general body ache | -72
    malaise | -72
    breathing difficulty | -48
    tachycardia (120 bpm) | 0
    tachypnea (36/min) | 0
    leukocytosis (white blood cell count > 52,000) | 0
    urinary tract infection (pus cell count - 12-15 cells) | 0
    antibiotics (meropenem, 500 mg thrice a day) | 0
    vasopressors | 0
    adequate fluid resuscitation | 0
    mechanical ventilation | 0
    deterioration with decreasing urine output | 0
    intubated | 4
    became anuric | 6
    sequential organ failure assessment (SOFA) score was 15 | 24
    MODS score was 10 | 24
    acute physiology and chronic health evaluation (APACHE II) score was 30 | 24
    septic shock (urosepsis) | 16
    low perfusion state | 16
    MODS (acute respiratory distress syndrome, acute kidney injury, arterial hypotension) | 16
    hemoadsorption column (CytoSorb®) added | 16
    continuous renal replacement therapy for 24 h | 16
    flow rate maintained at 250 ml/min | 16
    anticoagulated with heparin | 16
    activated partial thromboplastin time of 30-40 s | 16
    improved hemodynamically | 28
    inotropic support | 28
    intravenous hydrocortisone | 28
    other supportive measures along with CytoSorb | 28
    Noradrenalin stopped | 28
    vasopressors gradually weaned out | 28
    corticosteroids (intravenous hydrocortisone), 100 mg thrice daily | 28
    stabilized after 3 days | 72
    CytoSorb applied daily | 72
    urine output increased | 72
    improvement in ventilator parameters | 72
    SOFA score was 4 | 72
    MODS score was 5 | 72
    APACHE II score was 7 | 72
    laboratory parameters within normal range | 72
    
    
    36 years old | 0
    female | 0
    admitted to the hospital | 0
    diabetes mellitus type II | 0
    obstructive sleep apnea | 0
    hypertension | 0
    hypothyroidism | 0
    morbid obesity | 0
    general body ache | -72
    malaise | -72
    breathing difficulty | -48
    tachycardia (120 bpm) | 0
    tachypnea (36/min) | 0
    leukocytosis (white blood cell count > 52,000) | 0
    urinary tract infection (pus cell count - 12-15 cells) | 0
    antibiotics (meropenem, 500 mg thrice a day) | 0
    vasopressors | 0
    adequate fluid resuscitation | 0
    mechanical ventilation |? 0
    deterioration with decreasing urine output | 0
    intubated | 4
    became anuric | 6
    sequential organ failure assessment (SOFA) score was 15 | 24
    MODS score was 10 | 24
    acute physiology and chronic health evaluation (APACHE II) score was 30 | 24
    septic shock (urosepsis) | 16
    low perfusion state | 16
    MODS (acute respiratory distress syndrome, acute kidney injury, arterial hypotension) | 16
    hemoadsorption column (CytoSorb®) added | 16
    continuous renal replacement therapy for 24 h | 16
    flow rate maintained at 250 ml/min | 16
    anticoagulated with heparin | 16
    activated partial thromboplastin time of 30-40 s | 16
    improved hemodynamically | 28
    inotropic support | 28
    intravenous hydrocortisone | 28
    other supportive measures along with CytoSorb | 28
    Noradrenalin stopped | 28
    vasopressors gradually weaned out | 28
    corticosteroids (intravenous hydrocortisone), 100 mg thrice daily | 28
    stabilized after 3 days | 72
    CytoSorb applied daily | 72
    urine output increased | 72
    improvement in ventilator parameters | 72
    SOFA score was 4 | 72
    MODS score was 5 | 72
    APACHE II score was 7 | 72
    laboratory parameters within normal range | 72
    