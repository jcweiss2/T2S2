400 g | 0
male | 0
delivered by primary cesarean delivery | 0
small for gestational age | 0
signs of placental insufficiency | 0
clear amniotic fluid | 0
delayed newborn adaptation | 0
respiratory support by CPAP mask | 0
transferred to neonatal intensive care unit | 0
administration of surfactant | 0
caffeine citrate | 0
empirical antibacterial therapy with piperacillin | 0
spironolactone | 0
hydrochlorothiazide | 0
intracranial hemorrhages grade 1 (right side) | 0
intracranial hemorrhages grade 2 (left side) | 0
negative initial perianal smear | 0
colonization with multidrug-resistant Acinetobacter pittii on day 14 | 336
recovered appropriately | 336
age of 3 months | -2160
body weight 2620 g | 0
planned for open both-sided inguinal hernia repair | 0
monitored blood pressure | 0
monitored oxygen saturation | 0
monitored heart rate | 0
sedated with propofol | 0
positioned in left lateral position | 0
maintained spontaneous breathing | 0
caudal anesthesia performed | 0
skin disinfection with Braunoderm | 0
surgical face masks worn | 0
sterile gloves worn | 0
identified caudal space with ultrasound | 0
entered hiatus sacralis | 0
instilled ropivacaine | 0
negative aspiration for blood and CSF | 0
confirmed epidural spread | 0
confirmed sufficient analgesia | 0
started surgery | 10
finished surgery | 61
no further analgesics required | 61
adequate neurology | 61
no signs of spinal block | 61
developed fever up to 39°C | 12
elevated CRP 3 mg/dL | 12
elevated IL-6 1477 pg/dL | 12
increased CRP to 27.6 mg/dL | 72
increased IL-6 to 26105 pg/dL | 24
initiated empiric broad antibacterial therapy | 12
firm abdomen | 12
painful abdomen | 12
no signs of intestinal perforation | 12
performed explorative laparotomy | 36
general anesthesia for laparotomy | 36
no pathological findings | 36
brain sonography signs compatible with inflammatory process | 48
no spinal cord pathologies | 48
lumbar puncture with increased cell counts | 48
increased protein in CSF | 48
increased lactate in CSF | 48
Gram stain assay identified Gram-instable rods | 48
no bacterial growth in culture | 48
switched to meropenem and vancomycin | 48
repeated lumbar puncture | 72
high lactate 85.6 mg/dL | 72
decreased cell counts 450/µL | 72
decreased protein 674 mg/dL | 72
no bacterial growth in blood cultures | 72
presence of Clostridium perfringens in CSF | 72
administered dexamethasone | 72
deteriorated clinical condition | 120
cystic remodeling of brain tissue | 72
secondary brain edema grade 3 | 120
generalized epileptic seizures | 120
anticonvulsive therapy with diazepam | 120
anticonvulsive therapy with phenobarbital | 120
developed apnea | 168
severe disturbance of temperature homeostasis | 168
died | 240
fulminant bacterial meningoencephalitis | 240
multiorgan failure | 240
