severe headache | -24
generalized tonic–clonic seizures | -24
loss of consciousness | -24
measurement of arterial blood pressure showed a value of 195/110 mmHg | -24
heart rate of 120 beats/min | -24
provisional diagnosis of eclampsia | -24
treated with antihypertensive therapy | -24
given an intravenous infusion of magnesium sulphate | -24
given ebrantil | -24
given 20% manitol | -24
given diazepam | -24
bilateral vision loss | -12
complete blood count was normal | -12
liver function tests were normal | -12
clotting parameters were normal | -12
electrocardiogram was normal | -12
urine analysis revealed proteinuria 2+ | -12
seizures were not repeated | 0
headache was alleviated | 0
ophthalmological examination revealed significant bilateral loss of vision | 0
diagnosis to cortical blindness | 0
mild right-sided facial nerve paresis | 0
no other neurological disorders | 0
multislice computed tomography scan showed hypodensity of the posterior white matter | 0
magnetic resonance imaging showed hyperintense signals in the white matter | 0
general condition stabilized | 12
moved to an obstetrics clinic | 12
blood pressure was stabilized using oral antihypertensive medication | 12
human albumin was administered by IV | 12
follow-up ophthalmological examinations showed significant bilateral improvement of the visual function | 120
best-corrected visual acuity 1.0 | 120
visual field image showed bilaterally expressed peripheral relative scotoma | 120
depressed sensitivity of the paracentral left visual field | 120
neurologist confirmed the right-sided partial facial nerve paresis | 120
no other neurological disturbances | 120
follow-up magnetic resonance imaging showed a significant regression of the edema | 192
discrete residual changes over the posterior horns of the side ventricles | 192
discharged from the clinic | 216
recommendation to take oral antihypertensive therapy | 216
recommendation to continue with physical therapy for the paresis of the facial nerve | 216