72 years old | 0
male | 0
hypertension | -168
stage 3 chronic kidney disease | -168
several weeks of worsening abdominal discomfort | -504
several weeks of constipation | -504
several weeks of worsening oral intake | -504
abdominal pain | 0
somnolent | 0
afebrile | 0
tachypneic | 0
tachycardic | 0
white blood cell count 27.7 | 0
potassium 7.0 mmol/L | 0
metabolic acidosis CO2 11mmol/L | 0
acute kidney injury | 0
BUN 174 mg/dL | 0
creatinine 15.4 mg/dL | 0
microscopic urinalysis positive for >150 RBC | 0
microscopic urinalysis positive for >150 WBC | 0
