45 years old | 0
male | 0
admitted to the hospital | 0
general malaise | -336
fever | -336
purpura | -336
pancytopenia | 0
leukopenia | 0
anemia | 0
thrombocytopenia | 0
diffusely increased bone marrow concentration | 0
bone marrow aspiration | 0
bone marrow biopsy | 0
acute panmyelosis with myelofibrosis | 0
acute myeloid leukemia | 0
idarubicin hydrochloride | 8
cytosine arabinoside | 8
induction therapy | 8
febrile neutropenia | 2
cefozopran | 2
left cheek cellulitis | 20
meropenem | 29
vancomycin | 29
levofloxacin | 38
hematological complete remission | 38
consolidation therapy | 38
cytosine arabinoside | 38
febrile neutropenia | 49
cefozopran | 49
hyperthermia | 54
blood culture | 54
central venous catheter removal | 54
pneumonia | 56
meropenem | 56
amikacin | 56
S. maltophilia | 57
trimethoprim-sulfamethoxazole | 57
levofloxacin | 57
ceftazidime | 57
minocycline | 57
hematic tracheal aspirates | 60
intubation | 57
intravenous granulocyte-colony stimulating factor | 63
SMX-TMP | 63
neutropenia | 63
airway pressure-release ventilation | 66
intermittent prone positioning | 66
respiratory failure | 66
ARDS | 66
bronchoalveolar lavage | 66
catecholamines | 66
VV ECMO | 68
tracheotomy | 71
awakened | 71
lungs opened up | 71
spontaneous breathing | 71
active mobilization of bronchial secretions | 71
weaned off VV ECMO | 79
mechanical ventilation support | 79
bilateral pulmonary infiltration improved | 79
biphasic positive airway pressure | 88
oxygen supplementation discontinued | 131
discharged from the hospital | 145
consolidation chemotherapy | 145
allogenic hematopoietic stem cell transplantation | 145
complete remission | 145