22 years old | 0
female | 0
admitted to the hospital | 0
LRGB | -21168
weight loss | -21168
correction of metabolic disturbances | -21168
internal hernia | 0
acute abdomen | 0
pregnant | 0
sudden onset of upper abdominal pain | 0
gall bladder stones | 0
MRI scan | 0
severe pain | 0
open cholecystectomy | 0
trans-cystic balloon dilation of the papilla of Vater | 0
cholangiogram demonstrated poor drainage | 0
small gallstones in the common hepatic bile duct | 0
re-operated due to cholascos | 120
renewed cystic duct ligation | 120
drainage | 120
endoscopy due to hematamesis | 144
blood in the jejunum | 144
no specific bleeding site | 144
clinical condition worsened | 144
transferred to the ICU | 144
severe septicaemia | 144
acute respiratory distress syndrome | 144
laparotomy | 312
internal hernia through Petersen's space | 312
necrosis of 1 m jejunum | 312
vital premature girl delivered by caesarean | 312
necrotic intestine removed | 312
second look operation | 336
third look operation | 336
further small bowel resections | 336
saliva fistula | 336
jejunostomy | 336
blind closed ileum | 336
infectious complications | 336
pneumothorax | 336
thrombosis of the superior mesenteric vein | 336
thrombosis of the iliac veins | 336
exposed bowel parquet covered with split skin | 336
transferred to intestinal failure unit | 336
good appetite | 336
no absorption of food | 336
short fistula below pouch-enteric anastomosis | 336
Hickmann catheter inserted | 336
parenteral nutrition with SMOF Kabiven | 336
vitamins and trace elements added | 336
isotonic saline for fluid balance | 336
yeast infection with candida albicans | 336
Hickmann catheter removed | 336
PICCline inserted | 336
discharged with home parenteral nutrition | 2880
intestinal continuity reconstructed | 5832
defect in anterior abdominal wall closed | 5832
PICCline occluded | 6624
PICCline removed | 6624
patient tried without parenteral nutrition | 6624
weight increased 2 kg | 6624
1–2 bowel movements a day | 6624
blood values for haemoglobin increased | 6624
blood values for albumin increased | 6624
short bowel syndrome | 336
parenteral nutrition dependency | 336
re-established intestinal continuity | 5832
amount of parenteral nutrition reduced | 5832
weaned off parenteral nutrition | 6624
survived | 6624
maternal death cases reported | 0
severe complications (type 2 intestinal failure) | 336
rehabilitation period | 2880
type 3 intestinal failure | 2880
successful reconstruction | 6624
no previous reports of survival with massive bowel necrosis | 0
importance of extensive surgery | 0
importance of second and third look operations | 0
internal herniation during third trimester | 0
internal herniation postpartum | 0
growing uterus increases intra-abdominal pressure | 0
uterus decreases in size postpartum | 0
internal herniation in up to 16% of patients | 0
bariatric surgeries in women of reproductive age | 0
LRGB increases fertility | 0
complications during pregnancy expected | 0
changed anatomy disposes for herniation | 0
abdominal pain difficult to diagnose | 0
MRI or CT scans not postponed | 0
laparoscopy on wide indication | 0
laparotomy if anatomy unclear | 0
successful reconstruction literature examples | 0
younger age improves prognosis | 0
awareness of internal hernia | 0
surgery on wide indication | 0
bowel necrosis resection | 0
start parenteral nutrition | 0
evaluation in specialized centres | 0
