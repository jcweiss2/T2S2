39 years old | 0
male | 0
admitted to the hospital | -2160
confusion | -2160
intra-abdominal trauma | -2160
traffic accident | -2160
ventilator-associated pneumonia | -2160
A. baumannii | -2160
tigecycline | -120
fever | -168
pustular eruptions | -96
erythematous areas | -96
facial and neck region | -96
upper and lower extremity | -96
mild erupted lesions | -48
tigecycline stopped | -48
tigecycline restarted | 0
generalized erupted lesions | 96
erythema | 12
pustules | 24
dermatologic examination | 24
numerous pustules | 24
face | 24
neck | 24
legs | 24
erythematous areas | 24
follicular localization | 24
oral examination | 24
no pathologies | 24
psoriasis | 0
family history | 0
no known allergies | 0
fever | 24
leukocytosis | 24
culture | 24
negative | 24
punch biopsy | 24
histopathologic examination | 24
sub-corneal pustules | 24
intraepidermal pustules | 24
spongiosis | 24
neutrophil | 24
histiocyte infiltration | 24
exocytosis of eosinophils | 24
AGEP | 24
tigecycline stopped | 24
methylprednisolon | 24
local moisturizers | 24
topical steroids | 24
new pustules stopped | 72
healing | 72
exfoliation | 72
dermatologic pathologies | 360
sepsis | 2160
multiorgan failure | 2160
death | 2160