18 years old | 0
female | 0
admitted to the hospital | 0
increasing abdominal pain | -72
frequency and intensity of uterine contractions | -72
suprapubic pain | -72
urinary discomfort | -72
vaginal discharge | -72
abnormal vaginal discharge | -72
low abdominal pain | -72
positive fetal fibronectin test | -72
seizures as a child | -100000
depression | -100000
remote history of smoking | -100000
respiratory symptoms | -168
shortness of breath | -168
coughing | -168
rhinorrhea | -168
water damage | -168
utilizing a humidifier | -168
moved out of the location | -168
G1P0 | 0
34 weeks 6 days | 0
routine and consistent prenatal care | 0
non-completion of glucose tolerance test (GTT) | 0
normotensive | 0
appropriate fetal growth | 0
total weight gain of 14 pounds | 0
normal 20-week anatomy scan | 0
persistent productive cough | 0
shortness of breath | 0
intermittent nausea | 0
denies chest pain | 0
denies lower extremity swelling or pain | 0
tachycardia of 111 beats per minute | 0
rupture of membranes | 0
closed cervix | 0
lungs were clear to auscultation | 0
lower extremity edema 1+ | 0
urinary tract infection | 0
unknown group B streptococcus (GBS) status | 0
steroid prophylaxis | 0
GBS prophylaxis | 0
ampicillin intravenous (IV) | 0
cefazolin | 0
cesarean section | 72
fever of 40.2°C (104.3°F) | 96
tachycardia | 96
suspicion of sepsis | 96
gentamicin | 96
clindamycin | 96
endometritis | 96
portable chest x-ray (CXR) | 96
no acute cardiopulmonary disease | 96
blood cultures drawn | 96
influenza type A and B | 96
respiratory syncytial virus (RSV) | 96
urine Legionella antigen | 96
urine mycoplasma | 96
urine streptococcus antigen | 96
thyroid function tests | 96
lower extremity ultrasound (US) | 96
deep vein thrombosis (DVT) | 96
transaminitis | 96
right upper quadrant (RUQ) ultrasound | 120
normal liver and common bile duct (CBD) | 120
questionable mild gallbladder wall thickening | 120
ceftriaxone 1 gm IV | 120
azithromycin 500 mg IV | 120
urinary tract infection treatment | 120
levofloxacin | 144
recurrent fever | 144
tachycardia (heart rate up to 130 beats per minute) | 144
transferred to the Intensive Care Unit (ICU) | 144
computed tomography (CT) scan of the chest | 168
bilateral small basilar infiltrates | 168
ground glass opacity in the left upper lobe | 168
CT scan of the abdomen and pelvis | 168
hepatic steatosis | 168
hepatomegaly | 168
Infectious disease (ID) consultation | 168
oral azithromycin | 216
treated for endometritis with Zosyn | 216
condition steadily improved | 216
transferred out of the ICU | 288
discharged | 216
additional 4 days of therapy with azithromycin | 216
normal blood pressure | 0
transaminitis peaked | 288
aspartate amino-transferase (AST) | 288
alanine aminotransferase (ALT) | 288
international normalized ratio (INR) | 288
bilirubin | 288
gastroenterology service consulted | 288
extensive serologic evaluation | 288
hepatitis panel | 288
herpes simplex virus (HSV)-1 and HSV-2 IgM | 432
parvovirus B19 IgM | 432
ammonia level | 288
repeat US | 288
hepatic steatosis | 288
hepatomegaly | 288
edema adjacent to the gallbladder | 288
gallbladder itself and the common bile duct (2 mm) | 288
hepatic arterial and venous flow | 288
N-acetyl cysteine by mouth | 288
loading dose plus 15 out of 17 follow-up doses | 288
refused the last 2 doses | 288
repeat liver function tests (LFT) | 432
normalized | 432
mild thrombocytopenia | 96
anemia | 96
haptoglobin | 96
lactate dehydrogenase (LDH) | 96
sodium level | 0