52 years old | 0
female | 0
abdominal pain | 0
nausea | 0
vomiting | 0
increased level of liver enzyme alanine aminotransferase | -840
positive autoimmune antibody | -840
elevated immunoglobulin G | -840
coarse liver surface | -840
overlap syndrome predominantly with features of autoimmune hepatitis | -840
high dose of ursodeoxycholic acid | -840
prednisolone | -840
liver biopsy | -840
mild heartburn | -48
abdominal pain | -48
nausea | -24
vomiting | -24
diarrhea | -24
abdominal tenderness | 0
mild fever | 0
tachycardia | 0
tachypnea | 0
reduced white blood cells | 0
reduced platelets | 0
decreased neutrophil | 0
elevated C-reactive protein | 0
elevated aspartate aminotransferase | 0
elevated ALT | 0
elevated gamma glutamyl transferase | 0
elevated prothrombin time international normalized ratio | 0
huge stomach with layered wall thickening | 0
air in the stomach wall | 0
decrease of mucosal enhancement | 0
necrotizing gastritis | 0
septic shock | 0
intravenous hydration | 0
antibiotic treatment | 0
inotropics | 0.5
fluid treatment | 0.5
decreased blood pressure | 0.5
increased blood pressure | 2
severe stress-induced cardiomyopathy | 3
extracorporeal membrane oxygenation | 3
cardiac arrest | 3
death | 3