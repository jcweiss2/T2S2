36 years old | 0
woman | 0
cerebral palsy | 0
severe kyphoscoliosis | 0
admitted to respiratory intensive care unit | 0
severe respiratory failure | 0
pneumonia | 0
respiratory condition deteriorated | 24
orotracheal intubation | 24
invasive mechanical ventilation | 24
tracheotomy | 672
persistent type II respiratory failure | 672
continuous ventilatory support | 672
peristomal skin diastase | 1344
wide tracheocutaneous fistula | 1344
excessive cuff pressure | 1344
difficult ventilatory support management | 1344
size of fistula approximately 4 cm in diameter | 1344
surgical repair impossible | 1344
tracheotomy with suturing of distal stump | 1344
suturing of previous tracheotomy breach | 1344
careful dissection of trachea | 1344
anonymous artery protected by muscle flap | 1344
mechanical ventilation hindered | 1344
reduced length of residual trachea | 1344
cannula or endotracheal tube not secured | 1344
cuff securing system in two main bronchi | 1344
selectively intubated main bronchi | 1344
bronchoscopy guidance | 1344
two tubes (Portex Tracheal Tube) | 1344
inflating cuffs at both main stem bronchi inlets | 1344
Y-shaped bridge added | 1344
ventilator connection | 1344
adequate minute volume | 1344
correct blood gas levels | 1344
no significant leaks | 1344
ventilatory parameters stable | 1344
bronchoscopic examination | 1824
no evidence of alterations | 1824
died | 3456
sepsis | 3456
