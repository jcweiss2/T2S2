58 years old | 0
    female | 0
    hypertension | 0
    stage 3 chronic kidney disease | 0
    undiagnosed muscle spasticity | 0
    presented to the emergency department | 0
    worsening upper extremities tremors | -72
    paresthesia | -72
    limb weakness | -72
    pins and needle sensation | -72
    temperature of 103 F | 0
    tachycardia | 0
    hypertensive | 0
    tachypneic | 0
    oxygen saturation 97% | 0
    ill-appearing | 0
    coarse tremors | 0
    neurology examination | 0
    bilateral upper extremities strength 3/5 | 0
    bilateral lower extremities strength 4/5 | 0
    decreased sensation | 0
    lungs clear to auscultation | 0
    initial impression sepsis | 0
    initial impression fever of unknown origin | 0
    started on cefepime | 0
    started on vancomycin | 0
    started on metronidazole | 0
    non-significant WBC count | 0
    non-significant lactic acid | 0
    non-significant inflammatory markers | 0
    negative blood cultures | 0
    negative urine cultures | 0
    negative respiratory cultures | 0
    lumbar puncture | 0
    cerebrospinal fluid analysis | 0
    ruled out meningitis | 0
    chest x-ray unremarkable | 0
    abdominal ultrasound unremarkable | 0
    magnetic resonance imaging of head | 0
    magnetic resonance imaging of spine | 0
    ruled out intracranial pathology | 0
    ruled out osteomyelitis of spine | 0
    neurology consulted | 0
    electroencephalography | 0
    ruled out seizure disorder | 0
    ruled out Guillain Barre Syndrome | 0
    ruled out Alcohol withdrawal syndrome | 0
    toxicology consulted | 0
    ruled out anticholinergic toxicity | 0
    persistent fever | 96
    worsening mental status | 96
    visual hallucinations | 96
    hyperpyrexia | 96
    ocular clonus | 96
    profound muscle rigidity | 96
    somnolent | 96
    unable to follow command | 96
    continuous tremors | 96
    lorazepam 7 mg given | 96
    phenobarbital 250 mg given | 96
    no improvement | 96
    intravenous haloperidol | 96
    decline in condition | 96
    rapid response called | 96
    evaluated by ICU team | 96
    minimally responsive | 96
    tachypnea 40 breaths/minute | 96
    ABG pH 7.3 | 96
    ABG PCO2 28.6 | 96
    ABG PaO2 70 | 96
    intubated | 96
    respiratory distress | 96
    continued worsening mental status | 96
    transferred to ICU | 96
    possible diagnosis neuroleptic malignant syndrome | 96
    possible diagnosis baclofen withdrawal | 96
    normal serum creatinine kinase | 96
    normal lactic acid | 96
    bromocriptine started | 96
    no improvement of symptoms | 96
    home medications reviewed | 96
    oral baclofen 10 mg 3 times a day | 0
    stopped baclofen 3 days | 0
    baclofen restarted | 96
    resolution of fever | 144
    improvement in mental status | 144
    complete cessation of tremors | 144
    extubated | 192
    transferred to medical floor | 192
    discharged | 192
    