23 years old | 0
female | 0
presented to the Emergency Department | 0
painful right breast | -12
swollen right breast | -12
right breast entirely discoloured | 0
offensive nipple discharge | 0
breast pruritus near the inframammary fold | -72
dizziness | 0
nausea | 0
vomiting episodes | 0
denied trauma to the breast | 0
obesity | 0
BMI 34.7 | 0
polycystic ovarian syndrome | 0
alert | 0
oriented | 0
blood pressure 80/60 mmHg | 0
heart rate 130 beats/min | 0
saturations 95% on room air | 0
temperature 35.8 °C | 0
swollen right breast | 0
tender right breast | 0
discolouration | 0
erythema to the margins | 0
associated bullae | 0
left breast unremarkable | 0
severe sepsis | 0
end organ dysfunction | 0
white cell count 27.85 × 10^9/L | 0
neutrophilia 23.6 × 10^9/L | 0
C-reactive protein 400 mg/L | 0
metabolic acidosis | 0
pH 7.06 | 0
lactate 8.8 mmol/L | 0
creatinine 394 umol/L | 0
estimated glomerular filtration rate 13 mL/min | 0
international normalized ratio 1.8 | 0
activated partial thromboplastin time 44 s | 0
intravenous crystalloid resuscitation 5 L | 0
inotropic support | 0
metaraminol boluses 2 mg total | 0
adrenaline boluses 1.1 mg total | 0
anuric | 0
noradrenaline infusion | 0
central line | 0
peak pre-operative rate 1.5 mg/h | 0
vasopressin infusion 4 units/h | 0
possible penicillin allergy | 0
renal-adjusted doses of IV meropenem | 0
IV clindamycin | 0
IV vancomycin | 0
taken to operating theatre within 3 hours | 3
emergency right mastectomy | 3
debridement of all necrotic tissue | 3
preserving pectoralis major | 3
consulted haematologist | 3
coagulopathy | 3
fresh frozen plasma 2 units | 3
wound packed | 3
vacuum assisted closure dressing | 3
transferred to intensive care unit | 3
intubated | 3
sedated | 3
continuous renal replacement therapy commenced | 3
troponin-I rise to 20,203 ng/L | -18
ST elevation in inferior leads | -18
troponin-I peaked >40,000 ng/L | -18
adrenaline weaned | -18
vasopressin weaned | -18
packed cells transfused 2 units | -18
haemoglobin 83 g/L | -18
sepsis driven myocardial ischaemia | -18
aspirin commenced | -18
IV heparin infusion commenced | -18
noradrenaline infusion peaked at 3 mg/hour | 6
noradrenaline weaned from 6 hours post-operatively | 6
noradrenaline cessation on day 2 post-op | 48
CRRT ceased | 12
improving urine output | 12
improving renal function | 12
extubated on day 8 | 192
wound debridements | 24
VAC applications on days 1, 5, and 9 | 24
tissue culture positive for streptococcus pyogenes | 24
confirmed no allergies on day 5 | 120
antibiotic therapy changed to benzylpenicillin | 120
inflammatory markers improved | 120
afebrile on day 5 | 120
stepped down to oral amoxicillin | 456
resolving ST elevation | 192
transthoracic echocardiogram | 192
ejection fraction 55% | 192
normal systolic function | 192
small sized septal and inferior wall motion abnormality | 192
mild hypokinesis of segments | 192
CT coronary angiograms planned as outpatient | 192
transferred to tertiary hospital on day 16 | 384
further debridement | 384
skin grafting from left thigh | 384
all blood parameters normalised | 384
stable under plastics team | 384
discharged home | 432
necrotising fasciitis of the breast | 0
primary idiopathic necrotizing fasciitis of the breast | 0
streptococcal toxic shock syndrome | 0
myocardial infarction | -18
full recovery | 432
no further complications | 432
