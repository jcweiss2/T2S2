29 years old | 0
    Caucasian | 0
    diamniotic dichorionic twin pregnancy | 0
    24+1 weeks of gestation | 0
    admitted to the obstetric unit | 0
    preterm premature rupture of membranes (pPROM) | 0
    spontaneous abortion in the first trimester | -672
    hyperemesis gravidarum | -672
    chlorpromazine | -672
    amniocentesis | -336
    CGH array | -336
    discordant growth between the twins | -336
    35% discordance | -336
    first fetus small for gestational age | -336
    ARSA (aberrant right succlavian artery) | -336
    right ventriculum hypertrophy (first fetus) | -336
    double left renal artery (second fetus) | -336
    pPROM of one of two sacs | 0
    no fever | 0
    no signs of chorioamnionitis | 0
    WBC 12,970 | 0
    CRP 0.58 | 0
    PCT negative | 0
    no uterine contractions | 0
    cardiac activity (both fetuses) | 0
    cephalic presentation (both fetuses) | 0
    corticosteroids (betamethasone 12 mg i.m.) | 0
    intravenous atosiban | 0
    magnesium sulfate infusion | 0
    cefazoline 1 g i.v. | 0
    bemiparine 3500 IU s.c. | 0
    WBC 14,920 cells/microL | 96
    CPR 1.34 mg/dL | 96
    PCT negative (day 4) | 96
    no fever | 96
    no signs of infection | 96
    WBC 10,100 cells/microL | 168
    CPR negative | 168
    PCT negative (day 11) | 168
    uterine contractions | 192
    substantial discharge of amniotic fluid | 192
    no tocolytics | 192
    magnesium sulfate restarted | 192
    WBC 13,490 cells/microL | 192
    CPR negative | 192
    PCT negative (day 12) | 192
    delivered the first fetus | 336
    umbilical cord clamped and kept in uterus | 336
    newborn girl (330 g) | 336
    transferred to NICU | 336
    right ventricular hypertrophy confirmed | 336
    died after 7 days | 408
    mother intensively monitored | 336
    no fever | 336
    no clinical symptoms | 336
    WBC 10,320 cells/microL | 552
    tocolysis restarted with atosiban | 336
    bemiparine 3500 IU s.c. continued | 336
    cefazoline 3 g/day continued | 336
    fetus growth rate slowing | 336
    no anomalies on Doppler scans | 336
    pathological pattern of cardiotocography | 672
    low variability | 672
    late decelerations (ACOG III) | 672
    cesarean section | 672
    second baby girl (960 g) | 672
    Apgar score 7/10 at 5 min | 672
    intubated | 672
    admitted to NICU | 672
    external pulmonary support | 672
    surfactant treatment | 672
    received 3 blood units | 672
    erythropoietin for anemia | 672
    good heart morphology and activity | 672
    normal cerebral ultrasound scans | 672
    normal electroencephalograms | 672
    normal urinary function | 672
    normal gastroenterological function | 672
    started eating | 672
    parenteral feeding stopped | 672
    discharged after 2 months | 672
    weight 2050 g | 672
    no neurological defects at 6-month follow-up | 672
    no cardiac defects at 6-month follow-up | 672
    no other defects at 6-month follow-up | 672
    mother continued antibiotic (ceftriaxone) | 672
    anti-thrombotic (bemiparine) | 672
    uterotonic therapy (oxytocine) | 672
    no fever | 672
    no pain | 672
    no post-operative complications | 672
    blood exams returned to normal | 672
    discharged on day 32 | 672
    bemiparine 3500 IU for 15 days | 672
    cefuroxime 500 mg tablets | 672