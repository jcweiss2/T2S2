44 years old|0
male|0
Covid-19 infection|0
mildBingflu like syndrome|-144
fever|-144
chills|-144
headache|-144
myalgia|-144
cough|-144
fatigue|-144
RT-PCR positive|0
referred to emergency ward|0
respiratory failure|0
oxygen supply with cPAP|0
chest CT scan|0
denied other symptoms|0
diabetes mellitus type 2|0
obesity|0
mild cognitive impairment|0
psychotic disorder|0
transferred to intensive-care unit|0
acute renal failure|0
bacteric pulmonary sovrainfection|0
complete atelectasia of left lung|0
tracheostomy|0
systemic sepsis|0
urinary tract infection|0
high blood pressure levels|0
antihypertensive therapy|0
transferred to Rehabilitation ward|0
normal consciousness (GCS=15)|0
no cranial nerves abnormality|0
upper limbs strength (MRC scale)|0
lower limbs strength (MRC scale)|0
absent deep tendon reflexes|0
normal plantar response|0
no sensitivity alteration|0
good respiratory gas exchanges|0
axonal polineuropathy|0
absence of sural nerve SAP|0
absence of common peroneal nerve CMAP|0
decreased tibial nerve velocity|0
severely decreased tibial nerve CMAP amplitude|0
decreased ulnar nerve SAP amplitude|0
Motricity Index assessment|0
Timed Up and Go Test assessment|0
Barthel Index assessment|0
rehabilitation treatment|0
respiratory rehabilitation|0
motor rehabilitation|0
training program|0
sessions per week|0
duration of rehabilitation program|0
passive or active motion session|0
breathing exercises|0
coordination exercises|0
recovery of standing position|0
reconditioning of walking|0
functional activities|0
overground ambulatory training|0
prescription of orthosis|0
TUG test improvement (20.29 s)|0
upper extremities recovery (right side)|0
lower extremities impairment (left side)|0
lower extremities mild improvement (right side)|0
no ankle dorsiflexors activity|0
Barthel Index improvement (89)|0
self-care activities improvement|0
mobility improvement|0
needs two sticks|0
wears ankle-foot orthosis|0
partial recovery|0
