69 years old | 0
    woman | 0
    presented with general myalgia | -72
    presented with fever | -72
    presented with nausea | -72
    resided in urban area | -240
    picked ginkgo nuts | -240
    visited local hospital | -72
    right upper abdominal tenderness | -72
    referred to hospital | -72
    vital signs checked | 0
    blood pressure 110/90 mm Hg | 0
    pulse rate 78/min | 0
    respiratory rate 24/min | 0
    body temperature 38.5℃ | 0
    enlarged cervical lymph nodes | 0
    right upper abdominal tenderness | 0
    rebound tenderness | 0
    no eschar on trunk | 0
    white blood cell count 4,510/mm3 | 0
    segmented neutrophils 70.6% | 0
    hemoglobin 14.0 g/dL | 0
    platelet count 57 × 103/mm3 | 0
    C-reactive protein 17.51 mg/dL | 0
    aspartate aminotransferase 374 IU/L | 0
    alanine aminotransferase 254 IU/L | 0
    alkaline phosphatase 982 IU/L | 0
    lactate dehydrogenase 1,141 IU/L | 0
    total protein 7.0 g/dL | 0
    albumin 3.8 g/dL | 0
    total bilirubin 1.2 mg/dL | 0
    chest radiography no abnormalities | 0
    electrocardiogram no abnormalities |? 0
    abdominal CT edematous GB wall | 0
    GB stones | 0
    acute calculous cholecystitis suspected | 0
    ceftriaxone initiated | 0
    percutaneous cholecystostomy performed | 0
    sustained nausea | 0
    sustained abdominal pain | 0
    developed progressive shortness of breath | 96
    increased sputum production | 96
    hypoxemia | 96
    confusion | 96
    oxygen delivery 5 L/min | 96
    arterial blood gas analysis pH 7.45 | 96
    PaCO2 36 mm Hg | 96
    PaO2 67 mm Hg | 96
    HCO3- 25 | 96
    follow-up chest radiography airspace consolidation | 96
    endotracheal intubation | 96
    admitted to ICU | 96
    maculopapular rash on trunk | 120
    maculapapular rash on face | 120
    sputum culture negative | 120
    blood culture negative | 120
    scrub typhus suspected | 120
    acute cholecystitis | 120
    ARDS | 120
    doxycycline treatment | 120
    piperacillin treatment | 120
    serologic test positive | 120
    Orientia tsutsugamushi titer 1:5,120 | 120
    multi-organ function normal | 216
    mental alertness improved | 216
    follow-up chest radiography resolved | 216
    discharged | 312
    complete blood count normal | 312
    biochemistry normal | 312
    recovered | 312
    cholecystostomy catheter removed | ?
    elective cholecystectomy | ?
    stones three | ?
    black pigment stones | ?
    no complications | ?
    eschars | 0
    lymphadenopathy | 0
    maculopapular rash | 120
    fever | -72
    headache | ?
    anorexia | ?
    nausea | -72
    diffuse myalgias | -72
    abdominal pain | 0
    relative bradycardia | 0
    no septic shock | ?
    no meningoencephalitis | ?
    no acute renal failure | ?
    no hepatitis | ?
    no gastrointestinal bleeding | ?
    vasculitis | ?
    perivasculitis | ?
    leukocyte infiltration | ?
    pre-existing GB stones | -240
    symptoms of acute cholecystitis | -72
    ARDS | 96
    confusion | 96
    mechanical respiration | 96
    ICU admission | 96
    elderly patient | 0
    severe complications | 0
    relative bradycardia | 0
    pulse-temperature dissociation | 0
    history of exposure | -240
    symptoms present | -72
    clinical signs present | 0
    lab results present | 0
    endemic area | ?
    eschars not found | 0
    skin eruptions present | 120
    heart rate below 100 beats/min | 0
    pyrexia | -72
    prompt doxycycline treatment | 120
    clinical illness shortened | 312
    mortality reduced | 312
    