39 years old | 0
female | 0
height 155 cm | 0
weight 44.5 kg | 0
mild dyspnea | 0
adenoid cystic carcinoma in the carina | 0
carinal resection | 0
reconstruction | 0
chest computed tomography | -24
bronchoscopy | -24
mass in the left mainstem bronchus | -24
mass extended to the carina and right mainstem bronchus | -24
internal diameter of the RMB 11 mm | -24
length of the RMB 12 mm | -24
length of the distal LMB not involved by the mass 20 mm | -24
preoperative examinations normal findings | -24
moderate obstructive pattern of the pulmonary function test | -24
forced expiratory volume in one second 1.88 liter | -24
forced vital capacity 2.81 liter | -24
ratio of forced expiratory volume in one second to forced vital capacity 67% | -24
general anesthesia induced | 0
target-controlled infusion of propofol | 0
target-controlled infusion of remifentanil | 0
rocuronium administered | 0
tracheal intubation | 0
right-sided double-lumen tube | 0
patient moved to the right lateral position | 0
left bronchi and vasculature dissected | 0
thoracoscopic surgery under right OLV | 0
arterial oxygen tension 462 mmHg | 20
inspired oxygen fraction 1.0 | 20
right-sided double-lumen tube replaced with a single-lumen endotracheal tube | 20
bronchial blocker placed into the RMB | 20
patient moved to the left lateral position | 20
right thoracotomy | 20
peak airway pressure 28 cmH2O | 40
tidal volume 300 ml | 40
arterial oxygen tension 110 mmHg | 40
inspired oxygen fraction 1.0 | 40
carinal resection | 40
LMB resected | 40
sterile reinforced endotracheal tube inserted into the separated LMB | 40
airway pressure increased to 35 cmH2O | 40
oxygen saturation by pulse oximetry decreased to 70% | 40
RMB resected | 40
additional sterile endotracheal tube inserted into the separated right bronchus | 40
differential bilateral lung ventilation | 40
oxygen saturation by pulse oximetry restored to 100% | 42
carina removed | 42
lower trachea resected | 42
separated RMB anastomosed with the resected trachea | 42
no air leak in the anastomotic site | 42
left lung removed | 42
left endobronchial tube removed | 42
non-dependent right lung ventilated | 42
airway pressure lower than 20 cmH2O | 42
oxygen saturation by pulse oximetry decreased below 80% | 42
left endobronchial tube reinserted | 42
two-lung ventilation | 42
oxygen saturation by pulse oximetry maintained 100% | 47
right OLV reattempted | 47
oxygen saturation by pulse oximetry decreased below 90% | 50
left pulmonary artery clamped | 50
oxygen saturation by pulse oximetry maintained 100% | 50
left main pulmonary artery ligated | 50
left endobronchial tube removed | 50
right thoracotomy closed | 50
arterial oxygen tension 360 mmHg | 110
inspired oxygen fraction 1.0 | 110
patient moved to the right lateral position | 110
left thoracotomy | 110
left pulmonary artery and veins resected | 110
left pneumonectomy completed | 110
patient moved to the supine position | 110
chin tightly sutured to the chest | 110
tracheal extubation | 110
patient transferred to the intensive care unit | 110
discharged on the 13th postoperative day | 312