66 years old | 0
male | 0
diabetes mellitus | -672
obesity | -672
consumed rice wine | -672
colonoscopy | 0
polypectomy | 0
endoscopic mucosal resection | 0
preventive hemoclips | 0
discharged from endoscopy room | 0
right abdominal pain | 24
tenderness | 24
rebound tenderness | 24
severe infection | 24
white blood cell count elevated | 24
C-reactive protein elevated | 24
blood urea nitrogen elevated | 24
creatinine elevated | 24
lactic acid elevated | 24
total bilirubin elevated | 24
abdominopelvic CT | 24
multiple air bubbles in abdominal muscles | 24
broad-spectrum antibiotic therapy | 24
piperacillin/tazobactam | 24
emergency exploratory laparotomy | 44
laparoscopic right hemicolectomy | 44
multiple-organ failure | 44
metabolic acidosis | 44
diagnosis of necrotizing fasciitis | 48
surgical debridement | 48
drainage | 48
renal replacement therapy | 48
intensive care unit | 48
imipenem-resistant Acinetobacter baumannii | 72
extended spectrum beta-lactamase negative Escherichia coli | 72
septic shock | 840
multiple-organ failure | 840
death | 840