53 years old | 0
male | 0
admitted to hospital | 0
hydronephrosis | 0
urolithiasis | 0
ureteral stent placement | 0
hypertension | -672
hypercholesterolemia | -672
violent pain in epigastric region | -72
nausea | -72
afebrile | -72
pale | -72
sweaty | -72
cold | -72
sinus tachycardia | -72
hypotension | -72
distended abdomen | -72
moderate tenderness in epigastrium | -72
moderate tenderness in left hypochondrium | -72
anemia | -72
thrombopenia | -72
increased international normalized ratio | -72
increased activated partial thromboplastin time | -72
increased alanine aminotransferase | -72
decompensated metabolic acidosis | -72
rapid resuscitation | -72
free fluid in peritoneal cavity | -72
dilated left hepatic artery | -72
bleeding point | -72
aneurysm of 20 x 18 mm | -72
large intraperitoneal effusion | -72
heterogeneous hepatic enhancement | -72
hepatic hypoperfusion | -72
laparotomy | -48
massive hemoperitoneum | -48
ruptured aneurysm of hepatic arterial branch | -48
fresh blood clot | -48
diffused disruption of vascular wall | -48
clamping of aneurysm | -48
isolation of proximal stump | -48
aneurysmectomy | -48
intensive care unit | 0
correction of acidosis | 0
stabilization of hemodynamic conditions | 0
transfer to surgical ward | 48
noninfectious fever | 48
discharged from hospital | 360
good clinical condition | 360
asymptomatic | 360
liver function tests within normal reference ranges | 360