60 years old | 0
female | 0
impaired consciousness | -1
atrial fibrillation | -672
dilated cardiomyopathy | -672
oral warfarin | -672
biventricular pacing implantable cardioverter defibrillator | -672
found lying at home | -1
transported to hospital | -1
Japan Coma Scale score II-10 | 0
Glasgow Coma Scale score 14 | 0
no clear neurological deficits | 0
non-contrast head CT | 0
hemorrhage in third and fourth ventricles | 0
hemorrhage in bilateral lateral ventricles | 0
brain 3D-CTA | 0
spot enhancement on lateral wall of anterior horn of left lateral ventricle | 0
blood pressure control | 0
ventricular drainage not performed | 0
cerebral angiograph | 72
aneurysm at distal site of mLSA | 72
embolization | 72
endovascular treatment | 72
N-butyl-2-cyanoacrylate | 72
general anesthesia | 72
right femoral introducer replaced | 72
systemic heparinization | 72
guiding sheath navigated | 72
distal access catheter | 72
Marathon catheter advanced | 72
contralateral approach | 72
DeFrictor nano catheter | 72
TENROU S10 guide wire | 72
mLSA cannulation | 72
selective angiography | 72
NBCA-Lipiodol mixture injected | 72
aneurysm filled with NBCA | 72
postoperative head CT | 96
no hemorrhagic complications | 96
no cerebral infarction | 96
sepsis triggered by pneumonia | 120
decrease in muscle strength | 120
disuse | 120
rehabilitation | 720
discharged to home | 720
modified Rankin Scale 1 | 720
DRESS syndrome | -672 
fever | -672
rash | -672 
acne | -672 
minocycline | -672 
increased WBC count | 0
eosinophilia | 0
systemic involvement | 0
diffuse erythematous or maculopapular eruption | 0
pruritis | 0 
DRESS syndrome | 0 
fever persisted | 0
rash persisted | 0 
discharged | 24