32 years old | 0
    woman | 0
    family history of polycystic kidney disease | 0
    referred from a local hospital with a hemorrhagic left renal cyst | -24
    received one packed red blood cell | -24
    vital signs were stable | 0
    abdomen was distended | 0
    left kidney was palpable | 0
    abdomen was soft without signs of peritonitis | 0
    hemoglobin level of 9.6 g/dl | 0
    creatinine level of 64 μmol/l | 0
    enhanced CT of the abdomen demonstrated features of polycystic kidneys | 0
    enlarged left kidney | 0
    hemorrhagic component without associated extravasation | 0
    images discussed with intervention radiologist confirmed no signs of active bleeding | 0
    stability of the patient | 0
    discharged home | 0
    seen in the clinic 10 days later | 240
    still symptomatic with abdominal pain | 240
    abdomen was distended more | 240
    decision made to admit her electively for angioembolization | 240
    repeated enhanced CT showed a left complex renal cyst with thick septation | 240
    contrast extravasation suggesting active bleeding | 240
    angiogram showed no evidence of extravasation | 240
    significant tortuous arteries in the lower pole that were embolized | 240
    increasing abdominal distention | 240
    dropping of hemoglobin even after angioembolization | 240
    necessitated surgical intervention to evacuate the hematoma | 240
    intraoperatively, capsulated mass around 30 cm crossing the midline with bleeding around it | 240
    radical nephrectomy done without clear spillage of the tumor | 240
    bowel injury repaired primarily intraoperatively | 240
    postoperatively, chyle leak | 240
    chyle leak managed conservatively | 240
    histopathology revealed embryonal rhabdomyosarcoma | 240
    case discussed in the tumor board | 240
    planned for chemotherapy | 240
    multiple peritoneal metastatic deposits | 240
    liver metastasis | 240
    bone metastasis | 240
    received first cycle of Dactinomycin | 240
    received Vincristine | 240
    received Cyclophosphamide | 240
    complicated by sepsis | 240
    pulmonary embolism | 240
    profound neutropenia | 240
    intensive care unit admission | 240
    passed away 88 days post-operatively | 2112