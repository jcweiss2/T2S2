34 years old | 0
    pregnant | 0
    female | 0
    ITP | 0
    anemia | 0
    suspected hypoplastic anemia | 0
    blood transfusion during pregnancy | 0
    iron supplement | 0
    admitted to hospital | 0
    threatened preterm labor | 0
    low hemoglobin (7.1 g/dl) | 0
    low platelet count (27 × 10³/μl) | 0
    IVIG 0.5 g/kg/day for 4 days | 0
    hemoglobin increased to 8.3 g/dl | 6
    hemoglobin dropped to 7.8 g/dl | 96
    platelet count 22 × 10³/μl | 96
    hemoglobin 8.6 g/dl | 48
    platelet 25 × 10³/μl | 48
    IUGR diagnosis | 0
    elective cesarean section | 0
    oral dexamethasone 8 mg every 12 h | -72
    last dose completed 3.5 h before surgery | -3.5
    blood transfusion | 0
    blood products transfused | 0
    baby girl born | 0
    IUGR | 0
    weight 2235 g | 0
    Apgar scores 9 at 1 min | 1
    Apgar scores 10 at 5 min | 5
    mild grunting at 1 hour | 1
    supplemental oxygen 2 L/min for 1 hour | 1
    mild respiratory distress at 6 hours | 6
    admission to neonatal ward | 6
    grunting | 6
    equal air entry bilaterally | 6
    mild subcostal retraction | 6
    normal heart sounds | 6
    oxygen saturation 94-95% | 6
    respiratory rate 64/min | 6
    temperature 36.6°C | 6
    heart rate 148/min | 6
    blood pressure 65/35 mmHg | 6
    TTN suspected | 6
    nasal cannula 2 L/min for 1 day | 6
    weaned on third day | 72
    discontinued on third day | 72
    neonatal jaundice on second day | 48
    phototherapy for two days | 48
    feeding started on second day | 48
    full feed by third day | 72
    discharged on fourth day | 96
    chest X-ray suggestive of TTN | 6
    normal blood counts | 8
    normal serum electrolytes | 8
    negative blood culture | 8
    slightly hemolyzed potassium sample | 44
    