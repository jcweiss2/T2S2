68 years old| 0
woman | 0
jaundice | -72
jaundice developed 3 days before the visit | -72
general weakness | -72
fatigue | -72
decreased appetite | -72
icteric sclera | 0
no other abnormal findings on physical examination | 0
vital signs normal | 0
acute bronchitis | 0
tranexamic acid | 0
N-acetylcysteine | 0
dihydrocodeine | 0
azithromycin | 0
no history of allergic diseases | 0
denied alcohol consumption | 0
denied smoking | 0
white blood cell count 9,100/mm³ | 0
hemoglobin level 13.7 g/dL | 0
platelet count 149,000/mm³ | 0
aspartate aminotransferase level 1,631 IU/L | 0
alanine aminotransferase level 1,711 IU/L | 0
total bilirubin level 24.20 mg/dL | 0
direct bilirubin level 14.99 mg/dL | 0
alkaline phosphatase level 226 IU/L | 0
gamma-glutamyl transferase level 232 U/L | 0
total protein concentration 5.3 g/dL | 0
albumin level 3.1 g/dL | 0
blood urea nitrogen level 6.4 mg/dL | 0
creatinine level 0.5 mg/dL | 0
sodium concentration 142 mmol/L | 0
potassium concentration 3.7 mmol/L | 0
amylase level 29 IU/L | 0
lipase level 53 IU/L | 0
ammonia concentration 163 μMol/L | 0
prothrombin time extended to 37.5 seconds | 0
partial thromboplastin time extended to 55.9 seconds | 0
high sensitivity C-reactive protein level 0.932 mg/dL | 0
hepatitis A virus IgM antibody negative | 0
hepatitis B surface antigen negative | 0
anti-HCV negative | 0
Epstein-Barr virus IgM antibody negative | 0
cytomegalovirus IgM negative | 0
cytomegalovirus real-time PCR negative | 0
herpes simplex virus IgM positive | 0
herpes simplex virus IgG positive | 0
toxoplasma IgM negative | 0
human immunodeficiency virus serum tests negative | 0
antinuclear antibody negative | 0
anti-mitochondrial antibody negative | 0
anti-smooth muscle antibody negative | 0
liver kidney microsomal antibody negative | 0
IgG serum level 774.6 mg/dL | 0
CT showed normal liver before azithromycin treatment | 0
periportal edema | 0
gallbladder wall edema | 0
small amount of ascites | 0
clinically suspected azithromycin-induced liver injury | 0
medications discontinued | 0
RUCAM score for azithromycin 7 (probable) | 0
RUCAM scores for tranexamic acid, N-acetylcysteine, dihydrocodeine 4 (possible) | 0
R value more than 5 (hepatocellular type) | 0
diagnosis of azithromycin-induced liver injury | 0
diagnosis of acute liver failure | 0
medical treatment received | 0
laboratory test values worsened | 0
flapping tremor | 72
decreased consciousness to drowsiness | 72
hepatic encephalopathy | 72
consciousness deteriorated to semi-coma | 168
emergency living donor liver transplantation | 192
recovery of consciousness | 192
recovery of liver function | 192
discharged after 20 days of transplant | 480
alive | 480
asymptomatic | 480
adequate liver graft function | 480
fulminant hepatitis | 192
zone 3 necrosis | 192
extensive hepatocyte death | 192
jaundice developed 4 days after azithromycin prescription | 0
acute jaundice | 0
abdominal pain | 0
