79 years old | 0
male | 0
white | 0
admitted to the hospital | 0
laparoscopic cholecystectomy | -504
converted to open cholecystectomy | -504
gangrenous perforated gallbladder | -504
inability to obtain the critical view | -504
tubular structure | -504
ligated | -504
cystic artery | -504
cystic duct | -504
single drain | -504
persistent high-output bilious drainage | -504
discharged | -288
jaundice | -192
weakness | -192
fatigue | -192
pain | -192
CT scan | -192
nuclear cholescintigraphy scan | -192
biliary leak | -192
free intra-abdominal fluid | -192
biliary peritonitis | -192
broad spectrum antibiotics | -168
atrial fibrillation | -168
rapid ventricular response | -168
bilirubin level | -168
protein-calorie malnutrition | -168
albumin | -168
percutaneous cholangiogram | -168
hilar ligation | -168
hepatic duct | -168
inability to pass a wire | -168
inability to pass a catheter | -168
right posterior percutaneous cholangiogram catheter | -168
right anterior percutaneous cholangiogram catheter | -168
definitive biliary diversion | -168
high calorie | -168
high protein enteral nutrition | -168
nasogastric Dobhoff tube | -168
follow-up | 336
improved substantially | 336
repeat CT scan | 336
abdominal fluid collections | 336
bilirubin | 336
albumin | 336
prealbumin | 336
definitive biliary reconstruction | 504
porta dissection | 504
common hepatic arteries | 504
proper hepatic arteries | 504
identification of percutaneous biliary catheters | 504
transection of CBD | 504
removal of clips | 504
bile drainage | 504
identification of second tubular structure | 504
transection of second tubular structure | 504
identification of second extrahepatic bile duct | 504
anterior percutaneous catheter | 504
on-table cholangiogram | 504
fluoroscopy | 504
two separate extrahepatic biliary systems | 504
distal ducts ligation | 504
Roux limb | 504
anastomosis | 504
drain | 504
no evidence of bile leakage | 504
discharged | 510
normal hepatic function | 510
normal bilirubin | 510
no further complications | 510
follow-up cholangiogram | 672
normal intrahepatic ducts | 672
no evidence of stricture | 672
no evidence of leak | 672
successful repair | 672
cholangiogram catheters removal | 672
discharged from the clinic | 672