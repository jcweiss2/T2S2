52 years old | 0
female | 0
admitted to the emergency room | 0
abdominal pain | -120
nausea | -120
vomiting | -120
increased liver enzyme | -140
autoimmune antibody | -140
elevated immunoglobulin G | -140
chronic liver disease | -140
liver biopsy | -140
overlap syndrome | -140
ursodeoxycholic acid | -140
prednisolone | -140
mild heartburn | -168
abdominal pain | -168
mild fever | -168
tachycardia | -168
tachypnea | -168
abdominal tenderness | -168
elevated white blood cells | -168
elevated red blood cells | -168
elevated platelets | -168
elevated aspartate aminotransferase | -168
elevated alanine aminotransferase | -168
elevated gamma glutamyl transferase | -168
elevated C-reactive protein | -168
decreased neutrophil level | -168
contrast-enhanced abdominal CT | -168
necrotizing gastritis | -168
septic shock | -168
intravenous hydration | -168
antibiotic treatment | -168
systolic blood pressure decreased | -168
severe stress-induced cardiomyopathy | -168
extracorporeal membrane oxygenation | -168
cardiac arrest | -168
death | -168