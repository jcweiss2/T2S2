28 years old | 0
male | 0
history of peptic ulcer disease | 0
burning epigastric pain | -72
abdominal distention | -72
nausea | -72
vomiting | -72
bloody diarrhoea | -72
fevers | -72
blood pressure 90/60 | 0
heart rate 111 | 0
respiratory rate 34 | 0
oxygen saturation 91% on room air | 0
pale | 0
diaphoretic | 0
collapsing in triage | 0
weak pulses | 0
undetectable blood pressure | 0
respiratory rate 40 | 0
oxygen saturation 90% on ten litres of oxygen by face mask | 0
rigid abdomen | 0
distended abdomen | 0
absent bowel sounds | 0
decreased level of consciousness | 0
irregularly irregular wide complex tachycardia | 0
intravenous fluids bolused | 0
push dose of intravenous dextrose | 0
haemoglobin 15.8 g/dl | 0
haematocrit 50.1% | 0
white blood cell count 24 × 10³/mm³ | 0
segmented neutrophils 52.6% | 0
lymphocytes 17.4% | 0
platelets 175 × 10³/mm³ | 0
point-of-care echocardiogram | 0
large hyperechoic semisolid mobile mass within left ventricle | 0
abdominal ultrasound | 0
dilated loops of bowel | 0
thickened bowel | 0
absence of peristalsis | 0
echogenic foci in bowel wall suggesting pneumatosis intestinalis | 0
haemodynamic instability | 0
concern for mesenteric thromboembolism | 0
bowel ischaemia | 0
surgery consultation | 0
operating room mobilised | 0
exploratory laparotomy preparation | 0
antibiotics administration | 0
aggressive intravenous fluid resuscitation | 0
gangrenous necrosis of small bowel | 0
extension to cecum | 0
extension to ascending colon | 0
viable proximal jejunum | 0
viable transverse colon | 0
viable descending colon | 0
viable sigmoid colon | 0
normal pancreas | 0
palpable middle colic artery pulse | 0
absent distal superior mesenteric artery pulse | 0
evacuation of 600 mL haemorrhagic fluid from peritoneum | 0
lavage with warmed saline | 0
deferred bowel resection | 0
transfer to intensive care unit | 0
intubated | 0
broad spectrum antibiotics | 0
vasopressors | 0
overwhelming sepsis | 24
multi-organ failure | 24
cardiopulmonary arrest | 24
expired | 48
