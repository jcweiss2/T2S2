56 years old | 0
male | 0
admitted to the hospital | 0
end-stage renal disease | -8760
hemodialysis | -8760
coronary artery disease | -8760
type 2 diabetes mellitus | -8760
hypertension | -8760
chronic obstructive pulmonary disease | -8760
ischemic cardiomyopathy | -8760
hyperlipidemia | -8760
dyspnea | -144
coughing | -144
COVID-19 positive | 0
severe acute respiratory distress syndrome | 0
hypoxia | 0
oxygen saturation 85% | 0
required 3 liters of oxygen/min | 0
broad-spectrum antibiotics | -24
intubated | 0
tracheostomy | 600
vasopressor support | 0
heart rate 107/min | 0
blood pressure 140/50 mmHg | 0
oxygen saturation 94% | 0
fraction of inspired oxygen 90% | 0
positive end-expiratory pressure 14 cm H2O | 0
pupils round and reactive to light | 0
Glasgow coma scale 1T1 | 0
mild scleral icterus | 0
coarse breath sounds | 0
extensive anasarca | 0
elevated D-dimer | 0
inflammatory markers elevated | 0
procalcitonin level elevated | 0
thrombocytopenia | 0
normocytic anemia | 0
normal white cell counts | 0
lymphopenia | 0
chest X-ray showed multiple alveolar opacities | 0
COVID-19-induced pneumonia | 0
prothrombotic state | 0
ST elevations | 168
electrocardiogram consistent with inferior lead ST-segment elevations | 168
troponin I peaked at 5.5 ng/ml | 168
angiography findings showed a 40% proximal lesion in the right coronary artery | 168
percutaneous intervention with a drug-eluting stent | 168
thrombolysis in myocardial infarction flow 3 | 168
dual antiplatelet therapy | 168
tocilizumab | 168
failed extubation | 600
reintubation | 600
tracheostomy | 600
new unstageable decubitus ulcer | 600
discharged to a long-term care facility | 768
outpatient echocardiogram | 1056
followed up in an outpatient clinic | 1008
slightly improved physical strength | 1008
slightly improved nutritional status | 1008
no complications from the dual antiplatelet therapy | 1008