66 years old | 0
female | 0
recurrent fever | -672
history of Hashimoto’s disease | -672
history of pulmonary embolism | -672
admitted to the rheumatology department | 0
fever | -672
pneumonia | -672
urinary tract inflammation | -672
antibiotic therapy | -672
human immunodeficiency virus infection excluded | -672
hepatitis C virus infection excluded | -672
cytomegalovirus infection excluded | -672
toxoplasmosis excluded | -672
Lyme disease excluded | -672
tuberculosis excluded | -672
bone marrow biopsy | -672
no evidence of proliferative disease | -672
diagnosis of SLE confirmed | 0
methylprednisolone 80 mg/day initiated | 0
shortness of breath | 48
progressive decrease in blood pressure | 48
elevated procalcitonin serum concentration | 48
transferred to the Intensive Care Unit | 48
diagnosis of severe infection with risk of septic shock | 48
empirical antibiotic treatment | 48
glucocorticosteroid therapy | 48
atrial fibrillation | 48
amiodarone used | 48
improvement of general condition | 96
re-hospitalized in the rheumatology department | 96
GC therapy continued | 96
infusions of immunoglobulins | 96
flaccid four-limb weakness | 96
no abnormalities in brain imaging | 96
episode of unconsciousness | 120
left eye turning | 120
hypotension | 120
transthoracic echocardiography | 120
computed tomography of coronary arteries | 120
no significant deviations | 120
electroencephalography recording | 120
no irritation changes typical for epilepsy | 120
electromyography (EMG) | 120
features of generalized axonal damage of peripheral nerve motor fibers | 120
features of F wave disturbance | 120
limit values of conduction in sensory fibers | 120
recording from the muscles of the upper limbs and lower limbs | 120
features of depletion of exercise recording | 120
increased percentage of polyphasia | 120
critical illness polyneuropathy suspected | 120
follow-up EMG | 240
intensification of the lesions | 240
tendency to acute axonal polyneuropathy | 240
treatment with GCs continued | 240
methotrexate initiated | 240
hydroxychloroquine planned | 240
low molecular weight heparin | 240
transfer to the department of rehabilitation | 288
generalized weakness of trunk and limb muscle strength | 288
tetraparesis | 288
global paresis of the lower limbs | 288
abolition of tendon reflexes | 288
persistent lower limb allodynia | 288
treatment with pregabalin | 288
improvement rehabilitation program | 288
comprehensive improvement | 288
gradual verticalization | 288
increase of muscular strength | 288
isometric exercises | 288
learning to change position in the bed | 288
coordination exercises | 288
gradual improvement in muscle strength | 288
functional status | 288
change positions in bed independently | 432
cover a distance of several meters with a walker | 432
next cycle of rehabilitation | 504
gait improvement | 504
walk up the stairs | 504
technique of rising after a fall | 504
muscular strength and range of mobility of the left shoulder strengthened | 504
significant functional improvement | 504
discharge | 504
walk alone for short distances | 504
Barthel Index of Activities of Daily Living | 504