80 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
urinary tract infection | -120 | 0 | Possible
fever | -120 | 0 | Factual
dysuria | -120 | 0 | Factual
clean catch urine specimen | -120 | -120 | Factual
cephalexin | -120 | -96 | Factual
urine analysis | -120 | -120 | Factual
leukocyte esterase | -120 | -120 | Factual
bacteria | -120 | -120 | Factual
Escherichia coli | -120 | -120 | Factual
ampicillin resistance | -120 | -120 | Factual
levofloxacin resistance | -120 | -120 | Factual
trimethoprim resistance | -120 | -120 | Factual
sulfamethoxazole resistance | -120 | -120 | Factual
ampicillin/sulbactam sensitivity | -120 | -120 | Factual
cefazolin sensitivity | -120 | -120 | Factual
gentamicin sensitivity | -120 | -120 | Factual
nitrofurantoin sensitivity | -120 | -120 | Factual
cephalexin 500 mg | -96 | -48 | Factual
erythematous rash | -48 | 0 | Factual
sloughing of the skin | -24 | 0 | Factual
discontinued cephalexin | 0 | 0 | Factual
transferred to BICU | 0 | 0 | Factual
chronic obstructive pulmonary disease | 0 | 0 | Factual
type 2 diabetes mellitus | 0 | 0 | Factual
coronary artery disease | 0 | 0 | Factual
hypertension | 0 | 0 | Factual
hypothyroidism | 0 | 0 | Factual
depression | 0 | 0 | Factual
end-stage renal disease | 0 | 0 | Factual
hemodialysis | 0 | 0 | Factual
myocardial infarctions | 0 | 0 | Factual
ischemic cardiomyopathy | 0 | 0 | Factual
atrial fibrillation | 0 | 0 | Factual
hydrocodone/acetaminophen | 0 | 0 | Factual
levothyroxine | 0 | 0 | Factual
escitalopram | 0 | 0 | Factual
carvedilol | 0 | 0 | Factual
guaifenesin | 0 | 0 | Factual
docusate | 0 | 0 | Factual
calcitriol | 0 | 0 | Factual
albuterol | 0 | 0 | Factual
amiodarone | 0 | 0 | Factual
pulmonary infiltrates | 24 | 24 | Factual
respiratory failure | 24 | 24 | Factual
intubated | 24 | 24 | Factual
difficulty swallowing | 24 | 24 | Factual
endotracheal tube | 24 | 24 | Factual
toxic epidermal necrolysis syndrome | 0 | 0 | Factual
body surface area skin detachment | 0 | 0 | Factual
blood pressure | 0 | 0 | Factual
respiratory rate | 0 | 0 | Factual
temperature | 0 | 0 | Factual
white blood cell count | 0 | 0 | Factual
neutrophils | 0 | 0 | Factual
platelet count | 0 | 0 | Factual
serum creatinine | 0 | 0 | Factual
venous serum lactate | 0 | 0 | Factual
oxygen saturation | 0 | 0 | Factual
pain | 0 | 0 | Factual
peripheral blood cultures | 0 | 0 | Factual
skin surveillance cultures | 0 | 0 | Factual
urine culture | 0 | 0 | Factual
chest radiograph | 0 | 0 | Factual
right pleural effusion | 0 | 0 | Factual
right lower and left basilar opacities | 0 | 0 | Factual
norepinephrine | 0 | 0 | Factual
vasopressin | 0 | 0 | Factual
albumin | 0 | 0 | Factual
lactated Ringer’s | 0 | 0 | Factual
tetanus–diphtheria toxoids vaccine | 0 | 0 | Factual
gentamicin | 0 | 0 | Factual
fluconazole | 0 | 0 | Factual
WBC | 24 | 24 | Factual
SCr | 24 | 24 | Factual
venous serum lactate | 24 | 24 | Factual
random serum gentamicin level | 24 | 24 | Factual
gentamicin | 24 | 24 | Factual
fluconazole | 24 | 24 | Factual
supportive continuous renal replacement therapy | 24 | 24 | Factual
wide complex tachycardia | 96 | 96 | Factual
amiodarone | 96 | 96 | Factual
gentamicin | 96 | 96 | Factual
physical examination | 120 | 120 | Factual
sloughing of skin | 120 | 120 | Factual
culture and sensitivity results | 120 | 120 | Factual
Pseudomonas aeruginosa | 120 | 120 | Factual
gentamicin | 120 | 120 | Factual
expired | 144 | 144 | Factual
cardiac arrest | 144 | 144 | Factual
multisystem organ failure | 144 | 144 | Factual
autopsy | 144 | 144 | Factual
necrotizing bronchopneumonia | 144 | 144 | Factual
TEN | 144 | 144 | Factual
SCORTEN | 144 | 144 | Factual
predicted mortality | 144 | 144 | Factual