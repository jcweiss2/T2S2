56 years old | 0
male | 0
end-stage renal disease | -12768
hemodialysis (3 d/week) | -12768
coronary artery disease | -12768
type 2 diabetes mellitus | -12768
hypertension | -12768
chronic obstructive pulmonary disease | -12768
ischemic cardiomyopathy | -12768
hyperlipidemia | -12768
dyspnea | -144
coughing | -144
significant contact history for COVID-19 | -144
COVID-19-positive | 0
transferred due to worsening dyspnea | -144
hypoxia during hemodialysis | -144
oxygen saturation not improving | -144
intubated for 25 days before tracheostomy | -144
hypoxic with 85% oxygen saturation | 0
required 3 liters of oxygen/min | 0
received broad-spectrum antibiotics | -144
differential diagnosis of COVID-19 pneumonia | 0
differential diagnosis of acute bacterial pneumonia | 0
vasopressor support | 0
heart rate of 107/min | 0
blood pressure of 140/50 mmHg | 0
oxygen saturation of 94% | 0
fraction of inspired oxygen 90% | 0
positive end-expiratory pressure of 14 cm H2O | 0
pupils round and reactive to light | 0
Glasgow coma scale of 1T1 due to sedation | 0
mild scleral icterus | 0
coarse breath sounds | 0
extensive anasarca | 0
elevated D-dimer | 0
increased erythrocyte sedimentation rate | 0
increased ferritin | 0
increased C-reactive protein | 0
procalcitonin level falsely elevated | 0
thrombocytopenia | 0
normocytic anemia | 0
normal white cell counts | 0
lymphopenia | 0
chest X-ray showing multifocal pneumonia | 0
cultures negative | 0
diagnosis of COVID-19-induced pneumonia | 0
diagnosis of prothrombotic state | 0
started on broad-spectrum antibiotics | 0
prone positioning for severe ARDS | 0
ST elevations noted on telemetry | 168
electrocardiogram consistent with inferior lead ST-segment elevations | 168
troponin I peaked at 5.5 ng/ml | 168
angiography showing 40% proximal lesion in right coronary artery | 168
angiography showing 99% distal lesion in posterior descending artery | 168
thrombus localized in posterior descending artery | 168
catheterization showing mean aortic pressure of 80 mmHg | 168
catheterization showing left ventricular end-diastolic pressure of 18 mmHg | 168
percutaneous intervention with drug-eluting stent | 168
thrombolysis in myocardial infarction flow 3 | 168
started on dual antiplatelet therapy (clopidogrel and aspirin) | 168
started on tocilizumab | 168
failed extubation | 168
reintubation | 168
tracheostomy | 168
new unstageable decubitus ulcer | 168
managed conservatively for decubitus ulcer | 168
discharged after 32 days | 768
outpatient echocardiogram planned | 768
outpatient follow-up after 2 weeks | 1344
slightly improved physical strength | 1344
improved nutritional status | 1344
no complications from dual antiplatelet therapy | 1344
