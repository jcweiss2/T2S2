52 years old | 0
female | 0
Indian | 0
admitted to hospital | 0
one-week history of right-sided retro-orbital pain | -168
right-sided facial swelling | -168
no significant past medical history | 0
apyrexial | 0
pulse rate of 100 min–1 | 0
confused | 0
right-sided periorbital cellulitis | 0
decreased visual acuity in the right eye | 0
full range of extraocular muscle movements | 0
ipsilateral mild facial nerve weakness | 0
neutrophilic leukocytosis | 0
C-reactive protein of 456 mg/L | 0
random blood glucose of 56.1 mmol/L | 0
presence of ketones | 0
metabolic acidosis | 0
diabetic ketoacidosis | 0
treated with intravenous fluid replacement | 0
treated with intravenous antibiotics | 0
commenced on an insulin sliding scale | 0
CT head including both orbits | 0
right periorbital cellulitis | 0
stranding of the extraconal adipose tissue | 0
Chandler classification grade II | 0
no evidence of intra-orbital collection | 0
no evidence of intracranial extension | 0
complete opacification of the right nasal cavity | 0
complete opacification of the maxillary and frontal sinuses | 0
urgent endoscopic exploration | 12
necrotic mass in the right nasal cavity | 12
biopsies sent for histopathology | 12
histopathological assessment revealed fungal invasion | 24
fungal hyphae were seen to be broad and distorted | 24
branching at right angles | 24
surrounded by extensive necrotic debris | 24
no septae were present | 24
right nasal cavity and paranasal sinuses exenterated | 24
irrigated | 24
parenteral amphotericin B added to treatment | 24
initial transient improvement | 24
temperature improved | 24
conscious level improved | 24
cranial neuropathies persisted | 48
deteriorated | 48
becoming more confused | 48
losing vision completely from the right eye | 48
MRI scan of the head | 72
evidence of predominantly right frontal cerebritis | 72
early abscess formation | 72
re-accumulation of fluid | 72
thickening of the mucosa in the paranasal sinuses | 72
disease affecting the sphenoid and ethmoid sinuses | 72
further surgery | 96
right maxillectomy | 96
orbital exenteration | 96
frontal sinus opened | 96
mass extending into the dura | 96
dura opened | 96
necrotic cerebral parenchyma removed | 96
repeated irrigation | 96
transferred to ICU | 120
failed to recover | 120
died | 144
generalized seizure | 144