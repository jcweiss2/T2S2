53 years old | 0
    African American female | 0
    hypertension | -43200
    diabetes mellitus type 2 | -43200
    presented to the emergency department | 0
    altered mental status | 0
    feeling unwell | -72
    symptoms progressed | -72
    altered mentation | 0
    dyspnea | 0
    temperature 36.6 °C | 0
    heart rate 112 beats per minute | 0
    blood pressure 140/72 mm Hg | 0
    respiratory rate 28 breaths per minute | 0
    oxygen saturation 96% | 0
    confused | 0
    agitated | 0
    tachypneic | 0
    tachycardic | 0
    leukocytosis | 0
    white blood cell count 19.9 × 10^9/L | 0
    absolute neutrophils 89.3% | 0
    platelet count 507 × 10^9/L | 0
    sodium 131 mmol/L | 0
    potassium 6.2 mmol/L | 0
    chloride 104 mmol/L | 0
    total CO2 6 | 0
    glucose >38.8 mmol/L | 0
    BUN 25 mmol/L | 0
    creatinine 362.5 µmol/L | 0
    high anion gap 28 | 0
    acetone large | 0
    high anion gap metabolic acidosis | 0
    compensatory respiratory alkalosis | 0
    CT head unremarkable | 0
    intravenous fluids | 0
    insulin infusion | 0
    transferred to intensive care unit | 0
    DKA resolved | 72
    altered mentation improved | 72
    renal function progressively worsened | 72
    BUN trend up | 72
    serum creatinine trend up | 72
    oliguric | 72
    Udall catheter placed | 72
    creatinine 88 µmol/L | -1440
    BUN 3.6 mmol/L | -1440
    febrile | 96
    Tmax 39.1 °C | 96
    tachycardic | 96
    hemodynamically stable | 96
    septic workup performed | 96
    empiric broad-spectrum antibiotics | 96
    antipyretics | 96
    blood cultures grew K pneumoniae | 96
    CT abdomen and pelvis with oral contrast | 96
    hypoattenuating hepatic lesions | 96
    heterogeneous splenic hyperattenuation | 96
    splenic infarcts | 96
    MRI abdomen and pelvis | 96
    8 lesions in left hepatic lobe | 96
    largest lesion 3.9 × 3.2 × 3.7 cm | 96
    hepatic abscess | 96
    ill-defined splenic lesions | 96
    splenic abscesses | 96
    piperacillin/tazobactam de-escalated | 96
    ceftriaxone | 96
    metronidazole | 96
    percutaneous drainage of hepatic abscess | 96
    30 mL pus | 96
    K pneumoniae | 96
    repeat blood cultures negative | 168
    renal function stabilized | 168
    dialysis discontinued | 168
    repeat CT abdomen and pelvis | 168
    worsening splenic lesions | 168
    perisplenic fluid | 168
    percutaneous drainage of splenic abscesses | 168
    acute right femoral deep vein thrombosis | 168
    popliteal deep vein thrombosis | 168
    peroneal vein deep vein thrombosis | 168
    high-range heparin infusion | 168
    heparin discontinued | 192
    steep decline in hemoglobin | 192
    inferior vena cava filter inserted | 192
    colonoscopy | 192
    15-mm polyp in cecum | 192
    nonbleeding hemorrhoids | 192
    hemoglobin stabilized | 192
    blood transfusions | 192
    clinically improved | 192
    6-week course of antibiotics | 240
    discharged | 240
    follow-up outpatient | 240
    nephrology | 240
    infectious disease | 240
    primary care physician | 240
    