48 years old | 0
male | 0
peasant crop farmer | 0
admitted to the hospital | 0
generalised abdominal pains | -48
fever | -48
passing scanty urine | -48
painful irreducible right groin swelling | -120
absolute constipation | -120
vomiting | -120
reducible right groin swelling | -5280
occasional episodes of irreducibility | -5280
ill-looking patient | 0
pale | 0
jaundiced | 0
dehydrated | 0
febrile | 0
respiratory rate 25 breaths/min | 0
pulse rate 108 beats/min | 0
blood pressure 98/55 mmHg | 0
globally distended abdomen | 0
tense abdomen | 0
peritonism | 0
irreducible right inguinoscrotal swelling | 0
septic shock | 0
resuscitation | 0
intravenous fluid | 0
intravenous ciprofloxacin | 0
metronidazole | 0
intranasal oxygen | 0
adrenaline | 0
transfused 2 pints of blood | 0
nasogastric tube | 0
urethral catheter | 0
urine output >0.6 ml/kg/hour | 0
SPO2 -94% | 0
blood pressure 115/70 mmHg | 0
pulse rate 86 bpm | 0
respiratory rate 22 cycles | 0
Full Blood Count | 0
haemoglobin 7.4 g/dL | 0
leucocytosis | 0
differential neutrophilia | 0
decreased platelets level | 0
blood urea 11.2 mmol/L | 0
creatinine 162 μmol/L | 0
retroviral tested positive | 0
random blood sugar 6.1 mmol/L | 0
American Society of Anesthesiology score III | 0
counseled for surgery | 0
informed consent | 0
surgery | 0
extended midline incision | 0
free fluid with faecal matter | 0
herbal residue | 0
extensive exudate | 0
gangrenous perforated caecum | 0
mattered small bowel | 0
hernia sac contained redundant large bowel | 0
right hemicolectomy | 0
herniotomy | 0
nylon darn repair | 0
abdominal drain inserted | 0
Peritoneum lavage | 0
post-operative care | 0
transfused another pint of blood | 0
intravenous antibiotics | 0
intravenous fluids | 0
analgesia | 0
intravenous KCL | 0
intravenous omeprazole | 0
nil per oral route | 0
graded oral intake | 72
oral medications | 72
weight loss | 0
intravenous combine vitamins | 0
local formulated high carbohydrate diet | 0
wound care | 0
wound exposed | 48
cleaned with savlon | 48
normal saline | 48
dressed with povidone-soaked gauze | 48
discharging serosanguinous fluid | 72
draining offensive pus | 72
massive scrotal collection | 72
copious exudate | 72
cleaned twice daily | 72
irrigated with normal saline | 72
cavity packed with povidone-iodine-soaked gauze | 72
discharge subsided | 336
daily dressing | 336
granulation over nylon darn sutures | 360
secondary suturing | 432
discharged | 576
parts of abdominal wound healed | 576
wound dressing at primary facility | 576
methylated spirit | 576
further investigations | 576
treatment at Anti-Retroviral Clinic | 576
doing very well | 4380
no evidence of hernia recurrence | 4380