30 years old | 0
multigravida | 0
g3p2 | 0
repeated cesarean section | 0
32-weeks pregnant | 0
admitted to the hospital | 0
chills | -144
cough | -144
shortness of breath | -144
respiratory rate 26/min | 0
blood pressure 110/75 mm Hg | 0
oxygen-free saturation 84% | 0
body temperature 38.8 °C | 0
no uterine activity | 0
lymphopenia | 0
elevated liver enzymes | 0
low platelets | 0
increased Prothrombin Time (PT/INR) | 0
increased activated Partial Thromboplastin Time (aPTT) | 0
high D-dimer | 0
high total bilirubin | 0
high LDH | 0
normal hemoglobin | 0
normal kidney function tests | 0
COVID-19 diagnosis | 0
sepsis diagnosis | 0
HELLP syndrome diagnosis | 0
admitted to the 3rd level intensive care unit | 0
bilateral diffuse ground glass areas | 24
diffuse peripheral interstitial thickening | 24
bilateral mild pleural effusion | 24
viral pneumonia (COVID-19) | 24
positive COVID-19 PCR test | 24
hepatitis markers negative | 24
HIV test negative | 24
no growth in blood and urine cultures | 24
normal serum electrolytes | 24
normal cardiac markers | 24
Anti-Covid treatment started | 24
hypertensive | 48
oxygen-free saturation dropped below 80% | 48
change in consciousness level | 48
intubated | 48
antihypertensive treatment started | 48
magnesium sulfate started | 48
obstetrician consulted | 48
termination of pregnancy considered | 48
hemodynamic stabilization | 48
cesarean section performed | 72
singleton live baby boy delivered | 72
Apgar scores of two and six | 72
newborn intubated | 72
newborn chest X-ray normal | 72
newborn COVID-19 positive | 72
pancytopenia developed | 96
renal failure developed | 96
newborn died | 120
fluid resuscitation | 0
electrolyte resuscitation | 0
blood and blood products resuscitation | 0
antihypertensive treatment | 0
magnesium sulfate | 0
antibiotherapy | 0
hemodialysis | 0
brain MRI examination | 216
normal brain MRI findings | 216
extubation attempts unsuccessful | 240
mother patient died | 240