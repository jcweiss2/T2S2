14 years | 0
male | 0
fever | -96
abdominal pain | -72
cough | -24
chills | -96
sweating | -96
no rigors | -96
no recent travel | -96
no known sick contacts | -96
no medications for chronic illness | -96
no known allergies | -96
thinly built | 0
weight <3rd centile | 0
febrile | 0
tachypneic | 0
hypotension | 0
oxygen saturation maintained with 2L O2 per minute | 0
enlarged right inguinal lymph nodes | 0
non-tender lymph nodes | 0
abdomen soft and distended | 0
liver palpable 3 cm below the right subcostal margin | 0
liver span 12 cm | 0
fluid thrill present | 0
no splenomegaly | 0
decreased air entry on the right mammary area | 0
neutrophilia | 0
lymphopenia | 0
thrombocytopenia | 0
deranged liver function test | 0
elevated liver enzymes | 0
low serum albumin | 0
normal renal function test | 0
arterial blood gas analysis showed pH:7.43 | 0
Pco2- 27 | 0
Po2-135 | 0
HCO3-20 | 0
significant number of pus cells in urine | 0
no growth in urine culture | 0
tested negative for scrub typhus | 0
subtle diffuse coalescent opacities in bilateral lungs | 0
decrease in 4–7th intercostal space on the left side | 0
gross ascites | 0
minimal pleural effusion | 0
minimal pericardial effusion | 0
mild tricuspid regurgitation | 0
mild mitral regurgitation | 0
elevated white blood cell count with lymphocytosis in ascitic fluid | 0
high ADA in ascitic fluid | 0
no growth in ascitic fluid culture | 0
normal peripheral blood smear | 0
negative troponin marker | 0
CK-MB value 18IU/L | 0
admitted to pediatric ICU | 0
treated with intravenous antibiotics | 0
treated with intravenous fluids | 0
treated with vasopressors | 0
administered albumin | 0
CT scan of bilateral lung fields | 24
CT scan showed subpleural reticular opacities | 24
CT scan showed ground glass opacity | 24
abdominal CT scan showed grossly normal findings | 24
abdominal CT scan showed mild hepatomegaly | 24
tested positive for Covid-antibody | 24
treated with intravenous immunoglobulin | 24
treated with high dose of methylprednisolone | 24
diuretics added | 48
low molecular weight heparin added | 48
kept on BIPAP | 48
intravenous antibiotics upgraded | 96
troponin marker tested positive | 120
CK-MB value 26 IU/L | 120
condition improved | 120
inotropes tapered | 120
oxygen weaned off | 120
low molecular heparin stopped | 192
intravenous diuretics stopped | 192
oral rivaroxaban started | 192
oral diuretics started | 192
feeding initiated | 192
afebrile | 192
oxygen saturation maintained with oxygen at 3 L per minute | 192
shifted to pediatric ward | 312
oxygen saturation maintained in room air | 312
repeat echocardiography showed dilated and fixed IVC | 312
repeat echocardiography showed dilated left ventricle | 312
repeat echocardiography showed no diastolic dysfunction | 312
repeat echocardiography showed minimal pericardial effusion | 312
repeat echocardiography showed coronary artery diameter - 3mm | 312
repeat echocardiography showed ejection fraction of 65% | 312
repeat complete blood panel showed improvement in platelet count | 312
discharged | 336
oral antibiotics | 336
steroids | 336
anticoagulants | 336
diuretics | 336
multivitamins | 336
followed up in pediatric OPD | 504
doing fine | 504
chest x-ray normal | 672