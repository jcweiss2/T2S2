27 years old | 0
male | 0
presented to the emergency department | 0
fevers | -120
chills | -120
intermittent epigastric pain | -120
epigastric pain started acutely | -120
burning pain | -120
non-radiating pain | -120
pain lasted 20 minutes | -120
pain recurred several times | -120
subjective fevers | -48
chills (subjective) | -48
vomiting | -48
denied diarrhea | 0
denied sick contacts | 0
denied recent travel | 0
denied dysuria | 0
denied hematuria | 0
denied chest pain | 0
denied shortness of breath | 0
tachycardic | 0
afebrile | 0
normotensive | 0
diaphoretic | 0
jaundiced skin | 0
icteric sclera | 0
clear lungs | 0
negative cardiac exam | 0
normal extremities | 0
no edema | 0
no rash | 0
epigastric tenderness | 0
soft abdomen | 0
non-distended abdomen | 0
no rebound tenderness | 0
no involuntary guarding | 0
no Rovsing’s sign | 0
no Obturator sign | 0
no Murphy’s sign | 0
non-tender abdomen | 0
leukocytosis | 0
toxic granulations | 0
neutrophilic predominance | 0
thrombocytopenia | 0
elevated D-dimer | 0
elevated fibrinogen | 0
elevated total bilirubin | 0
elevated alkaline phosphatase | 0
normal chest radiograph | 0
normal electrocardiogram | 0
treated for severe sepsis | 0
treated for septic shock | 0
received normal saline boluses | 0
received broad-spectrum antibiotics | 0
responded to interventions | 0
normalized vital signs | 0
reported feeling better | 0
ordered abdominal ultrasound | 0
normal liver | 0
no ductal dilatation | 0
normal kidneys | 0
normal aorta | 0
normal spleen | 0
normal pancreas | 0
no gallbladder stones | 0
no gallbladder sludge | 0
thickened gallbladder wall | 0
no peri-cholecystic fluid | 0
surgical consult for cholecystitis/cholangitis | 0
no tenderness on surgical exam | 0
no distension on surgical exam | 0
abnormal lab findings | 0
gallbladder wall thickening | 0
possible atypical cholecystitis | 0
recommended CT abdomen/pelvis | 0
admitted to ICU | 0
continued antibiotic therapy | 0
standard infectious workup | 0
tested for influenza | 0
tested for viral hepatitis | 0
tested for HIV | 0
tested for malaria | 0
tested for tularemia | 0
blood cultures grew E. coli | 48
tailored antibiotics | 48
CT abdomen/pelvis obtained | 72
dilated retrocecal appendix | 72
thick-walled appendix | 72
adjacent inflammation | 72
free fluid | 72
acute appendicitis | 72
inflamed gallbladder wall | 72
secondary to appendicitis | 72
final CT confirmed appendicitis | 96
pylephlebitis | 96
laproscopic appendectomy | 96
procedure without complications | 96
continued IV antibiotics | 96
discharged | 144
no mention of pylephlebitis | 0
antibiotics discontinued | 144
elevated WBC count at discharge | 144
elevated total bilirubin at discharge | 144
follow-up in surgery clinic | 168
minimal pain | 168
able to eat and drink | 168
staples removed | 168
lost to follow-up | 168
Final Answer<|eot_id|>
negative cardiac exam |0
