38 years old | 0
male | 0
asthma | 0
acute onset fever | -144
chills | -144
cough | -144
bronchitis | -144
symptoms persisted | -144
left upper quadrant abdominal pain | -72
pain radiating to left shoulder | -72
severe hypotension | -72
malaria blood slide positive | -72
ultrasound showing fluid in abdomen | -72
artesunate administration | -72
referral for surgical review | -72
referral for infectious disease specialist review | -72
sick-looking appearance | 0
mild pallor | 0
jaundice | 0
tachycardia (122 bpm) | 0
normal blood pressure (121/59 mmHg) | 0
slightly distended abdomen | 0
mild generalized tenderness | 0
no acute peritonitis | 0
low hemoglobin (9.3 g/dl) | 0
normal red cell indices | 0
repeat malaria blood slide positive (4% parasitemia, P. falciparum) | 0
parenteral artemether administration | 0
oral doxycycline administration | 0
CT scan abdomen with IV contrast | 0
free peritoneal fluid | 0
no obvious splenic rupture | 0
no contrast extravasation | 0
monitored in ICU | 0
hemoglobin fell from 9.3 to 7.4 g/dl | 16
ongoing resuscitation with two pints whole blood | 16
normal vital signs | 16
worsening abdominal distension | 16
worsening abdominal pain | 16
exploratory laparotomy | 16
finding 2 liters frank blood | 16
enlarged spleen | 16
firm spleen | 16
circumferential upper pole laceration | 16
active bleeding after spleen mobilization | 16
splenectomy performed | 16
postoperative recovery without complications | 24
discharged home after 8 days | 192
fully recovered | 192
advised malaria prophylaxis with atovaquone/proguanil | 192
splenic rupture due to complicated P. falciparum malaria | 0
hypotension history | -72
positive Kehr's sign | -72
negative CT scan for splenic rupture | 0
tamponaded laceration | 16
ongoing splenic bleeding | 16
unsuccessful conservative management | 16
splenectomy necessitated | 16
histopathology showing enlarged spleen | 16
no trauma history | 0
no perisplenic adhesions | 0
no other spleen disease | 0
met Orloff and Peskins criteria for spontaneous splenic rupture | 16
intravenous fluids administration | 16
blood product use | 16
deterioration despite conservative management | 16
