53 years old | 0
    male | 0
    visited the emergency room | 0
    productive cough | -24
    fever | -24
    chills | -24
    30-pack/year history of cigarette smoking | 0
    consumed alcohol in moderation | 0
    treated for community-acquired pneumonia 2 years prior | -17520
    acutely ill appearance | 0
    blood pressure 82/46 mmHg | 0
    respiratory rate 22 breaths per minute | 0
    pulse rate 120 beats per minute | 0
    body temperature 40℃ | 0
    regular heart rhythm | 0
    coarse breathing sounds | 0
    crackles on the right lower lung field | 0
    white blood cell count 11,500/mm3 | 0
    neutrophils 86.1% | 0
    lymphocytes 11.5% | 0
    monocytes 1.9% | 0
    eosinophils 0.2% | 0
    hemoglobin 14.4 g/dL | 0
    platelet count 188,000/mm3 | 0
    C-reactive protein 1.28 mg/dL | 0
    pH 7.47 | 0
    pCO2 22.4 mmHg | 0
    pO2 52.5 mmHg | 0
    HCO3- 16 mmol/L | 0
    O2 saturation 89% | 0
    BUN/Cr 9/2.05 mg/dL | 0
    serum sodium 139 mmol/L | 0
    serum potassium 4.1 mmol/L | 0
    serum chloride 105 mmol/L | 0
    urine sodium 19 mmol/L | 0
    urine Cr 222.31 mg/dL | 0
    fractional excretion of sodium 0.1% | 0
    moderate patchy consolidation in the right lower lobe | 0
    presumptive diagnosis of sepsis caused by community-acquired pneumonia | 0
    septic shock | 0
    central line catheter insertion | 0
    fluid resuscitation | 0
    oxygen administered via nasal cannula | 0
    blood culture | 0
    sputum culture | 0
    urine culture | 0
    empiric piperacillin/tazobactam | 0
    ciprofloxacin injection | 0
    admission to intensive care unit | 0
    APACHE II score 25 | 0
    low blood pressure persisted | 0
    norepinephrine administration | 0
    vasopressin administration | 0
    respiratory distress worsened | 16
    acute respiratory failure | 16
    arterial blood gas analysis pH 7.085 | 16
    arterial blood gas analysis pCO2 61.4 mmHg | 16
    arterial blood gas analysis HCO3C 19 mmol/L | 16
    intubation | 16
    mechanical ventilation FiO2 1.0 | 16
    positive end expiratory pressure 14 cmH2O | 16
    hypoxia persisted | 16
    respiratory acidosis deteriorated | 16
    metabolic acidosis deteriorated | 16
    follow-up arterial blood gas analysis pH 7.096 | 24
    follow-up arterial blood gas analysis pCO2 63.7 mmHg | 24
    follow-up arterial blood gas analysis pO2 77.6 mmHg | 24
    follow-up arterial blood gas analysis HCO3C 20 mmol/L | 24
    follow-up arterial blood gas analysis O2 saturation 89% | 24
    exacerbated consolidation in the right lung field | 24
    patchy opacities in the left lower lobe | 24
    antibiotics switched to meropenem | 24
    antibiotics switched to teicoplanin | 24
    oliguria | 28
    acute kidney injury deteriorated | 28
    BUN/Cr 26/3.66 mg/dL | 28
    continuous renal replacement therapy | 28
    septic shock persisted | 36
    acute respiratory failure persisted | 36
    cardiac arrest | 36
    cardiopulmonary resuscitation | 36
    patient expired | 36
    Acinetobacter baumannii identified in sputum culture | 36
    Acinetobacter baumannii identified in blood cultures | 36
    bacterial susceptibility to piperacillin/tazobactam | 36
    bacterial susceptibility to ceftazidime | 36
    bacterial susceptibility to cefepime | 36
    bacterial susceptibility to imipenem | 36
    bacterial susceptibility to meropenem | 36
    bacterial susceptibility to gentamicin | 36
    bacterial susceptibility to tobramycin | 36
    bacterial tolerance to ampicillin | 36
    bacterial tolerance to amoxacillin/clavulanic acid | 36
    bacterial tolerance to cafalotin | 36
    bacterial tolerance to cefoxitin | 36
    bacterial tolerance to trimethoprim/sulfamethoxazole | 36
    bacterial moderate tolerance to cefotaxime | 36
    bacterial moderate tolerance to levofloxacin | 36