60 years old | 0
male | 0
dysphagia | -672
barium swallow study | 0
aspiration of barium | 0
dyspneic | 0
labored breathing | 0
respiratory rate >35 breaths/min | 0
tachycardia | 0
heart rate >120 beat/min | 0
blood pressure 160/100 mmHg | 0
SPO2 <90% | 0
oxygen flow 15lit/min by mask | 0
hypoxemia | 0
PO2 86.7 mmHg on oxygen flow 15 lit/min | 0
crepitation in both lung bases | 0
barium sulfate aspiration | 0
intubation | 0
positive pressure mechanical ventilation | 0
early bronchioalveolar lavage | 0
postural drainage techniques | 0
shock | 4
fluid resuscitation | 4
inotropic support | 4
infusion noradrenaline | 4
injection hydrocortisone 100 mg | 4
broad-spectrum antibiotics | 4
nebulization with N-acetylcystein | 4
stable hemodynamically | 24
extubation | 24
oxygen saturation of 99% on 5 litres of oxygen | 24
shifted to ward | 72
aspiration of oral feed and gastric contents | 144
shifted to ICU | 144
sepsis | 336
death | 336