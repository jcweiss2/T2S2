63 years old | 0
male | 0
smoking (20 packs/year) | -72
DVT in left leg | -72
rivaroxaban anticoagulant therapy | -72
hospitalized | -72
abrupt onset of dyspnea | -72
thoracic CT scan | -72
pulmonary thromboembolism (PTE) | -72
mass in lower lobe of right lung | -72
ipsilateral ilo?mediastinal lymph nodes | -72
infra-clavear pathological lymph nodes | -72
abdominal CT scan | -72
splenic infarctions | -72
renal infarctions | -72
right cerebellar signs | -72
confusion | -72
nystagmus | -72
ataxia | -72
dysmetria | -72
adiadochokinesia | -72
MRI of brain | -72
multiple diffuse bi-hemispheric cerebral areas | -72
cerebellar areas | -72
grey matter hyperintense | -72
occipital lobes | -72
deep cerebral white matter hyperintense | -72
diffusion restriction | -72
moderate patchy enhancement | -72
gyriform enhancement | -72
TTE | -72
TEE | -72
spontaneous rapid improvement | -72
complete resolution of confusion | -72
cerebellar symptoms resolved | -72
cardio embolic origin suspected | -72
PFO detected | -72
LMWH prescribed | -72
PET scan | -24
locally advanced disease (IIIB stage) | -24
EBUS-guided transbronchial needle aspiration | -24
large-cell carcinoma diagnosed | -24
immunohistochemistry positive for cytokeratin pool | -24
TTF-1 negative | -24
p40 negative | -24
chromogranin A negative | -24
synaptophysin negative | -24
CAM5.2 positive | -24
EGFR mutations absent | -24
ALK rearrangements absent | -24
PD-L1 55% | -24
candidate for pembrolizumab | -24
novel hospitalization | -24
diplopia | -24
gait impairment | -24
CT scan | -24
evolution of lesion | -24
substernal chest pain | -24
dyspnea | -24
regular body temperature | -24
regular blood pressure | -24
regular heart rate | -24
diastolic murmur | -24
aortic regurgitation | -24
sinus tachycardia | -24
ST segment elevation | -24
elevated serum troponin I | -24
reduced LVEF 45% | -24
mobile mass on mitral valve | -24
moderate aortic insufficiency | -24
acute pulmonary edema | -24
respiratory failure | -24
noninvasive ventilation | -24
coronary angiography | -24
reduced flow TIMI 2 | -24
embolus | -24
hemodynamic instability | -24
respiratory instability | -24
admitted to ICU | -24
aspirin therapy | -24
β-blockers therapy | -24
LMWH continued | -24
infective endocarditis suspected | -24
blood culture tests | -24
empiric antibiotic therapy | -24
linezolid | -24
daptomycin | -24
piperacillin/tazobactam | -24
petechiae on lower limbs | -24
peripheral embolization | -24
abdominal CT scan | -24
abdominal pain | -24
loss of blood in stool | -24
occlusion of superior mesenteric artery | -24
ileal loop thinning | -24
emergency ileo-cecal resection | -24
bowel infarction | -24
intubated | -24
TEE | -24
echogenic mass on mitral valve | -24
aortic insufficiency | -24
LVEF 40% | -24
negative blood cultures | -24
normal inflammatory markers | -24
NBTE diagnosed | -24
coma | 24
increased brain infarcts | 24
novel cerebral foci | 24
multi-organ failure | 24
passed away | 24
