35 years old | 0
female | 0
chronic pancreatitis | 0
alcoholic liver disease | 0
alcohol abuse | 0
admitted to the emergency department | 0
diffuse abdominal pain | -72
abdominal pain radiating to the thorax | -72
admitted | -168
discharged | -168
acute chronic pancreatitis | -168
pancreatic pseudocyst | -168
necrosis | -168
current smoker | 0
16-pack year history | 0
consuming 1 to 2 glasses of alcohol daily | 0
abstinent from alcohol ingestion | 0
denied illicit drug use | 0
blood pressure 91/55 | 0
pulse 114 bpm | 0
respiratory rate 18 | 0
temperature 98.1°F | 0
oxygen saturation 99% | 0
abdomen distended | 0
diffusely tender to palpation | 0
positive fluid wave | 0
voluntary guarding | 0
leukocytosis | 0
WBC 16.9 | 0
hemoglobin 10.3 | 0
sodium 130 | 0
lipase 149 | 0
liver function tests within normal limits | 0
CT abdomen and pelvis with contrast | 0
significant increase in ascites | 0
multiple pancreatic cysts | 0
10 mm fluid density lesion at the neck of the pancreas | 0
enlarged peripancreatic fluid | 0
paracentesis | 0
ascitic fluid removed | 0
WBC 8423 | 0
RBC 1570 | 0
PMN 82% | 0
protein 3.2 | 0
amylase 5507 | 0
LDH 478 | 0
SAAG 0.1 | 0
ERCP | 0
plastic stent placed | 0
clinical condition deteriorated | 0
transferred to ICU | 0
acute respiratory distress syndrome | 0
ABG pH 7.36 | 0
ABG PCO2 30 | 0
ABG PO2 50 | 0
ABG HCO3 18.8 | 0
100% FiO2 | 0
non-rebreathing mask | 0
vasopressor support | 0
MAP 65 | 0
septic shock | 0
leukocytosis 16.9 to 69.2K/µL | 0
ascitic fluid culture | 0
blood culture | 0
urine culture | 0
ET tube culture | 0
no microbial growth | 0
ceftriaxone 2000 mg | 0
SBP treatment | 0
switched to IV meropenem | 0
IV meropenem 1000 mg every 8 hours | 0
serial CT abdomen with contrast | 0
no postprocedure worsening of pancreatitis | 0
intubated | 0
acute respiratory failure | 0
tracheostomy | 0
PEG feeding tube inserted | 0
paracentesis procedures | 0
4 L ascitic fluid removed | 0
3 L ascitic fluid removed | 0
2 L ascitic fluid removed | 0
Jackson-Pratt drains placed | 0
CT abdomen | 0
pancreatic pseudocyst increased size 2.7 to 5.8 cm | 0
loculated mesenteric collections | 0
concern for serosal implants | 0
surgical consultation | 0
surgical intervention not advised | 0
hyperdense material in pseudocyst | 0
consistent decline in hemoglobin | 0
concern for hemorrhagic pancreatitis | 0
pseudocysts drained | 0
1.6 L dark purulent fluid | 0
no microorganism growth | 0
hemoglobin stabilized 8.5 g/dL | 0
CT scans showed resolving pseudocyst collections | 0
pancreatic edema | 0
bilateral pleural effusions | 0
thoracentesis | 0
600 mL fluid removed | 0
WBC 664/mm3 | 0
RBC 1580/mm3 | 0
PMN 62% | 0
glucose 81 mg/dL | 0
protein 2.2 g/dL | 0
LDH 232 µ/L | 0
Pseudomonas aeruginosa pneumonia | 0
IV meropenem course | 0
Clostridium difficile-associated diarrhea | 0
oral vancomycin 500 mg every 6 hours | 0
IV metronidazole 500 mg every 8 hours | 0
transferred to general medical ward | 0
weaned off ventilator | 51
trach collar | 51
significant improvement in symptoms | 0
tolerating oral feeds | 0
second ERCP | 0
CBD stent removal | 0
PEG tube removal | 0
discharged | 102
subacute rehabilitation facility | 102
1.5 LPM supplemental oxygen | 102
