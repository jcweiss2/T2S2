42 years old | 0
male | 0
admitted to the hospital | 0
dysuria | 0
right-sided loin pain | 0
blood pressure 140/80 mmHg | 0
pulse 80 beats/minute | 0
temperature 38.5°C | 0
white cell count 12.5 × 103/mm3 | 0
haemoglobin 9.5 g/L | 0
platelet count 568 × 103/mm3 | 0
albumin 32 g/L | 0
serum creatinine 258 μmol/L | 0
urea 15.8 mmol/L | 0
potassium 6.2 mmol/L | 0
bicarbonate 16 mmol/L | 0
intravenous co-amoxiclav | 0
E. coli sensitive to co-amoxiclav | 0
urine culture | 0
blood culture | 0
immunosuppression | 0
tacrolimus | 0
prednisolone | 0
clinical condition deteriorated | 168
antibiotic therapy | 168
stable graft function | 168
serum blood glucose level risen to 50 mmol/L | 168
transferred to the critical care unit | 168
antibiotics switched to piperacillin and tazobactam | 168
CT scan | 168
gas within both renal parenchyma | 168
bilateral emphysematous pyelonephritis | 168
intubated and ventilated | 168
inotropic support | 168
percutaneous drainage of the collection | 216
E. coli cultured from the minimal pus aspirated | 216
blood cultures grew E. coli | 216
Enterococcus | 216
Candida | 216
meropenem | 216
teicoplanin | 216
caspofungin | 216
repeat CT scan | 360
infection in both sides improved | 360
ventilatory and inotropic requirements reduced | 360
transplant graft function declined | 360
continuous veno-venous haemofiltration | 360
bilateral nephrectomies | 528
second operation for bleeding | 528
received 8 units of whole blood | 528
received 4 units of fresh frozen plasma | 528
received 2 units of cryoprecipitate | 528
patient’s condition improved | 576
transplant function recovered | 576
organ support not required | 576
histological examination of the kidneys | 576
inflammatory changes consistent with infection | 576
discharged home | 1440
serum creatinine 168 μmol/L | 1440
occasional urinary tract infections | 1440
diabetes mellitus well controlled on metformin | 1440
serum creatinine 200 μmol/L | 2592
renal failure | -5880
adult polycystic kidney disease | -5880
renal transplantation | -504
recurrent urinary tract infections | -504
established renal failure | -504
new diagnosis of diabetes mellitus | 168
post-transplant diabetes | 168