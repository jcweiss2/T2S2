48 years old | 0
male | 0
admitted to the hospital | 0
past medical history of intravenous drug abuse | -672
methadone treatment | -672
untreated chronic hepatitis C infection | -672
poorly controlled diabetes mellitus | -672
bilateral lower extremity pain | -2
severe and continuous pain | -2
no history of trauma | -2
no fever | -2
no chills | -2
no skin rashes | -2
no joint pain | -2
no atrial fibrillation | -2
no peripheral artery disease | -2
no blood clots | -2
no malignancies | -2
non-smoker | -2
last IV drug use was several months ago | -168
alert | 0
oriented | 0
afebrile | 0
hemodynamically stable | 0
BP 152/84 mm Hg | 0
heart rate 112/min | 0
temperature 97.9 F | 0
pale and cold feet | 0
normal range of motion | 0
bilateral femoral pulses were 2+ | 0
absent pedal pulses | 0
gross motor and sensory function intact | 0
white blood count of 12,900/µL | 0
hemoglobin of 10 g/dL | 0
platelet count of 144,000/µL | 0
blood glucose of 345 mg/dL | 0
normal renal function test | 0
normal liver function test | 0
normal thyroid function test | 0
normal coagulation profile | 0
sinus tachycardia | 0
prolonged QTc of 556 | 0
no atrial fibrillation | 0
multiple splenic and bilateral renal infarctions | 0
occlusion of left common iliac, left popliteal tibial, and right common femoral and right popliteal tibial arteries | 0
emergency embolectomy | 2
embolectomies involving multiple arteries | 2
intra-procedure hypoxemic respiratory failure | 2
ventilator support | 2
transthoracic echocardiogram | 4
large 1.2 cm highly mobile vegetation attached to the anterior mitral valve leaflet | 4
severe mitral regurgitation | 4
transesophageal echocardiogram | 6
small pulmonic valve vegetation | 6
patent foramen ovale | 6
broad spectrum antibiotics | 6
CT of the brain | 8
10-mm area suspicious for cerebral infarct in the right frontal lobe | 8
bilateral carotid duplex | 8
unremarkable | 8
HIV 1 and 2 antibodies non-reactive | 8
Rapid Plasma Reagin non-reactive | 8
Antiphospholipid and Beta-2 glycoprotein antibodies negative | 8
emergency cardiac catheterization | 10
100% embolic occlusion of the mid left posterior descending artery | 10
negative bacterial blood cultures | 10
embolectomy specimen examined histologically | 12
organizing blood clot with abundant fungal organisms | 12
fungal elements characterized by wide hyphae, lack of distinctive septa | 12
Mucorales | 12
empiric liposomal amphotericin B | 12
cardiothoracic surgery consulted | 12
mitral valve replacement | 12
pulmonic valve repair | 12
acute upper gastrointestinal bleeding | 14
urgent gastroenterology evaluation | 14
esophagogastroduodenoscopy | 14
3-cm friable pedunculated polypoid mass within the gastric antrum | 14
diffuse gastritis/gastropathy | 14
no active bleeding | 14
biopsy of the gastric mass | 14
negative for malignancy | 16
ventilator-dependent respiratory failure | 16
multi-organ dysfunction | 16
bacterial and fungal cultures negative | 16
aggressive medical management | 16
transiently weaned off ventilator support | 18
recurrent respiratory distress | 18
re-intubation | 18
repeat TTE | 18
increased mitral valve vegetation size | 18
additional vegetation on the posterior valve leaflet | 18
refractory shock | 18
multi-organ failure | 18
comfort care | 18
deterioration | 18
death | 432