11 years old | 0
female | 0
pallor of the lips | 0
low free T4 | 0
normal TSH | 0
uncomplicated full-term gestation | -13200
emergency cesarean section | -13200
fetal distress | -13200
maternal fever | -13200
2-week neonatal intensive care unit stay | -13200
phototherapy for hyperbilirubinemia | -13200
several urinary tract infections | -6570
septic shock | -4320
multi-organ dysfunction | -4320
nausea | -4320
vomiting | -4320
diarrhea | -4320
fever | -4320
abdominal pain | -4320
hypotension | -4320
tachycardia | -4320
tachypnea | -4320
hypoglycemia | -4320
unresponsive | -4320
intubated | -4320
broad-spectrum antibiotics | -4320
intravenous fluids | -4320
pressor support | -4320
acute renal failure | -4320
dialysis | -4320
high-dose intravenous glucocorticoids | -4320
febrile illness | -2190
sore throat | -2190
dry cough | -2190
temperature 102.5°F | -2190
blood pressure 114/69 mm Hg | -2190
empiric antibiotic therapy | -2190
episodic lip pallor | 0
dry skin | 0
denies cold intolerance | 0
denies constipation | 0
denies fatigue | 0
denies weakness | 0
denies recent change in weight | 0
well appearing | 0
weight at the 70th percentile | 0
height at the 60th percentile | 0
growth records showing a plateau | 0
mid-parental height at the 10th percentile | 0
mildly delayed deep tendon reflexes | 0
Tanner stage of B3PH1 | 0
thyroid gland not enlarged | 0
no proximal muscle weakness | 0
low free T4 | 0
mildly elevated TSH | 0
elevated TSH | 0
low IGF-binding protein-3 | 0
low IGF-1 | 0
low estradiol | 0
undetectable morning cortisol | 0
low peak cortisol on ACTH stimulation testing | 0
growth hormone deficiency | 0
gonadotropin deficiency | 0
hydrocortisone started | 24
thyroid hormone replacement initiated | 48
estrogen provided via oral contraceptive | 48
growth hormone treatment | 48
annualized growth velocity of 7.2 cm/year | 1560
first-year height gain of 6.8 cm | 8760
final height 5’7” | 26280
hypertension | 26280
low-dose lisinopril | 26280
septic shock due to adrenal crisis | -4320
adrenal insufficiency | -4320
high-dose glucocorticoids | -4320
hemodynamic instability | -4320
clinical deterioration | -4320
aggressive fluid resuscitation | -4320
empirical treatment | -4320
febrile illness | -2190
aggressively hydrated | -2190
no hypotension | -2190
no clinical decompensation | -2190
stress dosing for hydrocortisone | 0
Solu-Cortef provided for emergencies | 0