64 years old | 0
    male | 0
    multiple myeloma | 0
    admitted to the hospital | 0
    septic shock | 0
    febrile episode | 0
    lumargia | -144
    L1-2 compression fracture | -144
    vital signs at admission: blood pressure 82/60 mmHg | 0
    heart rate 78/min | 0
    body temperature 39.1℃ | 0
    respiration rate 20/min | 0
    SpO2 95% | 0
    physical examination revealed no clear focus of infection | 0
    did not complain of muscular pain | 0
    laboratory findings: massive myolysis | 0
    elevated creatinine kinase (3,582 U/L) | 0
    CK isotype analysis confirmed skeletal muscle origin (98.8%) | 0
    multiple myeloma diagnosed 5 years earlier | -43800
    IgG λ type | 0
    stage IIIA | 0
    treatment with melphalan | -43800
    prednisolone | -43800
    VAD chemotherapy | -43800
    BD chemotherapy | -43800
    thalidomide | -43800
    lenalidomide | -2160
    IgG gradually increased 6 months before current infection | -4320
    admission for sepsis caused by M. morganii | 0
    rehydration via central venous catheterization | 0
    dopamine infusion (3 mg/kg/h) | 0
    meropenem treatment (0.5 g three times a day) | 0
    cervical to pelvis CT on day of admission | 0
    no clear findings explaining massive myolysis | 0
    day 2: hypotension | 24
    day 2: oliguria | 24
    day 2: renal impairment | 24
    vital signs on day 2: blood pressure 61/45 mmHg | 24
    heart rate 87/min | 24
    body temperature 36.8℃ | 24
    hemodialysis initiated | 24
    endotoxin absorption | 24
    respiratory failure on night of day 2 | 24
    mechanical ventilation | 24
    rhabdomyolysis developed day-by-day | 24
    CK elevated to 19,790 U/L | 24
    M. morganii sensitive to broad spectrum beta-lactams | 0
    resistant to cefotiam, minomycin, ciprofloxacin | 0
    visited outpatient clinic 6 days before admission | -144
    death due to multi-organ failure | 72
    no clear focus of infection on CT | 0
    rhabdomyolysis caused by M. morganii | 0
    gram-negative bacillus rhabdomyolysis | 0
    no HIV | 0
    no Conflict of Interest (COI) | 0
    