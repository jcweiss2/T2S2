21 years old | 0
male | 0
admitted to emergency department | 0
recurrent generalized and pruritic skin lesions | -48
polymyalgia | -48
polyarthralgia | -48
no fever | -48
inflammatory syndrome | -48
hyperleukocytosis | -48
negativity of rheumatoid factor | -48
negative viral serology | -48
neurologically conscious | 0
well-oriented | 0
generalized papular cutaneous lesions | 0
erythematous pharynx | 0
no fever | 0
no headache | 0
no photophobia | 0
no neck stiffness | 0
cardiac frequency at 92/min | 0
blood pressure at 10.5/80 mm Hg | 0
saturation at 100% | 0
pulmonary examination normal | 0
cardiac examination normal | 0
abdomen soft and painless | 0
chest radiography normal | 0
leukocytosis | 0
relative polyneutrophilia | 0
elevated CRP | 0
no abnormalities of renal and hepatic functions | 0
no abnormalities of coagulation | 0
negative serologies | 0
dermatological opinion requested | 0
skin biopsy performed | 0
blood cultures performed | 0
blood cultures positive for Gram negative diplococci | 24
N. meningitidis identified by PCR | 24
intravenous treatment with Ceftriaxone | 24
transferred to intensive care unit | 24
lumbar puncture performed | 24
cerebrospinal fluid slightly turbid | 24
numerous leucocytes in cerebrospinal fluid | 24
protein in cerebrospinal fluid | 24
glucose in cerebrospinal fluid | 24
Gram staining examination negative | 24
CSF culture negative | 72
PCR positive for N. meningitidis serotype B | 72
regression of skin lesions | 72
decrease in leukocytosis | 72
decrease in CRP | 72
transferred to medical unit | 72
transesophageal ultrasound normal | 72
otolaryngology examination normal | 72
histologic examination of skin biopsy | 72
dermal ectatic lymph vessels and capillaries | 72
perivascular lymphocytic infiltration | 72
neutrophil granulocytes | 72
PAS and Gram staining negative | 72
PCR on skin biopsy positive for N. meningitidis | 72
no deficiency of classic and alternative pathway of hemolytic complement activity | 72
no deficiency of lectin pathways | 72
total IgG level slightly low | 72
IgG subclasses normal | 72
ceftriaxone treatment continued | 72
per oral quinolone treatment | 168
discharged | 168