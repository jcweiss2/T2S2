68 years old | 0
lady | 0
diagnosed with AML de novo | 0
FLT3-itd positive | 0
normal karyotype | 0
referred for allogeneic stem cell transplantation | 0
high-risk disease | 0
previously well | 0
no major comorbidities | 0
regular exercise | 0
swimming | 0
diagnosis | 0
fatigue | 0
pancytopenia | 0
blast count of 30% | 0
refractory to one course of DA-chemotherapy | 0
AML-17 | 0
excellent response to FLAG-IDA | 0
complete remission in the bone marrow | 0
1st cycle | 0
1 brother | 0
66 years old | 0
heavy smoker | 0
drinker | 0
not an ideal candidate for a potential donor | 0
unrelated donor search initiated | 0
tissue typing | 0
2nd course of FLAG-IDA | 0
complete remission | 0
underwent HLAmismatched reduced intensity-conditioned allogeneic transplant | 0
mismatch at HLA-A locus | 0
Fludarabine | 0
Busulphan for 2 days | 0
Alemtuzumab 50 mg over 2 days | 0
T-deplete | 0
matched unrelated donor | 0
day 0=13/9/14 | 0
allo-HCT | 0
first complete remission | 0
higher 3-5-year disease-free survival | 0
lower relapse risk | 0
chemotherapy | 0
auto- HCT | 0
CMV status negative (recipient) | 0
CMV positive (donor) | 0
blood groups A negative (recipient) | 0
blood groups A positive (donor) | 0
conditioning complicated by Enterobacter bacteremia | 0
E.coli bacteremia | 0
resolved following treatment with meropenem | 0
transplant well tolerated | 0
no major toxicities | 0
mild nausea | 0
diarrhea | 0
engrafted neutrophils on day +18 | 18
platelet engraftment on day +20 | 20
discharged on day +26 | 26
treated for febrile episode | 26
mild grade 1 skin GVHD | 1008
started 6 weeks post transplant | 1008
responded to topical steroids | 1008
clostridium difficile diarrhea | 1344
2 months post transplant | 1344
resolved with oral vancomycin | 1344
3-month bone marrow aspirate | 2160
trephine | 2160
100% donor chimerism in whole sample | 2160
99% donor chimerism in CD3+ T cells | 2160
ciclosporin tapered from January 2015 | 2160
ongoing diarrhea | 2160
3-4 episodes per day | 2160
flexible sigmoidoscopy | 2160
February 2015 | 2160
inflammation | 2160
no evidence of gut GVHD | 2160
ciclosporin stopped on 31st June 2015 | 4464
1-year post transplant | 8760
mild chronic skin GVHD | 8760
no sclerodermatous features | 8760
no mouth/eye/vaginal involvement | 8760
well-controlled with topical creams | 8760
stable pulmonary function | 8760
stable cardiac function | 8760
commenced on vaccination program | 8760
monthly monitoring | 8760
uneventful clinical course | 8760
attended clinic on 5/2/16 | 12528
18 months post transplant | 12528
significant reduction in Cher neutrophil count | 12528
viral screen sent | 12528
parvovirus | 12528
CMV | 12528
EBV | 12528
Adenovirus | 12528
HHV 6 | 12528
HHV 8 | 12528
urgent bone marrow arranged | 12528
relapsed disease confirmed | 12528
20% blasts detected | 12528
flt-3 ITD positive | 12528
normal cytogenetics | 12528
mixed chimerism | 12528
48% donor in whole sample | 12528
92% donor in CD3+ T cell fraction | 12528
2 months earlier | 12000
full chimera in whole blood | 12000
full chimera in T cells | 12000
commenced on azacitadine | 12528
75 mg/m2 for 7 days | 12528
1st donor lymphocyte infusion after 2 cycles | 12528
access to AC220 and Crenolanib applied for | 12528
compassionate access declined | 12528
tolerated 1st 2 cycles of azacitadine | 12528
chimerism post 2 cycles | 12528
53% donor in whole blood | 12528
91% donor in T cells | 12528
1st DLI on 14/4/16 | 13128
1×106 CD3+ cells/kg | 13128
cytopenic | 13128
required red cell transfusion | 13128
required platelet transfusion | 13128
proceeded with cycles 3 and 4 azacitadine | 13128
2nd DLI on 16/6/16 |?|
| 5x106 CD3 cells/kg | 13128
monthly cycles of azacitadine | 13128
3rd DLI on 26/8/16 |?|
| 1×107 CD3 cells/kg | 13128
attended clinic on 31st September 2016 | 16704
ongoing gastrointestinal symptoms | 16704
attributed to azacitadine | 16704
dose reduced by 50% | 16704
9th cycle started 1 week later | 16704
developed gram-negative sepsis | 16704
E.coli | 16704
brief intensive care admission | 16704
inotropic support | 16704
recovered well | 16704
bone marrow aspirate on 6/12/16 | 17136
trephine | 17136
complete morphological remission | 17136
FLT3-itd negativity | 17136
no further treatment | 17136
monitored monthly | 17136
regular blood chimerism monitoring | 17136
latest on 10/4/18 | 34320
100% donor chimerism in whole blood | 34320
100% donor chimerism in CD3+ T cells | 34320
