40 years old | 0 | 0 | Factual
African-American | 0 | 0 | Factual
female | 0 | 0 | Factual
chronic eczema | -672 | 0 | Factual
alcohol abuse | -672 | 0 | Factual
gout | -672 | 0 | Factual
hypothyroidism | -672 | 0 | Factual
worsening eruption | -720 | 0 | Factual
intermittent diarrhea | -720 | 0 | Factual
cutaneous eruption | -1440 | 0 | Factual
desquamation of the hands | -1440 | 0 | Factual
desquamation of the feet | -1440 | 0 | Factual
desquamation of the perioral skin | -1440 | 0 | Factual
desquamation of the perineal skin | -1440 | 0 | Factual
pain | -1440 | 0 | Factual
swelling | -1440 | 0 | Factual
hair loss | -1440 | 0 | Factual
increasing weakness | -2880 | 0 | Factual
fatigue | -2880 | 0 | Factual
unintentional weight loss | -2880 | 0 | Factual
weight loss 70 pounds | -2880 | 0 | Factual
drinking 1 to 2 glasses of wine a day | -672 | 0 | Factual
smoking | -672 | 0 | Factual
no significant family history | 0 | 0 | Factual
not on any medications | 0 | 0 | Factual
erythematous desquamative patches | 0 | 0 | Factual
erosions | 0 | 0 | Factual
crusted lesions | 0 | 0 | Factual
diffuse nonscarring alopecia | 0 | 0 | Factual
scaling patches on the vermillion lips | 0 | 0 | Factual
punch biopsy of the left medial thigh | 0 | 0 | Factual
psoriasiform epidermal spongiosis | 0 | 0 | Factual
superficial perivascular lymphohistiocytic infiltrate | 0 | 0 | Factual
diffuse hypogranulosis | 0 | 0 | Factual
broad overlying parakeratosis | 0 | 0 | Factual
ballooning degeneration of the spinous layer | 0 | 0 | Factual
methicillin-resistant Staphylococcus aureus sepsis | 0 | 24 | Factual
Escherichia coli sepsis | 0 | 24 | Factual
pneumonia | 0 | 24 | Factual
ventilator respiratory support | 0 | 24 | Factual
systemic antibiotics | 0 | 24 | Factual
low zinc levels | 0 | 0 | Factual
antitransglutaminase antibodies positive | 0 | 0 | Factual
antiendomysium antibodies positive | 0 | 0 | Factual
celiac disease | 0 | 0 | Factual
zinc deficiency | 0 | 0 | Factual
focal villi blunting | 0 | 0 | Factual
Brunner's gland hyperplasia | 0 | 0 | Factual
gluten-free diet | 0 | 672 | Factual
zinc sulfate | 0 | 672 | Factual
resolution of gastrointestinal symptoms | 672 | 672 | Factual
resolution of cutaneous symptoms | 672 | 672 | Factual