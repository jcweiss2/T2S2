26 years old | 0
male | 0
admitted to the hospital | 0
febrile illness | -168
involuntary movements | -168
hyperkinetic movements | -168
weakness of both upper and lower limbs | -168
autonomic dysfunction | -168
excessive sweating | -168
insomnia | -168
behavioral abnormalities | -168
auditory hallucinations | -168
resting pulse rate above 110 beats/min | 0
blood pressure elevated above 160/100 mm Hg | 0
wasting of muscles of all four limbs |> 0
hypokalemia (serum potassium: 3.2 mEq) | 0
hypoproteinemia (total protein: 5.8 g/dl) | 0
positive serum anti-CASPR2 antibody | 0
high-dose steroids | 0
intravenous immune globulin (IVIG) | 0
therapeutic plasma exchange (TPE) decision | 0
femoral line placement | 0
calcium infusion | 0
potassium correction | 0
FFP and saline replacement fluid | 0
TPE sessions | 0
hyperkinetic movements hindering flow | 0
limb restraining | 0
methyl prednisolone | 0
clonazepam | 0
allergic reaction to FFP | 0
rashes | 0
antihistamines | 0
elevated blood pressure | 0
tachycardia | 0
serum protein (5.2 g/dL) | 0
FFP transfusion | 0
total serum proteins (7.2 g/dL) | 0
hemodynamically stable | 0
improved sitting with support | 24
improved eating and walking with support | 24
mild occasional hyperkinetic movements | 24
autonomic dysfunction improvement | 24
pulse rate below 90 beats/min | 24
blood pressure below 140/90 mm Hg | 24
excessive sweating subsided | 24
restlessness subsided | 24
insomnia subsided | 24
no behavioral abnormalities | 24
anti-CASPR2 antibodies decline | 24
oral prednisolone | 0
remission | 24
