33 years old| 0
woman | 0
diagnosed with active methicillin-sensitive Staphylococcus aureus mitral valve acute bacterial endocarditis | 0
11th week of gestation | 0
high fever | 0
lower back pain | 0
admitted for intravenous antibiotic treatment for pyelonephritis | 0
platelet count decreased daily | 0
transferred to intensive care unit | 48
diagnosed with disseminated intravascular coagulation with sepsis | 48
body temperature 40°C | 48
tachycardia | 48
systolic murmur | 48
transthoracic echocardiography revealed severe mitral valve regurgitation without vegetation | 48
blood cultures grew MSSA | 0
intravenous gentamicin | 0
intravenous teicoplanin | 0
gradual improvement in inflammatory markers | 0
clinical condition worsened abruptly on hospital day 8 | 192
high-dose diuretic | 192
inotropic support | 192
noninvasive positive pressure ventilation | 192
exacerbation of mitral valve regurgitation | 192
heart failure due to mitral valve destruction | 192
minimally invasive thoracoscopic mitral valve repair | 240
fetal heart rate showed no abnormalities | 240
supine position | 240
rapid sequence induction of anesthesia | 240
tracheal intubation | 240
general anesthesia maintained with propofol | 240
oxygen-air mixture | 240
remifentanil | 240
fentanyl | 240
standard radial artery catheter | 240
Swan-Ganz catheter | 240
bispectral index monitoring | 240
cerebral oximetry monitoring | 240
intraoperative transesophageal echocardiography showed severe mitral valve regurgitation | 240
rupture of the chordae tendineae of the A3 segment | 240
other valves not affected | 240
hypothermic cardiopulmonary bypass at 32°C | 240
femoral artery cannula | 240
femoral vein cannula | 240
monitored maternal uteroplacental perfusion | 240
monitored fetus using Doppler flow ultrasound | 240
successful repair | 240
weaned off cardiopulmonary bypass with inotropic support | 240
total cardiopulmonary bypass duration 108 minutes | 240
aortic cross-clamp duration 70 minutes | 240
propofol used for sedation with dobutamine | 240
tracheal tube extubated | 240
postoperative condition favorable | 240
transvaginal ultrasound for fetal heart rate | 240
fetus diagnosed with hydrops fetalis | 312
dilation and curettage | 312
blood cultures did not detect bacterial growth | 120
antibiotics administered for 8 weeks | 0
