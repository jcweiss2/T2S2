27 years old | 0
female | 0
Filipino | 0
gravida 1 | 0
para 0 | 0
admitted to perinatology | 0
SEA heterozygote deletion | -672
partner is cis heterozygous carrier for SEA α-thalassemia deletion | -672
25% risk to fetus of having α-thalassemia major | -672
declined amniocentesis | -672
opted for expectant management | -672
initial ultrasound unremarkable | -504
follow-up ultrasound showed oligohydramnios | -336
shortened long bones | -336
severe cardiomegaly | -336
cardiothoracic circumference ratio of 0.65 | -336
Doppler velocimetry showed normal forward flow in umbilical artery | -336
middle cerebral artery peak systolic velocity of 1.49 multiples of the median | -336
referred to tertiary center for suspected Bart's hemoglobinopathy | -336
moderate hydrops | -336
informed of likely diagnosis of ATM | -336
discussed risks of IUT | -336
discussed need for chronic postnatal transfusion | -336
discussed possible bone marrow transplantation | -336
discussed increased risk for neurodevelopmental impairment | -336
elected to proceed with serial IUTs | -336
initial cordocentesis | -280
fetal hemoglobin level measured 7.9 g/dL | -280
fetal electrophoresis showed 35.3% Hb A1 and 62.5% Hb Bart | -280
IUT performed | -280
follow-up ultrasound showed resolving hydrops | -224
symmetric fetal growth restriction | -224
estimated fetal weight at 2.7th percentile | -224
hydrops and oligohydramnios resolved | -112
fetal weight at 29th percentile | -112
five IUTs performed | -112
intrauterine transfusions | -280
induced at 37 weeks' gestation | 0
delivered vaginally | 0
live, well-appearing, 2,984 g, female infant | 0
cord milking performed | 0
blow by oxygen | 0
face mask continuous positive pressure | 0
nasal CPAP for continued oxygen requirement | 0
empiric ampicillin and gentamicin started | 0
initial complete blood count significant for Hb of 19 g/dL | 0
hematocrit of 64% | 0
hypoxemic | 0
required high as 0.7 fraction inspired oxygen | 0
normal work of breathing | 0
no signs of respiratory distress | 0
chest X-ray showed mild ground glass opacities | 0
adequate lung expansion | 0
arterial blood gas unremarkable | 0
pH 7.38 | 0
PCO2 38 mm Hg | 0
PO2 95 mm Hg | 0
nasal CPAP with FiO2 at 0.67 | 0
pulse oximetry in lower extremities 5 to 10% lower than upper extremities | 0
oxygenation index calculated | 0
alveolar-arterial oxygen gradient | 0
echocardiogram showed evidence of elevated pulmonary vascular resistance | 0
estimated right ventricular systolic pressure of 65 mm Hg | 0
bidirectional shunts through patent ductus arteriosus and patent foramen ovale | 0
flattened interventricular septum | 0
no left heart obstructive lesion or myocardial dysfunction | 0
inhaled prostacyclin started | 0
immediate response demonstrated by 10 mm Hg decrease in estimated right ventricle pressure | 0
oxygen requirement decreased within 1 hour to 0.48 FiO2 | 1
weaned to 0.25 over next 24 hours | 24
inhaled PGI2 weaned off at 24 hours of life | 24
sustained improvement in oxygenation | 24
placed on high-flow nasal cannula on DOL 2 | 48
weaned to room air on DOL 5 | 120
desaturations into 80s necessitating oxygen therapy by low-flow nasal cannula on DOL 6 | 144
required oxygen between 0.21 and 0.3 FiO2 over next 14 days | 144
echocardiogram on DOL 12 demonstrated normalization of RV pressures | 288
primary pediatric hematologist consulted | 288
high hemoglobin precluded early transfusion of PRBCs | 288
hemoglobin electrophoresis from DOL 1 resulted as 45% Hb Bart, 50% Hb A, 1.3% Hb A2, and 3% Hb F | 24
partial volume exchange of 20 mL/kg with normal saline on DOL 18 | 432
transfused packed red blood cells | 432
Hb remained stable at 14.8 g/dL after transfusion | 432
oxygenation improved and weaned to room air on DOL 19 | 456
sepsis evaluation at birth | 0
initiation of empiric ampicillin and gentamicin | 0
antibiotics stopped with negative cultures at 48 hours | 48
bilirubin level reached peak of 13.6 mg/dL on DOL 2 | 48
phototherapy for 24 hours | 48
discharged 2 days after weaning to room air | 480
close follow-up with pediatric hematology within 2 weeks to set up future transfusions | 480
exhibited appropriate somatic growth for age and normal developmental milestones at 16 months | 11520
continues to receive chronic blood transfusions every 3 weeks | 11520
eczema | 11520
daily multivitamin | 11520
awaiting bone marrow transplantation | 11520