21 months old | 0
girl | 0
presented to a secondary care hospital | -720
isolated fever | -720
bacterial pulmonary infection | -720
discharged | -672
long-term course of oral antibiotics | -672
afebrile for 2 days | -672
presented to the health facility | -456
worsening abdominal pain | -456
fever | -456
no history of nausea | -456
no history of vomiting | -456
no history of any other associated sign | -456
abdominal ultrasound | -456
angio-computed tomography (CT) | -456
AAA measuring 40 mm in diameter | -456
referred to our hospital | -456
on admission | 0
hemodynamic shock | 0
pale | 0
tachycardic | 0
hypotensive | 0
admitted to the intensive care unit | 0
emergency CT scan | 0
ruptured infrarenal aortic aneurysm | 0
giant retroperitoneal hematoma measuring 93×54×92 mm3 | 0
underwent urgent surgery | 24
hemodynamic stabilization | 24
surgical exploration | 24
giant AAA compressing on approximate organs | 24
signs of inflammation | 24
signs of rupture | 24
aneurysm dissected firsthand | 24
aorta ligated below the origin of the renal arteries | 24
aorta ligated above the iliac bifurcation with 5-0 silk | 24
verifying collateral circulation on angio-CT | 24
remaining aortic aneurysm sac resected | 24
abdominal cavity rinsed | 24
closed after verifying local hemostasis | 24
put on intravenous (IV) antibiotics | 24
combination of amoxicillin | 24
combination of clavulanic acid | 24
combination of gentamicin | 24
anemia with hemoglobin at 10.5 mg/dL | 24
white blood cell count at 30,000 cells/µL | 24
erythrocyte sedimentation rate at 52 mm/hh | 24
C-reactive protein at 142.78 mg/L | 24
EKG normal | 24
echocardiography showed no signs of endocarditis | 24
postoperative angio-CT | 168
persistent retroperitoneal hematoma measuring 70×50 mm2 | 168
no signs of lower limb ischemia | 168
postoperative course remarkable for hypertension | 168
treated with combination of beta-blockers | 168
combination of ACE inhibitors | 168
combination of CCBs | 168
no other complications | 168
discharged home | 432
put on pain medication | 432
beta-blockers for 3 months | 432
pathologic examination of aortic tissue showed inflammatory signs | 432
suppuration | 432
conclusion of mycotic aneurysm | 432
microbiological cultures of aortic tissue sterile | 432
blood cultures sterile | 432
a year and a half of postoperative follow-up uneventful | 13200
no signs of lower limb ischemia | 13200
no exercise-induced fatigue | 13200
no growth retardation | 13200
long-term follow-up necessary | 13200
secondary reconstruction may be required | 13200
