31 years old| 0
male| 0
exposure to COVID-19-positive colleague| -672
COVID-19 nasal swab positive| 0
advised home quarantine/isolation| 0
acute severe left flank pain| 336
mild shortness of breath| 336
intermittent abdominal pain| 336
nausea| 336
occasional cough| 336
no fever| 336
no dehydration| 336
no vomiting| 336
no change in urinary/bowel habits| 336
mild tenderness in left lumbar region| 0
vitally stable| 0
elevated C-reactive protein| 0
elevated ferritin| 0
elevated lactate dehydrogenase| 0
mild leukocytosis| 0
deranged D-dimer| 0
deranged prothrombin time| 0
deranged INR| 0
COVID-19 nasal swab positive again| 0
normal creatinine| 0
normal eGFR| 0
no proteinuria| 0
negative thrombophilia work up| 0
negative lupus anticoagulant panel| 0
negative sickle hemoglobin| 0
negative paroxysmal nocturnal hemoglobinuria| 0
hypothyroidism| 0
treated with levothyroxine| 0
dyslipidemia| 0
treated with atorvastatin| 0
no personal/family history of hematological diseases| 0
sinus tachycardia| 0
rare premature atrial contractions| 0
rare premature ventricular contractions| 0
no intra-cardiac shunt| 0
multiple renal infarctions| 0
subpleural patchy ground glass opacities| 0
reticular opacities in lung bases| 0
COVID-19 pneumonia| 0
managed with enoxaparin| 0
replaced with warfarin| 120
injectable acetaminophen| 0
no specific treatment for COVID-19 pulmonary findings| 0
no intubation| 0
no ICU admission| 0
no supplementary oxygen| 0
focal scarring left kidney| 8784
poor compliance to warfarin| 8784
sub-therapeutic INR| 8784
advised lifelong warfarin| 8784
no supplementary oxygen|B0
