69 years old | 0
male | 0
white | 0
admitted to the hospital | 0
abdominal distension | 0
abdominal pain | 0
diabetes mellitus | -8760
hypertension | -8760
56 pack-year smoking | -8760
peritonitis | 0
severe abdominal tenderness | 0
rebound | 0
guarding | 0
white blood cell count: 9.4 × 10^9 cells/L | 0
hemoglobin: 10.9 g/dL | 0
platelets: 370 × 10^9 cells/L | 0
creatinine: 1.29 mg/dL | 0
thickening of the sigmoid colon | 0
pneumoperitoneum | 0
intraperitoneal free fluid | 0
multifocal liver lesions | 0
peritoneal and omental implants | 0
exploratory laparotomy | 2
perforated sigmoid | 2
multiple liver and omental lesions | 2
sigmoidectomy | 2
end colostomy | 2
partial omentectomy | 2
wedge resection of liver segment III | 2
admitted to the surgical intensive care unit | 2
routine postoperative care | 2
poorly differentiated SC carcinoma | 4
immunohistochemical staining | 4
primary pulmonary source | 4
tumor cells stained positive for CK5/6 | 4
tumor cells stained positive for p40 | 4
tumor cells negative for CK7 | 4
tumor cells negative for CK20 | 4
tumor cells negative for villin | 4
tumor cells negative for TTF1 | 4
right perihilar mass | 24
obstructing the right upper and middle lobe bronchi | 24
encasement of the right pulmonary artery branches | 24
extensive bulky mediastinal lymphadenopathy | 24
primary LC | 24
obstructive bronchopneumonia | 168 
died | 168