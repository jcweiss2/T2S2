45 years old | 0
female | 0
admitted to the hospital | 0
pain in abdomen | -48
vomiting | -48
caesarean section delivery | -4320
incisional hernia | -4320
LIHR | -336
ePTFE mesh placement | -336
conscious | 0
oriented | 0
pulse rate 120/min | 0
blood pressure 50mm Hg | 0
added sounds on chest auscultation | 0
mild distension | 0
tenderness | 0
rigidity | 0
guarding | 0
7cm fluctuant swelling in right lumbar quadrant | 0
blackish discoloration of overlying skin | 0
Hb 7.5 g/dl | 0
Total Leucocyte Count 5840 cells/cmm | 0
blood glucose 66 mg/dl | 0
serum creatinine 1.4 mg/dl | 0
serum albumin 1.3 g/dl | 0
serum sodium 142.6 meq/l | 0
serum potassium 3.1 meq/l | 0
loculated collection in pelvis | 0
parietal wall collection in right lower abdomen | 0
scar dehiscence | 0
patchy-confluent consolidation in bilateral lung fields | 0
admitted to ICU | 0
intravenous fluids | 0
inotropic drugs | 0
ventilatory support | 0
necrotising fasciitis of overlying abdominal wall | 0
infected mesh | 0
dense adhesions | 0
feculent fluid | 0
small bowel perforations | 0
liberal debridement | 0
resection of implanted mesh | 0
small bowel segmental resection | 0
exteriorisation of bowel ends | 0
multiorgan dysfunction syndrome | 72
expired | 72