42 years old | 0
male | 0
admitted to the hospital | 0
generalized weakness | -2160
fever | -2160
cough | -2160
12-kg weight loss | -2160
lived in Guatemala for five years | -8760
sought medical attention in Guatemala | -720
HIV-antibody test positive | -720
sputum AFB smear positive | -720
AIDS diagnosis | -720
came home to Seoul, South Korea | -720
HIV-1 Western blot test positive | -720
CD4 cell count 10/µL | -720
HIV RNA titer 18,000 copies/mL | -720
anti-tuberculosis medications started | -720
fluconazole started | -720
trimethoprim/sulfamethoxazole started | -720
generalized weakness persisted | 0
fever persisted | 0
oral thrush | 0
hepatosplenomegaly | 0
ascites | 0
hemoglobin 10.6g/dL | 0
white blood cell 2,700/µL | 0
platelet 58,000/µL | 0
total bilirubin 2.4mg/dL | 0
AST/ALT 131/48IU/L | 0
ALP 114IU/L | 0
GGT 133 IU/L | 0
costophrenic angle blunting | 0
fluid shifting in the right hemithorax | 0
mild pneumonic infiltration in left lung | 0
disseminated tuberculosis suspected | 0
Mycobacterium tuberculosis identified | 0
anti-tuberculosis medication continued | 0
anti-retroviral agents started | 24
pancytopenia progressed | 48
hemoglobin 7.4g/dL | 48
white blood cell 1,070/µL | 48
platelet 13,000/µL | 48
rifampin discontinued | 48
zidovudine discontinued | 48
trimethoprim/sulfamethoxazole discontinued | 48
new pulmonary infiltrates | 120
septic shock | 120
empirical antibiotic therapy started | 120
piperacillin/tazobactam started | 120
transferred to intensive care unit | 144
mechanical ventilator support | 144
Gram stain negative | 144
ordinary culture negative | 144
bone marrow aspiration and biopsy | 216
Histoplasma capsulatum identified | 216
disseminated histoplasmosis diagnosed | 216
died | 240