51 years old | 0
    male | 0
    end-stage renal disease | 0
    polycystic kidney disease | 0
    renal transplant (right lower quadrant, 2003) | 0
    renal transplant failure (right) due to malignant hypertension | 0
    renal transplant (left lower quadrant, 2015) | 0
    transferred from outside hospital | 0
    sepsis | 0
    E coli bacteremia | 0
    acute renal failure | 0
    hemodialysis | 0
    no history of recurrent infections | 0
    abdominal and pelvic CT scan | 0
    atrophic native kidneys | 0
    bilateral lower quadrant transplanted kidneys | 0
    right transplanted kidney appearing atrophic | 0
    intubation | 0
    pressors | 0
    broad-spectrum antibiotics | 0
    clinical status stabilized | 0
    weaned off pressor support | 144
    extubated | 144
    poor urine output | 144
    ongoing need for dialysis | 144
    transplant ultrasound performed | 144
    abdominal X-ray | 144
    development of new renal parenchymal gas | 144
    emphysematous pyelonephritis (EPN) | 144
    repeat CT confirmed diagnosis | 144
    management escalated | 144
    percutaneous drain placed | 144
    clinical picture declined | 168
    increasing pressor support required | 168
    re-intubated | 168
    taken emergently to OR for nephrectomy | 168
    nephrectomy performed | 168
    left lower quadrant modified Gibson incision | 168
    infected kidney soft and boggy | 168
    infarcted kidney | 168
    liquefaction necrosis | 168
    bed irrigated | 168
    drain left in situ | 168
    pathology indicated endarteritis | 168
    chronic transplant arteriopathy | 168
    arterial thrombi | 168
    cortical infarctions | 168
    thrombotic microangiopathy | 168
    micro abscess formation | 168
    extubated | 192
    pressor support discontinued | 192
    progressive ischemia | 192
    prolonged pressor use | 192
    peripheral artery disease | 192
    bilateral amputation | 192
    transmetatarsal amputation | 192
    bilateral knee amputation | 192
    worsening sepsis | 240
    lower limb extremity tissue necrosis | 240
    passed away | 240
    cardiopulmonary arrest | 240
    