42 years old | 0
female | 0
motorcycle accident | -720
fracture of the middle third of the right clavicle | -720
Allman's group I (AO 15-B1) | -720
deviation >2 cm | -720
right shoulder abrasions | -720
analgesics | -720
no sling use | -720
no therapeutic follow-up | -720
pain | -240
fever | -240
local hyperemia | -240
hospitalization | -240
febrile peaks | -216
local edema | -216
skin fluctuation on the right clavicle region | -216
drainage of a purulent secretion | -216
abscess drainage | -336
cleansing with 0.9% saline solution | -336
no material for culture | -336
leukogram WBC 12,000/mm3 | -336
eosinophilia (3% rods) | -336
ESR 25 mm/h | -336
CRP 11 mm/dl | -336
intravenous antibiotic therapy | -336
ceftriaxone 1 g 12/12 h | -336
metronidazole 500 mg 8/8 h | -336
clindamycin 600 mg 8/8 h | -336
admission to Salvador medical service | -600
extensive lesion of the right hemithorax | -600
toxemia | -600
sepsis | -600
HR 110 bpm | -600
RF 26 ripm | -600
Temp 38.5 °C | -600
clavicle bone exposure | -600
extensive necrosis of the skin | -600
no neurovascular alterations | -600
leukogram WBC 21,000/mm3 | -600
eosinophilia (5% rods) | -600
ESR 44 mm/h | -600
CRP 20 mm/dl | -600
creatinine 1.3 mg/dl | -600
urea 48 mg/dl | -600
CPK 900 u/l | -600
MRI thorax | -600
MRI neck | -600
ICU admission | -600
surgical debridement | -600
bone tissue culture | -600
antibiotic therapy modification | -600
meropenem 1 g 8/8 h | -600
vancomycin 1 g 12/12 h | -600
anti-tetanus prophylaxis | -600
osteolysis in the clavicle | -576
increase in necrotic area | -576
right clavicle resection | -576
aggressive debridement of devitalized tissue | -576
soft tissue culture | -576
bone culture | -576
clinical improvement | -576
discharged from ICU | -528
reduction of WBC | -528
reduction of inflammatory markers | -528
purulent secretion diminished | -528
special dressing every other day | -528
borders of lesion ceased necrosis | -528
raw area without purulent secretion | -528
granulation tissue | -528
negative bone culture | -528
negative soft tissue culture | -528
skin graft | -528
discharge from hospital | -528
complete wound healing | 1440
excellent upper limb functional score | 1440
healed wound | 4320
