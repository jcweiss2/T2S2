63 years old | 0
female | 0
168 cm height | 0
53 kg weight | 0
papillary thyroid carcinoma | -9720
resection | -9720
radiotherapy | -9720
stenosis of the esophagus | -8760
repeated aspiration | -8760
respiratory insufficiency | -8760
pneumonia | -8760
purulent pleurisy | -8760
pleurectomy | -8760
restrictive ventilation pattern | -8760
recurrent nerve palsy | -8760
percutaneous endoscopic gastrostomy | -7200
tracheostoma | -7200
home ventilation | -7200
decreased mobility | -8760
secondary depression | -8760
fixed mandible | -8760
limited mouth opening | -8760
stented left axis vertebralis | -4380
stenosis of the internal axis carotis | -4380
arterial hypertension | -4380
secondary lactase deficiency | -4380
esophageal stenosis dilation | -120
fistula between the esophagus and tracheal membrane | -120
decreasing general condition | 0
admitted to the University of Erlangen | 0
examined by chiefs and consultants | 0
deemed too unstable for open surgery | 0
inability to open the mouth | 0
recurrent nerve palsy | 0
referred to the surgical intensive care unit | 15
pneumonia by 4-multiresistente gramnegative Pseudomonas aeruginosa | 15
veno-venous extracorporeal membrane oxygenation | 15
partial thromboplastin time of 60 seconds | 15
preseptic status | 15
ventilated through a tracheostoma | 15
thoracic computed tomography | 16
big fistula of the tracheal membrane | 16
tracheal cannula ended shortly beneath the lower limit of the mediastinal fistula | 16
decision to try endobronchial stenting | 16
plan to close the fistula with a pedicled omentum majus replacement | 16
surgical plastic needed an abutment and a secured continuous airway replacement | 16
procedure performed on October 28, 2016 | 17
vv-ECMO began to be partly ineffective | 17
high volume input of physiological saline | 17
oral approach would only allow a small flexible bronchoscope | 17
approach for the upper part of the trachea had to be performed through the percutaneous tracheostoma | 17
retrograde stenting | 17
Dumon and one-hybrid self expandable metalic y-stent | 17
Freitag stent | 17
mandatory additional ventilation | 17
nasal jet catheter | 17
double-lumen endotracheal tube exchange catheter | 17
ventilation line introduced either orally or through the tracheostoma | 17
successful retrograde stenting performed in four steps | 17
Step I | 17
regular bronchoscopes, jagwires, jet-catheters, and DLETs | 17
manually compressed “y” of the FS pushed downward on the main carina | 17
Step II | 18
frontal surface of the stent cut with at least 1 cm opening | 18
stent surface reduced ~40% in the sagittal axis | 18
new stoma for a regular tracheal cannula created | 18
lower new edge of this stoma fixed subcutaneously | 18
Step III | 19
jagwire introduced through the mouth into the trachea | 19
jagwire running out of the new FS stoma | 19
DLET introduced for more stability | 19
distal jagwire introduced into the oral orifice of the FS | 19
FS flipped with its upper part over the soft-tip stiff DLET into the upper third of the trachea | 19
whole fistula bridged by the FS up to the level of the vocal cords | 19
upper edge of the new FS stoma fixed subcutaneously | 19
Step IV | 20
regular tracheal cannula introduced for ventilation | 20
lungs not aerated at that point of time | 20
spontaneous breathing work increased | 20
vv-ECMO support reduced | 20
lungs became re-aerated again | 20
patient woke up again | 20
could communicate with her family by writing and her eyes | 20
infections continued to be very severe | 20
spontaneous work of breathing never exceeded a tidal ventilation of 170 mL per breath | 20
reduction of intravenous saline injection limited | 20
vv-ECMO support mandatory but reduced | 20
patient and family decided to reduce vv-ECMO support | 20
patient died on 18 November 2016 | 30
pulmonary infection | 30