28 years old | 0
woman | 0
large left-to-right shunt through secundum ASD measuring 25 mm | 0
normal pulmonary venous drainage to the left atrium | 0
normal ventricular function on echocardiogram | 0
admitted for transcatheter closure | 0
negative RT-PCR for COVID-19 infection | 0
normal preprocedural blood investigations | 0
elevated right atrial pressure to 9 mmHg | 0
elevated left ventricular end-diastolic pressure to 12 mmHg | 0
normal pulmonary artery pressure | 0
placement of stiff guidewire and delivery sheath in the left upper pulmonary vein | 0
defect closure using 34 mm Cera septal occluder under transesophageal echocardiographic guidance | 0
LVEDP not rechecked after device closure | 0
brief postprocedural endotracheal bleeding delayed extubation by 48 hours | 0
managed with protamine to reverse the effect of heparin | 0
packed red cell transfusion for hemoglobin drop of 2 g/dl from baseline | 0
chest X-ray in baseline showed cardiomegaly with increased pulmonary flow | 0
chest X-ray postprocedure showed left upper zone infiltrates suggestive of lung bleed | 0
developed progressive respiratory distress after extubation | 48
hypoxia after extubation | 48
radiological evidence of acute respiratory distress syndrome | 48
pre-discharge chest X-ray showed resolution of radiological findings | 168
echocardiogram showed dilated right heart chambers | 72
significant biventricular systolic dysfunction | 72
mild pleural effusion | 72
mild pericardial effusion | 72
elevated right ventricular systolic pressures | 72
computed tomography excluded pulmonary thromboembolism | 72
computed tomography showed pleural effusion | 72
computed tomography showed lung collapse | 72
computed tomography showed features suggestive of pulmonary edema | 72
elevated inflammatory biomarkers | 72
CRP 24 mg/L | 72
d-Dimer 2335 ng/mL | 72
troponin I levels elevated to 0.075 ng/mL | 72
COVID RT-PCR repeatedly negative | 72
COVID total antibodies elevated to 209 units/ml | 72
unavailability of NT-proBNP | 72
unavailability of interleukin-6 | 72
unavailability of COVID antibody IgM fraction test | 72
differential diagnosis included infection | 72
differential diagnosis included pulmonary thromboembolism | 72
differential diagnosis included postA COVID inflammatory syndrome | 72
treated with supplemental oxygen | 72
treated with enoxaparin 40 units twice daily | 72
transitioned to warfarin | 72
treated with broad-spectrum antibiotic | 72
treated with aspirin | 72
treated with beta-blocker | 72
treated with sildenafil | 72
treated with diuretics | 72
responded well with reduction of biomarkers | 168
plan to start methylprednisolone abandoned due to clinical recovery | 168
discharged on day 7 postprocedure | 168
hemodynamically stable condition at discharge | 168
on aspirin at discharge | 168
on warfarin at discharge | 168
on weaning schedule of sildenafil at discharge | 168
echocardiogram before discharge showed reduction of right ventricular dimensions | 168
echocardiogram before discharge showed reduction of pleural effusion | 168
echocardiogram before discharge showed recovery of ventricular systolic function | 168
asymptomatic on 15-month follow-up | 1128
normal effort tolerance on 15-month follow-up | 1128
