2.980 Kg | 0
male | 0
admitted to the hospital | 0
perinatal asphyxia | 0
intubated | 0
transferred to NICU | 0
blood pressure 70/50 mmHg | 0
heart rate 144 beats/min | 0
breathing rate 66/min | 0
respiratory distress | 48
afebrile | 48
tachypnic | 48
no history of aspiration | 48
no lethargy | 48
no rash | 48
blood pressure 52/38 mmHg | 48
pulse rate 186/min | 48
S1 muffled | 48
S2 muffled | 48
lungs clear on auscultation | 48
ECG low voltage QRS complex | 48
ECG non-specific ST-T wave changes | 48
mild leucocytosis (13800/mm3) | 48
normal cardiac troponin | 48
normal CK | 48
normal CK-MB | 48
chest X-ray halo sign | 48
endotracheal tube deep in right main bronchus | 48
echocardiography air bubbles in pericardial sac | 48
diastolic collapse of right atrium | 48
diastolic collapse of right ventricular outflow tract | 48
normal bi-ventricular functions | 48
ruled out infection | 48
ruled out sepsis | 48
ruled out ARDS | 48
ruled out myocarditis | 48
hemodynamic instability | 48
tamponade physiology | 48
intravenous normal saline | 48
ceftriaxone 250 mg | 48
pericardiocentesis | 48
aspirated 40-50 ml air | 48
blood pressure 66/42 mmHg | 48
endotracheal tube repositioned | 48
ECG minimal air on anterior cardiac surface | 72
pericardial sheath removed | 72
repeated chest X-ray complete resolution of PPC | 72
weaned off mechanical ventilation | 168
discharged | 240
27-year-old mother | 0
primigravida | 0
primipara | 0
prolonged second stage of labour | 0
prolonged third stage of labour | 0
Apgar score 4 at 1 minute | 0
Apgar score 7 at 5 minutes | 0
Apgar score 10 at 10 minutes | 0
mechanical ventilation | 0
subcutaneous emphysema | -48
interstitial emphysema | -48
pneumomediastinum | -48
pneumothorax | -48
pneumoperitonium | -48
no fever | 48
normal blood count | 48
temporal course of events | 48
clear lung fields on auscultation | 48
normal chest X-ray (initially) | 0
pericardiocentesis under echocardiographic guidance | 48
informed consent obtained | 48
sub-costal area aseptically prepared | 48
skin infiltration with 2% xylocaine | 48
21-G needle inserted | 48
guide wires inserted | 48
4F radial angiographic sheath inserted | 48
underwater seal connected | 48
wire and dilator removed | 48
hemodynamic stability restored | 48
repeated ECG minimal air | 72
sheath in situ | 48
air aspiration | 48
endotracheal tube tip repositioned | 48
minimal air on anterior cardiac surface | 72
complete resolution of PPC | 72
gradual weaning off mechanical ventilation | 168
stable condition | 240
