23-week gestational age | 0
    female | 0
    born | 0
    HELLP syndrome | 0
    cesarean section | 0
    birthweight 485 grams | 0
    Apgar score 3 | 0
    Apgar score 8 | 0
    intubated | 0
    received surfactant | 0
    mechanical ventilation | 0
    transferred to neonatal intensive care unit | 0
    WBC 2.1×10^9/L | 0
    hematocrit 39.6% | 0
    hemoglobin 12.6 g/100 mL | 0
    platelet 186×10^3/mL | 0
    differential 9% segmental WBC | 0
    1% bands | 0
    60% lymphocytes | 0
    26% monocytes | 0
    603 nucleated red blood cells per 100 WBC | 0
    CRP less than 0.3 mg/dL | 0
    persistent neutropenia | 0
    thrombocytopenia | 0
    bandemia | 0
    hemodynamically significant hypotension | 0
    vasopressors | 0
    no definitive infection | 0
    ampicillin | 0
    gentamicin | 0
    early-onset sepsis | 0
    blood culture | 0
    anaerobic gram-positive branching rods | 0
    Actinomyces species | 0
    culture sent to reference laboratory | 0
    ampicillin switched to penicillin | 0
    Actinomyces bacteremia | 0
    ampicillin | 0
    gentamicin | 0
    penicillin | 0
    total antibiotic course 13 days | 0
    subsequent blood culture no growth | 0
    Actinomyces viscosus identified | 0
    16S ribosomal RNA gene sequencing | 0
    MALD-TOF unable to identify organism | 0
    clinically significant hypotension | 0
    vasopressor support | 0
    stress dose corticosteroid | 0
    persistent neutropenia | 0
    thrombocytopenia | 0
    disseminated intravascular coagulation | 0
    transient hypoglycemia | 0
    electrolyte imbalance | 0
    adrenal insufficiency | 0
    acute renal failure | 0
    endotracheal aspirate grew Staphylococcus aureus | 744
    urine culture grew Enterococcus faecalis | 744
    central line grew Staphylococcus epidermidis | 744
    clinical evidence of infection | 744
    vancomycin | 744
    ampicillin/sulbactam | 744
    discharged | 2160
    HELLP syndrome | -672
    preterm labor | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    maternal serology negative for HIV | -672
    hepatitis | -672
    chlamydia | -672
    syphilis | -672
    group B streptococcal status unknown | -672
    pregnancy complicated by HELLP syndrome | -672
    HELLP syndrome leading to cesarean section | -672
    respiratory distress requiring mechanical ventilation | 0
    sepsis at birth | 0
    persistent anemia | 0
    pulmonary hypertension | 0
    cardiac hypertension | 0
    cardiogenic pressor | 0
    stress dose corticosteroid | 0
    secondary infection at 30 days | 720
    Staphylococcus aureus oxacillin susceptible | 744
    Enterococcus faecalis | 744
    Staphylococcus epidermidis | 744
    no copious vaginal discharge | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    negative repeat blood culture | 168
    clinical instability | 0
    prolonged antibiotic therapy | 0
    risks of antibiotic resistance | 0
    microbiota alteration | 0
    impaired neutrophils | 0
    vulnerability to infection | 0
    contamination in neonatal blood culture | 0
    unnecessary antibiotic exposure | 0
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm illness of the mother | -672
    HELLP syndrome | -672
    extreme prematurity | -672
    preterm