29 years old| 0
pregnant | 0
female | 0
fever | -96
cough | -96
presented at emergency room | 0
second pregnancy | -20160
full-term cesarean delivery | -20160
regular antenatal visits | 0
body mass index 35 kg/m² | 0
anomaly scan at 20 weeks | -4032
glucose tolerance test at 24 weeks | -2016
last routine antenatal visit | -336
admitted to isolation ward | 0
X-ray showed patchy infiltrates | 0
nasopharyngeal swab confirmed COVID-19 | 0
prophylactic medication | 0
shifted to ICU | 72
intravenous piperacillin-tazobactam | 72
therapeutic dose of enoxaparin | 72
continuous positive airway pressure | 72
respiratory distress worsened | 72
intubated | 96
mechanical ventilation | 96
unable to maintain saturation | 96
synchronised intermittent mandatory ventilation | 96
pressure-regulated volume control | 96
multidisciplinary team decision | 96
ECMO insertion | 96
midazolam 5 mg/hour | 96
fentanyl 300 µg/hour | 96
cisatracurium 8 mg/hour | 96
effective anticoagulation | 96
activated partial thromboplastin time 53.2 seconds | 96
ECMO drainage cannula inserted | 96
ECMO return cannula inserted | 96
VVECMO circuit initiated | 96
fetal heart monitored | 96
transferred to Dubai Hospital | 96
monitored in surgical ICU | 96
daily fetal cardiotocography | 96
repeat COVID-19 swab negative | 168
condition improved | 168
weaned off ECMO | 168
haemodynamic stability | 168
monitored in general antenatal ward | 168
chest physiotherapy sessions | 168
fetal growth parameters normal | 168
umbilical artery Doppler studies normal | 168
white blood cell count 8.2 | 0
platelet count 145-198 | 0
D-dimer 1.03-1.23 | 0
blood sugar levels | 0
liver function tests | 0
renal function tests | 0
troponin T | 0
pro-brain natriuretic peptide | 0
ferritin 366-45 | 0
APTT levels 50-60 | 96
discharged | 552
advised to taper prednisolone | 552
enoxaparin once a day | 552
32-week outpatient antenatal visit | 1344
fetal growth parameters | 1344
transthoracic echocardiography | 1344
chest X-ray indicative of disease severity | 0
negative COVID-19 swab | 168
ECMO run for 5 days | 168
no significant bleeding | 168
no cannula dislodgement | 168
no haemolysis | 168
no superadded infections | 168
methylprednisolone 40 mg IV | 72
oral prednisolone 30 mg | 168
intramuscular betamethasone | 0
magnesium for neuroprotection | 0
enoxaparin started | 0
heparin infusion during ECMO | 96
enoxaparin continued after ECMO | 168
long-term follow-up | 1344
discharged home | 552
normal respiration | 552
obstetrical ultrasound Doppler studies | 552
ambulating | 552
maintaining saturation | 552
haemodynamically stable | 552
chest physiotherapy | 552
multivitamins | 552
pantoprazole | 552
ambroxol syrup | 552
ferritin increased | 336
D-dimer decreased | 336
lactate normal | 336
CKMB normal | 336
troponin normal | 336
chest X-ray improved | 336
patient perspective | 552
learning points | 552
multidisciplinary team | 552
counselling with relatives | 552
long-term outcome monitoring | 552
