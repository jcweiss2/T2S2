43 years old|0
male|0
admitted to the surgical ward|0
upper abdominal pain|-24
colic|-24
vomiting|-24
diarrhea|-24
history of similar attacks|0
afebrile|0
hemodynamically stable|0
right upper abdominal tenderness|0
positive Murphy's sign|0
leucocytosis (18 × 10³/mm³)|0
normal liver function tests|0
normal electrolytes|0
gall bladder stone|0
signs of acute cholecystitis|0
intravenous fluids|0
ceftriaxone|0
metronidazole|0
dalteparin|0
laparoscopic cholecystectomy|6
edematous gall bladder|6
single gall bladder stone|6
adhesions|6
normal other abdominal organs|6
perioperative period uneventful|6
intra-abdominal pressure 12-15 mmHg|6
acute cholecystitis on top of chronic cholecystitis|6
postoperative recovery well|6
scheduled discharge post-LC day 2|48
severe epigastric pain|48
afebrile|48
normal vital signs|48
severe leucocytosis (34 × 10³/mm³)|48
partial SMA obstruction|48
secondary small bowel ischemia|48
small bowel obstruction|48
dilatation proximal small bowel|48
ischemic terminal ileum|48
good SMA pulsation|48
ileum resection|48
anastomosis|48
Bogota bag closure|48
transfer to SICU|48
full heparinization|48
intubation|48
sedation|48
ventilation|48
second look laparotomy day 4|120
viable healthy bowel|120
no anastomosis leakage|120
abdominal wall closure|120
heparinization resumed|126
total parenteral nutrition started|120
normal echocardiogram|120
no embolism signs|120
no deep venous thrombus|120
sinus rhythm|120
no atrial fibrillation|120
increased abdominal distension day 12|288
intra-abdominal pressure 24 mmHg|288
hemoglobin 6.3 g/dl|288
blood transfusion|288
blood products received|288
abdominal collections day 13|312
deteriorated condition day 14|336
abdominal distension|336
full ventilatory support|336
oliguria|336
intra-abdominal pressure 25 mmHg|336
abdominal compartment syndrome diagnosis|336
decompressive laparotomy|336
old blood-stained fluid collection drained|336
Bogota bag closure|336
unstable condition|336
inotropic support|336
high fever (39.2°C) day 15|360
septic shock|360
renal failure|360
renal replacement therapy started|360
asystole day 16|384
death|384
