18 years old | 0
male | 0
admitted to the hospital | 0
fever | -24
vomiting | -24
generalized abdominal pain | -24
rash on palms and trunk | -24
no conjunctivitis | -24
severe drowsiness | -24
lethargic | -24
tender to palpation | -24
right lower quadrant | -24
negative meningeal signs | -24
tachycardic | -24
hypotension | -24
no associated murmurs | -24
white blood cell count of 13.5 × 103/μL | -24
segmented neutrophils, 94.5% | -24
erythrocyte sedimentation rate, 82 mm/h | -24
serum C-reactive protein, 298.5 mg/L | -24
procalcitonin concentrations, 18.45 mcg/L | -24
negative for SARS-CoV-2 by both rapid PCR and RT-PCR | -24
positive history of contact | -24
positive serology of SARS-CoV-2 (immunoglobulin G (IgG)) | -24
ferritin, IL6, high-sensitivity troponin, and D-dimer were all elevated | -24
enoxaparin, an anticoagulant | -24
IV immunoglobulin (IVIG; 2 g/kg) | -24
325 mg of aspirin per day | -24
red blood cell transfusion | -48
pulse dosage of systemic corticosteroids (30 mg/kg daily methylprednisolone) | -48
dobutamine | -48
favorable progression | -72
afebrile | -72
clinical symptoms improved | -72
arterial pressure was stable without inotropes | -72
histopathological examination resulted in the diagnosis of catarrhal appendicitis | -72
D-dimer showed a downward trend | -72
troponemia had resolved | -72
inflammatory parameters were normal | -72
LV function was improved, demonstrating normal biventricular function | -72
no aneurysms were observed in the proximal coronary artery system | -72
discharged | -72
follow-up outpatient visit after 2 weeks | -96
blood tests had normalized | -96
COV-2 IgG was elevated to 84 | -96
abdominal and cardiac ultrasounds were normal | -96