48 years old | 0
    male | 0
    hypertension | -720
    dyslipidemia | -720
    sudden onset of chest pain | -24
    ST-segment elevation on leads I, aVL, V1–V6 | -24
    ST-segment depression on leads II, III, aVF | -24
    severely impaired motion of the anterolateral wall of the left ventricle | -24
    white blood cell count of 19100/μL | -24
    lactase dehydrogenase level of 213 IU/L | -24
    creatinine kinase level of 77 mg/dL | -24
    C-reactive protein level of 0.6 mg/dL | -24
    D-dimer level of 1.85 μg/mL | -24
    AMI on the anterolateral wall of the left ventricle | -24
    emergent coronary angiography | -24
    severe narrowing of the LMT | -24
    PCI with IVUS guidance | -24
    intimal flap extending from the aortic wall of the ascending aorta to the ostium of the LMT | -24
    severe compression of the LMT ostium | -24
    critical AMI | -24
    pooling of blood in the false channel of the localized aortic dissection | -24
    collapsed with sustained ventricular tachycardia | -24
    resuscitated with tracheal intubation | -24
    recovered with normal sinus rhythm | -24
    drug-eluting stents placed from LMT ostium to LAD artery | -24
    severe hypotension persisted | -24
    VA-ECMO established | -24
    transferred to operating room for emergency surgery | -24
    exposed ascending aorta through median sternotomy | 0
    no signs of aortic dissection | 0
    localized hematoma on the posterior wall of the ascending aorta | 0
    trans-esophageal echocardiography showed localized dissection | 0
    CPB with tepid hypothermia (32°C) | 0
    cannulation of ascending aorta and right atrium | 0
    aortic cross clamping | 0
    antegrade and retrograde cardioplegia | 0
    distal side coronary artery bypass grafting to LAD and circumflex branch using SVGs | 0
    additional cardioplegic solution given selectively from SVGs | 0
    dissecting part of ascending aorta transversely opened | 0
    inside ascending aorta showed atherosclerotic changes | 0
    entry found at 15-mm distal site above LMT orifice | 0
    LMT dissected (Neri’s classification type B) | 0
    localized dissection encompassed one-third circumference of ascending aorta | 0
    localized at left Valsalva sinus and right Valsalva sinus | 0
    LMT compression | 0
    localized dissection repaired by obliterating false lumina | 0
    several mattress sutures of 4-0 Prolene with inside and outside felt strips | 0
    surgical glue (BioGlue) used | 0
    reinforced edges closed with horizontal mattress sutures | 0
    over-and-over sutures of 4-0 Prolene | 0
    proximal side coronary artery bypass grafting performed | 0
    CPB time 283 min | 0
    aortic cross clamping time 172 min | 0
    weaning from CPB unsuccessful | 0
    severely impaired left ventricle due to AMI | 0
    VA-ECMO and IABP support established | 0
    transferred to intensive care unit with VA.ECMO and IABP | 0
    maximum creatine kinase level of 7712 U/L | 0
    postoperative contrast-enhanced computed tomography showed successful repair | 0
    cardiac dysfunction persisted 5 days after operation | 120
    transferred to specialized hospital for left ventricular assist device | 120
    died of severe sepsis | 2880
    <|eot_id|>
    