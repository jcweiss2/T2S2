83 years old | 0\
male | 0\
admitted to the hospital | 0\
leg ecchymosis | 0\
anuric | 0\
rhabdomyolysis-induced AKI | 0\
septic state | 0\
syncope | -12\
fell to the ground | -12\
lying on the floor throughout the night | -12\
prostatic hypertrophy | -8760\
overactive bladder | -8760\
recurrent prostatitis | -8760\
statins | -8760\
volume expansion | 0\
diuretic | 0\
alpha-agonist | 0\
antibiotic treatment | 0\
furosemide | 0\
femoral central venous catheter | 0\
HFR-Supra | 0\
endogenous reinfusion | 0\
remove myoglobin | 0\
reduce the inflammatory status | 0\
maintain the fluid balance | 0\
ultrafiltration | 0\
adsorbent cartridge | 0\
low flux polyphenylene membrane | 0\
high-dose furosemide | 0\
intravenous fluids | 0\
24-h urine output 300 mL | 96\
24-h urine output 2,400 mL | 192\
furosemide tapered | 192\
oral administration | 192\
piperacillin/tazobactam | 0\
meropenem | 0\
E. coli resistant to piperacillin/tazobactam | 0\
myoglobin reduction | 120\
CPK reduction | 120\
LDH reduction | 120\
CRP reduction | 120\
PCT reduction | 120\
HFR-Supra sessions | 120\
femoral hemodialysis catheter removed | 168\
right jugular central venous catheter | 168\
on-line hemodiafiltration | 168\
high-flux hemodialysis | 168\
Phylter HF 17G dialyzer | 168\
dialysis no longer required | 504\
discharge | 504\
urea 96 mg/dL | 504\
creatinine 3.06 mg/dL | 504\
CRP 3.2 mg/dL | 504\
total bilirubin 0.81 mg/dL | 504\
ASL 27 IU/L | 504\
ALT 25 IU/L | 504\
PSA 61 ng/mL | 504\
white blood cells count 6,300 cells/µL | 504\
urea 89 mg/dL | 2160\
creatinine 2.41 mg/dL | 2160\
GFR 24 mL/min | 2160