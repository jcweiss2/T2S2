35 years old | 0
gravida 2 para 2 | 0
no previous history of chronic medical illnesses | 0
gestational diabetes | 0
presented at 16 weeks of gestation | 0
acute-onset excruciating headache | 0
tonic-clonic convulsions | 0
low Glasgow Coma Scores | 0
intubation | 0
computed tomography scan | 0
left frontal hematoma | 0
mild edema | 0
mass effect | 0
midline shift of 4 mm to the right | 0
bleeding spread to the left lateral ventricle | 0
third ventricle | 0
fourth ventricle | 0
left subdural hematoma | 0
open basal cisterns | 0
CT angiography of the brain | 0
frontal lobe bleeding | 0
carotid bifurcation aneurysm | 0
small subarachnoidal bleeding | 0
intraventricular bleeding | 0
possible hydrocephalus | 0
sent to the operating room | 0
trial of coiling of the aneurysm | 0
failed coiling | 0
admitted to the intensive care unit | 0
monitoring | 0
supportive measures | 0
remained sedated | 0
mechanical ventilation | 0
2 mm size midposition pupils | 0
sluggish reaction to light bilaterally | 0
second trial of endovascular coiling | 24
failed coiling | 24
sudden dilatation of the left pupil to 3 mm | 48
sluggish reaction to light | 48
right pupil remained 1 to 2 mm in size | 48
heart rate dropped to 55–59 beats/minute | 48
blood pressure of 110/60 mmHg | 48
managed with crystalloid and colloid therapy | 48
low doses of norepinephrine | 48
urgent CT of the brain | 48
modest subarachnoidal rebleeding | 48
spastic reaction of the vessels | 48
extended ischemia in the middle cerebral artery | 48
signs of mesotemporal herniation | 48
third ventricle well separated | 48
flow problem at the aqueduct level | 48
another trial of coiling | 72
difficult coiling | 72
occlusion of the left carotid system by a thrombus | 72
CT of the brain showed deterioration | 72
ischemic areas better demarcated | 72
midline shift increased | 72
increase in the effacement of gyri and sulci | 72
cerebral angiography | 72
thrombosis in the left internal cerebral artery | 72
thrombosis in the MCA | 72
no carotid artery aneurysm | 72
partial mechanical thrombectomy | 72
failed coiling | 72
pupils became fixed and dilated at 7 mm bilaterally | 72
decompressive craniotomy | 72
placement of external ventricular drains | 72
monitoring intracranial pressure | 72
ventilated and sedated | 72
fixed dilated pupils | 72
no cough or gag reflexes | 72
ICP monitor reading of less than 10 mmHg | 72
ICP started rising | 96
ICP reached up to 50 mmHg | 96
medical management for high ICP | 96
muscle relaxants | 96
mannitol | 96
hypertonic saline infusions | 96
thiopental coma | 96
ICP remained elevated | 96
removal of the monitor | 168
GCS of 3 | 168
no gag or cough reflexes | 168
pupils 5 mm dilated and fixed | 168
sedation stopped | 192
apnea test not done | 192
EEG not done | 192
diagnosis confirmation | 192
full ventilatory support | 192
nutritional support | 192
vasoactive drugs | 192
maintenance of normothermia | 192
supportive measures | 192
110-day hospital course | 0
severe hypotension | 0
managed with vasopressors | 0
hypertension | 0
treated with antihypertensives | 0
intranasal DDAVP | 0
water flushes through nasogastric tube | 0
diabetes insipidus | 0
hypernatremia | 0
episodes of sepsis | 0
pneumonia | 0
urinary tract infection | 0
line infection | 0
treated with antibiotics | 0
meningitis | 0
treated with meropenem | 0
treated with vancomycin | 0
panhypopituitarism | 0
thyroid hormone replacement | 0
steroids | 0
hypothermia | 0
managed with passive rewarming and blankets | 0
tracheostomy | 432
feeding through NG tube | 0
consensus of family | 0
multidisciplinary approach | 0
ethics committees involved | 0
decision to continue somatic support | 0
cesarean section planned at 32 weeks | 0
ultrasound scan revealed IUGR | 0
biometry corresponding to 25 weeks | 0
estimated fetal weight of 650 gm | 0
oligohydramnios | 0
no fetal anomalies | 0
intrauterine monitoring | 0
serial ultrasounds | 0
heart rate monitoring | 0
amniocentesis | 0
betamethasone therapy | 0
lower segment cesarean section | 2640
preterm male in breech presentation | 2640
Apgar score of 6/7/9 | 2640
average weight of 750 gm | 2640
transferred to NICU | 2640
nasal CPAP applied | 2640
apnea test done twice | 2640
positive apnea tests | 2640
death pronounced | 2640
