79 years old | 0
female | 0
presented to the Emergency Department | 0
slurred speech | 0
arm weakness | 0
deteriorating mobility | -2160
cognition | -2160
oral intake | -2160
radioactive iodine treatment for hyperthyroidism | -11640
iatrogenic hypothyroidism | -11640
stopped taking levothyroxine | -2880
temperature of 33.3°C | 0
heart rate of 45 bpm | 0
blood pressure of 170/99 mmHg | 0
oxygen saturations were 90% on room air | 0
GCS was 9/15 | 0
dry flaky skin | 0
coarse hair | 0
frontal balding | 0
globally depressed reflexes | 0
hoarse voice | 0
peripheral oedema | 0
no palpable goitre | 0
focal right cerebellar calcification | 0
Na+ 127 mmol/l | 0
CRP 19 mg/l | 0
creatine kinase (CK) 586 IU/l | 0
TSH 51 mU/l | 0
T4 2.6 pmol/l | 0
T3 <0.8 pmol/l | 0
cortisol 1,001 nmol/l | 0
re-warming initiated | 0
broad-spectrum intravenous antibiotics | 0
T4 25 μg via the nasogastric (NG) route | 0
T3 replacement three times a day | 0
hydrocortisone | 0
admitted to the critical care unit | 0
passed away | 672
recurrent hospital-acquired pneumonias | 672
non-ST-elevation myocardial infarction (NSTEMI) | 672
per rectum bleed | 672
raised CK secondary to thyroid myositis | 672