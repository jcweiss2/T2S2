19 years old | 0
male | 0
mild asthma | 0
admitted to the hospital | 0
scratched by a cat | -168
fever | -168
deep venous thrombosis | -168
fondaparinux treatment | -168
apixaban treatment | -161
macroscopic hematuria | -7
leg edema | -7
asthenia | -7
persistent fever | -7
lethargic | 0
Glasgow Coma Scale 15/15 | 0
blood pressure 100/66 mm Hg | 0
sinus tachycardia | 0
mitral murmur | 0
hemocultures taken | 0
piperacillin started | 0
ceftriaxone/gentamicin started | 0
Hb 6.3 g/dL | 0
red blood cells transfused | 0
anterograde amnesia | 0
cerebral computed tomography | 0
nuclear magnetic resonance scan | 0
large hematoma in left occipitoparietal region | 0
multiple bilateral microhemorrhage | 0
hematoma next to right cerebellum | 0
hematoma in right occipital region | 0
multiple ischemic microlesions | 0
left cerebellar ischemic stroke | 0
intracerebral mycotic aneurysm | 0
embolization of mycotic aneurysm | 0
transthoracic echocardiography | 0
large vegetation on mitral valve | 0
mitral valve prolapse | 0
septic shock | 0
intubated | 0
sedated | 0
norepinephrine started | 0
dobutamine started | 0
wake-up test | 12
obeying commands | 12
no neurological deficits | 12
emergency surgery | 48
minimal cardiopulmonary bypass | 48
in situ right radial arterial line | 48
left internal jugular central venous line | 48
intubated | 48
ventilated | 48
sedated | 48
hemodynamically supported | 48
tranexamic acid given | 48
MCPB primed | 48
retrograde priming technique | 48
Hb dropped to 7.8 g/dL | 48
red blood cells transfused | 48
mean arterial blood pressure maintained | 48
anterograde and retrograde cold cardioplegia | 48
central body temperature cooled | 48
transesophageal echocardiography | 48
surgical time kept to a minimum | 48
biological mitral valve replacement | 48
nonin cerebral oximeter | 48
tissue oxygen saturation monitored | 48
heparin administration | 48
activated clotting time monitored | 48
protamine given | 48
MCBP weaning | 48
atrioventricular pacemaker stimulation | 48
fresh frozen plasma transfused | 48
platelets transfused | 48
postoperative intensive care unit stay | 72
norepinephrine infusion | 72
reoperation to remove thromboemboli | 96
ventilation-acquired pneumonia | 96
tracheostomy | 96
percutaneous gastric feeding | 96
rehabilitation medicine | 432
good neurological recovery | 432
no loss in memory capacity | 432
no signs of neurological deficits | 432
discharged home | 432
residual bilateral claudication | 432
follow-up nuclear magnetic resonance | 432
resorption of occipital and left cerebellar hematoma | 432