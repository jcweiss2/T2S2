76 years old | 0
female | 0
Multiple Myeloma | -304
end-stage kidney disease | -304
fatigue | -304
bone pain | -304
weight loss | -304
hemodialysis | -304
Systemic Arterial Hypertension | -304
Glucose Intolerance | -304
International Staging System III | -304
Durie Salmon stage IIIB | -304
Myeloma Frailty Score: 3 | -304
Bortezomib | -168
Dexamethasone | -168
hypercalcemia | -168
anemia | -168
renal impairment | -168
lytic lesions | -168
admitted to emergency service | -72
confusion | -72
hip pain | -72
respiratory distress | -68
COVID-19 diagnosed | -68
plasmacytoma | -68
nasal swab real time polymerase chain reaction | -68
SARS-COV-2 | -68
computed tomography | -68
peripheral ground-glass opacities | -68
antibiotic therapy | -68
Ceftriaxone | -68
Vancomycin | -68
discharged | 0
RT-PCR test | 17
recovered symptoms | 17
delirium | 17
radiotherapy | 104
Daratumumab | 104
chills | 111
tremors | 111
hemodialysis | 111
negative blood culture | 111
dyspnea | 112
acute respiratory failure | 112
hypoxemia | 112
COVID-19 positive | 112
nasal swab RT-PCR | 112
SARS-COV-2 | 112
negative serology | 112
SARS-COV-2 IgG | 112
SARS-COV-2 IgM | 112
close family members infected | 112
Shilley catheter-related bloodstream infection | 112
Pseudomonas aeruginosa | 112
extended spectrum beta-lactamase | 112
blood culture | 112
Meropenen | 112
Vancomycin | 112
Dexamethasone | 112
catheter exchanged | 112
clinical stability | 119
Chest Computer Tomograph | 119
febrile event | 133
antibiotics escalated | 133
Polymixicin | 133
Linezolid | 133
RT-PCR SARS-COV-2 | 135
undetectable | 135
hemodynamic instability | 137
refractory septic shock | 137
Klebsiella pneumonia | 137
carbapenemase | 137
intensive care | 137
mechanical ventilation | 137
high-dose vasoactive drug | 137
death | 141