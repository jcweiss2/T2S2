50 years old | 0
female | 0
admitted to the Emergency Department | 0
continuous abdominal pain | -144
vomiting | -144
lactic acidosis | 0
thrombocytopenia | 0
rheumatic heart disease | -43296
aortic valve replacement | -43296
mitral valve replacement | -43296
chronic renal failure | -17280
anemia | -17280
palpitation | -672
fever | -672
endocarditis | -672
methicillin-resistant Staphylococcus intermedius | -672
neoplasm around the mechanical aortic valve | -672
serum creatinine 331 µmol/L | -672
estimated glomerular filtration rate 23 mL/min/1.73 m2 | -672
hemoglobin 78 g/L | -672
leukocytes 8.7×10^9/L | -672
polymorphonuclear neutrophils 7.57×10^9/L | -672
platelets 216×10^9/L | -672
LZD 600 mg intravenously every 12 hours | -672
warfarin 1.25 mg orally every 12 hours | -672
improved condition | -408
major symptoms disappeared | -408
body temperature returned to normal | -408
multiple blood culture results negative | -408
discharged | -408
drowsy | 0
dyspneic | 0
nausea | 0
vomiting | 0
persistent periumbilical pain | 0
no fever | 0
no chill | 0
no cough | 0
no diarrhea | 0
no expectoration | 0
no rash | 0
tachypneic (28 breaths/min) | 0
atrial fibrillation (83 beats/min) | 0
normotensive (112/50 mmHg) | 0
afebrile (36.5°C) | 0
microbiological investigations negative | 0
no sputum specimen collected | 0
severe lactic acidosis | 0
transferred to Emergency Intensive Care Unit | 24
worsening condition | 24
heart rate 115 beats/min | 24
atrial fibrillation | 24
blood pressure 70/35 mmHg | 24
respiratory rate 30 breaths/min | 24
hemodynamic support with norepinephrine | 24
mechanical ventilation | 24
continuous renal replacement therapy | 24
2U erythrocytes | 24
1U platelets | 24
shock | 24
multiple organ failure | 312
died | 312
D+25 admission | 600
D+26 | 624
D+27 | 648
D+28 | 672
PH 6.94 | 600
PCO2 <10 mmHg | 600
PO2 178 mmHg | 600
serum lactate >20 mmol/L | 600
Tot Bili 4.6 µmol/L | -48
serum creatinine 331 µmol/L | -48
platelet count 216×10^9/L | -48
leukocyte count 8.7×10^9/L | -48
red blood cell count 2.8×10^12/L | -48
PH 6.86 | 624
PCO2 14 mmHg | 624
PO2 118 mmHg | 624
serum lactate >20 mmol/L | 624
Tot Bili 5.4 µmol/L | 0
serum creatinine 333 µmol/L | 0
platelet count 271×10^9/L | 0
leukocyte count 8.45×10^9/L | 0
red blood cell count 3.04×10^12/L | 0
PH 7.09 | 648
PCO2 16.8 mmHg | 648
PO2 449.6 mmHg | 648
serum lactate >20 mmol/L | 648
Tot Bili 7.2 µmol/L | 120
serum creatinine 300 µmol/L | 120
platelet count 197×10^9/L | 120
leukocyte count 7.65×10^9/L | 120
red blood cell count 2.50×10^12/L | 120
PH 7.08 | 672
PCO2 24.5 mmHg | 672
PO2 100.3 mmHg | 672
serum lactate >20 mmol/L | 672
Tot Bili 7.1 µmol/L | 240
serum creatinine 316 µmol/L | 240
platelet count 143×10^9/L | 240
leukocyte count 5.50×10^9/L | 240
red blood cell count 2.71×10^12/L | 240
Tot Bili 8.1 µmol/L | 600
serum creatinine 496 µmol/L | 600
platelet count 12×10^9/L | 600
leukocyte count 4.15×10^9/L | 600
red blood cell count 2.02×10^12/L | 600
Tot Bili 7.6 µmol/L | 624
serum creatinine 467 µmol/L | 624
platelet count 15×10^9/L | 624
leukocyte count 3.36×10^9/L | 624
red blood cell count 2.46×10^12/L | 624
Tot Bili 9.9 µmol/L | 648
serum creatinine 322 µmol/L | 648
platelet count 59×10^9/L | 648
leukocyte count 3.06×10^9/L | 648
red blood cell count 2.04×10^12/L | 648
Tot Bili 10.5 µmol/L | 672
serum creatinine 291 µmol/L | 672
platelet count 40×10^9/L | 672
leukocyte count 2.41×10^9/L | 672
red blood cell count 2.76×10^12/L | 672
