22 years old | 0
male | 0
temporal lobe epilepsy | 0
mental retardation | 0
sodium valproate | 0
Levetiracetam | 0
generalized tonic clonic seizure | 0
three episodes within 15 minutes | 0
without returning to baseline consciousness between the seizures | 0
sedated | 0
intubated | 0
admitted to the Intensive Care Unit | 0
status epilepticus | 0
fever >38°c | 48
increased tracheobronchial secretions | 48
leukocyte count 18.3 x 109/mL | 48
culture tracheobronchial secretions showed Pseudomonas aeruginosa | 48
chest X-ray right lower lobe consolidation | 48
diagnosis of ventilator-associated pneumonia | 48
extubated | 96
stayed in ICU for 5 days | 96
transferred back to ward | 120
febrile | 144
hypotensive | 144
transferred back to ICU | 144
antibiotics modified to Piperacillin-Tazobactam and Vancomycin | 144
no mechanical ventilation | 144
improvement on second day of ICU stay | 168
afebrile | 192
transferred out of ICU to ward | 192
vital signs stable | 192
maintaining oxygen saturation on room air | 192
returned back to baseline condition | 192
progressive bulbar weakness | 336
ataxia | 336
pulse 48 beats per minute | 336
blood pressure 96/63 mmHg | 336
temperature 36.9°c | 336
ophthalmoplegia | 336
finger to nose dysmetria | 336
dysdiadochokinesia | 336
abnormal heel to shin test | 336
generalized areflexia | 336
difficulty in standing | 336
lumbar puncture | 336
CSF analysis proteins 100mg/dl | 336
white cell count 10 | 336
MRI brain and spine shows atrophic left hippocampus | 336
mesial temporal sclerosis | 336
anti-GD1b 198 | 336
anti-GD1a 175 | 336
anti-GM1 154 | 336
anti-GM2 41 | 336
anti-GQ1b <30 | 336
diagnosis of sero-negative MFS | 336
received 5 sessions of IVIG | 336
hemodynamic status improved | 360
blood pressure 113/67mmHg | 360
heart rate 68–75 beats per minutes | 360
neurologic symptoms did not improve | 360
hemodynamics stabilized | 360
rehabilitation team consulted | 360
written informed consent | 360
institutional approval not required | 360
