25 years old | 0
female | 0
admitted to the hospital | 0
epigastric pain | -144
intermittent low-grade fever | -144
multiple hospitalizations | -144
postprandial vomiting | -144
breathing difficulty on exertion | -144
orthopnoea | -144
loss of appetite | -144
weight loss | -144
severe shock | 0
tachycardia | 0
tachypnoea | 0
hypotension | 0
tenderness over the epigastric region | 0
left infrascapular crepts | 0
decreased breath sounds | 0
fluid resuscitation | 0
inotropes | 0
IV antibiotics | 0
Azithromycin | 0
Piperacillin/Tazobactam | 0
blood culture | 0
portable chest radiograph | 0
pneumopericardium | 0
2D-Echo | 0
cardiac tamponade | 0
echogenic materials in the pericardial space | 0
pericardiocentesis | 0
frank pus | 0
pyo-pneumopericardium | 0
IV Fluconazole | 0
intubation | 7
mechanical ventilation | 7
worsening metabolic acidosis | 7
deterioration of clinical condition | 13
death | 24
Hemoglobin | 0
total WBC | 0
Platelet count | 0
Total bilirubin | 0
direct bilirubin | 0
total protein | 0
albumin | 0
SGOT | 0
SGPT | 0
alkaline phosphatase | 0
Creatinine | 0
urea | 0
Sodium | 0
Potassium | 0
Bicarbonate | 0
Lipase | 0
Amylase | 0
Malarial parasite | 0
Procalcitonin | 0
Prothrombin time | 0
INR | 0
APTT | 0
Viral markers | 0
XPERT TB PCR test | 24
AFB smear | 24
Culture fungus | 24
Culture- aspirated pus | 24
Escherichia coli | 24
Serial arterial blood gas | 0
pH | 0
PCo2 | 0
PO2 | 0
Sodium | 0
Potassium | 0
Lactate | 0
Bicarbonate | 0
Chloride | 0
Glucose | 0
BEecf | 0
FIO2 | 0