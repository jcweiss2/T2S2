53 years old | 0  
    male | 0  
    long-standing left renal calculi | -2160  
    left-side pyelolithotomy | -2160  
    postoperative placement of a DJS | -2160  
    DJS placement not under fluoroscopy guidance | -2160  
    no postoperative imaging examinations | -2160  
    advised for stent removal after 5 months | -2160  
    KUB x-ray film showed abnormal DJS location | -2160  
    DJS appeared to enter into the IVC | -2160  
    transferred to our hospital | 0  
    moderate flank pain persisted | 0  
    normal leukocytes counts | 0  
    normal creatinine levels |3  
    increased leukocytes counts in urine | 0  
    increased erythrocyte counts in urine | 0  
    urine culture positive for Enterococcus faecalis | 0  
    CDFI showed small mural thrombus in IVC | 0  
    treated with anticoagulants | 0  
    treated with antibiotics | 0  
    next-day CTU performed | 24  
    CTU showed left-side hydronephrosis | 24  
    migration of DJS into IVC at left renal vein level | 24  
    proximal coil in IVC | 24  
    distal coil in left renal pelvis | 24  
    percutaneous nephroscope under C-arm guidance | 48  
    used 18G puncture needles | 48  
    used 20 Fr working sheaths | 48  
    distal coil of DJS visualized | 48  
    DJS removed successfully | 48  
    new DJS placed | 48  
    new DJS location confirmed by radiologic imaging | 48  
    transferred to ICU | 48  
    continued anticoagulants | 48  
    continued antibiotics | 48  
    CDFI showed no thrombus in IVC | 360  
    discharged | 384  
    symptom free | 384  
    follow-up uneventful | 384  
    