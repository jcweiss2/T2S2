47 years old | 0
    male | 0
    admitted to the emergency department | 0
    increasing weight loss over 6 weeks | -1008
    sudden onset dyspnea | 0
    chest pain | 0
    micro haemoptysis | 0
    low-grade fever | 0
    fatigue | 0
    fever | 0
    skin paleness | 0
    mild tachycardia | 0
    laterocervical lymphadenopathy | 0
    ECG sinus tachycardia | 0
    ECG right bundle branch block | 0
    ECG negative T waves in V1-V4, DIII, and aVF | 0
    chest-abdomen-pelvis CT pulmonary infarction | 0
    chest-abdomen-pelvis CT renal infarction | 0
    chest-abdomen-pelvis CT splenic infarction | 0
    chest-abdomen-pelvis CT bilateral pulmonary thromboembolism | 0
    brain CT hypodense lesion in right parietal lobe | 0
    TTE and TEE mobile echogenic mass on mitral valve | 0
    vascular Doppler ultrasonography no deep vein thrombosis | 0
    suspected bacterial endocarditis | 0
    admitted to Department of Cardiology | 0
    normal complete blood count | 0
    normal erythrocyte sedimentation rate | 0
    normal procalcitonin level |1
    normal C-Reactive Protein |1
    normal blood ion levels |1
    normal coagulation tests |1
    normal amylase |1
    normal urea |1
    normal creatinine |1
    elevated transaminase levels |1
    elevated D-dimers |1
    negative blood cultures |1
    intravenous cefuroxime |1
    intravenous gentamicin |1
    subcutaneous enoxaparin |1
    right-sided hemiparesis (4/5) |192
    severe motor aphasia |192
    brain MRI multiple embolic infarctions |192
    repeated TEE vegetation on mitral valve |192
    no mitral stenosis |192
    no mitral regurgitation |192
    negative hereditary thrombophilia panel |192
    normal antithrombin III |192
    normal protein C |192
    normal protein S |192
    normal Factor V Leiden |192
    normal methylenetetrahydrofolate reductase mutation screening |192
    negative autoimmune panel |192
    normal anti-cardiolipin IgG and IgM |192
    normal antinuclear antibodies |192
    negative lupus anticoagulant |192
    normal tumour markers (alpha-fetoprotein, carcinoembryonic antigen, prostate-specific antigen) |192
    elevated Cyfra 21-1 |192
    normochromic normocytic anemia |336
    decreased hemoglobin to 6.5 g/dl |336
    decreased haematocrit to 19.5% |336
    gastroscopy ulcerated gastric adenocarcinoma |336
    biopsy poorly differentiated gastric adenocarcinoma |336
    worsening neurological status |336
    tetraparesis |336
    left hemiplegia |336
    cerebral CT new right sylvian artery infarction |336
    impaired consciousness |336
    respiratory failure |336
    transfer to intensive care unit |336
    increased intracranial pressure |672
    transtentorial brain herniation |672
    death |672

    