38 years old | 0
female | 0
admitted to hospital | 0
bacteraemia | 0
fever | -48
nausea | -48
sepsis | 0
MSSA bacteraemia | 0
infection of CRT-D device | 0
intravenous antibiotics started | 0
vancomycin | 0
piperacillin-tazobactam | 0
cefazolin | 0
extraction of device generator and transvenous leads | 24
debridement of device pocket | 24
blood cultures negative for growth | 216
new device generator placed | 432
biventricular epicardial lead placement | 432
1st episode of cardiac tamponade | 600
pericardiocentesis | 600
colchicine | 600
2nd episode of cardiac tamponade | 672
repeat pericardiocentesis | 672
prednisone | 672
ibuprofen | 672
pericardial window with small-bore chest tube placement | 744
discharge home from hospital | 912
intravenous antibiotics completed | 1224
repeat echocardiogram showed no pericardial effusion | 1824
chest tube removed | 1824
repeat echocardiogram showed no pericardial effusion | 2928
permanent atrial fibrillation | 0
AVJ ablation | 0
heart failure with reduced ejection fraction | 0
non-ischaemic cardiomyopathy | 0
Type 2 diabetes | 0
obesity | 0
hyperlipidaemia | 0
lisinopril | 0
metformin | 0
metoprolol succinate | 0
rivaroxaban | 0
spironolactone | 0
torsemide | 0
left-sided CRT-D pocket infection | -672
device extraction and re-implantation | -672
MSSA bacteraemia | -672
dizziness | 600
diaphoresis | 600
malaise | 600
elevated leucocyte count | 600
stable haemoglobin | 600
elevated C-reactive protein | 600
elevated erythrocyte sedimentation rate | 600
normal anti-nuclear antibody | 600
normal C3 complement | 600
normal C4 complement | 600
normal thyroid-stimulating hormone | 600
AF with complete heart block | 600
100% ventricular pacing | 600
marked enlargement of cardiac silhouette | 600
pericardial effusion | 600
RV collapse | 600
diastolic RV collapse | 600
systolic right atrial collapse | 600
pericardial drain | 600
normal nucleated cell count | 600
neutrophilic predominance | 600
normal pericardial fluid protein | 600
serum protein | 600
no bacterial or fungal growth | 600
computed tomography scan | 600
appropriate position of epicardial electrodes | 600
re-accumulation of pericardial effusion | 672
elevated intracardiac filling pressures | 672
impending tamponade | 672
pericardial window | 744
small-bore chest tube | 744
drainage from chest tube | 912
transthoracic echocardiogram | 912
no significant pericardial effusion | 912
colchicine | 912
ibuprofen | 912
prednisone taper | 912
intravenous cefazolin | 912
stable condition | 912
asymptomatic | 1824
minimal drainage | 1824
no effusion recurrence | 1824
chest tube removed | 1824
feeling well | 2928
no pericardial effusion recurrence | 2928
epicardial lead settings | 2928