29 years old | 0
male | 0
admitted to the hospital | 0
cardiogenic shock | -720
biventricular failure | -720
ejection fraction 5-10% | -720
myopericarditis | -720
constrictive physiology | -720
PICC line placed | -720
discharged on milrinone | -720
fever | -24
chills | -24
septic shock | 0
PICC line removed | 0
IV vancomycin | 0
piperacillin/tazobactam | 0
vasopressor support | 0
Chryseobacterium indologenes | 48
ciprofloxacin | 48
pericardiectomy | 264
discharged from the hospital | 504
inotrope independent | 504
follow-up | 7440
no evidence of recurrent infection | 7440
NYHA Class I | 7440
non-ischaemic cardiomyopathy | -720
viral myopericarditis | -720
constrictive pericarditis | -720
atrial flutter | -720
radiofrequency ablation | -720
inotrope therapy | -720
home milrinone infusion | -720
peripherally inserted central catheter | -720
elective pericardiectomy | -24
fever of 38.7°C | -24
tachycardia | -24
hypotension | 0
elevated lactate level | 0
blood cultures drawn | 0
Gram-negative rods | 48
infectious disease team consulted | 48
susceptibility testing | 48
sensitivity to ciprofloxacin | 48
sensitivity to piperacillin | 48
sensitivity to trimethoprim/sulfamethoxazole | 48
resistance to meropenem | 48
improved clinically | 120
weaned off vasopressor support | 120
negative blood cultures | 120
interval echocardiogram | 168
left ventricular EF increased | 168
right ventricular systolic dysfunction improved | 168
inotrope independent | 504
guideline-directed medical therapy | 504
furosemide | 504
metoprolol succinate | 504
sacubitril-valsartan | 504
follow-up transthoracic echocardiogram | 7440
no evidence of valvular stenosis | 7440
no evidence of valvular regurgitation | 7440
no evidence of vegetations | 7440
simultaneous right and left heart catheterization | 168
discordance of right and left ventricular pressures | 168
diastolic equalization of pressures | 168
constrictive pericarditis | 168
dense areas of adhesions | 264
calcium laterally and towards the apex of the heart | 264
pericardiectomy | 264
complete removal of the pericardium | 264
left ventricular EF increased to 50-55% | 312
right ventricular systolic dysfunction improved | 312
intravenous piperacillin/tazobactam | 504
oral ciprofloxacin | 504
total of 14 days of antibiotics | 504
discharged following completion of antibiotic course | 504