87 years old | 0
    white | 0
    male | 0
    end-stage renal disease | 0
    atrial fibrillation | 0
    warfarin | 0
    maintenance home hemodialysis | 0
    NxStage machine | 0
    laparoscopic appendicectomy | 0
    intra-abdominal abscess | 0
    sepsis | 0
    tamponade | 0
    bloody pericardial effusion | 0
    emergent therapeutic pericardiocentesis | 0
    intensive care unit | 0
    warfarin discontinued | 0
    discharged home | 0
    heparin-free home hemodialysis | 0
    Fresenius machine | 0
    Optiflux 160 NR dialyzers | 0
    pump-delivered normal saline flushes | 0
    extracorporeal circuits clotting | 0
    filters clotting | 0
    high venous pressures | 0
    compromised home hemodialysis | 0
    heparin contraindicated | 0
    flushes with 250-500 mL normal saline | 0
    aliquots every 15-30 minutes | 0
    failed to prevent clotting | 0
    warfarin contraindicated | 0
    consideration to stop home hemodialysis | 0
    discussion of peritoneal dialysis switch | 0
    literature review failed | 0
    CAR-170-C NXSTAGE Chronic cartridge | 0
    early clot formation at 12-o'clock position | 0
    blood pooling | 0
    first signs of clotting | 0
    rotating filter 60 degrees clockwise | 0
    returning to neutral position | 0
    rotating filter 60 degrees counterclockwise | 0
    repeated cycles of rotations | 0
    resolved clotting problem | 0
    lines stopped clotting | 0
    no saline flushes needed | 0
    smooth heparin-free home hemodialysis | 0
    treatment sessions interrupted due to clotting | 0
    sessions lasting almost twice as long | 0
    sessions abandoned | 0
    observed fibrin formation at 12-o'clock position | 0
    Locke-Onuigbo Maneuver | 0
    reproducible results | 0
    heparin-free and saline-flush-free home hemodialysis | 0
    patient satisfaction | 0
    wife's detailed diary | 0
    December 2019 difficult month | 0
    January 2020 smooth treatments | 0
    hypothesis of antigravity effect | 0
    no air trap in CAR-170-C cartridge | 0
    novel method confirmed | 0
    electric motor proposal | 0

<|eot_id|>