42 years old | 0 | 0 
female | 0 | 0 
admitted to the hospital | 0 | 0 
altered mental status | 0 | 0 
low grade fevers | -120 | 0 
sudden deterioration in mental status | 0 | 0 
history of intravenous drug use | -8760 | -720 
extraction of all maxillary teeth | -2160 | -2160 
mandibular dental infection | -720 | -720 
treated with oral amoxicillin | -720 | -720 
temperature was 36.7 °C | 0 | 0 
heart rate was 98 beats/min | 0 | 0 
respiratory rate was 17 breaths/min | 0 | 0 
blood pressure was 131/66 mm Hg | 0 | 0 
oxygen saturation of 99% on room air | 0 | 0 
denies fevers | 0 | 0 
denies chills | 0 | 0 
denies chest pain | 0 | 0 
denies dyspnea | 0 | 0 
denies nausea | 0 | 0 
denies vomiting | 0 | 0 
denies diarrhea | 0 | 0 
denies skin lesions | 0 | 0 
denies numbness | 0 | 0 
denies tingling | 0 | 0 
denies weakness of the lower extremities | 0 | 0 
prominent holosystolic murmur at the apex | 0 | 0 
petechial rash scattered on the abdomen | 0 | 0 
petechial rash scattered on the palms | 0 | 0 
petechial rash scattered on the soles of the feet | 0 | 0 
encephalopathy | 0 | 0 
facial droop | 0 | 0 
slurred speech | 0 | 0 
admitted to the intensive care unit | 0 | 0 
started on empiric antibiotic treatment with vancomycin | 0 | 72 
started on empiric antibiotic treatment with meropenem | 0 | 72 
unresponsive to voice | 24 | 24 
minimally responsive to pain | 24 | 24 
left hemi-neglect | 24 | 24 
right gaze deviation | 24 | 24 
Glasgow Coma Scale (GCS) was 6 | 24 | 24 
intubated for airway protection | 24 | 24 
leukocytosis of 24.7 × 109/L | 0 | 0 
87.6% neutrophils | 0 | 0 
platelet count of 17 × 109/L | 0 | 0 
liver and kidney functions were within normal | 0 | 0 
declined a HIV test | 0 | 0 
innumerable acute to subacute embolic infarcts in both cerebral and cerebellar hemispheres | 0 | 0 
proximal right internal carotid artery T-shaped acute thrombus | 0 | 0 
occlusion of the right middle cerebral artery | 0 | 0 
subarachnoid hemorrhage in the right parietal region | 0 | 0 
subarachnoid hemorrhage around the posterior aspect of the midbrain | 0 | 0 
echo densities on the tricuspid valve | 0 | 0 
echo densities on the aortic valve | 0 | 0 
echo densities on the mitral valve | 0 | 0 
blood culture grew S. marcescens | 0 | 0 
antibiotic changed to cefepime | 72 | 72 
cardiothoracic surgery consulted | 72 | 72 
poor candidate for surgery | 72 | 72 
no cough or gag reflex | 144 | 144 
pupils were fixed and mid-dilated | 144 | 144 
withdraw care | 144 | 144 
discharged to hospice care | 144 | 144