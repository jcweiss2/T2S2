63 years old| 0
male | 0
alcoholic cirrhosis | -672
abdominal pain | -504
admitted to the hospital | 0
cachectic | 0
icteric |;0
holosystolic murmur | 0
abdomen diffusely tender | 0
abdomen distended | 0
erythematous macules | 0
purpuric macules | 0
papules scattered diffusely | 0
white blood cell count of 16.8 k/uL | 0
hemoglobin of 10 g/dl | 0
platelets of 292 k/uL | 0
prothrombin time 27.8 s | 0
sodium of 125 mEq/L | 0
potassium of 4.8 mmol/L | 0
urea of 54 mg/dL | 0
creatinine 3.3 mg/dL | 0
bilirubin 9.1 mg/dL | 0
alanine transaminase of 24 U/L | 0
aspartate transaminase of 76 U/L | 0
alkaline phosphatase of 93 U/L | 0
lactic acid dehydrogenase 829 U/L | 0
total protein of 7.4 g/dL | 0
albumin of 2.6 g/dL | 0
INR of 2.3 | 0
paracentesis | 0
ascitic fluid cell count of 2000 cells/mm3 | 0
polymorphonuclear cell count PMN of 700 cells/mm3 | 0
started on Piperacillin and Tazobactam | 0
blood culture revealed gram-positive cocci in clusters | 48
Vancomycin added | 48
final culture positive for MSSA | 72
paracentesis fluid culture positive for MSSA | 72
echocardiogram showed vegetation on the mitral valve 17 mm x 4 mm | 72
antibiotics changed to cefazolin | 72
no candidate for surgery | 72
kidney function continued to deteriorate | 72
urine studies showed UNa of 79 mEq/L | 72
U creatinine of 50.2 mg/dL | 72
FENa of 4.1% | 72
daily EKG did not show AV block | 72
no persistent fever | 72
no bacteremia | 72
hepatorenal syndrome | 72
started on octreotide | 72
started on midodrine | 72
started on albumin | 72
no response | 72
needed hemodialysis | 72
discharged to rehab | 216
long-term intravenous antibiotics for 6 weeks | 216
repeat echocardiogram showed improvement in valve function | 216
clearance of vegetation | 216
clinical course continued to deteriorate | 216
multiple admissions for refractory symptomatic ascites | 216
hepatic hydrothorax | 216
recurrent pleural effusion | 216
acute liver failure | 216
encephalopathy | 216
not a candidate for transplantation | 216
active alcohol abuse within last 6 months | 216
placement of palliative peritoneal drainage catheter | 216
transferred to tertiary care for TIPS | 216
pre-TIPS bilirubin of 2.6 mg/dL | 216
