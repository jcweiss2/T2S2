79 years old | 0
male | 0
septic shock | 0
urosepsis | 0
multi-organ failure | 0
acute on chronic renal failure | 0
acute respiratory distress syndrome | 0
Arterial hypotension | 0
drowsy mentation | 0
APACHE II score 32 | 0
started on CytoSorb therapy | 15
started on SLED | 15
standard surviving sepsis guidelines treatment | 15
improved hemodynamic parameters | 72
improved ventilator requirements | 72
increasing urine output | 72
APACHE II score 8 | 72
IL-6 levels 1356.3 pg/ml | 0
IL-6 levels 26.12 pg/ml | 72
deteriorated clinically | 120
CytoSorb hemadsorption | 15
SLED for 6 h every day | 15
immunosuppression | 120
removal of helpful anti-inflammatory cytokines | 120 
IL-1 | -1
IL-6 | -1
IL-8 | -1
tumor necrosis factor | -1
IL-10 | -1
tumor growth factor-β | -1