48 years old | 0
female | 0
brought to the emergency room | 0
shortness of breath | -3
headache | -3
nausea | -3
increased blood pressure | 0
painless loss of vision in both eyes | 0
no history of hypertension | 0
no other comorbidities | 0
no other significant history | 0
heart rate of 104/min | 0
blood pressure of 220/120 mm Hg | 0
basal crepitations | 0
drowsy | 0
arousable | 0
normal pupillary reflex | 0
normal extra-ocular movements | 0
normal fundoscopy | 0
no light perception | 0
no signs of meningeal irritation |+ 0
normal hemoglobin | 0
mild leukocytosis | 0
elevated C-reactive protein | 0
normal ESR | 0
normal liver function tests | 0
normal renal function tests | 0
normal other blood tests | 0
normal coagulation profile | 0
normal autoantibodies | 0
normal neoplastic markers | 0
cerebrospinal fluid protein increase | 0
chest radiography showing pulmonary edema | 0
normal arterial blood gas analysis | 0
MRI brain showing T2/FLAIR hyperintensities | 0
managed in intensive care unit | 0
nitroglycerin infusion | 0
furosemide | 0
calcium channel blockers | 0
telmisartan | 0
normal lipid profile | 0
normal thyroid profile | 0
electroencephalography diffuse theta/delta slowing | 0
electroencephalography bilateral temporal–occipital epileptiform discharges | 0
normal electrocardiogram | 0
normal echocardiogram | 0
normal ultrasound abdomen | 0
normal renal artery doppler | 0
normal neck vessel doppler | 0
reduced shortness of breath | 120
regaining vision completely | 120
blood pressure 160/90 mmHg on day 4 | 96
telmisartan 40 mg once daily | 96
cilnidipine 10 mg BID | 96
hydrochlorothiazide 12.5 mg once daily | 96
persistently high blood pressure | 96
anxiety | 96
metoprolol 25 mg BID added | 96
blood pressure increased to 180/100 mmHg | 96
paradoxical blood pressure increase | 96
serum cortisol normal | 96
parathormone normal | 96
calcium normal | 96
phosphorus normal | 96
urine VMA normal | 96
urine metanephrine elevated | 96
plasma metanephrine elevated | 96
CECT abdomen showing retroperitoneal mass | 96
PET scan no metastasis | 96
started on phenoxybenzamine | 96
other antihypertensives | 96
blood pressure normalized | 96
surgical resection of tumor | 168
biopsy confirmed neuroendocrine tumor | 168
discharged in stable condition | 168
normal blood pressure | 168
