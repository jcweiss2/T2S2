born | -2800
caesarean section | -2800
birth weight 2100 g | -2800
birth length 48 cm | -2800
prominent forehead | -2800
relative macrocephaly | -2800
limb asymmetry | -2800
5th finger clinodactyly of both hands | -2800
2/3 toe syndactyly of both legs feet | -2800
genetic examination | -16
hypomethylation of the 11p15 region of the paternal chromosome | -16
diagnosis of SRS | -16
delayed motor development | -14
walked independently | -14
hepatic dysfunction | -14
increased concentration of alanine aminotransferase | -14
increased concentration of aspartate aminotransferase | -14
increased creatine kinase level | -14
diagnosis of Duchenne muscular dystrophy | -14
genetic test | -9
mutation of the maternal DMD gene | -9
exon deletion 49–50 | -9
corticosteroids treatment | -6
prednisone treatment | -6
deflazacort treatment | -4
G-CSF treatment | -4
sepsis | -4
hypoglycaemia | -4
neurological symptoms | -4
glucose level of 14 mg/dl | -4
urological care | -4
hypospadias | -4
cardiological diagnostics | -2
episodes of sinus tachycardia | -2
heart murmur | -2
propranolol treatment | -2
growth hormone deficiency | -1
rhGH treatment | 0
height 115.9 cm | 0
weight 19.9 kg | 0
body mass index 14.8 kg/m2 | 0
target height 182.5 cm | 0
height velocity 4.3 cm/year | 0
glucose and insulin levels in oral glucose tolerance test | 0
IGF-1 and IGFBP-3 concentrations | 0
MRI of the hypothalamic-pituitary region | 0
transparent septum cyst | 0
rhGH therapy started | 0
height velocity increased | 3
height 118.6 cm | 6
height SDS –2.97 | 6
BMI 16.6 kg/m2 | 6
SDS-BMI –0.2 | 6
IGF-1 294 ng/ml | 6
IGFBP-3 5.76 µg/ml | 6
HbA1c 6.6% | 6
rhGH dose reduced | 6
behavioural treatment with lifestyle modification | 6
weight gain | 6
impaired glucose tolerance | 12
insulin resistance | 12
HOMA-IR 9.66 | 12
distance covered in 6MWT decreased | 12
abnormal gait | 12
rhGH therapy discontinued | 18
densitometry performed | 18
body mass composition examined | 18
bone density test of the lumbar spine | 18
Z-score –2.2 | 18