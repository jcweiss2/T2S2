61 years old | 0
female | 0
breathing difficulties | -48
vomiting | -48
diarrhea | -48
right hemithoracic pain | -48
arterial hypertension | -672
hypercholesterolemia | -672
arthritis | -672
type 2 diabetes | -672
allergy to molds | -672
metformin | -672
co-lisinopril | -672
tramadol | -672
atorvastatin | -672
allopurinol | -672
ranitidine | -672
quinine sulfate | -672
naproxen | -240
restless | 0
pale | 0
hypotensive | 0
sinus tachycardia | 0
marbled legs | 0
marbled thorax | 0
thirst | 0
admitted to ICU | 0
fluid resuscitation | 0
central venous pressure | 0
ScVO2 | 0
low urine output | 0
bradycardic | 2
cardiac arrest | 2
multiple organ failure | 2
respiratory failure | 2
renal failure | 2
liver failure | 2
coagulopathy | 2
inotropes | 2
broad-spectrum antibiotics | 2
amoxicillin-clavulanic acid | 2
amikacin | 2
meropenem | 2
vancomycin | 2
fluconazole | 2
SOFA score | 2
APACHE II score | 2
marbled skin pattern | 0
petechial lesions | 6
erythematous and bullous eruptions | 30
Nikolsky sign | 30
skin biopsy | 30
muscle biopsy | 30
extensive epidermal necrosis | 30
necrosis of striated muscle fibers | 30
necrosis of smooth muscle fibers | 30
elevated uric acid | 0
elevated creatine phosphokinase | 0
elevated C-reactive protein | 0
elevated D-Dimers | 0
lymphocyte transformation test | 24
discontinued naproxen | 24
intravenous methylprednisolone | 24
died | 48