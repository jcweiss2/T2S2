60 years old | 0
male | 0
motor-vehicle accident | -144
right side rib fractures | -144
bilateral pneumothorax | -144
left hip dislocation | -144
fractures of spinous processes of 5th to 8th thoracic vertebrae | -144
obese | 0
BMI 39 kg/m2 | 0
quit smoking | -105600
left lower lobectomy | -105600
carcinoid | -105600
initial regional hospital attendance | -144
thoracic cavity drained | -144
hip dislocation reduced under general anaesthesia | -144
mechanical ventilation dependence | -144
transferred to ICU | -96
respiratory insufficiency | -96
haemodynamic instability | -96
acute renal failure | -96
haemodialysis | -96
massive SE of face, neck, thoracic and abdominal wall | 0
CT scans showing persistent bilateral pneumothorax | 0
pneumomediastinum | 0
pneumoperitoneum | 0
subcutaneous emphysema extending to the pelvis | 0
thoracic drains replaced | 0
continuous venovenous haemodiafiltration initiated | 0
sepsis | 0
multi-resistant Acinetobacter baumanii isolated | 0
bilevel positive airway pressure (BPAP) mechanical ventilation | 0
high inspiratory airway pressure (Pinsp 30 mbar) | 0
high positive end-expiratory pressure (PEEP 10 mbar) | 0
low dynamic compliance (Cdyn 33–40 mL/mbar) | 0
respiratory status deterioration | 120
high inspired oxygen fraction (FiO2 100%) required | 120
control CT confirming thoracic drains position | 120
persistent massive SE | 120
surgical decompression | 120
subclavicular blowhole incisions | 120
NPWT dressing applied | 120
regression of SE | 132
improvement in ventilatory parameters | 132
transition to pressure support mode (PSV) | 132
NPWT dressing removed | 192
wounds sutured | 192
surgical tracheostomy performed | 192
weaned off ventilator | 192
renal function improved | 192
recovery | 192
