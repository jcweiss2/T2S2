72 years old | 0
female | 0
urinary incontinence | -672
ground-level fall | -672
right frontal meningioma | -672
dexamethasone | -672
neurosurgery | -672
outpatient surgery | -672
brain mass resection | -672
dyspnea | -72
nonproductive cough | -72
chest pain | -72
generalized weakness | -72
admitted to the hospital | 0
crackles in the right lung base | 0
consolidation in the right lung base | 0
elevated white blood cell counts | 0
elevated neutrophils | 0
thrombocytopenia | 0
normal renal function | 0
community-acquired pneumonia | 0
intravenous ceftriaxone | 0
azithromycin | 0
discontinued dexamethasone | -72
restarted on dexamethasone | 0
continued chest pain | 168
productive cough | 168
hemoptysis | 168
cavitary lesion | 168
computer tomography scan | 168
cavitary mass in the right middle lobe | 168
sputum samples for acid fast bacilli stain and culture | 168
negative acid fast bacilli stain and culture | 168
indeterminate serum QuantiFERON gold test | 168
negative repeat serum QuantiFERON gold test | 168
negative serum Aspergillus antigen enzyme immunoassay | 168
broadened antibiotic treatment | 168
vancomycin | 168
piperacillin-tazobactam | 168
large right-sided hydropneumothorax | 240
chest tube placement | 240
resolved pneumothorax | 240
pulmonary consult | 240
diagnostic bronchoscopy | 240
tissue sampling | 240
bronchoalveolar lavage | 240
negative AFB stain and culture | 240
grew Streptococcus viridians | 240
grew A. fumigatus | 240
cytology revealed acute-angle hyphae septate | 240
consistent with A. fumigatus | 240
started on voriconazole | 240
switched to isavuconazole | 288
thrombocytopenia | 288
rash | 288
continued pleural leak | 288
persistent and progressive pneumothorax | 288
prolonged ileus | 288
worsening renal function | 288
cardiothoracic surgery consult | 288
evaluation for lobectomy | 288
declined surgical intervention | 288
severe septic shock | 336
multiorgan failure | 336
died | 336