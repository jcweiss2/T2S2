66 years old | 0
morbid obesity | 0
hypertension | 0
hyperlipidemia | 0
non-insulin dependent diabetes mellitus | 0
coronary artery disease | 0
admitted to the hospital | 0
sepsis | 0
lower extremity ulceration | 0
osteomyelitis | 0
contacted family members | -336
immobilized | -336
collapsed floor | -336
without access to hydration | -336
squalid living condition | -336
refused outside assistance | -336
requested medical attention | -336
transported by emergency medical services | -336
anxious | 0
temperature 99.8o F | 0
pulse 109 beats per minute | 0
blood pressure 128/60 mm Hg | 0
respiratory rate 18 breaths per minute |## 数据结构：堆的应用
