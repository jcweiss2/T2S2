18 years old | 0
female | 0
SLE | 0
stage IV lupus nephritis | 0
prior stroke | 0
intravenous drug use | 0
cardiogenic shock | 0
mental status changes | 0
elevated jugular venous pressure | 0
prominent v wave | 0
fever | 0
blood pressure 95/66 mm Hg | 0
heart rate 94 beats/min | 0
hemoglobin 10.3 g/dL | 0
white blood cell count 18.9 × 10^9/L | 0
platelet count 64 × 10^9/L | 0
international normalized ratio 3.6 | 0
creatinine level 1.7 mg/dL | 0
narcotics positive | 0
cannabis positive | 0
negative antiphospholipid serology | 0
negative blood cultures | 0
mitral valve prosthesis dehiscence | 0
severe mitral regurgitation | 0
intervalvular fibrosa dehiscence | 0
cavity at the intervalvular fibrosa | 0
multiloculations | 0
bland fibrin thrombus and fibrous tissue with mild chronic inflammation | 0
destruction of the valves and the intervalvular fibrosa | 0
extensive reconstruction of the fibrous skeleton of the heart and atria | 0
mitral valve annulus reconstruction | 0
33-mm bioprosthesis | 0
bovine pericardium patch | 0
well-seated mitral valve bioprosthesis | 0
mean gradient 3 mm Hg | 0
no regurgitation | 0
left ventricular ejection fraction 25% | 0
sluggish flow in the left atrium | 0
extracorporeal membrane oxygenation | 0
multiple blood product transfusions | 0
layered thrombus in the left atrium | 5
surgical clot removal | 5
thrombus reaccumulation | 5
withdrawal of extracorporeal membrane oxygenation | 5
death | 5