52 years old | 0
woman | 0
presented with worsening shortness of breath | 0
treated as exacerbation of heart failure | 0
echocardiogram demonstrated 5.4 cm aortic root dilated ascending aorta | 0
bicuspid aortic valve | 0
moderate mixed aortic valve disease | 0
mild mitral regurgitation | 0
no prior medical history except penicillin allergy | 0
no known family history of aortopathy | 0
regular smoker | 0
denied illicit drug use | 0
Bentall’s procedure using 27 mm bio-integral valve aortic bio-conduit | -0
mitral valve annuloplasty | -0
no complications in postoperative period | -0
sternotomy wound healed | -8760
re-presented to cardiothoracic clinic with discharging sternal sinus | -30240
secondary to infection of sternal wires with Staphylococcus aureus (methicillin-sensitive) | -30240
chronic sternal osteomyelitis | -30240
sternal wound debridement | -30240
removal of superior infected sternal wires | -30240
antibiotics | -30240
negative pressure wound therapy | -30240
conventional dressings | -30240
co-trimoxazole advised | -30240
re-presented acutely to hospital complaining of chest pain | 0
dizziness | 0
multiple episodes of active bleeding from sternal wound | 0
hemodynamically stable | 0
swollen chronically infected sinus over previous sternotomy scar | 0
hematoma | 0
anemia | 0
hemoglobin of 95 g/L | 0
albumin 27 g/L | 0
raised inflammatory markers | 0
white cell count of 9 × 109/L | 0
platelet count of 613 × 109/L | 0
C-reactive protein 24 mg/L | 0
CT angiogram demonstrated pseudoaneurysm at distal anastomosis of ascending graft | 0
rim-enhancing soft tissue surrounding aorta | 0
sternal wound infection extended to ascending aortic bio graft forming pseudoaneurysm | 0
aorto-cutaneous fistula through osteomyelitic sternum and infected skin sinus | 0
discussed at aortic multidisciplinary team meeting | 0
definitive open repair contemplated | 0
radial surgical debridement | 0
removal of infective foreign material | 0
re-do Bentall’s proximal arch replacement | 0
or without removal of mitral ring under deep hypothermic circulatory arrest | 0
deemed high-risk | 0
not fit to tolerate re-do Bentall’s operation | 0
malnourishment | 0
low body mass index | 0
significant smoking history | 0
multiple psychosocial issues including nonadherence to medical advice | 0
consensus to exclude pseudoaneurysm with endovascular stent graft | 0
manage risk for exsanguination from repeat aorto-cutaneous fistula bleeding | 0
endovascular treatment intended as temporizing measure | 0
optimize patient before major cardiac revision surgery | 0
allow time for long-term antibiotics to suppress graft infection | 0
pseudoaneurysm located at distal anastomosis of ascending graft | 0
ascending graft proximal to pseudoaneurysm was 43 mm | 0
aorta distal to pseudoaneurysm was 42 × 38 mm | 0
distance between coronary arteries and proximal end of pseudoaneurysm was 53 mm | 0
distance from proximal end of brachiocephalic trunk to distal end of pseudoaneurysm was 30 mm | 0
46 mm × 46 mm 55-mm Valiant Navion stent graft selected | 0
flushed with rifampicin before insertion | 0
percutaneous femoral access used | 0
stent deployed under rapid pacing to 200 bpm | 0
dilated after placement | 0
completion angiogram confirmed exclusion of pseudoaneurysm | 0
CT angiogram performed 48 hours later demonstrated successful covering | 48
infectious disease team advised long-term antibiotics | 48
discharged 48 hours later | 48
follow-up plan included cardiothoracic and infectious disease clinic appointments at 2 weeks | 48
vascular clinic appointment at 6 weeks | 48
repeat CT angiography prior | 48
regular community nurse visits | 48
wound dressing changes | 48
regular dietician assessments | 48
regular blood tests | 48
red blood cell transfusions | 48
iron infusions | 48
psychological input | 48
psychiatric input | 48
social work input | 48
regular infectious disease follow-up | 48
community pharmacist visits | 48
re-presented acutely in septic shock | 1080
blood pressure 75/51 mm Hg | 1080
heart rate 127 | 1080
respiratory rate 27 | 1080
temperature 40 °C | 1080
white cell count 19.7 × 109/L | 1080
C-reactive protein 160 mg/L | 1080
lactate 2.2 mmol/L | 1080
CT angiogram demonstrated new infected pseudoaneurysm | 1080
intact ascending graft proximal to pseudoaneurysm | 1080
multidisciplinary meeting held | 1080
consensus to perform thoracic endovascular aortic repair | 1080
extension of graft to just distal to coronary arteries | 1080
intraoperative transesophageal echocardiogram performed | 1080
no signs of vegetation’s of aortic valve | 1080
second ascending stent graft performed percutaneously | 1080
SAFARI wire placed into left ventricle | 1080
pigtail catheter placed above aortic valve | 1080
Medtronic Valiant Navion 46 × 46 × 93 mm stent graft | 1080
flushed with rifampicin | 1080
deployed under rapid cardiac pacing | 1080
completion angiogram confirmed satisfactory stent position | 1080
CT angiogram day 6 after surgery demonstrated pseudoaneurysm covered | 1128
multiple admissions for red blood cell transfusions | 1128
iron infusions due to blood loss through sternotomy wound | 1128
regular dietician input | 1128
slow improvements in nutritional status | 1128
specialist cardiac input obtained | 1128
assessed for second opinion on surgical management | 1128
potential operative plan made | 1128
inpatient mortality risk over 50% | 1128
re-presented with sternal wound bleeding | 2160
hemoptysis | 2160
dizziness | 2160
hemoglobin 73 g/dL | 2160
required transfusion | 2160
CT angiography demonstrated extension of pseudoaneurysm superior to stent graft | 2160
up to level of brachiocephalic trunk | 2160
empyema | 2160
pseudoaneurysm compressing carina | 2160
abscess developing between airways | 2160
endovascular treatment as bridging therapy | 2160
patient decision not to proceed with further surgery | 2160
declined antibiotic therapy | 2160
palliated | 2160
died 7 months after first endovascular stent graft | 2160
no prior medical history except penicillin allergy |DONE
