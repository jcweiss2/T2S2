32 years old | 0
female | 0
no significant past medical history | 0
referred to a dermatologist | -72
diagnosed with Nicolau syndrome | -72
severe pain | -72
redness | -72
swelling | -72
left buttock | -72
surrounding back area | -72
intramuscular injection of methocarbamol | -72
musculoskeletal pain | -72
motor vehicle accident | -72
anxious | 0
severe distress | 0
discolored | 0
dusky appearance | 0
marked erythema | 0
edema | 0
necrotic tissue | 0
black | 0
eschar-like | 0
hypotension | 0
tachycardia | 0
leukocytosis | 0
left shift | 0
inflammatory response | 0
renal function normal | 0
hepatic function normal | 0
ultrasound | 0
computed tomography (CT) | 0
massive tissue necrosis | 0
impairment of peripheral perfusion | 0
aggressive resuscitation efforts | 0
broad-spectrum antibiotic therapy | 0
hemodynamic instability | 0
cardiac shock | 0
death | 144
autopsy | 144
external examination | 144
internal examination | 144
tissue samples | 144
histopathological analysis | 144
toxicological analysis | 144
mild fatty changes | 144
acute tubular necrosis | 144
acute kidney injury | 144
brain tissue normal | 144
therapeutic levels of metacarbamol | 144
skin integrity | -72
trauma | -72
infection | -72
pressure | -72
chronic diseases | -72
discomfort | -72
pain | -72
quality of life | -72
prevention | -72
injection technique | -72
patient-specific factors | -72
substance injected | -72
vasoconstriction | -72
tissue ischemia | -72
cytotoxic effect | -72
improper injection technique | -72
local ischemia | -72
necrosis | -72
compromised local circulation | -72
diabetes | -72
immunosuppression | -72
sepsis | 0
wound care | 0
debridement of necrotic tissue | 0
dressings | 0
surgical intervention | 0
skin grafting | 0
flap reconstruction | 0
pain control | 0
infection prevention | 0
discontinuing methocarbamol | 0