28 years old | 0
male | 0
admitted to a local hospital | 0
BMI of 70.1 kg/m2 | 0
gained approximately 80 kg in weight | -8760
worsening edema in both lower legs | -168
dyspnea on exertion | -168
transferred to our hospital | 0
respiratory failure | 0
super-obesity | 0
supplemental oxygen via face mask at 3 L/min | 0
arterial blood gas | 0
pH of 7.21 | 0
PaCO2 78 mmHg | 0
PaO2 105 mmHg | 0
HCO3− 30.7 mmol/L | 0
provisional diagnosis of acute cardiac failure | 0
obesity hypoventilation syndrome | 0
clinical examination | 0
chest X-ray | 0
elevated BNP level | 0
noninvasive positive-pressure ventilation therapy | 0
furosemide | 0
developed worsening hypercapnia | 24
impaired consciousness | 24
admitted to the ICU | 24
physical examination upon admission to the ICU | 24
GCS 14 | 24
blood pressure 128/74 mmHg | 24
heart rate 90 bpm | 24
SpO2 90% | 24
FIO2 0.45 | 24
expiratory positive airway pressure 6 cmH2O | 24
inspiratory positive airway pressure 18 cmH2O | 24
facial edema | 24
leg edema | 24
wheezing on expiration | 24
no heart murmur | 24
blood test | 24
mildly elevated inflammatory response | 24
elevated BNP level | 24
arterial blood gas analysis | 24
pH 7.236 | 24
PaCO2 94 mmHg | 24
PaO2 78 mmHg | 24
HCO3 39.1 mmol/L | 24
lactate 4.9 mmol/L | 24
respiratory acidosis | 24
chest radiograph | 24
marked cardiomegaly | 24
cardiothoracic ratio 66.2% | 24
enhanced pulmonary vasculature | 24
electrocardiogram | 24
heart rate 80 bpm | 24
sinus rhythm | 24
chest computed tomography | 24
no infiltrative shadow | 24
no pleural effusion | 24
no atelectasis | 24
contrast-enhanced CT | 24
no thrombus in the pulmonary artery | 24
intubated | 24
ventilator set to assist/control mode | 24
FIO2 0.6 | 24
ventilation frequency 16/min | 24
pressure control 16 cmH2O | 24
positive end-expiratory pressure 10 cmH2O | 24
PAC placed | 24
mean pulmonary artery pressure 49 mmHg | 24
central venous pressure 10 mmHg | 24
pulmonary artery wedge pressure 18 mmHg | 24
cardiac output 7.8 L/min | 24
cardiac index 2.8 L/min/m2 | 24
diagnosis of pulmonary hypertension | 24
transoesophageal echocardiography | 120
no abnormal left ventricular wall motion | 120
no significant valvular disease | 120
no patent foramen ovale | 120
positional changes | 120
tracheal aspiration | 120
systolic pulmonary artery pressure 80–90 mmHg | 120
systolic pressure 60–70 mmHg | 120
SpO2 <80% | 120
deep sedation management | 120
continuous administration of muscle relaxants | 120
catheter removed | 240
mean pulmonary artery pressure 31 mmHg | 240
rapid decrease in blood pressure | 240
SpO2 decrease | 240
suspicion of catheter infection | 240
septic shock | 240
noradrenaline continued | 240
muscle relaxants discontinued | 240
spontaneous respiration restored | 240
condition gradually improved | 240
hemodynamic stability | 360
NAd administration discontinued | 360
extubated | 552
discharged from the ICU | 672
discharged from the hospital | 2040
