52 years old | 0\
male | 0\
body mass index 23.6 kg/m2 | 0\
no comorbidities | 0\
referred to our institution for surgical consultation | 0\
chronic post-bariatric gastrocutaneous fistula | 0\
open modified Scopinaro procedure | -7200\
initial weight 216 kg | -7200\
BMI 57.4 kg/m2 | -7200\
weight reganance | -2400\
incisional hernia | -2400\
bariatric revisional surgery and hernia repair | -2400\
weight 170 kg | -2400\
BMI 45.1 | -2400\
gastric pouch leak | -2400\
multiple intra-abdominal collections | -2400\
sepsis | -2400\
conservative management with open abdomen | -2400\
negative wound pressure therapy | -2400\
parenteral nutrition | -2400\
intravenous antibiotics | -2400\
epithelized gastrocutaneous fistula | -1200\
controlled but persistent drainage | -1200\
proximal edge of his planned ventral hernia | -1200\
upper endoscopy | -1200\
fistulous orifice at the proximal edge of the vertical staple line | -1200\
just below the esophagogastric junction | -1200\
measuring approximately 8 mm | -1200\
extraluminal extravasation | -1200\
recurrent left subphrenic abscess | -1200\
endoscopic treatment | -1200\
poor nutritional status | -1200\
hostile abdomen | -1200\
multiple attempts at fistula closure | -1200\
argon plasma coagulation | -1200\
internal and external drainages | -1200\
clipping | -1200\
fibrin sealants | -1200\
e-vac therapy | -1200\
stenting | -1200\
multidisciplinary team discussion | -24\
decision to proceed with an innovative endoscopic technique | -24\
placement of a CSDO across the fistula orifice | -24\
Occlutech muscular VSD occluder | -24\
long funnel-shaped aspect of the defect | -24\
similar to a ventricular septal defect | -24\
braided nitinol disc | -24\
adapt to the shape of the defect | -24\
achieve immediate closure | -24\
patch material | -24\
matrix for subsequent tissue ingrowth and granulation | -24\
contribute to fistula closure | -24\
procedure performed in the catheterization laboratory | 0\
intravenous sedation | 0\
topic anesthesia | 0\
fistula cannulated from the esophagus | 0\
biliary stent deployment system | 0\
direct endoscopic guidance | 0\
extraluminal leakage | 0\
documented by contrast injection | 0\
Amplatz extra stiff guidewire | 0\
inserted through the fistula orifice | 0\
adequate position confirmed by fluoroscopy | 0\
delivery system introduced over the guidewire | 0\
CSDO deployed under endoscopic and fluoroscopic guidance | 0\
no immediate adverse events | 0\
contrast study after the CSDO placement | 0\
no extravasation of contrast material through the device | 0\
restricted oral intake for 24 h | 24\
liquid diet for 10 days | 240\
advanced to a regular diet on day 12 | 288\
10–15cc remaining daily drainage through the pigtail drain | 288\
pigtail drain positioned at his left subphrenic abscess | 288\
pigtail was accidentally displaced | 504\
systemic signs of sepsis | 504\
computed tomography and fluoroscopy | 504\
recurrence of the abscess | 504\
partial dislodgment of the 8-mm mVSD CSDO | 504\
device probably tore the friable tissue around the fistulous orifice | 504\
got stuck in the tunnel-shaped tract | 504\
not possible to see or snare the device by endoscopic view | 504\
second attempt with an oversized disc | 504\
Occlutech Figulla Flex II UNI 24-mm | 504\
sealing the fistulous orifice with the former device positioned between the two discs of the new one | 504\
6-month clinical and imaging follow-up | 2160\
upper endoscopy and contrast-enhanced CT scan | 2160\
device already engrafted | 2160\
significant reduction of the chronic abscess | 2160\
no signs of fistula recurrence | 2160\
pigtail was maintained in the subphrenic space | 2160\
monitor any sign of fistula recurrence | 2160\
occasionally drained debris from the chronic abscess | 2160\
finally removed after the follow-up imaging | 2160\
no drainage was observed from its insertion orifice or the previous cutaneous fistulous tract | 2160