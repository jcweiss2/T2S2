37 years old | 0
    man | 0
    admitted | 0
    fever | -96
    headache | -96
    myalgia | -96
    epigastralgia | -96
    nausea | -96
    diarrhoea | -96
    active smoking | 0
    no splenic disorders | 0
    no alcohol excess | 0
    no immunocompromised | 0
    no cardiac symptoms | 0
    dog bite (right hand) | -120
    temperature 38.2°C | 0
    heart rate 130 b.p.m. | 0
    blood pressure 118/72 mmHg | 0
    pulse oxygen saturation 100% | 0
    bite wound (right hand) | 0
    no rash | 0
    no sign of cellulitis | 0
    no soft tissue necrosis | 0
    C-reactive protein 417 mg/L | 0
    white blood cell count 9.45 G/L | 0
    neutrophils 91% | 0
    lymphocytes 3.5% | 0
    procalcitonin 8.42 μg/L | 0
    thrombocytopaenia (platelets 29 G/L) | 0
    acute kidney injury (creatinine 189 μmol/L) | 0
    abnormal liver enzymes (AST ×2, ALT ×3) | 0
    elevated high sensitivity-troponin T (peak 1129 ng/L) | 0
    N-terminal brain natriuretic peptide 1127 pg/mL | 0
    12-lead electrocardiogram (diffuse ST-segment elevation) | 0
    micro-Q waves (inferior and lateral leads) | 0
    transthoracic echocardiography (mild global LV hypokinesia) | 0
    LV ejection fraction 42% | 0
    preserved right ventricular function | 0
    no pericardial effusion | 0
    blood cultures drawn | 0
    parenteral cefotaxime (3 g/day) | 0
    Capnocytophaga canimorsus identified (blood cultures) | 47
    cefotaxime changed to amoxicillin (3 g/day for 7 days) | 47
    recovery of biological markers | 47
    coronary computed tomography angiography (normal coronary arteries) | 47
    cardiovascular magnetic resonance (Day 5) | 120
    non-dilated LV (87 mL/m²) | 120
    LV ejection fraction 56% | 120
    focal areas of subepicardial oedema (LV inferolateral wall) | 120
    early hyper-enhancement (LV inferolateral wall) | 120
    late gadolinium-enhancement (subepicardium of inferolateral and anterolateral walls) | 120
    increased T2 time (oedema) | 120
    increased extracellular volume (interstitial space) | 120
    no endomyocardial biopsy performed | 120
    no haemodynamic deterioration | 120
    no heart failure | 120
    no arrhythmias | 120
    Gram-negative rod bacteria covered with antibiotics | 120
    discharged | 168
    remains well at 1 year | 168
    no further symptoms | 168