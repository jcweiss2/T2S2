68 years old | 0
male | 0
admitted to the hospital | 0
decompressive laminectomy | -720
fatigue | -72
dyspnea | -72
cough | -72
chills | -72
fever (Tmax 101oF) | -72
hematuria | -72
hypoxia (SpO2 high 80s) | -72
tested positive for COVID-19 | -72
acute kidney injury | -72
started on hydroxychloroquine | 0
started on azithromycin | 0
progressive dyspnea | 24
hypoxia | 24
severe hypotension (blood pressures 60/40) | 24
intubated | 24
transitioned to intensive care unit | 24
increasing pressure requirements | 72
persistent fevers (Tmax 103.5oF) | 72
hypotension | 72
given Tocilizumab | 72
stabilized hemodynamically | 72
self-extubation | 168
placed on supplemental oxygen | 168
discharged to inpatient rehabilitation | 408
negative COVID-19 test result | 408
deep venous thrombosis | 408
transitioned to Enoxaparin sodium | 408
acute right knee pain | 600
limited range of motion | 600
could not bear weight | 600
swollen knee | 600
painful knee | 600
low-grade fever (100.8oF) | 600
warm knee | 600
erythematous knee | 600
knee arthrocentesis | 600
synovial fluid drained | 600
admitted back to the hospital | 648
started on Vancomycin | 648
started on Zosyn | 648
high white blood cell count | 648
high lymphocytes | 648
low monocytes | 648
elevated IL markers | 648
cloudy yellow synovial fluid | 648
neutrophilic predominance (87%) | 648
no crystals | 648
no bacterial culture growth | 648
transitioned to oral cephalexin | 648
started on Prednisone taper | 648
transferred back to inpatient rehabilitation | 648
transitioned to Apixaban | 648
discharged home | 1176
