18 years old | 0
female | 0
admitted to the hospital | 0
right lower quadrant abdominal pain | -336
nausea | -336
vomiting | -336
anorexia | -336
no fever | -336
eaten decayed wheat | -672
abdominal distension | 0
tenderness in the right lower quadrant | 0
fullness in the right lower quadrant | 0
CT scan of the abdomen and pelvis | 0
obstructing caecal mass | 0
colonoscopy | 24
necrotic caecal mass | 24
biopsies | 24
ulcerations | 48
necrosis | 48
microabscesses | 48
multinucleated giant cells | 48
fungal hyphae | 48
antifungal treatment with amphotericin B | 48
jaundice | 72
high fever | 72
per-rectal bleeding | 72
increased white cell count | 72
eosinophilia | 72
deranged liver function tests | 72
CT scan of the abdomen and pelvis | 72
anterior intra-abdominal collection | 72
right paracolic gutter collection | 72
panniculitis | 72
peritonitis | 72
multiple hypodense lesions in the liver | 72
septic shock | 96
exploratory laparotomy | 96
ileal perforation | 96
extensive white patches over the posterior abdominal wall | 96
small bowel | 96
liver | 96
bowel resection | 96
primary anastomosis | 96
histopathology | 120
fungal hyphae invading the bowel wall | 120
positive periodic acid-Schiff | 120
positive Gomori’s Methenamine Silver stain | 120
Splendore-Hoeppli phenomenon | 120
liver biopsies | 120
Basidiobolus species | 120
Candida | 120
Klebsiella pneumoniae | 120
voriconazole | 144
tigecycline | 144
meropenem | 144
enterocutaneous fistula | 168
vacuum-assisted closure device | 168
total parenteral nutrition | 168
inflammatory markers returned to normal | 240
white cell count returned to normal | 240
liver function tests returned to normal | 240
fever | 288
CT scan of the abdomen and pelvis | 288
enlargement of the right paracolic gutter collection | 288
common hepatic artery aneurysm | 288
large right pleural effusion | 288
ultrasound-guided drainage | 312
embolisation of the common hepatic artery pseudoaneurysm | 312
chest tube insertion | 312
liposomal amphotericin B | 336
posaconazole | 336
seizures | 360
MRI of the brain | 360
diffuse global brain oedema | 360
cortical laminar necrosis | 360
meningoencephalitis | 360
intubation | 384
high doses of inotropes | 384
multiple bilateral lung abscesses | 408
septic shock | 408
death | 432