spontaneous onset of labor | -1
fetal distress noted on cardiotocography | -0.5
ventouse-assisted delivery | 0
baby born with birth weight of 3940 grams | 0
immediate resuscitation with mask ventilation | 0
intubated at 8 minutes of age | 0.13
transferred to NICU | 0.13
commenced empirical antibiotics | 0.13
supported with SIPPV | 0.13
weaned from respiratory support | 12
extubated at 13.5 hours of age | 13.5
neutropenia with significant left shift | 18
elevated inflammatory markers | 18
lumbar puncture performed | 23
placental surface eSwab demonstrated light pure growth of an organism | 23
Gram-negative diplococci identified | 23
MALDI-TOF mass spectrometry identified Neisseria meningitidis | 23
molecular testing confirmed detection of meningococcus genogroup W CC11 | 23
blood cultures taken from newborn were negative | 0.48
heel-prick blood detected presence of N. meningitidis genogroup W DNA | 5.5
benzylpenicillin dosage decreased | 24
benzylpenicillin changed to cefotaxime | 24
completed 5-day course of β-lactam therapy | 120
maternal bloods showed elevated leucocyte count | -2.5
maternal bloods showed neutrophil count of 18.1×10^9/L | -2.5
mother remained well after birth | 0
baby remained well and discharged from NICU | 192
contact tracing identified staff members and family at risk | 192
chemoprophylaxis with ciprofloxacin provided | 192
vaccination with quadrivalent conjugate meningococcal vaccine provided | 192
placenta histopathology revealed acute funisitis and chorioamnionitis | 24
no shortness of breath | 0
denies chest pain | 0 
baby required immediate resuscitation | 0 
baby had poor respiratory effort | 0 
baby was intubated | 0.13 
baby was supported with SIPPV with minimal pressures | 0.13 
baby had no additional oxygen requirement | 0.13 
baby was weaned from respiratory support | 12 
baby was extubated | 13.5 
inflammatory markers were elevated | 18 
C-reactive protein was elevated | 18 
procalcitonin was elevated | 18 
lumbar puncture was negative for pathogens | 23 
lumbar puncture was negative for meningococcus | 23 
placental surface eSwab was performed | 23 
Gram-negative diplococci were identified | 23 
Neisseria meningitidis was identified | 23 
molecular testing was performed | 23 
molecular testing confirmed detection of meningococcus | 23 
blood cultures were taken from newborn | 0.48 
blood cultures were negative | 0.48 
heel-prick blood was taken | 5.5 
heel-prick blood detected presence of N. meningitidis | 5.5 
benzylpenicillin dosage was decreased | 24 
benzylpenicillin was changed to cefotaxime | 24 
β-lactam therapy was completed | 120 
maternal bloods were taken | -2.5 
maternal bloods showed elevated leucocyte count | -2.5 
maternal bloods showed neutrophil count | -2.5 
mother remained well | 0 
baby remained well | 192 
baby was discharged from NICU | 192 
contact tracing was performed | 192 
chemoprophylaxis was provided | 192 
vaccination was provided | 192 
placenta histopathology was performed | 24 
placenta histopathology revealed acute funisitis | 24 
placenta histopathology revealed chorioamnionitis | 24 
no shortness of breath | 0 
denies chest pain | 0 
baby required immediate resuscitation | 0 
baby had poor respiratory effort | 0 
baby was intubated | 0.13 
baby was supported with SIPPV | 0.13 
baby had no additional oxygen requirement | 0.13 
baby was weaned from respiratory support | 12 
baby was extubated | 13.5 
inflammatory markers were elevated | 18 
C-reactive protein was elevated | 18 
procalcitonin was elevated | 18 
lumbar puncture was negative for pathogens | 23 
lumbar puncture was negative for meningococcus | 23 
placental surface eSwab was performed | 23 
Gram-negative diplococci were identified | 23 
Neisseria meningitidis was identified | 23 
molecular testing was performed | 23 
molecular testing confirmed detection of meningococcus | 23 
blood cultures were taken from newborn | 0.48 
blood cultures were negative | 0.48 
heel-prick blood was taken | 5.5 
heel-prick blood detected presence of N. meningitidis | 5.5 
benzylpenicillin dosage was decreased | 24 
benzylpenicillin was changed to cefotaxime | 24 
β-lactam therapy was completed | 120 
maternal bloods were taken | -2.5 
maternal bloods showed elevated leucocyte count | -2.5 
maternal bloods showed neutrophil count | -2.5 
mother remained well | 0 
baby remained well | 192 
baby was discharged from NICU | 192 
contact tracing was performed | 192 
chemoprophylaxis was provided | 192 
vaccination was provided | 192 
placenta histopathology was performed | 24 
placenta histopathology revealed acute funisitis | 24 
placenta histopathology revealed chorioamnionitis | 24 
baby had neutropenia | 18 
baby had significant left shift | 18 
baby had elevated CRP | 18 
baby had elevated procalcitonin | 18 
baby had normal cell count | 23 
baby had negative lumbar puncture | 23 
baby had negative blood cultures | 0.48 
baby had positive heel-prick blood | 5.5 
mother had elevated leucocyte count | -2.5 
mother had elevated neutrophil count | -2.5 
mother had no symptoms | -2.5 
baby was treated with gentamicin | 0.13 
baby was treated with benzylpenicillin | 0.13 
baby was treated with cefotaxime | 24 
baby completed β-lactam therapy | 120 
staff members were at risk | 192 
family members were at risk | 192 
chemoprophylaxis was provided to staff members | 192 
chemoprophylaxis was provided to family members | 192 
vaccination was provided to staff members | 192 
vaccination was provided to family members | 192 
Neisseria meningitidis was detected in placental surface eSwab | 23 
Neisseria meningitidis was detected in heel-prick blood | 5.5 
Neisseria meningitidis was identified by MALDI-TOF | 23 
Neisseria meningitidis was identified by molecular testing | 23 
Neisseria meningitidis was serogroup W | 23 
Neisseria meningitidis was clonal complex 11 | 23 
baby had funisitis | 24 
baby had chorioamnionitis | 24 
mother had no symptoms after birth | 0 
baby had no symptoms after discharge | 192 
baby was discharged from NICU | 192 
contact tracing was performed | 192 
chemoprophylaxis was provided | 192 
vaccination was provided | 192 
placenta histopathology was performed | 24 
placenta histopathology revealed acute funisitis | 24 
placenta histopathology revealed chorioamnionitis | 24 
Neisseria meningitidis was detected in placental surface eSwab | 23 
Neisseria meningitidis was detected in heel-prick blood | 5.5 
Neisseria meningitidis was identified by MALDI-TOF | 23 
Neisseria meningitidis was identified by molecular testing | 23 
Neisseria meningitidis was serogroup W | 23 
Neisseria meningitidis was clonal complex 11 | 23 
baby had funisitis | 24 
baby had chorioamnionitis | 24 
mother had no symptoms after birth | 0 
baby had no symptoms after discharge | 192 
baby was treated with gentamicin | 0.13 
baby was treated with benzylpenicillin | 0.13 
baby was treated with cefotaxime | 24 
baby completed β-lactam therapy | 120 
staff members were at risk | 192 
family members were at risk | 192 
chemoprophylaxis was provided to staff members | 192 
chemoprophylaxis was provided to family members | 192 
vaccination was provided to staff members | 192 
vaccination was provided to family members | 192 
Neisseria meningitidis was detected in placental surface eSwab | 23 
Neisseria meningitidis was detected in heel-prick blood | 5.5 
Neisseria meningitidis was identified by MALDI-TOF | 23 
Neisseria meningitidis was identified by molecular testing | 23 
Neisseria meningitidis was serogroup W | 23 
Neisseria meningitidis was clonal complex 11 | 23 
baby had funisitis | 24 
baby had chorioamnionitis | 24 
mother had no symptoms after birth | 0 
baby had no symptoms after discharge | 192 
baby was discharged from NICU | 192 
contact tracing was performed | 192 
chemoprophylaxis was provided | 192 
vaccination was provided | 192 
placenta histopathology was performed | 24 
placenta histopathology revealed acute funisitis | 24 
placenta histopathology revealed chorioamnionitis | 24 
Neisseria meningitidis was detected in placental surface eSwab | 23 
Neisseria meningitidis was detected in heel-prick blood | 5.5 
Neisseria meningitidis was identified by MALDI-TOF | 23 
Neisseria meningitidis was identified by molecular testing | 23 
Neisseria meningitidis was serogroup W | 23 
Neisseria meningitidis was clonal complex 11 | 23 
baby had funisitis | 24 
baby had chorioamnionitis | 24 
mother had no symptoms after birth | 0 
baby had no symptoms after discharge | 192 
baby was treated with gentamicin | 0.13 
baby was treated with benzylpenicillin | 0.13 
baby was treated with cefotaxime | 24 
baby completed β-lactam therapy | 120 
staff members were at risk | 192 
family members were at risk | 192 
chemoprophylaxis was provided to staff members | 192 
chemoprophylaxis was provided to family members | 192 
vaccination was provided to staff members | 192 
vaccination was provided to family members | 192 
Neisseria meningitidis was detected in placental surface eSwab | 23 
Neisseria meningitidis was detected in heel-prick blood | 5.5 
Neisseria meningitidis was identified by MALDI-TOF | 23 
Neisseria meningitidis was identified by molecular testing | 23 
Neisseria meningitidis was serogroup W | 23 
Neisseria meningitidis was clonal complex 11 | 23 
baby had funisitis | 24 
baby had chorioamnionitis | 24 
mother had no symptoms after birth | 0 
baby had no symptoms after discharge | 192 
baby was discharged from NICU | 192 
contact tracing was performed | 192 
chemoprophylaxis was provided | 192 
vaccination was provided | 192 
placenta histopathology was performed | 24 
placenta histopathology revealed acute funisitis | 24 
placenta histopathology revealed chorioamnionitis | 24 
Neisseria meningitidis was detected in placental surface eSwab | 23 
Neisseria meningitidis was detected in heel-prick blood | 5.5 
Neisseria meningitidis was identified by MALDI-TOF | 23 
Neisseria meningitidis was identified by molecular testing | 23 
Neisseria meningitidis was serogroup W | 23 
Neisseria meningitidis was clonal complex 11 | 23 
baby had funisitis | 24 
baby had chorioamnionitis | 24 
mother had no symptoms after birth | 0 
baby had no symptoms after discharge | 192 
baby was treated with gentamicin | 0.13 
baby was treated with benzylpenicillin | 0.13 
baby was treated with cefotaxime | 24 
baby completed β-lactam therapy | 120 
staff members were at risk | 192 
family members were at risk | 192 
chemoprophylaxis was provided to staff members | 192 
chemoprophylaxis was provided to family members | 192 
vaccination was provided to staff members | 192 
vaccination was provided to family members | 192 
Neisseria meningitidis was detected in placental surface eSwab | 23 
Neisseria meningitidis was detected in heel-prick blood | 5.5 
Neisseria meningitidis was identified by MALDI-TOF | 23 
Neisseria meningitidis was identified by molecular testing | 23 
Neisseria meningitidis was serogroup W | 23 
Neisseria meningitidis was clonal complex 11 | 23 
baby had funisitis | 24 
baby had chorioamnionitis | 24 
mother had no symptoms after birth | 0 
baby had no symptoms after discharge | 192 
baby was discharged from NICU | 192 
contact tracing was performed | 192 
chemoprophylaxis was provided | 192 
vaccination was provided | 192 
placenta histopathology was performed | 24 
placenta histopathology revealed acute funisitis | 24 
placenta histopathology revealed chorioamnionitis | 24 
Neisseria meningitidis was detected in placental surface eSwab | 23 
Neisseria meningitidis was detected in heel-prick blood | 5.5 
Neisseria meningitidis was identified by MALDI-TOF | 23 
Neisseria meningitidis was identified by molecular testing | 23 
Neisseria meningitidis was serogroup W | 23 
Neisseria meningitidis was clonal complex 11 | 23 
baby had funisitis | 24 
baby had chorioamnionitis | 24 
mother had no symptoms after birth | 0 
baby had no symptoms after discharge | 192 
baby was treated with gentamicin | 0.13 
baby was treated with benzylpenicillin | 0.13 
baby was treated with cefotaxime | 24 
baby completed β-lactam therapy | 120 
staff members were at risk | 192 
family members were at risk | 192 
chemoprophylaxis was provided to staff members | 192 
chemoprophylaxis was provided to family members | 192 
vaccination was provided to staff members | 192 
vaccination was provided to family members | 192 
Neisseria meningitidis was detected in placental surface eSwab | 23 
Neisseria meningitidis was detected in heel-prick blood | 5.5 
Neisseria meningitidis was identified by MALDI-TOF | 23 
Neisseria meningitidis was identified by molecular testing | 23 
Neisseria meningitidis was serogroup W | 23 
Neisseria meningitidis was clonal complex 11 | 23 
baby had funisitis | 24 
baby had chorioamnionitis | 24 
mother had no symptoms after birth | 0 
baby had no symptoms after discharge | 192 
baby was discharged from NICU | 192 
contact tracing was performed | 192 
chemoprophylaxis was provided | 192 
vaccination was provided | 192 
placenta histopathology was performed | 24 
placenta histopathology revealed acute funisitis | 24 
placenta histopathology revealed chorioamnionitis | 24 
Neisseria meningitidis was detected in placental surface eSwab | 23 
Neisseria meningitidis was detected in heel-prick blood | 5.5 
Neisseria meningitidis was identified by MALDI-TOF | 23 
Neisseria meningitidis was identified by molecular testing | 23 
Neisseria meningitidis was serogroup W | 23 
Neisseria meningitidis was clonal complex 11 | 23 
baby had funisitis | 24 
baby had chorioamnionitis | 24 
mother had no symptoms after birth | 0 
baby had no symptoms after discharge | 192 
baby was treated with gentamicin | 0.13 
baby was treated with benzylpenicillin | 0.13 
baby was treated with cefotaxime | 24 
baby completed β-lactam therapy | 120 
staff members were at risk | 192 
family members were at risk | 192 
chemoprophylaxis was provided to staff members | 192 
chemoprophylaxis was provided to family members | 192 
vaccination was provided to staff members | 192 
vaccination was provided to family members | 192 
Neisseria meningitidis was detected in placental surface eSwab | 23 
Neisseria meningitidis was detected in heel-prick blood | 5.5 
Neisseria meningitidis was identified by MALDI-TOF | 23 
Neisseria meningitidis was identified by molecular testing | 23 
Neisseria meningitidis was serogroup W | 23 
Neisseria meningitidis was clonal complex 11 | 23 
baby had funisitis | 24 
baby had chorioamnionitis | 24 
mother had no symptoms after birth | 0 
baby had no symptoms after discharge | 192 
baby was discharged from NICU | 192 
contact tracing was performed | 192 
chemoprophylaxis was provided | 192 
vaccination was provided | 192 
placenta histopathology was performed | 24 
placenta histopathology revealed acute funisitis | 24 
placenta histopathology revealed chorioamnionitis | 24 
Neisseria meningitidis was detected in placental surface eSwab | 23 
Neisseria meningitidis was detected in heel-prick blood | 5.5 
Neisseria meningitidis was identified by MALDI-TOF | 23 
Neisseria meningitidis was identified by molecular testing | 23 
Neisseria meningitidis was serogroup W | 23 
Neisseria meningitidis was clonal complex 11 | 23 
baby had funisitis | 24 
baby had chorioamnionitis | 24 
mother had no symptoms after birth | 0 
baby had no symptoms after discharge | 192 
baby was treated with gentamicin | 0.13 
baby was treated with benzylpenicillin | 0.13 
baby was treated with cefotaxime | 24 
baby completed β-lactam therapy | 120 
staff members were at risk | 192 
family members were at risk | 192 
chemoprophylaxis was provided to staff members | 192 
chemoprophylaxis was provided to family members | 192 
vaccination was provided to staff members | 192 
vaccination was provided to family members | 192 
Neisseria meningitidis was detected in placental surface eSwab | 23 
Neisseria meningitidis was detected in heel-prick blood | 5.5 
Neisseria meningitidis was identified by MALDI-TOF | 23 
Neisseria meningitidis was identified by molecular testing | 23 
Neisseria meningitidis was serogroup W | 23 
Neisseria meningitidis was clonal complex 11 | 23 
baby had funisitis | 24 
baby had chorioamnionitis | 24 
mother had no symptoms after birth | 0 
baby had no symptoms after discharge | 192 
baby was discharged from NICU | 192 
contact tracing was performed | 192 
chemoprophylaxis was provided | 192 
vaccination was provided | 192 
placenta histopathology was performed | 24 
placenta histopathology revealed acute funisitis | 24 
placenta histopathology revealed chorioamnionitis | 24 
Neisseria meningitidis was detected in placental surface eSwab | 23 
Neisseria meningitidis was detected in heel-prick blood | 5.5 
Neisseria meningitidis was identified by MALDI-TOF | 23 
Neisseria meningitidis was identified by molecular testing | 23 
Neisseria meningitidis was serogroup W | 23 
Neisseria meningitidis was clonal complex 11 | 23 
baby had funisitis | 24 
baby had chorioamnionitis | 24 
mother had no symptoms after birth | 0 
baby had no symptoms after discharge | 192 
baby was treated with gentamicin | 0.13 
baby was treated with benzylpenicillin | 0.13 
baby was treated with cefotaxime | 24 
baby completed β-lactam therapy | 120 
staff members were at risk | 192 
family members were at risk | 192 
chemoprophylaxis was provided to staff members | 192 
chemoprophylaxis was provided to family members | 192 
vaccination was provided to staff members | 192 
vaccination was provided to family members | 192 
Neisseria meningitidis was detected in placental surface eSwab | 23 
Neisseria meningitidis was detected in heel-prick blood | 5.5 
Neisseria meningitidis was identified by MALDI-TOF | 23 
Neisseria meningitidis was identified by molecular testing | 23 
Neisseria meningitidis was serogroup W | 23 
Neisseria meningitidis was clonal complex 11 | 23 
baby had funisitis | 24 
baby had chorioamnionitis | 24 
mother had no symptoms after birth | 0 
baby had no symptoms after discharge | 192 
baby was discharged from NICU | 192 
contact tracing was performed | 192 
chemoprophylaxis was provided | 192 
vaccination was provided | 192 
placenta histopathology was performed | 24 
placenta histopathology revealed acute funisitis | 24 
placenta histopathology revealed chorioamnionitis | 24 
Neisseria meningitidis was detected in placental surface eSwab | 23 
Neisseria meningitidis was detected in heel-prick blood | 5.5 
Neisseria meningitidis was identified by MALDI-TOF | 23 
Neisseria meningitidis was identified by molecular testing | 23 
Neisseria meningitidis was serogroup W | 23 
Neisseria meningitidis was clonal complex 11 | 23 
baby had funisitis | 24 
baby had chorioamnionitis | 24 
mother had no symptoms after birth | 0 
baby had no symptoms after discharge | 192 
baby was treated with gentamicin | 0.13 
baby was treated with benzylpenicillin | 0.13 
baby was treated with cefotaxime | 24 
baby completed β-lactam therapy | 120 
staff members were at risk | 192 
family members were at risk | 192 
chemoprophylaxis was provided to staff members | 192 
chemoprophylaxis was provided to family members | 192 
vaccination was provided to staff members | 192 
vaccination was provided to family members | 192 
Neisseria meningitidis was detected in placental surface eSwab | 23 
Neisseria meningitidis was detected in heel-prick blood | 5.5 
Neisseria meningitidis was identified by MALDI-TOF | 23 
Neisseria meningitidis was identified by molecular testing | 23 
Neisseria meningitidis was serogroup W | 23 
Neisseria meningitidis was clonal complex 11 | 23 
baby had funisitis | 24 
baby had chorioamnionitis | 24 
mother had no symptoms after birth | 0 
baby had no symptoms after discharge | 192 
baby was discharged from NICU | 192 
contact tracing was performed | 192 
chemoprophylaxis was provided | 192 
vaccination was provided | 192 
placenta histopathology was performed | 24 
placenta histopathology revealed acute funisitis | 24 
placenta histopathology revealed chorioamnionitis | 24 
Neisseria meningitidis was detected in placental surface eSwab | 23 
Neisseria meningitidis was detected in heel-prick blood | 5.5 
Neisseria meningitidis was identified by MALDI-TOF | 23 
Neisseria meningitidis was identified by molecular testing | 23 
Neisseria meningitidis was serogroup W | 23 
Neisseria meningitidis was clonal complex 11 | 23 
baby had funisitis | 24 
baby had chorioamnionitis | 24 
mother had no symptoms after birth | 0 
baby had no symptoms after discharge | 192 
baby was treated with gentamicin | 0.13 
baby was treated with benzylpenicillin | 0.13 
baby was treated with cefotaxime | 24 
baby completed β-lactam therapy | 120 
staff members were at risk | 192 
family members were at risk | 192 
chemoprophylaxis was provided to staff members | 192 
chemoprophylaxis was provided to family members | 192 
vaccination was provided to staff members | 192 
vaccination was provided to family members | 192 
Neisseria meningitidis was detected in placental surface eSwab | 23 
Neisseria meningitidis was detected in heel-prick blood | 5.5 
Neisseria meningitidis was identified by MALDI-TOF | 23 
Neisseria meningitidis was identified by molecular testing | 23 
Neisseria meningitidis was serogroup W | 23 
Neisseria meningitidis was clonal complex 11 | 23 
baby had funisitis | 24 
baby had chorioamnionitis | 24 
mother had no symptoms after birth | 0 
baby had no symptoms after discharge | 192 
baby was discharged from NICU | 192 
contact tracing was performed | 192 
chemoprophylaxis was provided | 192 
vaccination was provided | 192 
placenta histopathology was performed | 24 
placenta histopathology revealed acute funisitis | 24 
placenta histopathology revealed chorioamnionitis | 24 
Neisseria meningitidis was detected in placental surface eSwab | 23 
Neisseria meningitidis was detected in heel-prick blood | 5.5 
Neisseria meningitidis was identified by MALDI-TOF | 23 
Neisseria meningitidis was identified by molecular testing | 23 
Neisseria meningitidis was serogroup W | 23 
Neisseria meningitidis was clonal complex 11 | 23 
baby had funisitis | 24 
baby had chorioamnionitis | 24 
mother had no symptoms after birth | 0 
baby had no symptoms after discharge | 192 
baby was treated with gentamicin | 0.13 
baby was treated with benzylpenicillin | 0.13 
baby was treated with cefotaxime | 24 
baby completed β-lactam therapy | 120 
staff members were at risk | 192 
family members were at risk | 192 
chemoprophylaxis was provided to staff members | 192 
chemoprophylaxis was provided to family members | 192 
vaccination was provided to staff members | 192 
vaccination was provided to family members | 192 
Neisseria meningitidis was detected in placental surface eSwab | 23 
Neisseria meningitidis was detected in heel-prick blood | 5.5 
Neisseria meningitidis was identified by MALDI-TOF | 23 
Neisseria meningitidis was identified by molecular testing | 23 
Neisseria meningitidis was serogroup W | 23 
Neisseria meningitidis was clonal complex 11 | 23 
baby had funisitis | 24 
baby had chorioamnionitis | 24 
mother had no symptoms after birth | 0 
baby had no symptoms after discharge | 192 
baby was discharged from NICU | 192 
contact tracing was performed | 192 
chemoprophylaxis was provided | 192 
vaccination was provided | 192 
placenta histopathology was performed | 24 
placenta histopathology revealed acute funisitis | 24 
placenta histopathology revealed chorioamnionitis | 24 
Neisseria meningitidis was detected in placental surface eSwab | 23 
Neisseria meningitidis was detected in heel-prick blood | 5.5 
Neisseria meningitidis was identified by MALDI-TOF | 23 
Neisseria meningitidis was identified by molecular testing | 23 
Neisseria meningitidis was serogroup W | 23 
Neisseria meningitidis was clonal complex 11 | 23 
baby had funisitis | 24 
baby had chorioamnionitis | 24 
mother had no symptoms after birth | 0 
baby had no symptoms after discharge | 192 
baby was treated with gentamicin | 0.13 
baby was treated with benzylpenicillin | 0.13 
baby was treated with cefotaxime | 24 
baby completed β-lactam therapy | 120 
staff members were at risk | 192 
family members were at risk | 192 
chemoprophylaxis was provided to staff members | 192 
chemoprophylaxis was provided to family members | 192 
vaccination was provided to staff members | 192 
vaccination was provided to family members | 192 
Neisseria meningitidis was detected in placental surface eSwab | 23 
Neisseria meningitidis was detected in heel-prick blood | 5.5 
Neisseria meningitidis was identified by MALDI-TOF | 23 
Neisseria meningitidis was identified by molecular testing | 23 
Neisseria meningitidis was serogroup W | 23 
Neisseria meningitidis was clonal complex 11 | 23 
baby had funisitis | 24 
baby had chorioamnionitis | 24 
mother had no symptoms after birth | 0 
baby had no symptoms after discharge | 192 
baby was discharged from NICU | 192 
contact tracing was performed | 192 
chemoprophylaxis was provided | 192 
vaccination was provided | 192 
placenta histopathology was performed | 24 
placenta histopathology revealed acute funisitis | 24 
placenta histopathology revealed chorioamnionitis | 24 
Neisseria meningitidis was detected in placental surface eSwab | 23 
Neisseria meningitidis was detected in heel-prick blood | 5.5 
Neisseria meningitidis was identified by MALDI-TOF | 23 
Neisseria meningitidis was identified by molecular testing | 23 
Neisseria meningitidis was serogroup W | 23 
Neisseria meningitidis was clonal complex 11 | 23 
baby had funisitis | 24 
baby had chorioamnionitis | 24 
mother had no symptoms after birth | 0 
baby had no symptoms after discharge | 192 
baby was treated with gentamicin | 0.13 
baby was treated with benzylpenicillin | 0.13 
baby was treated with cefotaxime | 24 
baby completed β-lactam therapy | 120 
staff members were at risk | 192 
family members were at risk | 192 
chemoprophylaxis was provided to staff members | 192 
chemoprophylaxis was provided to family members | 192 
vaccination was provided to staff members | 192 
vaccination was provided to family members | 192 
Neisseria meningitidis was detected in placental surface eSwab | 23 
Neisseria meningitidis was detected in heel-prick blood | 5.5 
Neisseria meningitidis was identified by MALDI-TOF | 23 
Neisseria meningitidis was identified by molecular testing | 23 
Neisseria meningitidis was serogroup W | 23 
Neisseria meningitidis was clonal complex 11 | 23 
baby had funisitis | 24 
baby had chorioamnionitis | 24 
mother had no symptoms after birth | 0 
baby had no symptoms after discharge | 192 
baby was discharged from NICU | 192 
contact tracing was performed | 192 
chemoprophylaxis was provided | 192 
vaccination was provided | 192 
placenta histopathology was performed | 24 
placenta histopathology revealed acute funisitis | 24 
placenta histopathology revealed chorioamnionitis | 24 
Neisseria meningitidis was detected in placental surface eSwab | 23 
Neisseria meningitidis was detected in heel-prick blood | 5.5 
Neisseria meningitidis was identified by MALDI-TOF | 23 
Neisseria meningitidis was identified by molecular testing | 23 
Neisseria meningitidis was serogroup W | 23 
Neisseria meningitidis was clonal complex 11 | 23 
baby had funisitis | 24 
baby had chorioamnionitis | 24 
mother had no symptoms after birth | 0 
baby had no symptoms after discharge | 192 
baby was treated with gentamicin | 0.13 
baby was treated with benzylpenicillin | 0.13 
baby was treated with cefotaxime | 24 
baby completed β-lactam therapy | 120 
staff members were at risk | 192 
family members were at risk | 192 
chemoprophylaxis was provided to staff members | 192 
chemoprophylaxis was provided to family members | 192 
vaccination was provided to staff members | 192 
vaccination was provided to family members | 192 
Neisseria meningitidis was detected in placental surface eSwab | 23 
Neisseria meningitidis was detected in heel-prick blood | 5.5 
Neisseria meningitidis was identified by MALDI-TOF | 23 
Neisseria meningitidis was identified by molecular testing | 23 
Neisseria meningitidis was serogroup W | 23 
Neisseria meningitidis was clonal complex 11 | 23 
baby had funisitis | 24 
baby had chorioamnionitis | 24 
mother had no symptoms after birth | 0 
baby had no symptoms after discharge | 192 
baby was discharged from NICU | 192 
contact tracing