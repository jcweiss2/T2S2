29 years old | 0
woman | 0
presented 3 weeks post-partum | 0
right hip pain | 0
right flank pain | 0
right flank bruising | 0
pain started 4 months prior | -2880
6-months pregnant | -2880
uncomplicated spontaneous vaginal delivery | 0
healthy son | 0
severe right flank pain continued post-delivery | 0
past medical history: 5-year opioid addiction | -672
Methadone use | -672
Crohn’s disease diagnosed at 17 years old | -672
Azathioprine 100 mg twice daily | -672
acute flares started 2 years prior | -17520
severe abdominal pain | -17520
vomiting | -17520
bloody diarrhea | -17520
Infliximab infusions monthly | -17520
stopped Infliximab 6 months prior | -4320
financial concerns | -4320
mild acute flares continued | -4320
discharged from 2 GI practices due to noncompliance | -4320
treated flares with oral prednisone 80 mg | -4320
copper intrauterine device | -672
no history of sexually transmitted diseases | -672
fever 100.9°F (38.3°C) | 0
pulse 177 bpm | 0
blood pressure 106/62 mmHg | 0
white blood cell count 50,000 cells/mm3 | 0
elevated platelet count 717 mcL | 0
hemoglobin 6.0 g/dL | 0
lactic acid 5.2 mmol/L | 0
elevated alkaline phosphatase 207 unit/L | 0
chest X-ray no acute abnormalities | 0
CT scan: large complex air-fluid collection | 0
diagnosed with severe sepsis due to retroperitoneal abscess | 0
taken to operating room (OR) | 0
colonic intramural retroperitoneal fistula | 0
incision, drainage, debridement of necrotizing infection | 0
ileal perforation | 0
ileal resection | 0
transferred to ICU intubated | 0
OR cultures: Escherichia coli | 0
OR cultures: Beta Hemolytic Group C Streptococcus | 0
IV Meropenem 500 mg daily | 0
IV Vancomycin 1000 mg daily | 0
IV Clindamycin 900 mg TID | 0
post-op day 1: additional debridement | 24
irrigation of necrotizing infection | 24
wound VAC device placed | 24
sepsis improved | 24
transferred to medical floor on day 4 | 96
hospital day 7: worsening sepsis | 168
tachycardia | 168
tachypnea | 168
fever | 168
leukocytosis 62,000 cells/mm3 | 168
acute respiratory failure | 168
4 liters oxygen via nasal cannula | 168
hospital day 9: exploratory laparotomy | 216
intraperitoneal abscess | 216
transverse colon staple line leak | 216
drainage of abscess | 216
repair of leak with omental patch | 216
pathology: transmural chronic inflammation | 216
serosal fibrous adhesions with granulation | 216
peri-colonic abscesses | 216
cultures: Enterococcus faecalis | 216
cultures: Candida albicans | 216
Vancomycin continued | 216
Micafungin 100 mg daily | 216
blood cultures: no growth | 216
transferred to medical floor on day 11 | 264
discharged on day 14 | 336
long-term acute care | 336
IV antibiotic therapy | 336
aggressive wound management | 336
left long-term care 4 weeks later | 1344
no shortness of breath | 0
denies chest pain | 0
