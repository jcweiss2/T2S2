13 years old|0
    male|0
    admitted to the pediatric department|24
    fever|0
    limping|-24
    left-sided knee pain|-24
    knee pain|0
    tenderness at the infrapatellar ligament|0
    passive flexion|0
    radiography of the knee and leg|0
    elevated leucocytes|0
    elevated CRP|0
    sent home|0
    febrile|24
    IV vancomycin treatment|72
    red and swollen knee|72
    cutaneous micro&dash;ulcerations|72
    MRI synovitis|72
    knee joint effusion|72
    medullary osteomyelitis in the proximal tibia|72
    subperiostal fluid accumulation|72
    elevated CRP|72
    elevated sedimentation rate|72
    acute arthroscopy|72
    synovectomy|72
    lavage of the knee joint|72
    MRSA cultured from blood|72
    MRSA cultured from nasal swabs|72
    MRSA cultured from biopsy materials|72
    PVL-positive|72
    pain increased|168
    CRP and leucocytes continued to rise|168
    MRI progression of infection|168
    renewed surgical debridement|168
    IV vancomycin continued|168
    condition deteriorated|168
    sepsis|168
    multiple bilateral pulmonary infiltrates|168
    respiratory distress|168
    admitted to ICU|168
    necrotizing pneumonia|168
    oral linezolid added|168
    ICU discharge after 4 days|192
    returned to orthopedic ward|192
    clinical improvement|192
    biochemical improvement|192
    CRP rose again|504
    MRI new subperiostal abscess|504
    osteomyelitis progression|504
    edema and enhancement in medullary canal|504
    cortical destruction of the tibia|504
    renewed surgery|504
    condition improved|504
    discharged after 49 days|1176
    IV antibiotics for 7 weeks|1176
    outpatient follow-up|1176
    clinical controls|1176
    biochemical controls|1176
    radiological controls|1176
    progression of osteomyelitis radiologically|1176
    MRI|1176
    CT|1176
    bone scintigraphy|1176
    leukocyte scintigraphy|1176
    no active infection|1176
    radiography normal tibia after 22 months|1584
    fever persisted for 51 days|1224
    elevated CRP for 23 weeks|3864
    elevated SR for 23 weeks|3864
    surgical scar tissue|1176
    plastic surgery|1176
    bilateral pneumonia|168
    necrotizing pneumonia|168
    pleural effusion|168
    atelectasis|216
    linezolid stopped|432
    IV clindamycin|432
    IV rifampicin|432
    progression of osseous changes|1008
    active osteomyelitis|1176
    sequestrum|1176
    irregular osteomyelitis changes|1176
    vital bone uptake|1176
    no pathological leucocyte accumulation|1176
    regression of osteomyelitis|1176
    healed tibia|1584

