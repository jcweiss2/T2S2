23 years old | 0
    female | 0
    presented in the emergency room | -72
    C-section delivery | -72
    pseudotumor cerebri | 0
    acetazolamide | 0
    transferred to the operation room | 0
    emergent laparotomy | 0
    diffuse abdominal rebound tenderness | 0
    guarding | 0
    small bowel gangrene | 0
    gangrened bowel segments resected | 0
    stoma created | 0
    septic shock | 0
    gangrene of the stoma | 0
    transferred to our center | 0
    remnant of the small intestine resected | 0
    gastrodouodenostomy tube inserted | 0
    transferred to the intensive care unit | 0
    admitted to the intestinal rehabilitation unit | 0
    parenteral nutrition | 0
    listed on the waiting list for small intestinal transplantation | 0
    AB+ blood group | 0
    negative flow panel reactive assay | 0
    anti-human leukocyte antigen antibodies | 0
    two time positive bacterial culture from central venous catheters | 0
    pulmonary thromboembolism | 0
    small intestine transplantation | 0
    donor found | 0
    16-year-old brain-dead patient | 0
    O+ blood group | 0
    operation lasted 210 min | 0
    bled 200 cc | 0
    no RBC transfusion | 0
    cold phase 30 min | 0
    weaned from the ventilator | 6
    methylprednisolone 1 gr for 3 days | 0
    60 mg daily dose of thymoglobulin for 5 days | 0
    500 mg of rituximab | 0
    rituximab repeated on the 5th POD | 120
    immunosuppressive maintenance regimen | 0
    tacrolimus | 0
    mycophenolate mofetil | 0
    prednisolone | 0
    small bowel biopsy done | 120
    no rejection | 120
    oral nutrition started | 120
    hemoglobin 9 g/dL | 120
    hemoglobin level dropped to 7.2 g/dL | 240
    hypotension | 240
    tachycardia | 240
    received two units of AB+ RBC transfusion | 240
    hemoglobin level reached 6.2 g/dL | 264
    received another AB+ RBC transfusion | 264
    hemoglobin corrected to 8 g/dL | 264
    hemoglobin dropped to 6 g/dL | 288
    acute jaundice | 288
    total bilirubin level 22 mg/dL | 288
    transferred to the operation room for exploratory laparotomy | 288
    small intestinal hernia observed | 288
    reduced hernia | 288
    bowel intact | 288
    no internal bleeding | 288
    Lactate dehydrogenase (LDH) 935 U/L | 288
    reticulocyte count 10% | 288
    haptoglobin level 0.149 g/L | 288
    total bilirubin 34.9 mg/dL | 288
    indirect bilirubin 18 mg/dL | 288
    2+ bilirubin in urine | 288
    peripheral blood smear fragmented RBCs | 288
    mean corpuscular volume 97 fL | 288
    hemolysis | 288
    medications reviewed | 288
    no medication causing hemolysis | 288
    no preexisting hemolytic disease | 288
    no infection causing hemolysis | 288
    normal G6PD enzyme | 288
    normal hemoglobin electrophoresis | 288
    kidney function tests normal | 288
    platelet count normal | 288
    PLS suspected | 288
    direct coombs test demanded on 12th POD | 288
    direct coombs test negative | 288
    ongoing hemolysis | 312
    received RBC transfusion O+ | 312
    second direct coombs test done on 14th POD | 336
    direct coombs test positive | 336
    total bilirubin decreasing to 11 mg/dL | 432
    IVIG transfusion | 432
    7 cycles of plasmapheresis | 432
    severity of hemolysis decreased | 432
    discharged on 43rd POD | 1032
    episode of cytomegalovirus infection | 1032
    acute rejection | 1032
    discharged with hemoglobin 8.7 g/dL | 1032
    admitted a month later | 1776
    neck soft tissue abscess | 1776
    died of sepsis | 1776
    