76 years old | 0
    woman | 0
    transferred to Daegu Catholic University Medical Center | 0
    worsening dyspnea | 0
    inability to ambulate effectively | -8760
    cerebrovascular disease | -8760
    hypertension | -157248
    type 2 diabetes mellitus | -157248
    subarachnoid hemorrhage | -157248
    endobronchial tuberculosis | -131328
    intracerebral hemorrhage | -35040
    pneumonia episodes | various
    crackle breathing sounds | 0
    no skin lesions | 0
    indwelling urinary catheter | 0
    white blood cell count 361,000/µL | 0
    neutrophils 95.8% | 0
    lymphocytes 1.1% | 0
    monocytes 2.5% | 0
    hemoglobin level 7.2 g/dL | 0
    platelet count 76×103/µL | 0
    C-reactive protein level 41.7 mg/L | 0
    blood urea nitrogen 61 mg/dL | 0
    creatinine 0.8 mg/dL |' 0
    Na 130 mEq/L | 0
    total protein 3.4 g/dL | 0
    albumin 2.2 g/dL | 0
    pro B-natriuretic peptide 3,669 pg/mL | 0
    arterial pH 7.3999 | 0
    arterial carbon dioxide partial pressure 53.1 mmHg | 0
    arterial oxygen partial pressure 61.9 mmHg | 0
    peripheral oxygen saturation 99% | 0
    Candida tropicalis in blood culture | 0
    Candida tropicalis in urine culture | 0
    Klebsiella pneumoniae in sputum culture | 0
    chest radiography findings | 0
    chest CT findings | 0
    pneumonia diagnosis | 0
    acute respiratory failure diagnosis | 0
    candidemia diagnosis | 0
    meropenem treatment | 0
    colistimethate sodium treatment | 0
    fluconazole treatment | 0
    high-flow nasal cannula oxygen therapy | 0
    flexible bronchoscopy on day 2 | 48
    narrowing of the right main bronchus | 48
    anthracotic pigmentation | 48
    bronchial washing | 48
    no infected cells in bronchial washing cytology | 48
    worsening hypoxia | 57
    worsening dyspnea | 57
    endotracheal intubation | 57
    mechanical ventilation | 57
    microscopic hematuria | 72
    urine cytology test | 72
    HSV IgM negative | 72
    HSV IgG positive | 72
    HSV titers 27.9 index value | 72
    weaning failure | 168
    percutaneous dilatational tracheostomy | 168
    bronchoscopy | 168
    bronchial washing cytology | 168
    HSV type 1-positive cells | 168
    intranuclear inclusions | 168
    multinucleation | 168
    RT-PCR positive for HSV type 1 | 168
    HSV type 1-infected cells in urine cytology | 72
    acyclovir treatment | 168
    subsequent urine cytology absence of HSV | 216
    repeat bronchoscopy not performed | 168
    vital signs stable without fever | 168
    white blood cell count 4,400/µL | 168
    neutrophils 88.7% | 168
    lymphocytes 7.5% | 168
    monocytes 2.4% | 168
    hemoglobin level 8.6 g/dL | 168
    platelet count 65×103/µL | 168
    C-reactive protein level 78.1 mg/L | 168
    chest radiography stable | 168
    vancomycin-resistant Enterococci in urine culture | 480
    vancomycin-resistant Enterococci in stool culture | 480
    sepsis | 480
    linezolid treatment | 480
    urine output decrease | 480
    acute renal failure | 480
    refusal of hemodialysis | 480
    refusal of cardiopulmonary resuscitation | 480
    patient death | 672
    