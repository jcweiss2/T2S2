Here is the extracted table of clinical events and timestamps:

Hodgkin lymphoma | -7200
mantle field RT | -7200
chemotherapy | -7200
splenectomy | -7200
DLBCL | -480
denosumab | -480
rituximab | -480
cyclophosphamide | -480
doxorubicin | -480
vincristine | -480
prednisone | -480
dizziness | -480
ataxia | -480
memory loss | -480
brain MRI | -480
whole brain radiation therapy | -480
intrathecal cytarabine | -480
coronary artery disease | 0
hypertension | 0
hypothyroidism | 0
gastroesophageal reflux disease | 0
mini-stroke | 0
coronary artery bypass grafting | 0
right carotid endarterectomy | 0
appendectomy | 0
aortic valve replacement | 0
neck mass | 0
CT scan | 0
biopsy | 0
EMC | 0
resection | 0
revision surgery | 24
adjuvant chemoradiation | 24
xerostomia | 168
fibrosis | 168
restaging PET scan | 168
neuroendocrine tumor | 168
bronchoscopy | 168
biopsy | 168
Hurthle cell adenoma | 168
thyroid ultrasound | 168
fine needle aspiration | 168
hemithyroidectomy | 240
follow-up CT scan | 360
interval growth | 360
PET scan | 360
stereotactic body radiation therapy | 420
epistaxis | 480
supratherapeutic international normalized ratio | 480
warfarin | 480
fall | 480
altered mental status | 480
hypoxic respiratory failure | 480
intubation | 480
pneumonia | 480
sepsis | 480
vasopressor requirement | 480
bilateral pleural effusions | 480
therapeutic thoracentesis | 480
flow cytometry | 480
CD10-positive lambda-skewed B cell population | 480
small B cell lymphoma | 480
palliative care | 504
inpatient hospice | 504
death | 504