74 years old | 0
female | 0
admitted for bilateral total knee replacement arthroplasty | 0
degenerative osteoarthritis | -8760
angina | -8760
hypertension | -8760
isosorbide-5-mononitrate | -8760
atenolol | -8760
blood and biochemistry tests within normal ranges | 0
cardiomegaly | 0
sinus bradycardia | 0
first degree atrioventricular block | 0
T wave inversion in leads V2-3 | 0
ejection fraction 60% | 0
combined spinal epidural anesthesia | 0
bupivacaine | 0
levobupivacaine | 0
epidural catheter | 0
surgery began | 0
oxygen administered via face mask | 0
vital signs stable | 0
pulse oxygen saturation 100% | 0
arterial blood gas analysis within normal ranges | 0
operation time 3 hours 5 minutes | 0
anesthesia period 4 hours 25 minutes | 0
estimated blood loss 1100 ml | 0
urine volume 850 ml | 0
hydroxyethyl starch | 0
Hartmann solution | 0
packed red blood cells | 0
recovery room | 205
oxygen supply 6 L/min | 205
pain controlled by epidural catheter | 205
stable vital signs | 205
arterial blood gas analysis within normal ranges | 205
transported to ward | 210
oxygen supply 2 L/min | 210
pulse oxygen saturation 90% | 210
oxygen supply 5 L/min | 210
drowsy mental state | 9
unresponsive to calling | 9
blood pressure within normal range | 9
heart rate within normal range | 9
respiratory rate 20 times/min | 9
pulse oxygen saturation 90% | 9
oxygen supply 7 L/min | 9
simple chest radiography | 9
brain computed tomography | 9
bilateral pulmonary effusion | 9
no abnormal findings on brain CT | 9
brain magnetic resonance imaging | 24
3D pulmonary arteriography | 24
high signal intensity lesions in cerebral and cerebellar cortices | 24
reduced apparent diffusion coefficient | 24
fat embolism | 24
transferred to stroke unit | 24
breathing shallow and irregular | 24
pulse oxygen saturation 84% | 24
eyeball deviation | 24
nystagmus | 24
unresponsive to stimulation | 24
stuporous | 24
intubated | 24
mechanical ventilator | 24
blood pressure 95/60 | 24
fever 38 | 24
low molecular weight heparin | 24
hemoglobin 8.3 g/dl | 24
platelets 34,000/µl | 24
coagulation time increased | 24
packed RBCs and platelets transfused | 24
inotropics and diuretics administered | 24
ischemic colitis | 72
petechial rash | 72
low molecular weight heparin administered | 96
conscious state still stuporous | 120
neurological symptoms unimproved | 120
electroencephalogram | 120
moderate to severe diffuse cerebral dysfunction | 120
weaned off mechanical ventilator | 168
endotracheal tube removed | 312
respiratory and neurological symptoms improved | 312
transferred to general ward | 408
brain MRI revealed multiple brain infarctions | 624
discharged | 1056