32 years old| 0
male | 0
admitted to the hospital | 0
abdominal pain | -4320
recurrent ascites | -4320
paracentesis procedures | -4320
albumin therapy | -4320
difficulty ambulating | -4320
nausea | -4320
dizziness | -4320
sodium level of 120 mEq/L | -4320
ceftriaxone | -4320
dyspnea | -4320
increased oxygen requirements | -4320
pleural fluid analysis positive for Cryptococcal antigen | -4320
IV fluconazole (400 mg) | -4320
cryptogenic cirrhosis | 0
right hypothalamic juvenile pilocytic astrocytoma status-post resection | 0
radiation (20 years prior) | 0
bilateral occipital ventriculoperitoneal (VP) shunt placement | 0
panhypopituitarism | 0
oral hydrocortisone (30 mg/daily) | 0
desmopressin (DDVAP) | 0
hypernatremic | 0
afebrile | 0
normal white blood cell (WBC) count | 0
blood cultures initially negative | 0
HIV test negative | 0
ALT 28 units/L | 0
AST 35 units/L | 0
viral hepatitis panel negative | 0
stress-dose steroids (IV hydrocortisone 50 mg q8) |A0
symptomatic relief of dyspnea after thoracentesis | 24
thoracentesis removed 1.5 L transudative fluid | 24
paracentesis performed | 36
206 nucleated cells/μL | 36
ceftriaxone discontinued | 36
CT thorax revealed massive left-sided pleural effusion | 24
atypical pneumonia | 24
reactive lymphadenopathy | 24
serum Cryptococcal Ag positive | 72
liposomal amphotericin B (3 mg/kg q24h) | 72
flucytosine (25 mg/kg q6h) | 72
flucytosine toxicities monitored | 72
pleural fluid Cryptococcal Ag positive | 96
blood cultures grew C. neoformans | 120
pleural fluid cultures grew C. neoformans | 120
abdominal fluid cultures grew C. neoformans | 120
transthoracic echo showed no vegetation | 120
CT head no ventriculitis | 120
lumbar puncture completed | 96
CSF positive for Cryptococcal Ag | 96
CSF culture positive | 168
VP shunt removed | 120
external ventricular drain (EVD) placed | 120
CSF remained positive for Cryptococcal Ag | 264
therapeutic thoracentesis revealed exudative fluid | 264
serosanguinous fluid | 264
pleural fluid grew three Cryptococcus colonies | 264
lethargic | 264
altered mental status | 264
EEG consistent with non-convulsive status epilepticus | 264
levetiracetam | 264
lacosamide | 264
intubated | 264
midazolam drip | 264
ketamine | 264
pressor support | 264
anuric AKI | 264
acute tubular necrosis | 264
continuous veno-venous hemofiltration (CVVH) | 264
flucytosine renally adjusted | 264
worsening septic shock | 312
negative repeat blood cultures | 312
piperacillin/tazobactam | 312
vancomycin | 312
meropenem | 312
daptomycin | 312
five pressors | 312
sodium bicarbonate infusion | 312
increase in stress steroids | 312
shock liver | 336
disseminated intravascular coagulopathy (DIC) | 336
bleed from nasogastric tube | 336
transfusions of blood | 336
transfusions of platelets | 336
transfusions of fresh frozen plasma | 336
transfusions of cryoprecipitate | 336
comfort care measures | 360
died | 360
