64 years old | 0
male | 0
admitted to the emergency room | 0
exertional dyspnea | 0
history of alcohol consumption | -672
liver cirrhosis | -672
productive cough | -48
fever | -48
temperature of 36 °C | 0
blood pressure 100/60 mmHg | 0
heart rate 78 bpm | 0
respiratory rate 19 bpm | 0
oxygen saturation of 96% | 0
round opacity in the right upper lobe | 0
antibiotic therapy started | 0
intravenous ceftriaxone | 0
oral clarithromycin | 0
sputum culture positive for E. hormaechei | 24
bacterium sensitive to levofloxacin | 24
therapy modified | 24
levofloxacin | 24
systemic respiratory distress syndrome | 48
intubated | 48
transferred to the intensive care unit | 48
mechanical ventilation | 48
lung-protective strategy | 48
hemodynamic instability | 72
additional blood cultures drawn | 72
antibiotic therapy escalation | 72
imipenem/cilastatin | 72
septic shock | 96
died | 96