47 years old | 0
male | 0
admitted to the hospital | 0
COVID-19 diagnosis | -144
shortness of breath | -144
fever | -144
non-productive cough | -144
dyspnea | -144
hypertension | 0
anginal pain | 48
typical anginal pain | 48
oxygen desaturation | -96
thorax CT | -96
diffuse bilateral infiltrates | -96
ground glass opacities | -96
crazy paving with thickened interlobular septa | -96
consolidation in lower lobes | -96
enoxaparin sodium treatment | -96
prednisolon treatment | -96
moxifloksasin treatment | -96
amlodipin treatment | -96
favirapiravir treatment | -240
ceftriaxone treatment | -144
high-flow nasal oxygen | 48
blood pressure 135/68 mmHg | 48
heart rate 73 bpm | 48
oxygen saturation 88-93% | 48
body temperature 36.7°C | 48
cardiac examination | 48
inferior STEMI | 48
acetylsalicylic acid treatment | 48
ticagrelor treatment | 48
heparin treatment | 48
cardiac symptoms decreased | 48
emergency coronary angiography | 48
30-40% stenosis in left anterior descending artery | 48
left main coronary artery normal | 48
left circumflex artery normal | 48
right coronary artery normal | 48
ST segment elevation regressed | 48
high sensitivity troponin 0.012 ng/mL | 48
troponin 0.056 ng/mL | 48
kidney function tests normal | 48
liver function tests normal | 48
d-dimer 520 ng/mL | 48
fibrinogen 589 mg/dL | 48
ferritin 1693 ng/mL | 48
lactate dehydrogenase 466 U/L | 48
C-reactive protein 4.1 mg/dL | 48
pro-brain natriuretic peptide 20 pg/mL | 48
computed tomographic pulmonary angiography | 48
no pulmonary embolism | 48
MINOCA diagnosis | 48
cardiogoniometry | 72
septal inferior myocardial ischemia | 72
medical treatment | 72
clinical improvement | 120
hemodynamic improvement | 120
transferred to normal medical ward | 120
discharged | 264