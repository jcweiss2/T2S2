72 years old | 0
    man | 0
    history of clinically quiescent Crohn's disease | 0
    presented to the emergency department | 0
    fever | -96
    fatigue | -96
    altered mental status | -96
    nausea | -96
    vomiting | -96
    new diagnosis of acute myelogenous leukemia | -96
    tumor lysis syndrome | -96
    acute kidney injury | -96
    hyperleukocytosis | -96
    intensive care unit admission | 0
    initial diagnostic uncertainty | 0
    multi-organ failure | 0
    treated empirically with ceftazidime | 0
    treated empirically with vancomycin | 0
    possible septic shock | 0
    blood cultures were sterile | 0
    urine cultures were sterile | 0
    computed tomography of chest | 0
    computed tomography of abdomen | 0
    computed tomography of pelvis | 0
    became neutropenic | 0
    cytoreductive therapy with hydroxyurea | 0
    cytoreductive therapy with cytarabine | 0
    defervesced | 0
    received dose-reduced G-CLAM | 0
    ceftazidime continued for neutropenic prophylaxis | 0
    vancomycin stopped | 0
    lack of evidence for active infection | 0
    fevered | 120
    reported mild abdominal pain | 144
    reported new diarrhea | 144
    febrile neutropenia | 144
    enteric pathogen panel obtained | 144
    rapid PCR using Biofire FilmArray GI panel | 144
    blood agar plate | 144
    no pathogens detected by PCR | 144
    loperamide started | 144
    blood agar plate showed 4+ MRSA | 168
    reduced normal fecal flora | 168
    profound immunocompromised status | 168
    oral vancomycin started | 168
    possible MRSA enterocolitis | 168
    gram-negative coverage broadened to piperacillin-tazobactam | 168
    anaerobic coverage broadened to piperacillin-tazobactam | 168
    developed respiratory distress | 192
    intubated | 192
    recurrence of acute kidney injury | 192
    recurrence of shock | 192
    vancomycin IV added | 192
    computed tomography of abdomen | 192
    computed tomography of pelvis | 192
    diffuse small bowel wall edema | 192
    diffuse small bowel wall thickening | 192
    diffuse small bowel wall dilatation | 192
    pneumatosis | 192
    no pneumoperitoneum | 192
    no surgical interventions available | 192
    transitioned to comfort care | 192
    expired | 192
    postmortem evaluation | 192
    gross dilatation of duodenum | 192
    gross dilatation of jejunum | 192
    dusky discoloration | 192
    mucosal erythema | 192
    congestion | 192
    gram positive cocci | 192
    focal mucosal erosions in stomach | 192
    focal mucosal erosions in cecum | 192
    no pseudomembranes found | 192
    cause of death attributed to septic shock | 192
    multiorgan failure | 192
    secondary to MRSA enterocolitis | 192