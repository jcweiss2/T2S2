18 years old | 0
male | 0
unrestrained driver in a rollover motor vehicle accident | -1
prolonged extrication | -1
positive blood alcohol screen | -1
intubated at the scene | -1
taken to a Level-1 trauma center | -1
multiple fractures | 0
open book pelvic fracture | 0
complete disruption of the posterior sacroiliac complex | 0
vertical and rotational instability of the left hemipelvis | 0
pubic symphysis diastasis | 0
left greater than right sacroiliac joint disruption | 0
left open comminuted femoral shaft fracture | 0
left distal tibia shaft fracture | 0
systolic blood pressure in the 80s | 0
tachycardic | 0
focused assessment with sonography for trauma scan was positive | 0
pelvis bound with a sheet and secured using hemostats | 0
pulses detected with Doppler ultrasound in the bilateral lower extremities | 0
poor response to initial fluid bolus | 0
sustained tachycardia | 0
taken to the angiography suite | 0
significant slowing of flow within the left superior gluteal and left internal pudendal arteries | 0
radiographic blush | 0
vasospasm versus distal arterial injury | 0
empiric Gelfoam embolization of the left internal iliac artery | 0
hypotension and tachycardia subsequently stabilized | 0
hemodynamic instability began to respond to resuscitation | 0
pelvic fractures temporarily stabilized through an external fixator | 0
left femoral shaft fracture stabilized | 0
definitive fixation of the pelvis and both sacroiliac joints | 48
definitive fixation of the left femur | 96
definitive fixation of the left tibia | 48
remained intubated post-operatively | 0
transferred out of the Intensive Care Unit | 192
transferred to a transitional care unit | 192
wounds followed throughout hospital course | 0
incisions remained clean and dry | 0
intermittently febrile | 0
increasing lymphocyte count | 240
computed tomography of the pelvis | 240
evidence of a 15cm diameter simple-appearing fluid collection | 240
scant gas collection located lateral to the left hip | 240
managed with observation | 240
discharged to a rehabilitation center | 360
continued to have drainage from the left buttock area | 528
developed early signs of wound margin epidermolysis | 528
readmitted to the hospital | 528
evidence of increasing drainage | 528
marginal erythema | 528
induration | 528
epidermolysis | 528
early signs of sepsis | 528
started on intravenous vancomycin | 528
underwent local debridement of his left hip/buttock wound | 528
cavitation extending posterior to the greater trochanter | 528
significant fat necrosis | 528
epidermolysis | 528
scheduled for repeat debridement | 528
repeat CT scan | 528
questionable intramuscular abscess formation | 528
ill-defined collection of fluid and gas in the left gluteal musculature | 528
underwent aggressive repeat surgical debridement of left hip | 576
massive gluteal muscle necrosis identified | 576
wound and tissue cultures positive for Proteus mirabilis | 528
wound and tissue cultures positive for Serratia marcescens | 528
wound and tissue cultures positive for Klebsiella pneumoniae | 528
underwent a third surgical debridement of the left hip wound | 600
drain placed | 600
continued on vancomycin | 528
piperacillin/tazobactam added | 528
wound noted to have no erythema or drainage | 696
significant decrease in swelling | 696
continued induration of the abductor compartment | 696
progressed with physical therapy | 696
recovered from traumatic injuries | 696
seen for 4-month follow-up | 1056
significant gluteal fold asymmetry | 1056
necrosis and atrophy | 1056
ambulated with a Trendelenburg gait | 1056
orthopedic fractures healed | 1056
unable to return to competitive football | 1056