12 years old | 0
abdominal lymphoma removal | -120
open drainage site on abdomen | -120
MRSA infection | 0
admission | 0
isolation | 0
scheduled chemotherapy | 0
local antiseptic (octenidin) treatment | 0
no improvement | 12
Medihoney™ application | 12
wound free of bacteria | 24
chemotherapy started | 24
MRSA infection |D0
isolation |D0
scheduled chemotherapy |D0
local antiseptic (octenidin) treatment |D0 (start)
no improvement |D+12 (288 hours)
Medihoney™ application |D+12 (288 hours)
wound free of bacteria |D+14 (336 hours)
chemotherapy started |D+14 (336 hours)
