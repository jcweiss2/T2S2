22 years old | 0
male | 0
admitted to the hospital | 0
fatigue | -360
chest tightness | -360
shortness of breath | -360
cold | -72
inability to walk | -72
aggravation of shortness of breath | -96
hospitalized in 2016 | -2160
muscle weakness | -2160
chest tightness | -2160
shortness of breath | -2160
electromyography | -2160
myogenic changes | -2160
methylprednisolone | -2160
family history of muscle weakness | -4320
family history of tachycardia | -4320
pseudohypertrophic muscular dystrophy | -4320
hereditary muscular dystrophy | -4320
progressive shortness of breath | 0
respiratory rate 32/min | 0
SpO2 96% | 0
sinus tachycardia | 0
pCO2 65 mmHg | 0
blood pressure 16.7/9.04 Kpa | 0
body temperature 36.8 °C | 0
muscle strength grade 4 | 0
abnormal breath sounds | 0
lactate 25 mmol/L | 0
creatinine phosphokinase-MB 385 U/L | 0
N-terminal pro-brain natriuretic peptide 1622 pg/mL | 0
white blood cell count 1.88 × 10^10/L | 0
procalcitonin 5.6 ng/mL | 0
interleukin-6 32 pg/mL | 0
global heart enlargement | 0
mild mitral and tricuspid valve regurgitation | 0
pulmonary artery pressure 3.86 Kpa | 0
pericardial effusion | 0
mitochondrial crisis | 0
hyperlactic acidemia | 0
respiratory failure | 0
multiple organ failure | 0
limb muscle weakness | 0
intravenous methylprednisone | 0
intravenous immunoglobulin | 0
high-dose B vitamins | 0
coenzyme Q10 | 0
L-carnitine | 0
adenosine triphosphate | 0
fat emulsion | 0
amino acids | 0
hormones | 0
traditional Chinese medicine | 0
mitochondrial myopathy | 0
myasthenia | 0
stroke | 0
epilepsy-like symptoms | 0
hyperlactatemia | 0
severe shock | 0
multiple visceral failures | 0
poor microcirculation | 0
organ support | 0
mitochondrial TRNL1 3243A>G mutation | 0
sepsis | 0
hyperlactatemia | 0
respiratory insufficiency | 0
circulatory failure | 0
mechanical ventilation | 24
veno-arterial extracorporeal membrane oxygenation | 24
continuous renal replacement therapy | 24
antibiotics | 24
nutrition | 24
regained consciousness | 48
severe respiratory muscle weakness | 48
severe limb muscle weakness | 48
diaphragmatic pacing | 168
rehabilitation training | 168
muscle strength training | 168
disengaged from ventilator | 720
standing training | 720
walking with assistance | 1440
walking independently | 2160
discharged | 2160