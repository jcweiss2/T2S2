62 years old | 0
male | 0
admitted to hospital | 0
lumbar back pain | -168
fever | -168
chronic congestive heart failure | 0
hypertension | 0
diabetes mellitus | 0
peripheral arterial disease | 0
atrial fibrillation | 0
hemodynamically stable | 0
no acute signs of worsening cardiac or lung function | 0
abdomen diffusely tender on palpation | 0
no signs of peritoneal inflammation | 0
non-contrast computed tomography scan | 0
confluent mass of periaortic soft tissue | 0
retroperitoneal fibrosis | 0
aortic calcifications | 0
abnormal acute phase inflammatory markers | 0
leukocytes 12.280/mmc | 0
neutrophils 96% | 0
C-reactive protein 225 mg/L | 0
magnetic resonance imaging of dorsal and lumbar spine | 0
no spondylodiscitis | 0
transthoracic echocardiogram | 0
no cardiac vegetations | 0
intravenous meropenem | 0
intravenous vancomycin | 0
blood cultures positive for methicillin-sensitive Staphylococcus aureus | 0
treatment changed to intravenous cloxacillin | 0
new onset syncope | 168
shock | 168
progressively worsening lumbar pain | 168
repeat abdominal CT scan | 168
retroperitoneal collection of blood | 168
aortic rupture at the level of the left renal artery | 168
angiography | 168
aortic balloon inflated above the superior mesenteric artery | 168
endovascular aortic cuff placed at the level of the renal arteries | 168
transferred to Intensive Care Unit | 168
repeat abdominal and pelvis CT scan | 192
small leak to the right renal artery | 192
patency of celiac trunk | 192
patency of SMA | 192
patency of right renal artery | 192
patency of inferior mesenteric artery | 192
operated on again | 216
right colon ischemia | 216
transverse colon ischemia | 216
left colon ischemia | 216
resection performed | 216
repeat abdominal CT scan | 240
no endoleak | 240
patency of all splachnic arteries except the left renal | 240
dependent on vasopressor and inotropic support | 168
mechanical ventilation | 168
hemodialysis | 168
intravenous vancomycin and cloxacillin continued post-operatively | 168
persistence of MSSA bacteremia | 168
expired 17 days after admission | 408
autopsy | 408
mycotic thrombosed abdominal aneurysm | 408
necrosis of left aortic wall | 408
thrombosis of the left renal artery | 408
no aortic rupture | 408
aortic wall heavily infiltrated with neutrophils | 408
gram positive cocci present in the sections | 408
no endocardial or valvular vegetations | 408
no fibrotic tissue found on peritoneum | 408
multiple abscess of peritoneal fat with bacterial and yeast | 408
vascular invasion | 408