66 years old | 0
male | 0
diabetes mellitus | 0
obesity | 0
body mass index 25.3 kg/m2 | 0
consumed rice wine thrice a week | 0
admitted for colonoscopy | 0
positive fecal immunochemical test result | -24
colonoscopy | 0
endoscopic mucosal resection | 0
15 polyps resected | 0
preventive hemoclips applied | 0
discharged from endoscopy room | 0
visited emergency department | 24
complained of right abdominal pain | 24
tenderness and rebound tenderness | 24
severe infection | 24
white blood cell count 21460/mm3 | 24
C-reactive protein level 17.8 mg/dL | 24
blood urea nitrogen level 28 mg/dL | 24
creatinine 2.13 mg/dL | 24
lactic acid 2.4 mmol/L | 24
total bilirubin 1.7 mg/dL | 24
abdominopelvic computed tomography | 24
multiple air bubbles in right lateral abdominal muscles | 24
intensive medical treatments | 24
broad-spectrum antibiotic therapy | 24
piperacillin/tazobactam 4.5 g/day | 24
emergency exploratory laparotomy | 44
laparoscopic right hemicolectomy | 44
no perforation found | 44
condition aggravated | 44
multiple-organ failure | 44
metabolic acidosis | 44
diagnosis of necrotizing fasciitis | 48
urgent surgical debridement and drainage | 48
extensive broad-spectrum antibiotic therapy | 48
renal replacement therapy | 48
intensive care unit | 48
two more surgical debridements and drainages | 72
imipenem-resistant Acinetobacter baumannii | 72
extended spectrum beta-lactamase negative Escherichia coli | 72
septic shock | 840
multiple-organ failure | 840
death | 840