40 years old | 0
male | 0
admitted to the Haematology Clinic of ‘Attikon’ Hospital | 0
recurrent acute lymphoblastic leukaemia (ALL) | 0
allogeneic bone marrow transplantation | 0
extensive maculopapular skin rash | 2160
widespread hyperpigmentation of the skin | 2160
clinical diagnosis of GVHD | 2160
confirmed histologically with a skin biopsy | 2160
systemic corticosteroids | 2160
no observed change in mental and emotional state | 2160
treatment with systemic steroids on a gradually reducing regime | 2160
monitored as an outpatient | 2160
remained fairly stable clinically | 2160
unexplained fever | 10800
admitted to the Haematology Clinic | 10800
intravenous antibiotics | 10800
became apyrexial | 10800
no changes in mental state | 10800
mood remained euthymic | 10800
non-specific, vague abdominal disturbance | 10824
acute onset of depressive effect | 10824
low mood | 10824
stopped eating | 10824
severely disturbed night sleep | 10824
stopped communicating | 10824
no evidence of frank aphasia | 10824
reluctant to see wife and children | 10824
markedly reduced motivation | 10824
markedly reduced energy | 10824
fear of death | 10824
jovial | 10824
hopeful | 10824
sociable | 10824
no report of depressive symptoms in recent past | 10824
extensive investigations | 10824
abdominal CT scans | 10824
liaison with other medical specialties | 10824
no specific cause for abdominal disturbance | 10824
ALL remained in remission | 10824
mood continued to deteriorate | 10824
consultation by Liaison Psychiatric team requested | 10824
profoundly low in mood | 10824
pronounced anhedonia | 10824
biological symptoms of severe depression | 10824
significantly reduced energy | 10824
severely disturbed sleep | 10824
lack of reduced appetite | 10824
marked weight loss | 10824
hopelessness | 10824
helplessness | 10824
passive death wishes | 10824
suicidal thoughts | 10824
no suicidal plan | 10824
well-orientated | 10824
MMSE score 30/30 | 10824
excluded hypoactive delirium | 10824
excluded organic brain cause | 10824
severe depressive episode without psychotic symptoms | 10824
HAM-D score 25 | 10824
treatment with duloxetine initiated | 10824
duloxetine titrated up to 60 mg daily | 10824
partial response | 10824
death wishes subsided | 10824
remained very low in mood | 10824
continued biological symptoms of depression | 10824
HAM-D score 17 | 10824
vague abdominal disturbance | 10824
no definite organic cause | 10824
localized abdominal pain in lower left quadrant | 10896
repeat abdominal CT scan | 10896
intestinal leakage | 10896
explorative laparotomy | 10896
sepsis | 10896
passed away | 10944
no marked change in mental state | 10944
remained severely depressed | 10944
