35 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
pregnant | 0 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
fever | -240 | 0 | Factual
cough | -240 | 0 | Factual
dyspnoea | -120 | 0 | Factual
chest distress | -240 | 0 | Factual
shortness of breath | -240 | 0 | Factual
yellow viscous sputum | -240 | 0 | Factual
no chills | -240 | 0 | Negated
cyanosis of the lip | 0 | 0 | Factual
thick breathing sounds in both lungs | 0 | 0 | Factual
dry and wet rales in the right lower lung | 0 | 0 | Factual
heart rate of 130 beats/min | 0 | 0 | Factual
respiratory rate of 20 times/min | 0 | 0 | Factual
gestational age of 34 + 4 wk | 0 | 0 | Factual
G2P1 | 0 | 0 | Factual
left occiput anterior | 0 | 0 | Factual
maternal lower weight | 0 | 0 | Factual
oligohydramnion | 0 | 0 | Factual
premature live baby | 0 | 0 | Factual
electrolyte disturbance | 0 | 0 | Factual
hypoproteinaemia | 0 | 0 | Factual
pH 7.472 | 0 | 0 | Factual
partial pressure of carbon dioxide 34.0 mmHg | 0 | 0 | Factual
partial pressure of oxygen 56 mmHg | 0 | 0 | Factual
sulfur dioxide 88.6% | 0 | 0 | Factual
C-reactive protein (CRP): 186.33 mg/L | 0 | 0 | Factual
erythrocyte sedimentation rate: 69.00 mm/h | 0 | 0 | Factual
procalcitonin (PCT): 2.24 ng/mL | 0 | 0 | Factual
White blood cell (WBC) 18.29 × 10^9/L | 0 | 0 | Factual
neutrophil % 90.10% | 0 | 0 | Factual
lymphocyte 0.97 × 10^9/L | 0 | 0 | Factual
Alkaline phosphatase 232 U/L | 0 | 0 | Factual
total bilirubin 23.1 μmol/L | 0 | 0 | Factual
albumin (ALB) 33.9 g/L | 0 | 0 | Factual
K+ 2.93 mmol/L | 0 | 0 | Factual
sodium 129 mmol/L | 0 | 0 | Factual
chloride 89 mmol/L | 0 | 0 | Factual
D-dimer 3.50 mg/L | 0 | 0 | Factual
multiple plaques, miliary foci, nodular foci with partial consolidation and cavities in the upper and lower lobes of both lungs | 0 | 0 | Factual
single viable foetus | 0 | 0 | Factual
head presentation | 0 | 0 | Factual
oligohydramnios | 0 | 0 | Factual
caesarean section | 24 | 24 | Factual
oxyhemoglobin saturation increased to 95%-98% | 24 | 48 | Factual
assisted ventilation by endotracheal intubation | 24 | 48 | Factual
empirical antibiotic therapy | 24 | 120 | Factual
symptomatic treatment of fluid and ALB infusion | 24 | 120 | Factual
irrigation solution collected and tested for metagenomic next-generation sequencing (mNGS) | 24 | 48 | Factual
S. aureus combined with novel coronavirus infection | 24 | 48 | Factual
no acid-fast bacilli in the sputum tuberculosis smear | 48 | 48 | Negated
tubercle bacillus-polymerase chain reaction (TB-PCR) and nontuberculosis mycobacterium-PCR were negative | 48 | 48 | Negated
galactomannan experiments were normal | 48 | 48 | Negated
vancomycin and meropenem | 48 | 120 | Factual
anticoagulant therapy | 48 | 120 | Factual
treatments to relieve the cough and reduce the amount of sputum | 48 | 120 | Factual
nasal tube oxygen with a flow rate of 3-4 L/min | 48 | 120 | Factual
multiple areas of inflammation in both lungs, mildly enlarged mediastinal lymph nodes and a small amount of bilateral pleural effusion | 96 | 96 | Factual
CRP was 38.54 mg/L | 96 | 96 | Factual
WBC count was 8.25 × 10^9/L | 96 | 96 | Factual
PCT was 0.129 ng/mL | 96 | 96 | Factual
potassium was 4.04 mmol/L | 96 | 96 | Factual
D-dimer was 2.44 mg/L | 96 | 96 | Factual
TB-PCR was negative | 96 | 96 | Negated
inflammatory lesions were gradually absorbed and improved | 216 | 216 | Factual
sitafloxacin 50 mg twice daily | 216 | 240 | Factual
discharged from the hospital | 240 | 240 | Factual
multiple lung inflammation was absorbed slightly | 336 | 336 | Factual
multiple lung inflammation was apparently absorbed | 744 | 744 | Factual