70 years old | 0
male | 0
BMI 31.14 | 0
smoker | 0
hypertensive | 0
endovascular aortic aneurysm repair | -52560
nephrectomy for kidney cancer | -52560
incisional hernia | -52560
laparoscopic multilayered mesh repair (Proceed®) | -52560
CT scan showed endoleak | -672
recurrent incisional hernia | -672
admitted to our hospital | 0
aorto-bi-iliac bypass | 0
abdominal wall sublay prosthetic repair with composite mesh (Parietex™) | 0
partial resection of ileum | 0
postoperative course uneventful | 0
discharged after twenty-eight days | 672
US scan showed large periprosthetic haematoma | 792
percutaneous drain placement under radiological guidance | 792
drains removed after seven days | 960
fever | 1200
leakage of enteric material from previous drain path | 1200
CT scan demonstrated xifo-pubic fluid collection | 1200
jejunal fistula (iatrogenic lesion from drain placement) | 1200
US guided positioning of two drains | 1200
evacuation of 1800 cc enteric material | 1200
nasogastric tube | 1200
total parenteral nutrition tailored to caloric and nutrient demands | 1200
intravenous octreotide | 1200
antibiotics | 1200
supervening sepsis | 1200
surgical treatment | 1200
infected mesh removed | 1200
open abdomen with thick granulation tissue | 1200
jejunal perforation confirmed | 1200
Kehr drain inside open fistula connected to vacuum-assisted system | 1200
Negative Pressure Wound Treatment (NPWT) (V.A.C. ULTA™) | 1200
baby bottle nipple of soft silicone over fistula | 1200
absorbable stitches (PDS®) | 1200
biologic glue (BioGlue-Levibiotech) | 1200
NPWT with low pressure (25 mmHg) | 1200
stitches and glue dissolved by enteric enzymes | 1200
subsequent unsuccessful efforts with Hyalomatrix® | 1200
platelet gel | 1200
non-cross-linked biologic implant (Tutomesh®) | 1200
biologic glue (Tisseel-Baxter) | 1200
NPWT | 1200
handmade “fistula patch” system | 1200
10 cm silastic drain placed across fistula as tutor | 1200
anchored to surface | 1200
replaced by smaller caliber drains | 1200
released into intestinal lumen | 1200
device effective to narrow fistula and protect surrounding tissue | 1200
