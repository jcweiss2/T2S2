generalized malaise | -168
shortness of breath | -168
lower extremity swelling | -168
subjective fever | -168
denies chest pain | -168
denies orthopnea | -168
denies paroxysmal nocturnal dyspnea | -168
blood pressure of 79/54 mmHg | 0
oral temperature of 38.3°C | 0
heart rate of 55 beats/min | 0
crackles up to the mid-lung fields bilaterally | 0
irregularly, irregular heart rhythm | 0
2+ pitting edema up to the knees | 0
congestion in the bilateral lower lung fields | 0
cardiomegaly | 0
sodium level of 126 | 0
potassium of 5.2 | 0
blood urea nitrogen of 33 | 0
creatinine of 2.77 | 0
white blood count of 4.9 | 0
INR of 2.8 | 0
signs of digoxin toxicity | 0
peak troponin level of 0.20 ng/mL | 0
digoxin level of 3.6 ng/mL | 0
admitted to the Cardiac Intensive Care Unit | 0
given digoxin immune fab | 1
echocardiogram showed ejection fraction of 45% to 49% | 2
possible vegetation on the mitral valve | 2
severe eccentric mitral and tricuspid regurgitation | 2
transesophageal echocardiogram showed mitral valve vegetation | 4
severe biatrial enlargement | 4
left atrium volume of 101.40 mL/m2 | 4
right atrium volume of 233.80 mL/m2 | 4
blood cultures positive for Pasteurella multocida | 6
started ceftriaxone for Pasteurella septicemia | 6
head computed tomography showed numerous chronic infarctions | 12
patient owned 4 cats | 12
evaluated for multi-valve replacement surgery | 24
chose conservative treatment | 24
condition stabilized | 72
discharged to a skilled nursing facility | 72
started 6-week course of ceftriaxone | 72
readmitted for congestive heart failure exacerbation | 720
elected for hospice care | 720