75 years old | 0
male | 0
admitted to the hospital | 0
high fever | -24
cough | -24
sore throat | -24
upper respiratory tract infection | -24
dyspnea | 0
mental fog | 0
blood pressure 140/100 mm Hg | 0
pulse 109/min | 0
temperature 38.4 C° | 0
drowsiness | 0
PA chest x-ray | 0
Thorax CT | 0
arterial blood gas analysis | 0
PaO2 30 mmHg | 0
PaCO2 60 mmHg | 0
pH 7.27 | 0
FiO2 40% | 0
rapid-sequence intubation | 0
mechanical ventilation | 0
assist control mode | 0
tidal volume 600 mL | 0
FiO2 100% | 0
trigger 0.2 lit/min | 0
PEEP 5 mmHg | 0
antibiotic treatment | 0
leukocytosis 23000/μL | 0
CRP 50 mg/L | 0
ventilator mode changed to SIMV + PS | 24
tidal volume 550 mL | 24
respiratory rate 10/min | 24
FiO2 0.4-0.6 | 24
PEEP 5 mmHg | 24
PS 15 mmHg | 24
trigger 2 lit/min | 24
PS and respiratory rate decreased | 48
ventilator mode changed to PSV | 48
PS 8 mmHg | 48
blood gases normal | 72
disconnected from mechanical ventilator | 72
extubated | 72
non-invasive ventilation | 72
PaCO2 increased | 96
intubated again | 96
mechanical ventilator support | 96
neurology consultation | 96
anamnesis | 96
physical examination | 96
bilateral hemiptosis | 96
minimal restriction in eye movements | 96
complaints of weakness | -6720
inability | -6720
easy exhaustibility | -6720
occasional diplopia | -6720
chewing difficulty | -6720
diagnosed with COPD | -6720
COPD treatment discontinued | -6720
Neostigmine Methylsulphate administered | 96
spontaneous respiratory activity | 96
mechanical ventilator assisted inspiration | 96
tidal volumes increased | 96
spontaneous respiratory activity stopped | 141
mechanical ventilator controlled inspiration | 141
electromyoneurography | 141
motor and sensory nerve conductions normal | 141
muscle responses normal | 141
AChR Ab level 205 nmol/L | 141
pyridostigmine bromide administered | 141
IVIG administered | 141
serial blood gas analysis | 141
weaning process | 141
pyridostigmine bromide 180 mg/day | 168
azathioprine 100 mg/day | 168
complaints disappeared | 168
discharged | 168