67 years old | 0
man | 0
hypertension | 0
degenerative joint disease | 0
bilateral knee replacement | -109680
substance abuse | 0
recent history of trauma to his face | 0
recent history of trauma to his chest wall | 0
presented for new-onset lightheadedness | 0
presented for new-onset fatigue | 0
leukocytosis | 0
hemoglobin | 0
venous lactic acid | 0
noncontrast computerized tomography of chest/abdomen/pelvis | 0
intramuscular hematoma | 0
subpectoral hematoma | 0
acute right second through fifth anterior rib fractures | 0
bilateral lower lobe bronchopneumonia | 0
blood cultures obtained | 0
started on empiric antibiotics with intravenous piperacillin-tazobactam | 0
afebrile | 0
hypotensive | 0
blood pressure | 0
admitted to intensive care unit | 0
suspected septic shock | 0
initiation of vasopressors | 0
antibiotics broadened to intravenous vancomycin | 24
antibiotics broadened to intravenous cefepime | 24
antibiotics broadened to intravenous metronidazole | 24
repeat blood cultures obtained | 24
repeat urine cultures obtained | 24
repeat sputum cultures obtained | 24
blood cultures negative | 24
urine cultures negative | 24
sputum cultures grew methicillin-resistant Staphylococcus aureus | 24
antibiotics narrowed to intravenous vancomycin | 96
complained of left knee pain | 120
notable swelling on physical exam | 120
sterile left knee aspiration performed | 120
synovial fluid cloudy | 120
synovial fluid amber colored | 120
white blood cells | 120
calcium pyrophosphate crystals | 120
underwent complete washout and debridement of the joint | 144
retention of the prosthesis | 144
infected knee with purulence | 144
five cultures obtained | 144
joint specimen | 144
tissue specimen | 144
fluid specimen | 144
antibiotic regimen transitioned to intravenous cefazolin | 168
two sets of cultures grew Clostridium bifermentans | 192
antibiotic regimen transitioned to intravenous ampicillin-sulbactam | 192
oral suppression with amoxicillin-clavulanic acid | 192
contrast computerized tomography scan of abdomen | 192
human immunodeficiency virus screening | 192
discharged to rehabilitation facility | 384
referral to gastroenterology for outpatient colonoscopy | 384
recovered full range of motion of left knee | 2304
no signs of lingering joint infection | 2304
no signs of systemic infection | 2304
continued taking Augmentin | 2304
medication adherence | 2304
had not undergone colonoscopy | 2304
DAIR procedure | 144
intravenous antibiotics | 192
oral antibiotics | 192
risk of treatment failure | 2304
risk of recurrence | 2304
close follow-up | 2304
possible two-stage arthroplasty | 2304
