16 years old| 0
female | 0
syncope | -144
malaise | -144
fever | -144
fatigue | -144
chest pain | -144
shortness of breath | -144
presyncopal episode | -144
dizziness | -144
vision changes | -144
sweating | -144
true syncopal episode | -144
chipping tooth | -144
hypotension | 0
sinus tachycardia | 0
tachypnea | 0
admitted | 0
telemetry | 0
serial troponins | 0
troponin I elevation | 0
fluid refractory hypotension | 24
transferred to cardiac intensive care unit | 24
vasopressor support | 24
dopamine | 24
milrinone | 24
myocarditis | 24
viral sepsis | 24
influenza A positive | 24
peramivir | 24
increased pericardial effusion | 48
tamponade physiology | 48
pericardiocentesis | 48
pericardial drain placement | 48
increased respiratory effort | 48
hypoxemia | 48
biphasic positive airway pressure | 48
intravenous immunoglobulin | 48
improved | 120
weaned from intravenous infusions | 120
weaned from supplemental oxygen | 120
increased ejection fraction | 168
persistent concentric LVH | 168
symptoms resolved | 168
resolving LVH | 168
discharged | 168
normal biventricular chamber sizes | 2880
normal biventricular systolic function | 2880
normal LV mass | 2880
no LVH | 2880
no late gadolinium enhancement | 2880
resolution of LVH | 2880
