severe pain | -12
shortness of breath | -12
worsening pain over right thigh | -12
drowsy | -12
tachypneic | -12
oxygen saturation of 56% on room air | -12
tachycardia with a pulse of 121 bpm | -12
afebrile at 36 °C | -12
unrecordable blood pressure | -12
hypotensive with a blood pressure of 56/30 mmHg | -12
noradrenaline infusion started | -12
IV heparin 5000 units given | -12
IV amoxicillin-clavulanate given | -12
electively intubated | 0
metabolic and lactic acidosis | 0
worsening respiratory distress | 0
120 mL/kg of crystalloid given | 0
persistently hypotensive post-intubation | 0
adrenaline, vasopressin and dobutamine added | 0
grossly swollen right thigh with extensive blistering ecchymotic patches | 0
necrotizing fasciitis of the right thigh | 0
septicemic shock | 0
acute kidney injury | 0
rhabdomyolysis | 0
coagulopathy with thrombocytopenia | 0
ischemic hepatitis | 0
IV meropenem, IV clindamycin and IV vancomycin started | 0
high vaginal swab for culture and sensitivity taken | 0
CT pulmonary angiography done | 0
bedside echocardiography showed good contractility | 0
intravenous immunoglobulin given | 0
continuous veno-venous hemofiltration started | 0
lactic acidosis | 0
elevated creatinine kinase | 0
skin lesion spread over bilateral upper and lower limbs | 12
bluish discoloration | 12
blistering of bilateral lower limbs | 12
lesion on right upper limb | 12
high vaginal swab culture revealed Gram positive cocci in chains | 24
blister fluid culture revealed Gram positive cocci in chains | 24
blood culture positive for group A beta hemolytic streptococcus | 24
IV clindamycin restarted | 48
high dose of IV crystalline penicillin G given | 48
CVVH continued | 48
multidisciplinary discussion held | 48
diagnosis of group A streptococcal toxic shock syndrome with necrotizing fasciitis | 48
death | 72