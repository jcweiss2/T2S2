50 years old | 0
female | 0
relapsing idiopathic membranous nephropathy | 0
presented to hospital in August 2016 | 0
maculopapular rash | -168
received rituximab | -168
IMN first diagnosed in 2000 | -138240
complete remission with cyclophosphamide and prednisolone | -138240
remission maintained with methotrexate | -138240
intolerance to cyclosporine | -138240
presented with nephrotic syndrome in July 2016 | -288
intact renal function | -288
renal biopsy confirmed relapse | -288
new nodular changes consistent with early diabetic nephropathy | -288
serum antiphospholipase-A2 receptor antibody negative | -288
cumulative cyclophosphamide exposure concerns | -288
treatment with rituximab (two doses of 1000 mg a fortnight apart) | -288
trimethoprim-sulfamethoxazole started for Pneumocystis jirovecii pneumonia prophylaxis | -288
metformin for diabetes | -288
widespread maculopapular rash on admission | 0
rash involving face, torso, peripheries | 0
haemodynamically stable | 0
presumptive diagnosis of allergic urticaria | 0
commenced on prednisolone 30 mg | 0
commenced on cetirizine 10 mg | 0
commenced on promethazine 25 mg | 0
became hypotensive (systolic BP 70 mmHg) | 24
febrile (38.1°C) | 24
tachycardic (heart rate 110 bpm) | 24
developed generalized myalgias | 24
developed arthralgias | 24
developed cervical lymphadenopathy | 24
did not respond to fluid resuscitation | 24
admission to ICU | 24
inotropic support | 24
empirical antibiotics commenced | 24
intravenous hydrocortisone for anaphylactic shock | 24
leucocytosis (WBC 24.9 ×10^9/L) | 24
lymphocytosis (7.2 ×10^9/L) | 24
serum eosinophils normal (0.0 ×10^9/L) | 24
neutrophils normal (6.4 ×10^9/L) | 24
blood film demonstrated non-specific reactive leucocytosis | 24
C-reactive protein elevated (3581 nmol/L) | 24
C3 low (0.63 g/L) | 24
C4 normal (0.20 g/L) | 24
septic workup negative | 24
lactic acidosis (lactate 15 mmol/L; pH 7.12) | 24
acute kidney injury (creatinine 339 µmol/L) | 24
urine microscopy showed 36 ×10^6 red cells | 24
no pyuria | 24
procalcitonin levels not tested | 24
symptoms resolved within 48 hours | 72
inotropic support weaned within 24 hours | 72
renal function normalized | 72
Rituximab-induced serum sickness diagnosis | 72
antibiotics ceased | 72
hydrocortisone changed to prednisolone weaning course | 72
rechallenged with trimethoprim-sulfamethoxazole | 72
no issues with rechallenge | 72
arrangements for outpatient skin allergen testing | 72
discharged home | 72
no recurrence of symptoms over 3 months | 720
rash involving face, torso, peripheries |>
presented with nephrotic syndrome in July 2016 | -672
intact renal function | -672
renal biopsy confirmed relapse | -672
new nodular changes consistent with early diabetic nephropathy | -672
serum antiphospholipase-A2 receptor antibody negative | -672
cumulative cyclophosphamide exposure concerns | -672
treatment with rituximab (two doses of 1000 mg a fortnight apart) | -672
trimethoprim-sulfamethoxazole started for Pneumocystis jirovecii pneumonia prophylaxis | -672
metformin for diabetes | -672
symptoms resolved within 48 hours | 48
