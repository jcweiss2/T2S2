58 years old | 0
African American | 0
male | 0
admitted to the hospital | 0
alcohol abuse | -672
hepatitis C | -672
left hand swelling | -36
left hand pain | -36
malaise | -36
catfish injury | -48
nausea | -48
progressive nausea | -48
edema of the dorsum of the hand | 0
edema of the thenar eminence | 0
mild pain on active motion | 0
altered mental status | 0
compartment pressures measured | 4
duplex of the left upper extremity | 4
antibiotics initiated | 0
blood cultures obtained | 0
hand swelling increased | 4
digit flexion limited | 4
digit extension limited | 4
hypotensive | 8
intubation | 8
high-dose vasopressor support | 8
blood cultures revealed ET | 8
infectious disease consultation | 8
multiorgan failure | 36
significant swelling of entire upper extremity | 36
bullae formation | 36
epidermolysis | 36
ischemia to the fingertips | 36
bullae and swelling over the remaining extremities | 36
plastic surgery team consulted | 48
surgical exploration | 48
dorsal hand incised | 48
flexor/extensor compartments of the forearm incised | 48
serous fluid found | 48
normal muscle and soft tissue appearance | 48
skin and muscle biopsies | 48
no evidence of tissue necrosis | 48
intraoperative cultures negative | 48
multiorgan failure progressed | 72
severe acidosis | 72
hemodynamic instability | 72
expired | 120
history of catfish bone injury | -48
exposure to catfish | -48
fulminant tissue necrosis | 48
cellulitis | 36
skin changes | 36
broad-spectrum antibiotic treatment | 0
involvement of an infectious disease specialist | 8
early aggressive surgical exploration | 48
multiple premorbid conditions | -672
high potential for mortality | 0