19 years old | 0
asymptomatic | 0
gravida 4 | 0
para 3 | 0
Syrian | 0
preterm premature rupture of the membranes | 0
admitted to hospital | 0
white blood cell count within normal range | 0
C-reactive protein levels elevated | 0
ampicillin | 0
erythromycin | 0
amoxicillin | 48
dexamethasone | 48
delivered a female infant | 168
spontaneous vaginal delivery | 168
Apgar scores 6 and 8 | 168
intubated | 168
severe respiratory depression | 168
surfactant administered | 168
transferred to neonatal intensive care unit | 168
mechanical ventilation initiated | 168
temperature 36.9°C | 168
heart rate 127 beats per min | 168
weight 1.085g | 168
head circumference 26cm | 168
length 38cm | 168
hypotensive | 168
dobutamine infusion started | 168
high-frequency ventilation initiated | 168
early-onset sepsis suspected | 168
blood specimens for cultures obtained | 168
ampicillin | 168
gentamicin | 168
high WBC count | 168
neutrophils 48.8% | 168
attempt to extubate failed | 48
re-intubated | 48
Gram-negative coccobacilli detected | 144
Rose Bengal test positive | 144
ampicillin stopped | 144
rifampin started | 144
gentamicin continued | 144
serum agglutination test positive | 192
B. melitensis | 192
B. abortus | 192
ciprofloxacin added | 288
gentamicin discontinued | 408
meropenem added | 408
general condition improved | 408
nasal cannula | 408
total parenteral nutrition | 408
meropenem withdrawn | 576
ciprofloxacin continued | 576
rifampin continued | 576
nasal cannula removed | 840
preterm milk formula | 840
discharged | 912
intermittent headaches | -672
anorexia | -672
malaise | -672
profuse sweating | -672
abdominal pain | -672
urinary tract infection | -504
antibiotics for UTI | -504
frequent visits to family farm | -1008
consumed unpasteurized sheep milk | -1008
grandfather had brucellosis | -1008
grandfather received treatment for brucellosis | -1008