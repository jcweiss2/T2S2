60 years old | 0
male | 0
Honduran | 0
admitted to hospital | 0
acute delirium | 0
alcohol abuse | -672
hypertension | -672
hydrochlorothiazide | -672
MSSA bacteremia | 0
aortic valvular endocarditis | 0
disseminated septic emboli | 0
MSSA meningitis | 0
C6-7 osteomyelitis | 0
spinal abscess | 0
sternoclavicular joint abscess | 0
septic emboli infarcts in brain | 0
septic emboli infarcts in liver | 0
septic emboli infarcts in spleen | 0
septic emboli infarcts in kidneys | 0
aortic valve replacement | 0
upper GI bleeding | 24
duodenal ulcers | 24
visible vessels | 24
endoscopy | 24
epinephrine injection | 48
BICAP cauterization | 48
endoclipping of vessels | 48
hemospray with procoagulant | 48
argon plasma coagulation | 48
IR embolization of gastroduodenal artery | 72
IR embolization of superior pancreaticoduodenal arteries | 72
IR embolization of inferior pancreaticoduodenal arteries | 72
duodenal resection | 168
Whipple procedure | 168
total pancreatectomy | 168
splenectomy | 168
gastrojejunostomy | 192
hepaticojejunostomy | 192
CMV duodenitis | 168
viral cytopathic changes | 168
intranuclear inclusion bodies | 168
immunohistochemical stains for CMV | 168
CMV IgM antibodies nonreactive | 168
CMV IgG antibodies reactive | 168
DNA quantitative PCR for CMV negative | 168
HIV immunologic assay normal | 168
hepatitis B immunologic assay normal | 168
hepatitis C immunologic assay normal | 168
intravenous ganciclovir | 192
oral valganciclovir | 216
discharged | 720