36 years old | 0
    woman | 0
    subarachnoid haemorrhage | -6480
    right-sided middle cerebral artery aneurysm rupture | -6480
    secondary vasospastic malignant infarction of the right middle cerebral artery territory | -6480
    haemicraniectomy | -6480
    posthaemorrhagic cerebrospinal fluid circulatory dysfunction | -6480
    ventriculoperitoneal shunt implantation | -6480
    coma | -6480
    left-sided hemiparesis | -6480
    basic communication ability | -6480
    simple actions (e.g., drinking from a feeding cup) | -6480
    condition deterioration over several weeks | -6480
    unresponsive to external stimuli | -6480
    vegetative dysfunction (vomiting, extreme sweating, tachypnoea, tachycardia) | -6480
    correction of suspected overdrainage of ventriculoperitoneal shunt | -6480
    cranioplastic skull reconstruction | -6480
    unresponsive wakefulness syndrome | -6480
    weaned from respirator | -6480
    breathing spontaneously through tracheal cannula | -6480
    infected decubiti | -6480
    upper limb phlegmon | -6480
    pneumothorax | -6480
    anaemia | -6480
    anovesical fistula | -6480
    multiple infections (pneumonia, urinary tract infection, catheter-associated sepsis) | -6480
    prolonged ICU stay | -6480
    rhythmic myoclonus of right upper and lower limbs | -6480
    rhythmic myoclonus of mandible muscles and tongue | -6480
    tremor (differential diagnosis) | -6480
    levetiracetam 4 g/day | -6480
    valproic acid 300 mg/day | -6480
    clonazepam 1.5 mg/day | -6480
    no seizures | -6480
    no epileptic activity in EEGs | -6480
    transfer to university hospital for second opinion | 0
    cranial CT (no over/underdrainage of ventriculoperitoneal shunt) | 0
    brain MRI (superficial siderosis, laminar necrosis, temporal, frontal, opercular atrophies) | 0
    spinal MRI (no structural abnormalities) | 0
    FDG-PET (normal glucose metabolism except infarction area) | 0
    cerebrospinal fluid examination (normal cell counts, lactate, glucose, protein; negative autoimmune antibodies) | 0
    spasticity (50% movement restriction) | 0
    fixed contractions (50% movement restriction) | 0
    baclofen 30 mg/day (no effect) | 0
    intrathecal baclofen (no effect) | 0
    levetiracetam discontinuation | 0
    valproic acid discontinuation | 0
    clonazepam discontinuation | 0
    lamotrigine treatment | 0
    amantadine therapy (initiated with 100 mg/day, increased to 300 mg/day) | 0
    improvement in revised coma recovery scale (5 to 23 points) | 24
    speaking valve use | 24
    speech apraxia | 24
    retrograde amnesia | 24
    full orientation | 24
    adequate communication (2-6 word sentences) | 24
    active movements with muscle power 4/5 | 24
    reduced spasticity | 24
    resolved myoclonus (except rare agitated situations) | 24
    transfer to neurorehabilitation centre | 24
    fully oriented at 3 months follow-up | 2160
    improved general condition | 2160
    mild cognitive deficits | 2160
    decannulation | 2160
    autonomous eating of precut food | 2160
    ability to stand with help | 2160
    difficulty walking due to fixed contractions | 2160
    <|eot_id|>
    