73 years old | 0
    female | 0
    left nasal obstruction | -480
    left side facial pain | -480
    headache | -480
    COVID-19 infection | -720
    home isolation treatment | -720
    no steroid use | -720
    black mucopurulent secretion in the nose | 0
    oroantral ulcer perforating through the left side of the palate | 0
    histopathological examination revealing fungal hyphae | 0
    MRI showing maxillary sinusitis with erosive lesions and left oroantral fistula | 0
    endoscopic surgical debridement planned | 0
    AmB 5 mg/kg/day initiated | 0
    bronchial asthma | 0
    hypertension | 0
    uncontrolled diabetes mellitus | 0
    regular treatment | 0
    normal airway examination | 0
    total leucocyte count 14,000/μL | 0
    fasting blood sugar 246 mg/dL | 0
    HbA1c 10.9% | 0
    ECG normal | 0
    chest roentgenogram normal | 0
    echocardiography normal | 0
    pulmonary function test normal | 0
    preoperative optimisation with regular insulin | 0
    nebulisation with budesonide and salbutamol | 0
    antifungal (AmB) | 0
    antibiotics | 0
    blood sugar control | 0
    COVID-19 negative RT-PCR test | 0
    surgery with informed consent | 0
    intravenous fluid via right subclavian central line | 0
    standard monitoring (ECG, NBP, pulse oximetry) | 0
    glycopyrrolate 0.2 mg | 0
    fentanyl 100 μg | 0
    propofol induction | 0
    vecuronium | 0
    endotracheal tube placement | 0
    anaesthesia maintained with oxygen, nitrous oxide, isoflurane | 0
    capnography monitoring | 0
    neuromuscular monitoring | 0
    urine output monitoring | 0
    stable intraoperative condition | 0
    extubation after surgery | 0
    postoperative ICU management | 0
    monitoring renal parameters | 0
    monitoring blood sugar | 0
    no residual shortness of breath | 0
    no deranged PFTs | 0
    no stress cardiomyopathy | 0
    no myocardial injury | 0
    no hypercoagulable state | 0
    no prolonged corticosteroid use | 0
    no adrenal suppression | 0
    no perioperative hypotension | 0
    no succinylcholine use | 0
    no difficult mask ventilation | 0
    no endotracheal intubation difficulties | 0
    no epiglottitis | 0
    no supraglottic oedema | 0
    no blood transfusion needed | 0
    no inotropic support needed | 0
    no AmB-induced nephrotoxicity | 0
    no AmB-induced hypotension | 0
    no hypokalaemia | 0
    no hypomagnesemia | 0
    no arrhythmias | 0
    no fever | 0
    successful anaesthetic management | 0
    postoperative recovery | 0
    