53 years old|0
male|0
hospitalized with worsening diarrhea|0
hematochezia|0
weight loss|0
abdominal pain|0
petechial rash of the trunk|0
petechial rash of the arms|0
petechial rash of the neck|0
petechial rash of the face|0
petechial rash of the eyelids|0
reported 6 months of chronic diarrhea|-4320
intermittent hematochezia|-4320
13.5-18 kg weight loss|-4320
two weeks prior to presentation at our institution|-336
presented to an outside community hospital's emergency department|-336
underwent colonoscopy|-336
colonoscopy showed edematous, friable mucosa|-336
pathology report noted acute and chronic inflammation|-336
preserved glandular architecture|-336
suspicious for Crohn disease|-336
discharged from outside hospital|-336
scheduled follow-up for presumed Crohn disease|-336
worsening symptoms of nausea|-336
worsening symptoms of vomiting|-336
worsening symptoms of diarrhea|-336
worsening symptoms of dyspnea|-336
worsening symptoms of rash|-336
presented to emergency department at our institution|0
ill-appearing|0
diffusely tender abdomen|0
new petechial rash|0
lungs clear to auscultation bilaterally without wheezing|0
heart in regular rhythm with increased rate|0
no murmur|0
hypotensive|0
tachycardic|0
afebrile|0
non-hypoxic on room air|0
blood pressure dropped to 87/50 mmHg|0
required intravenous fluid resuscitation|0
anemia|0
Hgb 9.1 g/dL|0
Hct 27.9%|0
RDW 15.4%|0
MCV 80.9 fL|0
platelet count 233 k/μL|0
acute kidney injury|0
Cr 1.57 mg/dL|0
low calcium|0
Ca 7.7 mg/dL|0
elevated BUN|0
BUN 21 mg/dL|0
low albumin|0
albumin 1.9 g/dL|0
C-reactive protein 0.80 mg/dL|0
high stool lactoferrin|0
lactoferrin 332.15 μg/mL|0
high pro-BNP|0
pro-BNP 10212 pg/mL|0
low folate|0
low thiamine|0
proteinuria|0
protein 100 mg/dL|0
presence of numerous hyaline casts|0
presence of coarse granular casts|0
CT chest showed moderate pericardial effusion|0
CT chest showed trace pleural effusions|0
CT abdomen/pelvis showed moderate wall thickening of the small bowel loops|0
CT abdomen/pelvis showed moderate wall thickening of the colon|0
echocardiogram showed normal left ventricular ejection fraction|0
echocardiogram showed small to moderate sized circumferential pericardial effusion|0
no tamponade|0
suspected diagnosis of Crohn disease|0
dermatology evaluation of petechial skin rash|0
fat pad biopsy performed|0
esophagogastroduodenoscopy|0
colonoscopy with biopsies|0
biopsies from esophagus|0
biopsies from stomach|0
biopsies from duodenum|0
biopsies from terminal ileum|0
biopsies from colon|0
pink amorphous material in abdominal fat pad biopsy|0
pink amorphous material in gastrointestinal tract biopsies|0
elevated IgG|0
IgG 3412 mg/dL|0
low IgA|0
IgA 33 mg/dL|0
quantitative kappa 1090 mg/dL|0
quantitative lambda 22 mg/dL|0
kappa/lambda ratio 49.55|0
serum protein electrophoresis showed M-spike|0
immunofixation showed IgG kappa monoclonal gammopathy|0
abnormal kappa free light chain present|0
24-hour urine protein elevated|0
urine protein 745 mg/d|0
bone marrow biopsy|0
kappa-restricted plasma cell neoplasm|0
30%-40% cellularity|0
negative for amyloid|0
plasma cell FISH detected duplication of chromosome 1q|0
plasma cell FISH detected gain of chromosomes 5|0
plasma cell FISH detected gain of chromosomes 9|0
plasma cell FISH detected gain of chromosomes 15|0
peripheral blood smear identified early rouleaux formation|0
Congo red staining showed apple green birefringence|0
diagnosis of amyloidosis|0
amyloid typing confirmed kappa light chain type amyloidosis|0
received IV fluid|0
admitted to ICU|0
started on empiric antibiotics|0
antibiotics discontinued after negative blood cultures|0
received midodrine|0
hemoglobin dropped to 6.7 g/dL|0
required multiple blood product transfusions|0
received electrolyte supplementation|0
received folate supplementation|0
received thiamine supplementation|0
scheduled outpatient follow-up with hematology and oncology|0
stabilized and discharged|0
returned to emergency department with worsening shortness of breath|24
worsening nausea|24
worsening vomiting|24
worsening diarrhea|24
worsening fatigue|24
hypotensive to 83/53 mmHg|24
admitted to ICU|24
work up for bacteremia|24
work up for septic shock|24
started on cyclophosphamide|24
started on bortezomib|24
started on dexamethasone|24
stabilized and discharged|24
continued treatment outpatient|24
seven months prior presented to outpatient clinic|-5040
new onset diarrhea|-5040
intermittent scant hematochezia|-5040
denied dyspnea|-5040
denied weight loss|-5040
denied fatigue|-5040
denied rash|-5040
differential diagnosis of hemorrhoids|-5040
differential diagnosis of diverticulosis|-5040
differential diagnosis of malignancy|-5040
stable vital signs|-5040
Hgb 13.6 g/dL|-5040
caseinomacropeptide within normal limits|-5040
elevated total protein 8.6 g/dL|-5040
referred for colonoscopy|-5040
colonoscopy not completed|-5040
elevated immunoglobulin G|0
low immunoglobulin A|0
quantitative kappa and lambda imbalance|0
serum protein electrophoresis with M-spike|0
immunofixation confirmed IgG kappa monoclonal gammopathy|0
bone marrow biopsy showing plasma cell neoplasm|0
Congo red positive biopsies|0
final diagnosis of AL amyloidosis|0
initial diagnosis of Crohn disease|-336
hypotension requiring IV fluids|0
anemia requiring transfusions|0
electrolyte supplementation|0
petechial rash leading to fat pad biopsy|0
presence of pericardial effusion|0
pleural effusions|0
wall thickening of small bowel and colon|0
high pro-BNP indicating cardiac involvement|0
proteinuria indicating renal involvement|0
malabsorption suggested by low folate and thiamine|0
outpatient amyloidosis treatment initiation|24
admission to ICU|0
discharge home|24
return to emergency department|24
septic shock management|24
ongoing treatment with cyclophosphamide|24
ongoing treatment with bortezomib|24
ongoing treatment with dexamethasone|24
outpatient follow-up continuation|24
