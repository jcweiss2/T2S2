46 years old | 0
male | 0
chronic bilateral hip and leg pain | 0
left sacral fracture | -time unknown
sacro-iliac joint separation | -time unknown
tingling sensation | -time unknown
lancinating pain | -time unknown
pain intensity 8 mm | 0
motor weakness of the lower extremities | 0
sensory weakness of the lower extremities | 0
electromyography | -time unknown
nerve conduction velocity | -time unknown
left lumbosacral plexopathy | -time unknown
right chronic L5-S1 radiculopathy | -time unknown
acetaminophen/tramadol | -time unknown
imipramine | -time unknown
divalproate | -time unknown
pregabalin | -time unknown
lumbar sympathetic ganglion block | -time unknown
pethidine HCl | -time unknown
patient-controlled continuous epidural morphine infusion | -time unknown
satisfactory catheter placement | -time unknown
epidurogram | -time unknown
preservative free morphine | -time unknown
basal rate 0.5 ml/h | -time unknown
on-demand bolus dose 4.0 ml | -time unknown
lock out interval 30 minutes | -time unknown
20% pain reduction | -time unknown
basal rate increased to 1.0 ml/h | -time unknown
no further improvement in pain intensity | -time unknown
neuromodulation | 0
spinal cord stimulation | 0
implantation of an intrathecal morphine pump | 0
epidural PCA stopped | 0
lateral decubitus position | 0
skin preparation | 0
spinal needle insertion | 0
cerebrospinal fluid flow | 0
intrathecal morphine administration | 0
0.3 mg morphine sulfate | 0
60% pain reduction | 1
respiratory rate 17/min | 1
pain recurred | 8
VAS 7 | 8
tramadol 50 mg | 15
dysarthria | 15
drowsiness | 15
unresponsive | 21
respiratory rate 15/min | 25
blood pressure 88/54 mmHg | 25
pulse oximetry 69-71% | 25
oxygen mask | 25
transferred to intensive care unit | 25
naloxone 0.4 mg | 25
no improvement in mental state | 25
chest radiograph | 25
multifocal patchy consolidation | 25
aspiration pneumonia | 25
conservative therapy | 25
antibiotic therapy | 25
ventilation care | 25
blood gas within normal range | 72
mentally alert | 72
extubation | 72
chest radiograph improved | 72
discharged | 72
previous medication | 72
VAS score 7 | 72