33 years old | 0
    male | 0
    admitted to the hospital (First Affiliated Hospital of Sun Yat-sen University) | -72
    fever | -2160
    diarrhea | -2160
    unexplained anemia | -2160
    splenomegaly | -2160
    mechanical ventilation | -72
    respiratory failure | -72
    antibiotic treatment for suspected pneumonia | -72
    antibiotic treatment for suspected cholecystitis | -72
    diarrhea with watery stool | -62
    itraconazole | -62
    norvancomycin | -62
    colonoscopy | -56
    inflammatory colitis | -56
    CMV in colon biopsy | -56
    ganciclovir treatment | -56
    abdominal pain | -56
    bloating | -56
    body temperature returned to normal | -56
    diarrhea persisted | -56
    CMV negative in peripheral blood | -28
    bone marrow aspiration | -28
    no hemophagocytosis | -28
    improved total bilirubin | -28
    improved conjugated bilirubin | -28
    improved γ-GT | -28
    decreased fibrinogen | -28
    discharged from First Affiliated Hospital of Sun Yat-sen University | -3
    presented to First Affiliated Hospital of Guangzhou University of Chinese Medicine | 0
    fever (41.0°C) | 0
    jaundice | 0
    distended lower abdomen | 0
    hepatomegaly | 0
    splenomegaly | 0
    normal chest X-ray | 0
    nutritional support | 0
    anemia (hemoglobin 36 g/l) | 0
    hyperbilirubinemia | 0
    fever persisted (40°C) | 0
    transferred to ICU | 10
    CMV IgM negative | 10
    CD3+ 79.2% | 10
    CD4+ 38.2% | 10
    CD8+ 35.3% | 10
    T helper/suppressor ratio 1.08 | 10
    hemoglobin 39 g/l | 10
    red blood cell count 1.61×10^12/l | 10
    leukocyte count 2.67×10^9/l | 10
    platelet count 57×10^9/l | 10
    ferritin 7931.21 mg/l | 10
    total bilirubin 299.5 mmol/l | 10
    conjugated bilirubin 215.7 mmol/l | 10
    occult blood (++) in urinalysis | 10
    urinary bilirubin (++) | 10
    erythrocytes 10/HPF | 10
    splenomegaly on abdominal CT | 10
    gall bladder stones | 10
    inflammatory changes in gall bladder | 10
    hemophagocytosis in bone marrow | 10
    whole-body PET/CT scan negative | 10
    peripheral blood culture | 10
    bone marrow culture | 10
    L. pseudomesenteroides identified | 14
    stool culture negative for C. difficile | 14
    vancomycin-resistant | 14
    clindamycin-sensitive | 14
    clindamycin therapy | 14
    red blood cell transfusion | 14
    frozen plasma transfusion | 14
    parenteral nutrition | 14
    fever subsided (37.0°C) | 14
    afebrile | 21
    repeat blood culture positive for L. pseudomesenteroides | 24
    improved hemoglobin (77 g/l) | 19
    improved red blood cell count (3.05×10^12/l) | 19
    improved platelet count (139×10^9/l) | 19
    improved total bilirubin (71.5 mmol/l) | 19
    improved conjugated bilirubin (45.2 mmol/l) | 19
    normal body temperature (36.5°C) | 19
    reduced stool volume (350 ml/day) | 19
    repeat blood culture negative for L. pseudomesenteroides | 28
    discharged due to financial concern | 35
    telephone follow-up | 49
    negative blood culture | 49
    visited hospital 8 months later | 5040
    anemia (hemoglobin 89 g/l) | 5040
    no other complaints | 5040

    33 years old | 0
    male | 0
    admitted to the hospital (First Affiliated Hospital of Sun Yat-sen University) | -72
    fever | -2160
    diarrhea | -2160
    unexplained anemia | -2160
    splenomegaly | -2160
    mechanical ventilation | -72
    respiratory failure | -72
    antibiotic treatment for suspected pneumonia | -72
    antibiotic treatment for suspected cholecystitis | -72
    diarrhea with watery stool | -62
    itraconazole | -62
    norvancomycin | -62
    colonoscopy | -56
    inflammatory colitis | -56
    CMV in colon biopsy | -56
    ganciclovir treatment | -56
    abdominal pain | -56
    bloating | -56
    body temperature returned to normal | -56
    diarrhea persisted | -56
    CMV negative in peripheral blood | -28
    bone marrow aspiration | -28
    no hemophagocytosis | -28
    improved total bilirubin | -28
    improved conjugated bilirubin | -28
    improved γ-GT | -28
    decreased fibrinogen | -28
    discharged from First Affiliated Hospital of Sun Yat-sen University | -3
    presented to First Affiliated Hospital of Guangzhou University of Chinese Medicine | 0
    fever (41.0°C) | 0
    jaundice | 0
    distended lower abdomen | 0
    hepatomegaly | 0
    splenomegaly | 0
    normal chest X-ray | 0
    nutritional support | 0
    anemia (hemoglobin 36 g/l) | 0
    hyperbilirubinemia |9
    fever persisted (40°C) | 0
    transferred to ICU | 10
    CMV IgM negative | 10
    CD3+ 79.2% | 10
    CD4+ 38.2% | 10
    CD8+ 35.3% | 10
    T helper/suppressor ratio 1.08 | 10
    hemoglobin 39 g/l | 10
    red blood cell count 1.61×10^12/l | 10
    leukocyte count 2.67×10^9/l | 10
    platelet count 57×10^9/l | 10
    ferritin 7931.21 mg/l | 10
    total bilirubin 299.5 mmol/l | 10
    conjugated bilirubin 215.7 mmol/l | 10
    occult blood (++) in urinalysis | 10
    urinary bilirubin (++) | 10
    erythrocytes 10/HPF | 10
    splenomegaly on abdominal CT | 10
    gall bladder stones | 10
    inflammatory changes in gall bladder | 10
    hemophagocytosis in bone marrow | 10
    whole-body PET/CT scan negative | 10
    peripheral blood culture | 10
    bone marrow culture | 10
    L. pseudomesenteroides identified | 14
    stool culture negative for C. difficile | 14
    vancomycin-resistant | 14
    clindamycin-sensitive | 14
    clindamycin therapy | 14
    red blood cell transfusion | 14
    frozen plasma transfusion | 14
    parenteral nutrition | 14
    fever subsided (37.0°C) | 14
    afebrile | 21
    repeat blood culture positive for L. pseudomesenteroides | 24
    improved hemoglobin (77 g/l) | 19
    improved red blood cell count (3.05×10^12/l) | 19
    improved platelet count (139×10^9/l) | 19
    improved total bilirubin (71.5 mmol/l) | 19
    improved conjugated bilirubin (45.2 mmol/l) | 19
    normal body temperature (36.5°C) | 19
    reduced stool volume (350 ml/day) | 19
    repeat blood culture negative for L. pseudomesenteroides | 28
    discharged due to financial concern | 35
    telephone follow-up | 49
    negative blood culture | 49
    visited hospital 8 months later | 5040
    anemia (hemoglobin 89 g/l) | 5040
    no other complaints | 5040