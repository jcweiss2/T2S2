31 years old | 0
male | 0
Caucasian | 0
alcohol use disorder | 0
admitted to the hospital | 0
generalized fatigue | -168
weakness | -168
myalgias | -168
throat pain | -672
GAS pharyngitis | -672
azithromycin | -672
severe penicillin allergy | -672
fever | -168
chills | -168
nausea | -168
vomiting | -168
arthralgias | -168
febrile | 0
tachycardic | 0
neutrophilic leukocytosis | 0
thrombocytopenia | 0
hyponatremia | 0
abnormal liver enzymes | 0
elevated Nt-ProBNP | 0
negative HIV | 0
elevated troponin T | 0
COVID-19 test negative | 0
hepatic steatosis | 0
acute viral hepatitis panel negative | 0
bilateral striated nephrograms | 0
perinephric fat stranding | 0
bilateral pyelonephritis | 0
mild hepatosplenomegaly | 0
alcoholic hepatitis | 0
alcohol withdrawal | 0
high fevers | 24
worsening myalgias | 24
nausea | 24
vomiting | 24
leukocytosis | 24
thrombocytopenia | 24
acute hypoxic respiratory failure | 48
desaturation | 48
SpO2 78 % | 48
extensive diffuse and bilateral interstitial and alveolar markings | 48
ground-glass airspace consolidations | 48
GAS bacteremia | 48
erythromycin resistance | 48
inducible clindamycin resistance | 48
vancomycin | 48
cefepime | 48
doxycycline | 48
broad spectrum antibiotics | 48
non-invasive positive pressure ventilation | 72
transferred to hospital | 72
evaluated by pulmonary medicine | 72
evaluated by infectious diseases teams | 72
transthoracic echocardiogram | 72
left ventricular ejection fraction 55–60 % | 72
mildly thickened aortic valve | 72
severe aortic regurgitation | 72
Janeway lesions | 96
splinter hemorrhages | 96
conjunctival hemorrhages | 96
desquamative rash | 96
cardiac intensive care unit | 96
urgent valve surgery | 120
aortic root abscess | 120
partial aortic valve annuloplasty reconstruction | 120
incision and drainage of root abscess | 120
partial root repair | 120
intraoperative culture of the aortic valve | 120
gram positive cocci | 120
GAS | 120
recovered well | 168
repeat blood cultures sterile | 168
discharged home | 168
ceftriaxone | 168