18 years old | 0
female | 0
65 years old | 0
chief complaint of recurrent fever for more than 1 month | 0
nausea | 0
vomiting for 1 week | 0
no obvious induction of fever | -1 month
highest body temperature 38 ℃ | -1 month
no obvious clinical signs | -1 month
neutrophil count 6.96×10^9/L ↑ | 0
monocyte count 0.86×10^9/L ↑ | 0
lymphocyte percentage 14.9% ↓ | 0
red blood cell count 3.17×10^12/L ↓ | 0
hemoglobin content 87 g/L ↓ | 0
hematocrit 0.28 L/L ↓ | 0
average red blood cell hemoglobin concentration 312 g/L ↓ | 0
platelet count 363×10^9/L ↑ | 0
platelet distribution width 8.3 fl ↓ | 0
C-reactive protein (CRP) 52.01 mg/L ↑ | 0
megakaryocyte maturation disorder | 0
Klebsiella pneumoniae sepsis | 0
admitted to the hematology department | 0
diagnosed with secondary infectious thrombocytopenia, gram-negative bacilli septicemia (Klebsiella pneumoniae), liver abscess, bilateral lung inflammation, type 2 diabetes, and hypertension grade 3 (extremely high risk) | 0
vancomycin, caspofungin, dexamethasone, and posaconazole oral suspension for therapy | 0
liver abscess puncture and drainage treatment | 0
inflammatory indexes tested by laboratory tests decreased significantly after treatment | 0
light perception disappeared in the left eye | 0
eyelid redness and pain | 0
purulent secretion | 0
repeated fever | 0
left-sided headache | 0
endogenous endophthalmitis (left), orbital cellulitis (left), rubeosis iridis (left), exudative retinal detachment (left), and diabetic retinopathy (right) | 0
intravitreal injection with vancomycin and ceftazidime | 0
symptoms were relieved | 0
patient’s current systemic infection was under control | 0
left eyeball enucleation | 7
fever again after the operation | 7
anti-infection medicine including moxifloxacin and sulperazon | 7
temperature elevated again | 7
inflammation of both lungs, pericardial effusion, bilateral pleural thickening and effusion, and atelectasis in right inferior lobe | 12
liver cyst and liver abscess, right renal cyst, and myoma of the uterus | 12
hypertension for more than 10 years | -10 years
highest blood pressure 180/100 mmHg | -10 years
oral valsartan was applied to control blood pressure at 140/80 mmHg | -10 years
sepsis | 0
secondary thrombocytopenia | 0
liver abscess | 0
gram-negative bacilli sepsis (Klebsiella pneumoniae) | 0
infection of lumbar vertebrae | 0
mesenteric panniculitis | 0
pelvic effusion | 0
pericardial effusion | 0
suppurative endophthalmitis (left) | 0
orbital cellulitis (left) | 0
retinal detachment (left) | 0
choroidal detachment (left) | 0
type 2 diabetes retinopathy (right) | 0
cortical senile cataract (right, immature stage) | 0
type 2 diabetes | 0
type 2 diabetes nephropathy stage I | 0
type 2 diabetic peripheral neuropathy | 0
hypertension, grade 3 (extremely high risk) | 0
hepatic cyst | 0
renal cyst | 0
hypoproteinemia | 0
coronary atherosclerotic heart disease | 0
lacunar cerebral infarction | 0
moderate anemia | 0
risk of malnutrition | 0
convulsion with unconsciousness | 20
transferred to the respiratory intensive care unit with pharmaceutical care | 20
emergency CT examination revealed the lacunar infarction and encephalomalacia | 20
bilateral pleural effusion, and the lower lobe of the right lung was insufficiently inflated | 20
intracranial infection | 20
lumbar puncture was performed | 20
cerebrospinal fluid (CSF) was sent for biochemistry analysis and microbial metagenomic next-generation sequencing (mNGS) | 20
biochemistry analysis on 21 April | 21
glucose <1.1 mmol/L ↓ | 21
chlorine 108 mmol/L ↓ | 21
CSF protein >3,000 mg/L ↑ | 21
microbial mNGS results showed a high sequence of Klebsiella pneumoniae with drug-resistant gene SHV-type beta-lactamases (blaSHV) | 21
2 g meropenem every 8 hours (q8h) prolonged for 3 hours to treat intracranial infection | 21
body temperature, blood routine, and CRP were gradually improved | 21
CT examination on 18 May | 18
pulmonary edema and pleural effusion were gradually dissipated and absorbed | 18
CSF analyses performed on 23 May | 23
chlorine 119 mmol/L ↓ | 23
micro amount of proteins 1,107 mg/L ↑ | 23
microalbumin 816.3 mg/L ↑ | 23
immunoglobulin G 308.5 mg/L ↑ | 23
α2-macroglobulin 18.5 mg/L ↑ | 23
β2-microglobulin 2.67 mg/L ↑ | 23
discharged from the hospital | 31