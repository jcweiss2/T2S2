12 years old | 0
female | 0
cerebral palsy | 0
admitted to ICU | 0
decreased level of consciousness | 0
sepsis | 0
respiratory distress | 0
gastrointestinal bleeding | 0
hypoglycemia | 0
noninvasive ventilation | 0
wide spectrum antibiotics | 0
hypertonic glucose | 0
improved general condition | 0
larva escaped from nose | 240
nasal myiasis | 240
L. sericata | 240
pancytopenia | 0
Klebsiella pneumoniae | 0
larva collected | 240
larva preserved | 240
larva identified | 240
Ivermectin treatment | 240
no other worm detected | 336
discharged | 336 
nosocomial myiasis | 240 
L. sericata identified | 240 
third instar larva | 240 
larva length | 240 
larva width | 240 
body segments | 240 
spine band | 240 
pseudocephalon | 240 
anterior spiracles | 240 
posterior spiracles | 240 
L. sericata diagnosis | 240 
Ivermectin dose | 240 
Ivermectin repeated | 432 
informed consent | 0 
ethics committee approval | 0 
Research Center of Pediatric Infectious Diseases | 0 
Iran University of Medical Sciences | 0 
Tehran | 0 
Firoozabadi Hospital | 0 
Intensive Care Unit | 0 
nosocomial infection | 240 
myiasis | 240 
Diptera | 240 
Calliphoridae | 240 
Lucilia | 240 
L. sericata | 240 
L. cuprina | 240 
Chrysomyia | 240 
Cochliomyia | 240 
Sarcophagidae | 0 
Wohlfartia magnifica | 0 
L. illustris | 0 
L. caesar | 0 
L. richardsi | 0 
Klebsiella pneumoniae infection | 0 
sepsis | 0 
respiratory distress | 0 
gastrointestinal bleeding | 0 
hypoglycemia | 0 
pancytopenia | 0 
nosocomial myiasis rate | 0 
mortality rate | 0 
larval feeding stage | 0 
egg laying | 0 
larval stage | 0 
instar stage | 0 
larva development | 0 
temperature | 0 
detection of larva | 240 
ICU admission | 0 
ICU stay | 240 
hospital stay | 336 
discharge | 336 
treatment outcome | 336 
follow-up | 336 
L. sericata infestation | 240 
nosocomial infestation | 240 
myiasis diagnosis | 240 
L. sericata identification | 240 
larva morphology | 240 
larva identification | 240 
species identification | 240 
dipterans | 0 
myiasis species | 0 
Calliphoridae family | 0 
Sarcophagidae family | 0 
Lucilia species | 0 
L. sericata species | 0 
Cochliomyia species | 0 
Chrysomyia species | 0 
Wohlfartia species | 0 
L. illustris species | 0 
L. caesar species | 0 
L. richardsi species | 0 
Klebsiella pneumoniae species | 0 
bacterial infection | 0 
sepsis | 0 
respiratory distress | 0 
gastrointestinal bleeding | 0 
hypoglycemia | 0 
pancytopenia | 0 
nosocomial infection rate | 0 
mortality rate | 0 
larval development | 0 
egg laying | 0 
larval stage | 0 
instar stage | 0 
temperature | 0 
detection of larva | 240 
ICU admission | 0 
ICU stay | 240 
hospital stay | 336 
discharge | 336 
treatment outcome | 336 
follow-up | 336 
L. sericata infestation | 240 
nosocomial infestation | 240 
myiasis diagnosis | 240 
L. sericata identification | 240 
larva morphology | 240 
larva identification | 240 
species identification | 240 
dipterans | 0 
myiasis species | 0 
Calliphoridae family | 0 
Sarcophagidae family | 0 
Lucilia species | 0 
L. sericata species | 0 
Cochliomyia species | 0 
Chrysomyia species | 0 
Wohlfartia species | 0 
L. illustris species | 0 
L. caesar species | 0 
L. richardsi species | 0 
Klebsiella pneumoniae species | 0 
bacterial infection | 0 
sepsis | 0 
respiratory distress | 0 
gastrointestinal bleeding | 0 
hypoglycemia | 0 
pancytopenia | 0 
nosocomial infection rate | 0 
mortality rate | 0 
larval development | 0 
egg laying | 0 
larval stage | 0 
instar stage | 0 
temperature | 0 
detection of larva | 240 
ICU admission | 0 
ICU stay | 240 
hospital stay | 336 
discharge | 336 
treatment outcome | 336 
follow-up | 336 
L. sericata infestation | 240 
nosocomial infestation | 240 
myiasis diagnosis | 240 
L. sericata identification | 240 
larva morphology | 240 
larva identification | 240 
species identification | 240 
dipterans | 0 
myiasis species | 0 
Calliphoridae family | 0 
Sarcophagidae family | 0 
Lucilia species | 0 
L. sericata species | 0 
Cochliomyia species | 0 
Chrysomyia species | 0 
Wohlfartia species | 0 
L. illustris species | 0 
L. caesar species | 0 
L. richardsi species | 0 
Klebsiella pneumoniae species | 0 
bacterial infection | 0 
sepsis | 0 
respiratory distress | 0 
gastrointestinal bleeding | 0 
hypoglycemia | 0 
pancytopenia | 0 
nosocomial infection rate | 0 
mortality rate | 0 
larval development | 0 
egg laying | 0 
larval stage | 0 
instar stage | 0 
temperature | 0 
detection of larva | 240 
ICU admission | 0 
ICU stay | 240 
hospital stay | 336 
discharge | 336 
treatment outcome | 336 
follow-up | 336 
L. sericata infestation | 240 
nosocomial infestation | 240 
myiasis diagnosis | 240 
L. sericata identification | 240 
larva morphology | 240 
larva identification | 240 
species identification | 240 
dipterans | 0 
myiasis species | 0 
Calliphoridae family | 0 
Sarcophagidae family | 0 
Lucilia species | 0 
L. sericata species | 0 
Cochliomyia species | 0 
Chrysomyia species | 0 
Wohlfartia species | 0 
L. illustris species | 0 
L. caesar species | 0 
L. richardsi species | 0 
Klebsiella pneumoniae species | 0 
bacterial infection | 0 
sepsis | 0 
respiratory distress | 0 
gastrointestinal bleeding | 0 
hypoglycemia | 0 
pancytopenia | 0 
nosocomial infection rate | 0 
mortality rate | 0 
larval development | 0 
egg laying | 0 
larval stage | 0 
instar stage | 0 
temperature | 0 
detection of larva | 240 
ICU admission | 0 
ICU stay | 240 
hospital stay | 336 
discharge | 336 
treatment outcome | 336 
follow-up | 336 
L. sericata infestation | 240 
nosocomial infestation | 240 
myiasis diagnosis | 240 
L. sericata identification | 240 
larva morphology | 240 
larva identification | 240 
species identification | 240 
dipterans | 0 
myiasis species | 0 
Calliphoridae family | 0 
Sarcophagidae family | 0 
Lucilia species | 0 
L. sericata species | 0 
Cochliomyia species | 0 
Chrysomyia species | 0 
Wohlfartia species | 0 
L. illustris species | 0 
L. caesar species | 0 
L. richardsi species | 0 
Klebsiella pneumoniae species | 0 
bacterial infection | 0 
sepsis | 0 
respiratory distress | 0 
gastrointestinal bleeding | 0 
hypoglycemia | 0 
pancytopenia | 0 
nosocomial infection rate | 0 
mortality rate | 0 
larval development | 0 
egg laying | 0 
larval stage | 0 
instar stage | 0 
temperature | 0 
detection of larva | 240 
ICU admission | 0 
ICU stay | 240 
hospital stay | 336 
discharge | 336 
treatment outcome | 336 
follow-up | 336 
L. sericata infestation | 240 
nosocomial infestation | 240 
myiasis diagnosis | 240 
L. sericata identification | 240 
larva morphology | 240 
larva identification | 240 
species identification | 240 
dipterans | 0 
myiasis species | 0 
Calliphoridae family | 0 
Sarcophagidae family | 0 
Lucilia species | 0 
L. sericata species | 0 
Cochliomyia species | 0 
Chrysomyia species | 0 
Wohlfartia species | 0 
L. illustris species | 0 
L. caesar species | 0 
L. richardsi species | 0 
Klebsiella pneumoniae species | 0 
bacterial infection | 0 
sepsis | 0 
respiratory distress | 0 
gastrointestinal bleeding | 0 
hypoglycemia | 0 
pancytopenia | 0 
nosocomial infection rate | 0 
mortality rate | 0 
larval development | 0 
egg laying | 0 
larval stage | 0 
instar stage | 0 
temperature | 0 
detection of larva | 240 
ICU admission | 0 
ICU stay | 240 
hospital stay | 336 
discharge | 336 
treatment outcome | 336 
follow-up | 336 
L. sericata infestation | 240 
nosocomial infestation | 240 
myiasis diagnosis | 240 
L. sericata identification | 240 
larva morphology | 240 
larva identification | 240 
species identification | 240 
dipterans | 0 
myiasis species | 0 
Calliphoridae family | 0 
Sarcophagidae family | 0 
Lucilia species | 0 
L. sericata species | 0 
Cochliomyia species | 0 
Chrysomyia species | 0 
Wohlfartia species | 0 
L. illustris species | 0 
L. caesar species | 0 
L. richardsi species | 0 
Klebsiella pneumoniae species | 0 
bacterial infection | 0 
sepsis | 0 
respiratory distress | 0 
gastrointestinal bleeding | 0 
hypoglycemia | 0 
pancytopenia | 0 
nosocomial infection rate | 0 
mortality rate | 0 
larval development | 0 
egg laying | 0 
larval stage | 0 
instar stage | 0 
temperature | 0 
detection of larva | 240 
ICU admission | 0 
ICU stay | 240 
hospital stay | 336 
discharge | 336 
treatment outcome | 336 
follow-up | 336 
L. sericata infestation | 240 
nosocomial infestation | 240 
myiasis diagnosis | 240 
L. sericata identification | 240 
larva morphology | 240 
larva identification | 240 
species identification | 240 
dipterans | 0 
myiasis species | 0 
Calliphoridae family | 0 
Sarcophagidae family | 0 
Lucilia species | 0 
L. sericata species | 0 
Cochliomyia species | 0 
Chrysomyia species | 0 
Wohlfartia species | 0 
L. illustris species | 0 
L. caesar species | 0 
L. richardsi species | 0 
Klebsiella pneumoniae species | 0 
bacterial infection | 0 
sepsis | 0 
respiratory distress | 0 
gastrointestinal bleeding | 0 
hypoglycemia | 0 
pancytopenia | 0 
nosocomial infection rate | 0 
mortality rate | 0 
larval development | 0 
egg laying | 0 
larval stage | 0 
instar stage | 0 
temperature | 0 
detection of larva | 240 
ICU admission | 0 
ICU stay | 240 
hospital stay | 336 
discharge | 336 
treatment outcome | 336 
follow-up | 336 
L. sericata infestation | 240 
nosocomial infestation | 240 
myiasis diagnosis | 240 
L. sericata identification | 240 
larva morphology | 240 
larva identification | 240 
species identification | 240 
dipterans | 0 
myiasis species | 0 
Calliphoridae family | 0 
Sarcophagidae family | 0 
Lucilia species | 0 
L. sericata species | 0 
Cochliomyia species | 0 
Chrysomyia species | 0 
Wohlfartia species | 0 
L. illustris species | 0 
L. caesar species | 0 
L. richardsi species | 0 
Klebsiella pneumoniae species | 0 
bacterial infection | 0 
sepsis | 0 
respiratory distress | 0 
gastrointestinal bleeding | 0 
hypoglycemia | 0 
pancytopenia | 0 
nosocomial infection rate | 0 
mortality rate | 0 
larval development | 0 
egg laying | 0 
larval stage | 0 
instar stage | 0 
temperature | 0 
detection of larva | 240 
ICU admission | 0 
ICU stay | 240 
hospital stay | 336 
discharge | 336 
treatment outcome | 336 
follow-up | 336 
L. sericata infestation | 240 
nosocomial infestation | 240 
myiasis diagnosis | 240 
L. sericata identification | 240 
larva morphology | 240 
larva identification | 240 
species identification | 240 
dipterans | 0 
myiasis species | 0 
Calliphoridae family | 0 
Sarcophagidae family | 0 
Lucilia species | 0 
L. sericata species | 0 
Cochliomyia species | 0 
Chrysomyia species | 0 
Wohlfartia species | 0 
L. illustris species | 0 
L. caesar species | 0 
L. richardsi species | 0 
Klebsiella pneumoniae species | 0 
bacterial infection | 0 
sepsis | 0 
respiratory distress | 0 
gastrointestinal bleeding | 0 
hypoglycemia | 0 
pancytopenia | 0 
nosocomial infection rate | 0 
mortality rate | 0 
larval development | 0 
egg laying | 0 
larval stage | 0 
instar stage | 0 
temperature | 0 
detection of larva | 240 
ICU admission | 0 
ICU stay | 240 
hospital stay | 336 
discharge | 336 
treatment outcome | 336 
follow-up | 336 
L. sericata infestation | 240 
nosocomial infestation | 240 
myiasis diagnosis | 240 
L. sericata identification | 240 
larva morphology | 240 
larva identification | 240 
species identification | 240 
dipterans | 0 
myiasis species | 0 
Calliphoridae family | 0 
Sarcophagidae family | 0 
Lucilia species | 0 
L. sericata species | 0 
Cochliomyia species | 0 
Chrysomyia species | 0 
Wohlfartia species | 0 
L. illustris species | 0 
L. caesar species | 0 
L. richardsi species | 0 
Klebsiella pneumoniae species | 0 
bacterial infection | 0 
sepsis | 0 
respiratory distress | 0 
gastrointestinal bleeding | 0 
hypoglycemia | 0 
pancytopenia | 0 
nosocomial infection rate | 0 
mortality rate | 0 
larval development | 0 
egg laying | 0 
larval stage | 0 
instar stage | 0 
temperature | 0 
detection of larva | 240 
ICU admission | 0 
ICU stay | 240 
hospital stay | 336 
discharge | 336 
treatment outcome | 336 
follow-up | 336 
L. sericata infestation | 240 
nosocomial infestation | 240 
myiasis diagnosis | 240 
L. sericata identification | 240 
larva morphology | 240 
larva identification | 240 
species identification | 240 
dipterans | 0 
myiasis species | 0 
Calliphoridae family | 0 
Sarcophagidae family | 0 
Lucilia species | 0 
L. sericata species | 0 
Cochliomyia species | 0 
Chrysomyia species | 0 
Wohlfartia species | 0 
L. illustris species | 0 
L. caesar species | 0 
L. richardsi species | 0 
Klebsiella pneumoniae species | 0 
bacterial infection | 0 
sepsis | 0 
respiratory distress | 0 
gastrointestinal bleeding | 0 
hypoglycemia | 0 
pancytopenia | 0 
nosocomial infection rate | 0 
mortality rate | 0 
larval development | 0 
egg laying | 0 
larval stage | 0 
instar stage | 0 
temperature | 0 
detection of larva | 240 
ICU admission | 0 
ICU stay | 240 
hospital stay | 336 
discharge | 336 
treatment outcome | 336 
follow-up | 336 
L. sericata infestation | 240 
nosocomial infestation | 240 
myiasis diagnosis | 240 
L. sericata identification | 240 
larva morphology | 240 
larva identification | 240 
species identification | 240 
dipterans | 0 
myiasis species | 0 
Calliphoridae family | 0 
Sarcophagidae family | 0 
Lucilia species | 0 
L. sericata species | 0 
Cochliomyia species | 0 
Chrysomyia species | 0 
Wohlfartia species | 0 
L. illustris species | 0 
L. caesar species | 0 
L. richardsi species | 0 
Klebsiella pneumoniae species | 0 
bacterial infection | 0 
sepsis | 0 
respiratory distress | 0 
gastrointestinal bleeding | 0 
hypoglycemia | 0 
pancytopenia | 0 
nosocomial infection rate | 0 
mortality rate | 0 
larval development | 0 
egg laying | 0 
larval stage | 0 
instar stage | 0 
temperature | 0 
detection of larva | 240 
ICU admission | 0 
ICU stay | 240 
hospital stay | 336 
discharge | 336 
treatment outcome | 336 
follow-up | 336 
L. sericata infestation | 240 
nosocomial infestation | 240 
myiasis diagnosis | 240 
L. sericata identification | 240 
larva morphology | 240 
larva identification | 240 
species identification | 240 
dipterans | 0 
myiasis species | 0 
Calliphoridae family | 0 
Sarcophagidae family | 0 
Lucilia species | 0 
L. sericata species | 0 
Cochliomyia species | 0 
Chrysomyia species | 0 
Wohlfartia species | 0 
L. illustris species | 0 
L. caesar species | 0 
L. richardsi species | 0 
Klebsiella pneumoniae species | 0 
bacterial infection | 0 
sepsis | 0 
respiratory distress | 0 
gastrointestinal bleeding | 0 
hypoglycemia | 0 
pancytopenia | 0 
nosocomial infection rate | 0 
mortality rate | 0 
larval development | 0 
egg laying | 0 
larval stage | 0 
instar stage | 0 
temperature | 0 
detection of larva | 240 
ICU admission | 0 
ICU stay | 240 
hospital stay | 336 
discharge | 336 
treatment outcome | 336 
follow-up | 336 
L. sericata infestation | 240 
nosocomial infestation | 240 
myiasis diagnosis | 240 
L. sericata identification | 240 
larva morphology | 240 
larva identification | 240 
species identification | 240 
dipterans | 0 
myiasis species | 0 
Calliphoridae family | 0 
Sarcophagidae family | 0 
Lucilia species | 0 
L. sericata species | 0 
Cochliomyia species | 0 
Chrysomyia species | 0 
Wohlfartia species | 0 
L. illustris species | 0 
L. caesar species | 0 
L. richardsi species | 0 
Klebsiella pneumoniae species | 0 
bacterial infection | 0 
sepsis | 0 
respiratory distress | 0 
gastrointestinal bleeding | 0 
hypoglycemia | 0 
pancytopenia | 0 
nosocomial infection rate | 0 
mortality rate | 0 
larval development | 0 
egg laying | 0 
larval stage | 0 
instar stage | 0 
temperature | 0 
detection of larva | 240 
ICU admission | 0 
ICU stay | 240 
hospital stay | 336 
discharge | 336 
treatment outcome | 336 
follow-up | 336 
L. sericata infestation | 240 
nosocomial infestation | 240 
myiasis diagnosis | 240 
L. sericata identification | 240 
larva morphology | 240 
larva identification | 240 
species identification | 240 
dipterans | 0 
myiasis species | 0 
Calliphoridae family | 0 
Sarcophagidae family | 0 
Lucilia species | 0 
L. sericata species | 0 
Cochliomyia species | 0 
Chrysomyia species | 0 
Wohlfartia species | 0 
L. illustris species | 0 
L. caesar species | 0 
L. richardsi species | 0 
Klebsiella pneumoniae species | 0 
bacterial infection | 0 
sepsis | 0 
respiratory distress | 0 
gastrointestinal bleeding | 0 
hypoglycemia | 0 
pancytopenia | 0 
nosocomial infection rate | 0 
mortality rate | 0 
larval development | 0 
egg laying | 0 
larval stage | 0 
instar stage | 0 
temperature | 0 
detection of larva | 240 
ICU admission | 0 
ICU stay | 240 
hospital stay | 336 
discharge | 336 
treatment outcome | 336 
follow-up | 336 
L. sericata infestation | 240 
nosocomial infestation | 240 
myiasis diagnosis | 240 
L. sericata identification | 240 
larva morphology | 240 
larva identification | 240 
species identification | 240 
dipterans | 0 
myiasis species | 0 
Calliphoridae family | 0 
Sarcophagidae family | 0 
Lucilia species | 0 
L. sericata species | 0 
Cochliomyia species | 0 
Chrysomyia species | 0 
Wohlfartia species | 0 
L. illustris species | 0 
L. caesar species | 0 
L. richardsi species | 0 
Klebsiella pneumoniae species | 0 
bacterial infection | 0 
sepsis | 0 
respiratory distress | 0 
gastrointestinal bleeding | 0 
hypoglycemia | 0 
pancytopenia | 0 
nosocomial infection rate | 0 
mortality rate | 0 
larval development | 0 
egg laying | 0 
larval stage | 0 
instar stage | 0 
temperature | 0 
detection of larva | 240 
ICU admission | 0 
ICU stay | 240 
hospital stay | 336 
discharge | 336 
treatment outcome | 336 
follow-up | 336 
L. sericata infestation | 240 
nosocomial infestation | 240 
myiasis diagnosis | 240 
L. sericata identification | 240 
larva morphology | 240 
larva identification | 240 
species identification | 240 
dipterans | 0 
myiasis species | 0 
Calliphoridae family | 0 
Sarcophagidae family | 0 
Lucilia species | 0 
L. sericata species | 0 
Cochliomyia species | 0 
Chrysomyia species | 0 
Wohlfartia species | 0 
L. illustris species | 0 
L. caesar species | 0 
L. richardsi species | 0 
Klebsiella pneumoniae species | 0 
bacterial infection | 0 
sepsis | 0 
respiratory distress | 0 
gastrointestinal bleeding | 0 
hypoglycemia | 0 
pancytopenia | 0 
nosocomial infection rate | 0 
mortality rate | 0 
larval development | 0 
egg laying | 0 
larval stage | 0 
instar stage | 0 
temperature | 0 
detection of larva | 240 
ICU admission | 0 
ICU stay | 240 
hospital stay | 336 
discharge | 336 
treatment outcome | 336 
follow-up | 336 
L. sericata infestation | 240 
nosocomial infestation | 240 
myiasis diagnosis | 240 
L. sericata identification | 240 
larva morphology | 240 
larva identification | 240 
species identification | 240 
dipterans | 0 
myiasis species | 0 
Calliphoridae family | 0 
Sarcophagidae family | 0 
Lucilia species | 0 
L. sericata species | 0 
Cochliomyia species | 0 
Chrysomyia species | 0 
Wohlfartia species | 0 
L. illustris species | 0 
L. caesar species | 0 
L. richardsi species | 0 
Klebsiella pneumoniae species | 0 
bacterial infection | 0 
sepsis | 0 
respiratory distress | 0 
gastrointestinal bleeding | 0 
hypoglycemia | 0 
pancytopenia | 0 
nosocomial infection rate | 0 
mortality rate | 0 
larval development | 0 
egg laying | 0 
larval stage | 0 
instar stage | 0 
temperature | 0 
detection of larva | 240 
ICU admission | 0 
ICU stay | 240 
hospital stay | 336 
discharge | 336 
treatment outcome | 336 
follow-up | 336 
L. sericata infestation | 240 
nosocomial infestation | 240 
myiasis diagnosis | 240 
L. sericata identification | 240 
larva morphology | 240 
larva identification | 240 
species identification | 240 
dipterans | 0 
myiasis species | 0 
Calliphoridae family | 0 
Sarcophagidae family | 0 
Lucilia species | 0 
L. sericata species | 0 
Cochliomyia species | 0 
Chrysomyia species | 0 
Wohlfartia species | 0 
L. illustris species | 0 
L. caesar species | 0 
L. richardsi species | 0 
Klebsiella pneumoniae species | 0 
bacterial infection | 0 
sepsis | 0 
respiratory distress | 0 
gastrointestinal bleeding | 0 
hypoglycemia | 0 
pancytopenia | 0 
nosocomial infection rate | 0 
mortality rate | 0 
larval development | 0 
egg laying | 0 
larval stage | 0 
instar stage | 0 
temperature | 0 
detection of larva | 240 
ICU admission | 0 
ICU stay | 240 
hospital stay | 336 
discharge | 336 
treatment outcome | 336 
follow-up | 336 
L. sericata infestation | 240 
nosocomial infestation | 240 
myiasis diagnosis | 240 
L. sericata identification | 240 
larva morphology | 240 
larva identification | 240 
species identification | 240 
dipterans | 0 
myiasis species | 0 
Calliphoridae family | 0 
Sarcophagidae family | 0 
Lucilia species | 0 
L. sericata species | 0 
Cochliomyia species | 0 
Chrysomyia species | 0 
Wohlfartia species | 0 
L. illustris species | 0 
L. caesar species | 0 
L. richardsi species | 0 
Klebsiella pneumoniae species | 0 
bacterial infection | 0 
sepsis | 0 
respiratory distress | 0 
gastrointestinal bleeding | 0 
hypoglycemia | 0 
pancytopenia | 0 
nosocomial infection rate | 0 
mortality rate | 0 
larval development | 0 
egg laying | 0 
larval stage | 0 
instar stage | 0 
temperature | 0 
detection of larva | 240 
ICU admission | 0 
ICU stay | 240 
hospital stay | 336 
discharge | 336 
treatment outcome | 336 
follow-up | 336 
L. sericata infestation | 240 
nosocomial infestation | 240 
myiasis diagnosis | 240 
L. sericata identification | 240 
larva morphology | 240 
larva identification | 240 
species identification | 240 
dipterans | 0 
myiasis species | 0 
Calliphoridae family | 0 
Sarcophagidae family | 0 
Lucilia species | 0 
L. sericata species | 0 
Cochliomyia species | 0 
Chrysomyia species | 0 
Wohlfartia species | 0 
L. illustris species | 0 
L. caesar species | 0 
L. richardsi species | 0 
Klebsiella pneumoniae species | 0 
bacterial infection | 0 
sepsis | 0 
respiratory distress | 0 
gastrointestinal bleeding | 0 
hypoglycemia | 0 
pancytopenia | 0 
nosocomial infection rate | 0 
mortality rate | 0 
larval development | 0 
egg laying | 0 
larval stage | 0 
instar stage | 0 
temperature | 0 
detection of larva | 240 
ICU admission | 0 
ICU stay | 240 
hospital stay | 336 
discharge | 336 
treatment outcome | 336 
follow-up | 336 
L. sericata infestation | 240 
nosocomial infestation | 240 
myiasis diagnosis | 240 
L. sericata identification | 240 
larva morphology | 240 
larva identification | 240 
species identification | 240 
dipterans | 0 
myiasis species | 0 
Calliphoridae family | 0 
Sarcophagidae family | 0 
Lucilia species | 0 
L. sericata species | 0 
Cochliomyia species | 0 
Chrysomyia species | 0 
Wohlfartia species | 0 
L. illustris species | 0 
L. caesar species | 0 
L. richardsi species | 0 
Klebsiella pneumoniae species | 0 
bacterial infection | 0 
sepsis | 0 
respiratory distress | 0 
gastrointestinal bleeding | 0 
hypoglycemia | 0 
pancytopenia | 0 
nosocomial infection rate | 0 
mortality rate | 0 
larval development | 0 
egg laying | 0 
larval stage | 0 
instar stage | 0 
temperature | 0 
detection of larva | 240 
ICU admission | 0 
ICU stay | 240 
hospital stay | 336 
discharge | 336 
treatment outcome | 336 
follow-up | 336 
L. sericata infestation | 240 
nosocomial infestation | 240 
myiasis diagnosis | 240 
L. sericata identification | 240 
larva morphology | 240 
larva identification |