80 years old | 0
female | 0
admitted to the hospital | 0
right femur fracture | 0
5-year history of hypertension | -43800
antihypertensive agent | -43800
aspirin | -43800
obesity | 0
depression | 0
delirium symptoms | 0
brain computerized tomography (CT) | 0
severe stenosis of the middle cerebral artery (MCA) | 0
old localized infarction of the basal ganglia | 0
diffuse atrophy of the brain | 0
cardiomegaly | 0
1 degree A-V block | 0
ejection fraction of 65% | 0
preoperative PT/PTT | 0
INR | 0
arterial blood gas analysis (ABGA) | 0
scheduled to undergo total hip replacement surgery | 96
aspirin maintained | -72
aspirin discontinued | 72
spinal anesthesia administered | 96
unresponsive | 96
BP 70/40 mmHg | 96
HR 40-45 beats/min | 96
ephedrine administration | 96
epinephrine administration | 96
endotracheal intubation | 103
norepinephrine administration | 103
dopamine administration | 103
IV epinephrine administration | 103
ABGA | 103
central venous catheterization | 103
emergent TEE | 103
enlargement of the right atrium (RA) and right ventricle (RV) | 103
straightening of the interventricular septum | 103
hypokinesia | 103
IV heparine administration | 103
milrinone administration | 103
operation postponed | 103
transported to the ICU | 103
cardiopulmonary resuscitation | 123
chest 3 dimensional PTCA | 123
non-contrast brain CT | 123
low density ovoid thromboembolism | 123
enlargement of the right atrium and ventricle | 123
low density large acute infarct | 123
gyral swelling of the right insula and temporal lobe | 123
heart rate decreased to 30 beats/min | 215
resuscitation ineffective | 215
death | 215