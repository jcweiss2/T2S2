87 years old | 0
man | 0
presented to the emergency department | 0
epigastric discomfort | -12
burning sensation radiating to chest | -12
burning sensation radiating to left upper quadrant | -12
nausea | -12
watery, nonbloody emesis | -12
hiccupping | -12
denied chest pain | 0
denied fever | 0
denied diarrhea | 0
denied constipation | 0
denied sneezing | 0
denied coughing | 0
denied Valsalva maneuvers | 0
coronary artery disease | 0
angina | 0
valvular heart disease | 0
hypertension | 0
hyperlipidemia | 0
gout | 0
gastroesophageal reflux disease | 0
recent hospital admission for constipation | 0
denied autoimmune disease | 0
denied connective tissue disorder | 0
denied upper gastrointestinal endoscopy | 0
denied esophageal biopsy | 0
furosemide | 0
atenolol | 0
doxazosin | 0
nifedipine | 0
simvastatin | 0
nitroglycerin PRN | 0
omeprazole | 0
oxybutynin | 0
denied current smoking | 0
denied alcohol usage | 0
hypertension (170/74 mm Hg) | 0
afebrile | 0
slight abdominal distention | 0
sluggish bowel sounds | 0
soft abdomen | 0
nontender abdomen | 0
negative cardiac enzymes | 0
no acute electrocardiogram changes | 0
unremarkable laboratory studies | 0
contrast-enhanced CT of abdominal and pelvis | 0
diffuse dilation of small bowel | 0
diffuse dilation of stomach | 0
diffuse dilation of mid-to-distal esophagus | 0
esophageal pneumatosis | 0
no pneumomediastinum | 0
no pneumoperitoneum | 0
no other sites of pneumatosis | 0
upper gastrointestinal ileus | 0
small bowel ileus | 0
attempted esophagram | 0
nondiagnostic esophagram | 0
decompensate | 0
admitted to surgical intensive care unit | 0
nasogastric tube placement | 0
decompression of 1700 ccs nonbloody fluid | 0
bowel rest | 0
intravenous fluids | 0
close observation | 0
esophagram performed through NG tube | 4
negative for perforation | 4
unremarkable esophagram | 4
additional nasogastric tube decompression | 4
repeat CT examination | 11
complete resolution of esophageal pneumatosis | 11
interval improvement of upper gastrointestinal ileus | 11
septic on hospital day 2 | 48
started broad-spectrum antibiotics | 48
tracheal aspirates grew Klebsiella pneumoniae | 48
acute kidney injury | 48
adjusted antibiotic regimen | 48
resolved acute kidney injury | 48
discharged home | 288
tolerating regular oral diet | 288
