81 years old | 0
female | 0
admitted to the hospital | 0
hypertension | -672
dyslipidemia | -672
asthma | -672
degenerative valve disease | -672
acute precordial pain | 0
dyspnea | 0
nausea | 0
vomiting | 0
fever | 0
respiratory distress | 0
hypoxemia | 0
aspiration pneumonia | 0
amoxicillin | 0
clavulanate acid | 0
blood cultures | 0
elevated troponin level | 24
type 2 myocardial infarction | 24
transthoracic echocardiography | 24
degenerative valve disease | 24
moderate to severe aortic disease | 24
mitral valve calcification | 24
moderate insufficiency | 24
worsening dyspnea | 96
worsening hypoxia | 96
chest pain | 96
chest computed tomography | 96
extensive parenchymal consolidation | 96
meropenem | 96
azithromycin | 96
mechanical ventilation | 120
intensive care unit | 120
noradrenalin | 120
circulatory shock | 120
bilateral infiltrates | 192
bronchofibroscopy | 192
bronchial lavage | 192
sputum collection | 192
corticosteroids | 192
excessive post-infectious inflammatory process | 192
interstitial lung disease | 192
febrile | 216
progressive lung infiltrates | 216
steroids suspended | 216
transesophageal echocardiography | 384
P-MAIVF | 384
important degenerative valve disease | 384
severe aortic stenosis | 384
expansibility | 384
solution of continuity | 384
severe mitral regurgitation jet | 384
mass in the tricuspid valve | 384
infection | 384
death | 480