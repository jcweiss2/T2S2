51-year-old | 0
    male | 0
    admitted to the hospital | 0
    right chest pain | -1464
    back pain | -1464
    inactive condition | -1464
    no family history | 0
    no medical history | 0
    biopsy (needle aspiration) | -1464
    right lower pulmonary pseudotumor diagnosis | -1464
    wedge resection of the right lower lobe | -2088
    CT scan showing right lung mass | 0
    bone destruction of thoracic vertebrae 7, 8, 9 | 0
    suspected metastasis | 0
    multiple enlarged lymph nodes in right hilar | 0
    bilateral pleural hypertrophy | 0
    fibre cord signs in both lungs | 0
    lesions after resection of inflammatory pseudotumor | 0
    thoracic spine space diagnosis | 0
    previous conservative treatment deemed invalid | -168
    thoracic vertebral lesions removal | -168
    right lung lesions needle aspiration | -168
    acute and chronic purulent inflammations | -168
    inflammatory granulation | -168
    granuloma | -168
    tuberculosis exclusion | -168
    negative sputum culture | -168
    neutrophils in lung tissues | -168
    lymphocytes in lung tissues | -168
    monocytes in lung tissues | -168
    scattered eosinophils | -168
    multinucleated giant-cell infiltration | -168
    fibrinous exudation | -168
    organization in alveolar cavity | -168
    significant focal necrosis in thoracic vertebrae | -168
    neutrophil aggregation | -168
    abscesses | -168
    special infectious disease | -168
    non-caseating necrosis | -168
    tuberculosis exclusion | -168
    increased plasma cells | -168
    myeloma exclusion | -168
    sudden high fever (40°C) | 24
    antibiotics administration | 24
    antipyretic treatment | 24
    symptom improvement | 24
    left upper arm pain | 384
    CT imaging showing rib destruction | 384
    suspected malignant tumors | 384
    small right pleural effusion | 384
    left upper lobe solitary nodule | 384
    striped high-density shadows in right lung | 384
    multiple enlarged mediastinal lymph nodes | 384
    suspected malignant bone tumors in left humerus | 384
    left humeral tumor lesion removal | 576
    osteoma-like hyperplasia | 576
    hemorrhaging in bone marrow cavity | 576
    inflammatory granulation tissues | 576
    granulomas | 576
    no bacterial growth in culture | 576
    postoperative CT scan suggesting peripheral lung cancer | 672
    inflammatory pseudotumor suspected | 672
    soft tissue density mass in right lung | 672
    pain related to right lower lobe lesion | 672
    right lower lobe resection attempted | 720
    extensive adhesions | 720
    significant bleeding | 720
    suspected lung inflammatory pseudotumor | 720
    postoperative recovery | 720
    discharge after incision healing | 720
    second hospital admission | 1344
    enlarged left upper lobe nodules | 1344
    patched high-density shadows in right lung | 1344
    lung inflammatory pseudotumor diagnosis | 1344
    severe left humerus pain | 1344
    radiation therapy (20 Gy/10 F) | 1440
    reduced CT scan shadows | 1464
    prednisone acetate administration | 1464
    percutaneous puncture biopsy | 1584
    argon-helium knife ablation | 1584
    chronic inflammation of fibrous tissues | 1584
    compound cyclophosphamide administration | 2376
    bone marrow suppression | 2376
    discontinued cyclophosphamide | 2376
    hemoglobin drop (91 g/L to 71 g/L) | 2376
    discharge after symptom improvement | 2376
    third hospital admission | 2160
    postoperative inflammatory pseudotumor diagnosis | 2160
    lung infection | 2160
    perianal abscess | 2160
    enlarged left upper lobe tumor | 2160
    enlarged right lower lobe tumor | 2160
    absorbed interstitial lesions | 2160
    reduced pleural effusion | 2160
    3 cm perianal mass | 2160
    perianal abscess incision and drainage | 2208
    acute purulent inflammation | 2208
    necrosis | 2208
    granulation tissues | 2208
    Klebsiella pneumoniae sputum culture | 2208
    levofloxacin treatment | 2208
    negative sputum culture | 2208
    symptom improvement | 2208
    discharge after treatment | 2208
    fourth hospital admission | 2472
    severe anemia diagnosis | 2472
    red-blood cell transfusion | 2472
    nutritional support | 2472
    symptomatic treatment | 2472
    rhGCSF administration | 2472
    pulmonary infection treatment | 2472
    improved anemia | 2472
    discharge after treatment | 2472
    fifth hospital admission | 10560
    left humerus pain | 10560
    MRI indicating chronic osteomyelitis | 10560
    peripheral inflammatory pseudotumor with infection | 10560
    antibiotic treatment | 10560
    debridement of osteomyelitis | 10560
    broken gray soft tissue | 10560
    inflammatory granulation | 10560
    purulent necrosis | 10560
    supportive treatments | 10560
    lung infection | 10560
    urinary tract infection | 10560
    antibiotic therapy | 10560
    discharge after improvement | 10560
    sixth hospital admission |"10768
    breathing difficulties | 10768
    unconsciousness | 10768
    severe pneumonia diagnosis | 10768
    septic shock | 10768
    multiple organ dysfunction syndromes | 10768
    metabolic acidosis | 10768
    type II respiratory failure | 10768
    osteomyelitis of left humerus | 10768
    soft tissue infection | 10768
    urinary system infection | 10768
    hypoalbuminemia | 10768
    incomplete paralysis | 10768
    postoperative right pulmonary pseudotumor | 10768
    chest tightness | 10768
    intensive care admission | 10768
    active treatments | 10768
    no significant improvement | 10768
    death | 10776
    septic shock as cause of death | 10776
    