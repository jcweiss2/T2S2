79 years old | 0
woman | 0
abdominal pain | -672
nausea | -672
weight loss | -672
postprandial abdominal pain | -288
femoral-tibial bypass | -288
emergency department presentation | -168
constipation treatment | -168
discharge | -168
hemodynamic compromise | -24
imaging studies | -24
distal superior mesenteric artery occlusion | -24
mucosal wall changes | -24
acute bowel ischemia | -24
peripheral vascular disease | 0
coronary artery disease | 0
asthma | 0
rheumatoid arthritis | 0
hypertension | 0
hyperlipidemia | 0
type 2 diabetes | 0
hypothyroidism | 0
breast cancer | 0
smoking history | -182760
quit smoking | -182760
septic shock | 0
abdominal peritonitis | 0
hypoxemia | 0
hypotension | 0
electrocardiogram ST-segment elevations | 0
troponin level elevated | 0
SMA embolectomy | 0
resuscitation | 0
thromboembolectomy | 0
necrotic jejunum resection | 0
pathologic examination | 0
transesophageal echocardiography | 0
pulmonary vein thrombus | 0
left atrium thrombus | 0
biventricular dysfunction | 0
intensive care unit admission | 0
vasopressor support | 0
cardiac catheterization | 0
right coronary artery stenosis | 0
saphenous vein bypass graft stenosis | 0
additional abdominal surgeries | 24
bowel resection | 24
spindle cell carcinoma diagnosis | 336
right upper lobe mass | 336
pulmonary vein thrombus burden | 336
left atrium thrombus burden | 336
postoperative complications | 504
palliative measures | 504
hypothyroidism |# Updated Table
rheumatrial arthritis | 0
