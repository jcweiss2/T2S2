71 years old | 0
woman | 0
admitted to the emergency department | 0
painful abdominal mass | 0
malnourished | 0
poor hygiene | 0
febrile | 0
temperature of 38℃ | 0
pulse rate of 106 beats per minute | 0
no heart murmur | 0
no lung crackles | 0
clear breath sounds | 0
no abdominal tenderness | 0
no rebound tenderness | 0
large tender mass in the abdominal left upper quadrant | 0
hemoglobin 8.3 g/dl | 0
white blood cell count 17,510/ml | 0
89.3% neutrophils | 0
blood urea nitrogen 27.5 mg/dl | 0
creatinine 0.38 mg/dl | 0
sodium 142 mEq/L | 0
chloride 105 mEq/L | 0
potassium 3.2 mEq/L | 0
C-reactive protein 304 mg/L | 0
normal urinalysis | 0
no chest radiography abnormalities | 0
computed tomography abdomen showing large abscess pocket | 0
incised the mass | 0
drained large abscess | 0
diagnostic laparotomy | 0
midline incision | 0
observed huge gastric cancer invading abdominal wall | 0
no distant metastasis | 0
peritoneal cavity not contaminated | 0
dissection impossible due to cancer penetration into abdominal wall | 0
total gastrectomy | 0
resection of involved abdominal wall | 0
no remaining muscle or subcutaneous layer on left upper quadrant | 0
overlying skin not viable | 0
wet gauze packing of the wound | 0
D1 lymph node dissection | 0
patient hypotensive | 0
patient septic | 0
R1 status expected | 0
admitted to intensive care unit | 24
postoperative care | 24
resuscitation | 24
vital signs stable | 24
febrile | 24
temperature 38.8℃ | 24
chest radiography showing diffuse haziness | 24
pneumonia suspected | 24
intensive treatment | 24
broad-spectrum antibiotics | 24
parenteral nutrition | 24
observation for anastomosis leakage | 24
resumed oral intake | 72
chest radiography improvement of pneumonia | 168
moved to general ward | 192
resumed ambulation | 192
wet dressing of the wound continued | 192
abdominal binder used | 192
planned chemotherapy | 192
cancer growth progressed rapidly | 960
wound filled with growing cancer | 960
prognosis expected to deteriorate | 960
conservative management | 960
analgesics | 960
sedatives | 960
nutrition for palliation | 960
oral intake impossible | 1440
intestinal obstruction | 1440
died | 1968
multiorgan failure | 1968
sepsis | 1968
pneumonia | 1968
poorly differentiated adenocarcinoma | 1968
5 of 13 lymph nodes cancer-cell positive (N2) | 1968
T stage suspected T4a | 1968
cancer stage IIIB | 1968
