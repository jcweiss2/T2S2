37 weeks of gestation | 0  
    male neonate | 0  
    born via caesarean section | 0  
    breech presentation | 0  
    Apgar score 8 at 1st minute | 0  
    Apgar score 9 at 5th minute | 0  
    admitted to NICU | 0  
    chest retractions | 0  
    fever (38.5°C) | 0  
    pale | 0  
    moderate tachypnoea | 0  
    dyspnoea | 0  
    bilateral fine gasps | 0  
    accentuated bronchovascular markings | 0  
    WBC count 11.9 × 109/L | 0  
    polymorphonuclear cells 59.4% | 0  
    normal C-reactive protein | 0  
    sterile blood culture | 0  
    RSV type A identified | 0  
    nasopharyngeal samples negative for bacteria | 0  
    penicillin 150,000 IU/kg/die | 0  
    gentamicin 5 mg/kg/die | 0  
    nCPAP started | 0  
    increasing fraction of oxygen required | 0  
    i.v. systemic corticosteroids | 0  
    chest X-ray opacities upper right and hilar-perihilar left lung regions | 24  
    antibiotics discontinued | 96  
    clinical improvement | 96  
    sterile blood culture | 96  
    RSV detection in nasopharyngeal samples | 96  
    normal procalcitonin levels | 96  
    nCPAP replaced with high-flow nasal cannula | 96  
    clinical conditions worsened | 168  
    severe hypotension | 168  
    i.v. fluids | 168  
    catecholamine support | 168  
    septic shock | 168  
    chest X-ray massive opacification right upper and left lower lobes | 168  
    hypertrophic interventricular septum | 168  
    ampicillin 150 mg/kg/die | 168  
    gentamicin 5 mg/kg/die | 168  
    cefotaxime 100 mg/kg/die | 168  
    nCPAP re-started | 168  
    WBC count 23.2 × 109/L | 168  
    polymorphonuclear cells 77.7% | 168  
    C-reactive protein 15.2 mg/dL | 168  
    S. pneumoniae serotype 3 in blood culture | 168  
    sterile CSF culture | 168  
    i.v. cefotaxime for 10 days | 168  
    C-reactive protein normal | 408  
    procalcitonin normal | 408  
    nCPAP discontinued | 312  
    discharged home | 312  
    uneventful clinical course | 312  
    normal neurodevelopmental outcome at 18 months | 312  

