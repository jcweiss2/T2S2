57 years old | 0
    Hispanic man | 0
    coronary artery disease | -77760
    myocardial infarction | -77760
    ischemic dilated cardiomyopathy | -77760
    cardiac resynchronization therapy defibrillator | 0
    implanted 9 years ago | -77760
    generator change 6 months ago | -4320
    2-month history of erythema | -1440
    discomfort around left upper chest implant site | -1440
    edema | -1440
    serosanguinous drainage | -1440
    oral amoxicillin treatment | -1440
    nonbacteremic | 0
    afebrile | 0
    laboratory investigations within normal limits | 0
    echocardiography: reduced left ventricular systolic function | 0
    ejection fraction 20%–25% | 0
    global hypokinesis of left ventricle | 0
    no vegetations | 0
    preoperative computed tomography: leads scarred to lateral wall of superior vena cava | 0
    transvenous lead extraction | 0
    pocket capsule dissected out | 0
    device removed | 0
    coronary sinus lead extracted with gentle traction | 0
    right atrial leads extracted with laser assistance | 0
    16F laser sheath passed first coil of right ventricular lead | 0
    hypotensive | 0
    transesophageal echocardiography: large pericardial effusion | 0
    emergency midsternotomy performed | 0
    pericardium opened | 0
    significant blood obscuring operative field | 0
    bleeding manually controlled with pressure | 0
    cardiopulmonary bypass instituted | 0
    5-mm tear in superior cavoatrial junction | 0
    perforation in right atrium | 0
    oozing hematoma at innominate vein | 0
    lesions repaired with polypropylene sutures | 0
    right ventricular lead capped and abandoned | 0
    intra-aortic balloon pump placed through left femoral artery | 0
    hemodynamic instability | 0
    multiple blood transfusions | 0
    coagulopathy developed | 0
    cryoprecipitate transfusions | 0
    platelet transfusions | 0
    fresh frozen plasma transfusions | 0
    factor VII transfusions | 0
    bleeding under control | 0
    chest closed | 0
    26 units of blood products given | 0
    postoperative transfer to ICU | 24
    critical condition | 24
    severe cardiogenic shock | 24
    multiorgan failure | 24
    hypotensive (79/48 mm Hg) | 24
    pulse 99 beats/min | 24
    vasopressin required | 24
    epinephrine required | 24
    norepinephrine required (50 mcg/h) | 24
    hypoxic respiratory failure | 24
    mechanical ventilation dependent | 24
    liver failure managed with albumin | 24
    blood products given for coagulopathy | 24
    broad-spectrum antibiotics adjusted | 24
    oliguric | 24
    continuous venovenous hemodialysis for acute renal failure | 24
    bilateral symmetrical cyanotic changes to digits | 216
    vasopressor administration stopped | 216
    marked surface pallor | 216
    coldness in affected areas | 216
    upper-digit ischemia progressed to dry gangrene | 216
    lower-digit ischemia progressed to dry gangrene | 216
    dull pain | 216
    no ability to move fingers and toes | 216
    bilateral stiffness | 216
    2+ pitting edema | 216
    nonexistent capillary refill time | 216
    2+ peripheral pulses | 216
    Doppler study: flat waveforms on digits and toes | 216
    no proximal occlusion or stenosis | 216
    intra-aortic balloon pump removed | 168
    endotracheal tube removed | 168
    albumin discontinued | 264
    liver enzymes returned to normal | 264
    kidney function improved | 984
    hemodialysis stopped | 984
    mental status improved | 984
    sedation weaned | 984
    necrotic lesions treated with povidone; iodine dressings | 648
    debridement on POD 27 | 648
    negative-pressure wound therapy | 648
    continued drainage of purulent material | 648
    foul-smelling material from left infraclavicular site | 648
    stabilized | 1296
    transferred to our facility on POD 54 | 1296
    preoperative transesophageal echocardiography: ejection fraction 10%–15% | 1296
    laser extraction of retained lead on POD 58 | 1392
    60 mL pus drained from subfascial area | 1392
    antibiotic regimen started | 1392
    Enterobacter cloacae culture | 1392
    Staphylococcus epidermidis culture | 1392
    failed screening for subcutaneous implantable cardioverter-defibrillator | 1536
    transvenous implantable cardioverter-defibrillator implanted on POD 64 | 1536
    no signs of local infection | 1536
    no wet gangrene | 1536
    black skin changes | 1536
    demarcation lines | 1536
    frank mummification of digits and toes | 1536
    discharged on POD 77 | 1848
    amputation and debridement of necrotic feet on POD 106 | 2544
    amputation of fingers scheduled | 2544
    <|eot_id|>
    