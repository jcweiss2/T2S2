64 years old | 0
male | 0
hypertension | 0
hiatal hernia | 0
osteoarthritis | 0
admitted to the hospital | 0
acute worsening of chronic lower back pain | -336
progressive weakness in lower extremities | -336
subjective fevers | -336
temperature of 100.1°F | 0
leukocytosis of 25,500 | 0
neutrophils 89% | 0
sedimentation rate of 44 | 0
lactic acid 1.6 | 0
anion gap 18 | 0
crepitus in both knees | 0
limping gait | 0
Kernig’s sign and Brudzinski’s sign obscured | 0
chronic bilateral knee pain | 0
congenital deformation of right knee | 0
smoker of 40 pack-years | 0
occasional user of alcohol and marijuana | 0
denies intravenous drugs | 0
toxicology positive for oxycodone | 0
thoracic and lumbar spine CT scan | 0
multilevel central canal and bilateral neural foraminal compromise | 0
cavitary lesion in left lower lobe | 0
left inferior renal pole abnormalities | 0
blood cultures grew S. aureus | 0
started empirically on vancomycin | 0
TTE performed | 0
ejection fraction of 65% | 0
normal valves and no vegetations | 0
altered mental status | 48
nuchal rigidity | 48
lumbar puncture | 48
cerebrospinal fluid leukocytosis | 48
culture positive for S. aureus | 48
testing for HIV, HSV, and PPD | 48
negative results | 48
spine MRI | 48
osteomyelitis at T12-L1 | 48
renal infarcts | 48
continued to be febrile | 96
tachypnea | 144
hypoxia | 144
new systolic 2/6 murmur | 144
bilateral respiratory crackles | 144
new right hemiparesis | 144
upgoing babinski reflex | 144
switched to nafcillin | 72
head MRI | 144
multiple infarcts in non-vascular pattern | 144
TEE | 144
severe mitral and tricuspid regurgitations | 144
1.5 cm mobile vegetation on mitral valve | 144
transferred to intensive care unit | 144
nafcillin continued | 144
resolution of leukocytosis and fever | 240
mental status improved | 240
indications for emergent mitral valve replacement | 240
mitral and tricuspid valve replacements | 672
completed 8 weeks of nafcillin | 1344
discharged home | 1344
dual-chamber pacemaker | 1344