58 years old | 0
hypertensive | 0
male | 0
admitted with acute pancreatitis | 0
biliary etiology not established | 0
toxonutritive etiology not established | 0
laboratory values at admittance | 0
ultrasonography not beneficial | 0
CT showed mass in head of pancreas | 0
oncomarkers without pathological values | 0
PET-CT confirmed lesion in head of pancreas | 0
diagnosis of tumor of pancreatic head | 0
preoperative T2N0M0 | 0
surgical resection recommended | 0
standard pylorus-preserving Traverso-Longmire pancreatoduodenectomy performed | 0
pancreatic duct thin | 0
pancreas fine structure | 0
blood loss perioperatively 400 ml | 0
antibiotic prophylaxis administered | 0
postoperative hyperamylasemia | 0
octreotide administered for 5 days | 0
began nutrition p.o. on day 5 | 120
secretion from drains minimal volume | 120
drains removed on day 6 | 144
histology findings described moderately differentiated ductal adenocarcinoma | 0
discharged on day 11 | 264
postoperative complications grade II | 264
blood count before discharge | 264
outpatient follow-up on day 16 | 384
felt good | 384
realimented | 384
proton pump inhibitor initiated | 264
exocrine secretion substitution initiated | 264
sudden upper abdominal pain on day 18 | 432
chills | 432
shivers | 432
nausea | 432
came to emergency room | 432
laboratory tests showed HGB 112 | 432
melena appeared | 432
esophagogastroduodenoscopy revealed subcardial erosions | 432
digested blood in stomach | 432
coagula | 432
stagnation fluid | 432
acute bleeding not seen | 432
blood transfusions administered | 432
antiulcer therapy administered | 432
CT revealed mass adjoining stump of gastroduodenal artery | 432
CT angiography performed | 432
pseudoaneurysm discovered | 432
angiography confirmed bleeding | 432
implantation of stent graft selected | 432
stent graft implantation confirmed | 432
under observation at ICU | 432
no signs of continued hemorrhage | 432
stable vital signs | 432
melena ceased | 432
follow-up endoscopy showed no hemorrhage | 432
antiaggregation therapy initiated | 432
clopidogrel added | 432
7 blood transfusions administered within 48 hours | 432
completed postoperative radiochemotherapy | 12960
oncomarkers without pathological values |3
