28 years old | 0  
    male | 0  
    attended a health center with symptoms of fatigue | -24  
    anosmia | -24  
    dyspnea for progressively shorter efforts | -24  
    SpO2 levels were 55% | -24  
    improved to 75% with nasal cannula oxygen therapy | -24  
    hospitalized | -24  
    evaluated at an emergency department | -24  
    chest radiography ordered | -24  
    bilateral lung infiltrates | -24  
    RT-PCR swab tested positive for SARS-CoV-2 infection | -24  
    admitted in a COVID-19 infirmary unit | -24  
    non-invasive ventilation support was unsuccessful | -24  
    intubation | -24  
    invasive mechanical ventilation with ventral decubitus positioning | -24  
    Escherichia coli detected on sputum culture | 48  
    methicillin-sensitive Staphylococcus aureus detected on sputum culture | 48  
    confirmed superinfection | 48  
    prescription of an 8-day regimen of amoxicillin | 48  
    blood culture revealed methicillin-resistant Staphylococcus aureus | 48  
    dismissed | 48  
    steady clinical improvement | 48  
    extubated | 48  
    discharged | 48  
    attended the emergency department of our hospital | 168  
    complaints of retrosternal thoracalgia irradiating to the left upper limb | 168  
    started shortly after transfer from the intensive care unit to the infirmary in the previous hospital | 168  
    abduction limited due to pain complaints | 168  
    external rotation limited due to pain complaints | 168  
    soft tissue swelling of the shoulder | 168  
    soft tissue swelling of the arm | 168  
    fever | 168  
    increased levels of C-reactive protein | 168  
    hemoculture proved negative | 168  
    urine culture proved negative | 168  
    chest radiograph performed | 168  
    thoracic CT performed | 168  
    bilateral peripheral ground glass opacities | 168  
    greater involvement of the lower lobes | 168  
    admitted for further investigation and treatment planning | 168  
    previous blood culture had been dismissed | 168  
    gentamicin prescribed | 168  
    gentamicin administered throughout the whole length of hospital stay | 168  
    thoracic CT with intravenous contrast administration performed | 312  
    scapulohumeral synovitis | 312  
    multiple intra-muscular collections | 312  
    continuity with the glenohumeral joint | 312  
    scapulohumeral synovitis on the right shoulder | 312  
    less pronounced joint fluid on the right shoulder | 312  
    bilateral shoulder magnetic resonance imaging (MRI) with intravenous contrast administration performed | 384  
    persistent shoulder pain | 384  
    persistent shoulder weakness | 384  
    infraspinatus fossa collections on the left shoulder | 384  
    subscapular fossa collections on the left shoulder | 384  
    extending and communicating with the glenohumeral joint | 384  
    capsular thickening | 384  
    increased signal intensity post-gadolinium administration | 384  
    similar changes on the right shoulder | 384  
    less pronounced changes on the right shoulder | 384  
    suggestive of septic arthritis | 384  
    rotator cuff collections | 384  
    possibly associated with myonecrosis | 384  
    aspiration of the infraspinatus fossa collection performed | 384  
    20 cc of seropurulent fluid sent for analysis | 384  
    8,5 Fr drainage catheter left on the left infraspinatus collection | 384  
    removed the day after due to patient complaints of discomfort | 432  
    direct tests for Mycobacterium tuberculosis | 384  
    culture tests for Mycobacterium tuberculosis | 384  
    anaerobic bacteria tests | 384  
    aerobic bacteria tests | 384  
    negative tests | 384  
    improvement of left shoulder range of motion | 384  
    physical rehabilitation exercises | 384  
    transferred to another hospital | 432  
    indication to continue physical therapy | 432  
    rehabilitation exercises | 432  
    prolonged immobilization | 0  
    mechanical ventilation | 0  
    muscle atrophy | 0  
    risk factor for development of heterotopic ossification around the shoulder | 0  
    delirium | 0  
    lung damage | 0  
    muscle weakness | 0  
    long-term rehabilitation process | 0  
    rhabdomyolysis | 0  
    myalgia | 0  
    fatigue | 0  
    pigmenturia | 0  
    acute renal failure | 0  
    enlargement of the affected muscles | 0  
    heterogeneous and hypodense on CT | 0  
    hyperintense signal on fluid-sensitive sequences | 0  
    heterogeneous enhancement following intravenous contrast administration | 0  
    rim enhancement | 0  
    myonecrosis | 0  
    arthritis associated with COVID-19 infection | 0  
    muscle pain | 0  
    arthralgia | 0  
    chronic rheumatologic diseases triggered by COVID-19 infection | 0  
    serological tests | 0  
    joint fluid tests | 0  
    no known arthropathy | 0  
    no previous shoulder problems | 0  
    no episodes of arthritis reported | 0  
    no causative agent detected | 0  
    under an antibiotic regimen | 0  
    lab results may have been affected | 0  
    cause of bilateral shoulder arthritis remained unknown | 0  
    presumed of septic nature | 0  
    treated accordingly | 0  

    <|eot_id|>
    