19 years old | 0
male | 0
newly recruited army officer | 0
fever | -120
arthralgia | -120
myalgia | -120
headache | -120
intermittent productive cough | -120
yellowish sputum | -120
chest heaviness | -120
dyspnea | -120
diarrhea | -120
reducing oral intake | -120
denies history of travelling | -120
denies recent jungle activities | -120
stayed in the military base camp | -120
no past medical illness | -120
no previous hospitalization | -120
no previous medical treatment | -120
conscious | -120
dehydrated | -120
cold peripheries | -120
febrile | -120
hypotensive | -120
tachycardic | -120
tachypnoeic | -120
oxygen saturation 75-80% | -120
coarse crepitation | -120
tenderness at epigastric region | -120
palpable liver | -120
no cervical lymph nodes | -120
no inguinal lymph nodes | -120
no axillary lymph nodes | -120
haemoglobin 11.3 g/dL | -120
low white blood cell 0.5×10^6/L | -120
neutrophil predominance | -120
platelet count 80×10^6/L | -120
C-reactive protein 28.28 mg/dL | -120
acute kidney injury | -120
serum sodium 137 mmol/L | -120
potassium 3.7 mmol/L | -120
urea 14 mmol/L | -120
creatinine 206 μmol/L | -120
normal liver function tests | -120
serum albumin 22 g/dL | -120
creatinine kinase 351 IU/L | -120
negative Dengue NS-1 Antigen | -120
negative Dengue IgG | -120
negative Dengue IgM | -120
consolidation of right upper lobe | -120
consolidation of left lower lobe | -120
severe community acquired pneumonia | -120
acute kidney injury | -120
resuscitated with normal saline | -120
non-invasive ventilation | -120
hypotensive | -120
inotropic support | -120
ceftriaxone | -120
azithromycin | -120
intubation | -120
mechanical ventilation | -120
type 2 respiratory failure | -120
bronchoscopy | -120
copious amount of haemoserous and greenish secretion | -120
worsening consolidation | -120
abscess formation | -120
meropenem | -120
cloxacillin | -120
oseltamivir | -120
continuous venous-venous haemofiltration | -120
severe metabolic acidosis | -120
oliguric acute kidney injury | -120
persistent spiking of temperature | -120
worsening of septic parameters | -120
refractory hypotension | -120
succumbed | 72
MDR Acinetobacter baumannii | 72
positive for MDR Acinetobacter baumannii | 72
susceptible to polymyxin B | 72
minimum inhibitory concentration (MIC) 0.5 μg/ml | 72
tested resistance to penicillin group | 72
tested resistance to ampicillin/sulbactam | 72
tested resistance to third generation cephalosporins | 72
tested resistance to fluoroquinolone | 72
tested resistance to carbapenem group | 72
negative blood cultures | 72
negative atypical bacterial serologies | 72
negative Leptospiral serologies | 72
negative Hepatitis B/C serologies | 72
negative HIV serologies | 72
negative respiratory viruses screening | 72
tracheal aspiration positive for MDR Acinetobacter baumannii | 72
bronchoalveolar lavage positive for MDR Acinetobacter baumannii | 72