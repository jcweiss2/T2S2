11 years old | 0
female | 0
admitted to the hospital | 0
fever | 0
vomiting | 0
generalized abdominal pain | 0
rash on palms and trunk | 0
severe drowsiness | 0
lethargy | 0
no conjunctivitis | 0
no lymphadenopathy | 0
respiratory rate 25/min | 0
oxygen saturation 93% | 0
tachycardic | 0
hypotension | 0
abdomen tender to palpation | 0
right lower quadrant tenderness | 0
white blood cell count 13.5 × 10^3/μL | 0
red blood cell count 3.5–5.8 × 10^6/mm^3 | 0
erythrocyte sedimentation rate 82 mm/h | 0
C-reactive protein 298.5 mg/L | 0
procalcitonin 18.45 mcg/L | 0
abdominal ultrasound showing enlarged appendix | 0
appendectomy | 0
postoperative course toxic | 0
tachycardia | 0
hypotension | 0
fractional shortening | 0
oxygen therapy | 0
chest X-ray showing bronchopneumonia | 0
treatment with ceftriaxone and amikacin | 0
switched to imipenem | 0
positive history of contact with COVID-19 | 0
grandfather diagnosed with COVID-19 | -720
serologic test positive for SARS-CoV-2 IgG | 0
ferritin elevated | 0
IL6 elevated | 0
high-sensitivity troponin elevated | 0
D-dimer elevated | 0
enoxaparin initiated | 0
IV immunoglobulin administered | 24
aspirin administered | 24
condition worsened | 24
febrile | 24
anemic | 24
red blood cell transfusion | 48
pulse dosage of systemic corticosteroids | 48
re-evaluation of emerging shock | 48
aggravation of heart dysfunction | 48
echocardiogram showing decreased LV function | 48
septal hypokinesia | 48
ejection fraction 30% | 48
dobutamine added | 48
vasoactive drugs discontinued | 72
afebrile | 96
clinical symptoms improved | 96
arterial pressure stable | 96
no pathogenic agents detected | 96
histopathological examination showing catarrhal appendicitis | 96
D-dimer downward trend | 96
troponemia resolved | 96
inflammatory parameters normal | 96
LV function improved | 96
normal biventricular function | 96
no aneurysms observed | 96
discharged | 288
follow-up outpatient visit | 336
blood tests normalized | 336
COV-2 IgG elevated | 336
abdominal and cardiac ultrasounds normal | 336