7 years old | 0
boy | 0
referred to the University Children's Hospital Tuebingen | 0
second relapse of pre-B-ALL | 0
first relapse treated with allogeneic HSCT | -672
hemoglobin 8.5 g/dl | 0
thrombocytes 13.000/μl | 0
WBC 940/μl | 0
neutrophils 50/μl |.0
CRP 6.83 mg/dl | 0
ferritin 182 μg/dl | 0
chronically reduced general condition | 0
cachexia | 0
dry skin | 0
pallor | 0
multiple hematomas | 0
hepatosplenomegaly | 0
antibiotic chemoprophylaxis | 0
ceftriaxone | 0
teicoplanin | 0
acyclovir | 0
antifungal chemoprophylaxis | 0
caspofungin | 0
pain in the left flank | 0
continuous infusion of morphine | 0
pain aggravated | 120
ultrasound scan | 120
no pathology apart from hepatosplenomegaly | 120
day +5 of blinatumomab treatment | 120
somnolent | 144
sleepy | 144
overdose of morphine assumed | 144
dose reduction | 144
reacted with delay | 144
opened eyes when addressed | 144
cerebral side effect of blinatumomab presumed | 144
neurological condition worsened | 168
cerebral CT scan | 168
MRI scan | 168
multiple cerebral hemorrhages | 168
cardio-respiratory decompensation | 168
transferred to intensive care unit | 168
mechanical ventilation | 168
catecholamine therapy | 168
blinatumomab treatment stopped | 168
hemoglobin 6.7 g/dl | 168
thrombocytes 49.000/μl | 168
WBC 120/μl | 168
neutrophils 20/μl | 168
CRP 23.13 mg/dl | 168
ferritin 1439 μg/dl | 168
echocardiography | 168
multiple thrombi in left and right ventricle | 168
thromboembolic events presumed | 168
endocarditis with multiple septic embolisms suspected | 168
antibiotic regimen intensified | 168
meropenem | 168
teicoplanin | 168
gentamicin | 168
antimycotic treatment continued | 168
caspofungin 50 mg/day | 168
CT scans of thorax | 180
CT scans of abdomen | 180
CT scans of pelvis | 180
multiple systemic thromboembolic lesions | 180
ischemia | 180
bleeding | 180
infarction | 180
lungs | 180
heart | 180
kidneys | 180
liver | 180
intestines | 180
muscles | 180
bone marrow aspiration | 180
bone marrow aplasia | 180
lymphatic blasts | 180
cerebral pressure rising | 180
etiology unknown | 180
cerebral herniation | 192
died | 192
autopsy | 192
invasive mycosis | 192
R. pusillus | 192
macroscopic examination | 192
microscopic examination | 192
systemic fungal infection | 192
PCR-based identification | 192
cerebral lesions | 168
septic embolic infarctions | 168
bleeding | 168
right ventricular thrombi | 180
left ventricular thrombi | 180
coronary artery occlusion | 180
fungal hyphae in coronary artery | 180
multiple infarcts in left kidney | 180
tubular necrosis | 180
hemorrhagic infarct | 180
occluded artery | 180
fungal hyphae in vessel | 180
ulcerations in colon | 180
neutropenia | 0
disseminated disease | 180
disseminated mucormycosis | 180
fungal infection | 180
cerebral infiltration | 168
pulmonary mucormycosis | 180
systemic thromboembolic lesions | 180
septic embolic infarctions in multiple organs | 180
death | 192
autopsy findings | 192
PCR confirmation of R. pusillus | 192
no detection in tracheal secretion | 192
proof of R. pusillus in lungs | 192
other organs | 192
original location of infection unclear | 180
health care-related infection not excluded | 180
caspofungin prophylaxis | 0
lack of amphotericin B treatment | 168
delay in diagnosis | 168
active malignancy | 0
cytopenia | 0
fulminant mucormycosis | 180
blinatumomab treatment | 0
targeted therapy | 0
reduced immunocompetence after HSCT | -672
increased vulnerability to infections | 0
lack of prospective studies | 0
antifungal prophylaxis | 0
need for amphotericin B prophylaxis | 0
