76 years old| 0
male | 0
admitted to the hospital | 0
history of bladder cancer | 0
regional lymph node involvement | 0
Clostridium difficile infection | 0
vomiting | -72
watery diarrhea | -72
anorexia | -72
mild odynophagia | -72
recurrent CDI | -72
oral vancomycin | -72
minimal symptomatic improvement | -72
hypotensive | 0
blood pressure 80/40 mm Hg | 0
acute renal dysfunction | 0
lactic acidosis | 0
leukocytosis | 0
bandemia | 0
basilar atelectasis | 0
diffuse colonic wall-thickening | 0
peri-colonic fat-stranding | 0
normal saline boluses | 0
lactated ringers boluses | 0
norepinephrine titration | 0
broad-spectrum intravenous antibiotics | 0
clinical improvement | 0
admitted to medical ICU | 0
septic shock secondary to fulminant CDI | 0
excellent mental status | 0
urine output >0.5 mL/kg/hr | 0
resolving lactic acidosis | 0
unexplained back pain | 6
worsening shock | 6
multi-organ failure | 6
five vasopressors | 6
emergent endotracheal intubation | 6
orogastric tube placement | 6
bilateral hydropneumothorax | 6
pneumomediastinum | 6
bilateral chest tube placement | 6
dark fluid from pleural spaces | 6
suspected esophageal perforation | 6
pleural fluid amylase 2,238 units/L | 6
Gram-positive cocci and rods | 6
aerobic Gram-positive organisms | 6
shock complicated by progressive renal impairment | 6
mixed refractory acidemia | 6
continuous veno-venous hemodiafiltration | 6
mechanical ventilation | 6
vasopressor support | 6
condition stabilized | 6
CT chest suggestive of esophageal perforation | 24
air communicating from pleural spaces to distal esophagus | 24
orogastric tube penetrating into lesser sac of stomach | 24
extensive esophageal necrosis | 72
complete separation of lower esophagus from stomach | 72
endoscopic intervention | 72
unsutured metal stent deployment | 72
parental nutrition | 72
chest tubes maintained | 72
vasopressors titrated off | 168
dialysis discontinued | 168
extubated | 168
mediastinitis | 264
recurrent respiratory failure | 264
comfort-focused approach | 264
passed away | 264
resolving lactic acidosis |,0
