28 years old | 0
male | 0
admitted to the hospital | 0
hepatomegaly | 0
splenomegaly | 0
leukopenia | 0
thrombocytopenia | 0
Gilbert’s syndrome | 0
slightly elevated activity of aminotransferases | 0
increased total bilirubin level | 0
fever | 0
persistent dry cough | 0
Escherichia coli in urine culture | 0
Chlamydophila pneumoniae antigen in urine | 0
increased lactate dehydrogenase (LDH) activity | 0
recurrence of fever | -24
worsening of neutropenia | -24
steroid therapy initiated | -24
fever subsided | -24
leukocyte count increased | -24
persistent elevated activity of aminotransferases | -24
liver biopsy performed | -72
fever recurred | -72
severe abdominal pain | -72
enlargement of the liver | -72
enlargement of the spleen | -72
free fluid in the abdominal cavity | -72
rapid drop in hemoglobin concentration | -72
subcapsular rupture of spleen | -72
retroperitoneal enlarged lymph nodes | -72
splenectomy performed | -72
histopathological examination of lymph nodes | -72
transfusions required | -72
hematoma found | -72
laparotomy performed | -72
hemophagocytes present in aspiration biopsy | -72
significant increase in ferritinemia | -72
met HLH 04 criteria | -72
HScore evaluation | -72
treatment initiated with dexamethasone, etoposide, cyclosporine A | -72
multiple-organ failure | -72
died | 0
PTCL-NOS diagnosis confirmed | 0
