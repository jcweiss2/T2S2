52 years old | 0
male | 0
admitted to the hospital | 0
sore throat | -240
right laterocervical swelling | -240
diabetes | 0
no pharmacological allergies | 0
no psychosocial problems | 0
no family genetic disease | 0
inflammatory right laterocervical swelling | 0
indurated painful right laterocervical swelling | 0
marked trismus | 0
raised tongue | 0
right peritonsillar swelling | 0
very bad dentition | 0
early signs of sepsis | 0
low-grade temperature of 38.5 °C | 0
mild tachycardia | 0
hemoglobin 13,2 g/dl | 0
WBC: 13120/mm3 | 0
Absolute neutrophils 22530/mm3 | 0
C-reactive protein, 441.9 mg/l | 0
creatinine 76.5 mg/L | 0
urea: 0.69 g/L |,<|eot_id|>
mild tachycardia |' 0
urea: 0.69 g/L | 0
ASAT: 585 UI/l | 0
ALAT 607 UI/l | 0
PT: 48% | 0
fasting blood glucose: 3.05 g/L | 0
multidrug-resistant streptococcus intermedius | 0
right IJV thrombosis | 0
right tonsil abscess | 0
bilateral submandibular lymph nodes abscesses | 0
narrowing adjacent pharyngeal lumen | 0
emphysematous cervical cellulitis | 0
hospitalized | 0
multidisciplinary management | 0
no bacteremia | 0
no metastatic infectious lesions | 0
broad-spectrum antibiotic therapy | 0
intravenous amoxicillin/clavulanic acid | 0
intravenous metronidazole | 0
intravenous gentamycin | 0
daily puncture of right tonsil abscess | 0
anticoagulant therapy with Enoxaparin | 0
endobucal adenophlegmon incision | 0
drainage of pus | 0
improvement of trismus | 0
increase in lateral cervical tumefaction | 0
emphysematous cervical facial cellulitis | 0
drain collections under general anesthesia | 0
sebileau incision | 0
cervical facial collections | 0
communication with oral cavity | 0
necrosis of submandibular gland | 0
delbet drain placement | 0
closure of communications | 0
good tolerance to surgery | 0
post-operative antibiotics | 0
local care | 0
no complications postoperatively | 0
anticoagulated with heparin | 0
negative echocardiogram for endocarditis | 0
discharged | 288
