43 years old|0
male|0
diagnosed with grade II hepatocellular carcinoma|0
admitted to Zhongnan Hospital's organ transplant center|0
allogeneic liver transplantation|0
sent to the center's intensive care unit|0
treated with Tacrolimus FK506|0
treated with Mycophenolate mofetil|0
treated with prednisone|0
peripheral T cell count 181.68/μL|0
peripheral B cell count 59.57/μL|0
peripheral NK cell count 70.66/μL|0
P. sputorum bacteremia detected|0
blood samples collected on July 17|0
blood samples collected on July 20|0
serum procalcitonin 0.56 ng/mL|0
C-reactive protein 61.00 mg/L|0
peripheral neutrophil granulocyte percentage 96.8%|0
imipenem administered|0
ceftriaxone/tazobactam administered|0
infection controlled|336
very low serum PCT levels|336
normal peripheral Neu% 73.67%|336
liver cancer due to chronic hepatitis B virus infection|0
undergone allogeneic liver transplantation|0
immunosuppressive treatment|0
compromised immune function|0
severe underlying disease|0
surgery|0
immunosuppressive therapy|0
very low levels of peripheral T lymphocytes|0
very low levels of peripheral B lymphocytes|0
very low levels of peripheral NK lymphocytes|0
multi-drug resistant P. sputorum isolates|0
resistant to aztreonam|0
resistant to cefepime|0
resistant to ceftazidime|0
resistant to gentamicin|0
resistant to meropenem|0
resistant to tobramycin|0
susceptible to ceftriaxone|0
susceptible to ciprofloxacin|0
susceptible to imipenem|0
susceptible to levofloxacin|0
susceptible to minocycline|0
susceptible to piperacillin|0
susceptible to piperacillin-tazobactam|0
susceptible to tetracycline|0
susceptible to ticarcillin/clavulanic acid|0
susceptible to tigecycline|0
susceptible to trimethoprim|0
intermediate to amikacin|0
improved clinical condition|336
chronic hepatitis B virus infection|0
P. sputorum bacteremia|0
pro-inflammatory response|0
inflammatory response|0
lung dysfunction|0
pronounced pro-inflammatory response|0
overwhelming inflammatory response|0
compromised immune function contributes to bacteremia|0
multi-drug resistance|0
characteristic resistance profiles|0
successfully eliminated P. sputorum|336
improved after treatment|336
