60 years old | 0
female | 0
hepatitis C-related cirrhosis | -6720
recurrent hepatic encephalopathies | -6720
chronic portal vein thrombosis | -6720
liver transplantation | 0
construction of an end-to-side anastomosis | 0
end-to-end bile duct anastomosis | 0
massive venous bleeding | 0
iliac conduit construction | 0
normal liver graft function | 0
stenosis of the bile duct anastomosis | -720
biliary leakage | -720
elevated liver enzymes | -720
pigtail treatment | -720
FCSCEMS insertion | -360
persisting leakage | -360
stent extraction | -120
hepatitis C reinfection | -120
recurrent stenosis of the biliary anastomosis | -120
ERCP | -120
balloon dilatations | -120
pigtail placements | -120
stent placements | -120
biopsy-proven significant fibrosis | -6240
treatment with pegylated interferon and ribavirin | -6240
elective ERCP | 0
recovery of 3 plastic double-pigtails | 0
cholangiogram | 0
large portobiliary fistula | 0
hemobilia | 0
FCSEMS placement | 0
prophylactic antibiotic treatment with ciprofloxacin | 0
septic shock | 48
admission to the intensive care unit | 48
hemodynamic support | 48
empiric broad-spectrum antibiotic treatment | 48
computed tomography | 48
angiography | 48
chronic obliteration of the iliac conduit | 48
partial perfusion of the hepatic artery | 48
anuric kidney failure | 48
continuous venovenous hemofiltration | 48
intermittent hemodialysis | 48
evaluation for liver re-transplantation | 4032
FCSEMS replacement | 4032
extraction of the lying FCSEMS | 4032
no evidence of persisting leakage | 4032
no relevant stenosis | 4032
no further endoscopic intervention | 7200