25 years old | 0
Hispanic female | 0
presented to emergency center | 0
sudden onset severe neck pain | 0
headache | 0
fever of 101.4°F | 0
history of sacral myofibroblastic sarcoma | -336
underwent remote sacrectomy | -336
lumbopelvic fixation | -336
complicated course involving multiple hardware revisions | -336
hardware revisions at L2–L4 levels | -336
wound breakdown | -336
two weeks prior to presentation | -336
underwent iliac screw revision | -336
placement of intrathecal pain pump | -336
somnolent | 0
without focal motor deficits | 0
developed new-onset seizure | 0
given lorazepam 2 mg/mL IV | 0
given levetiracetam 1,500 mg IV | 0
head CT revealed nonspecific hypodensities | 0
hypodensities in right frontal lobe | 0
hypodensities in left parietal lobe | 0
hypodensities in left cerebellum | 0
lumbar puncture performed | 0
broad-spectrum antibiotics initiated | 0
suspected bacterial meningitis | 0
admitted to intensive care unit | 0
intubated | 0
depressed level of consciousness | 0
electroencephalogram showed mild generalized slowing | 0
left temporal dysfunction | 0
no epileptiform discharges | 0
CSF WBC count of 5,781 mm3 | 0
CSF protein 578 mg/dL | 0
CSF glucose <30 mg/dL | 0
Gram-negative rods seen on stains | 0
CSF multiplexed NAAT positive for E. coli | 0
BioFire CNS multiplex panel detected K1 strain of E. coli | 0
corticosteroids not administered | 0
underwent intrathecal pump removal | 0
wound culture around pump insertion revealed E. coli | 0
wound culture around pump insertion revealed Candida parapsilosis | 0
treated with fluconazole | 0
MRI brain with and without contrast obtained one day after admission | 24
MRI demonstrated multifocal bilateral cerebral cortically based nonenhancing diffusion restricting lesions | 24
bilateral cerebellar cortically based nonenhancing diffusion restricting lesions | 24
lesions consistent with cortical infarcts | 24
MR susceptibility within cortical infarcts compatible with microhemorrhage | 24
no leptomeningeal enhancement | 24
stroke workup pursued | 24
CT angiogram of head/neck showed no arterial occlusion | 24
no stenosis | 24
no dissection | 24
no vasospasm of circle of Willis vessels | 24
transthoracic echocardiogram unremarkable | 24
transesophageal echocardiogram not pursued | 24
MRI brain venogram revealed no dural venous sinus thrombosis | 24
cortical infarcts determined secondary to E. coli K1 meningitis-induced vasculopathy | 24
day 4 of admission | 96
successfully extubated | 96
neurologically intact | 96
mild encephalopathy | 96
no focal findings | 96
meropenem changed to ceftriaxone | 96
ceftriaxone at meningeal doses for 14 days | 96
suppressive therapy with 400 mg cefpodoxine twice daily | 96
discharged on day 16 after admission | 384
phenytoin | 384
ceftriaxone | 384
cefpodoxime | 384
four days later | 480
phenytoin stopped | 480
good recovery | 480
no neurological deficits | 480
septic emboli considered | 0
no cardiac abnormalities | 0
no carotid abnormalities | 0
infarction patterns atypical for septic emboli | 0
diagnosis followed IDSA guidelines | 0
standard treatment antimicrobial therapy | 0
given meropenem 2 g | 0
given fluconazole 800 mg IV | 0
meropenem switched to ceftriaxone 2 g | 96
no corticosteroid therapy | 0
no meningeal biopsy | 0
no delay in diagnosis and therapy | 0
successfully treated with appropriate antibiotic course | 384
no chronic neurological sequelae | 384
