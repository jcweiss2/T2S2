41 years old | 0
female | 0
Caucasian | 0
admitted to the hospital | 0
intermittent headaches | -504
dizziness | -504
visual disturbance | -504
weight loss | -168
epilepsy | -13200
Carbamazepine | -13200
headaches localized around the occipital cortex | -336
dizziness | -336
visual blurriness | -336
morning emesis | -336
unintentional weight loss | -168
initial presenting symptoms | -504
provisional diagnosis of occipital neuralgia | 0
Pregabalin | 0
discharged | 0
re-admitted | 504
worsening headache | 504
nausea | 504
vomiting | 504
bilateral double vision | 504
dry cough | 504
shortness of breath | 504
bilateral abducens nerve palsy | 504
community acquired pneumonia | 504
ceftriaxone | 504
doxycycline | 504
increased C-reactive protein | 504
chest radiograph | 504
right middle lobe consolidation | 504
inpatient MRI scan | 504
neurological opinion | 504
meningioma | 504
meningitis | 504
lumbar puncture | 504
high opening pressure | 504
high protein | 504
low glucose | 504
high white cell count | 504
positive cryptococcal titer | 504
Cerebrospinal fluid culture | 504
C. neoformans | 504
AmBisome liposomal | 504
5-fluorocytosine | 504
induction therapy | 504
fluconazole | 504
chest CT scan | 504
cryptoccoma | 504
bronchoscopy | 504
bronchial lavage | 504
lumbar percutaneous drainage | 504
Methicillin-resistant Staphylococcus aureus infection | 1008
vancomycin | 1008
rifampicin | 1008
removal of the drain | 1008
source control | 1008
initial presenting symptoms began to improve | 1008
cryptococcal clearance | 1008
transferred to the rehabilitation ward | 1008
Fluconazole | 1008
external ventricular drain | 1008
ventriculoperitoneal shunt | 1008
fever | 1512
worsening vision | 1512
confusion | 1512
non-localized headache | 1512
septic screen | 1512
repeated CSF analysis | 1512
MRI brain | 1512
gyro hyper-intensity | 1512
IV cefepime | 1512
IV vancomycin | 1512
endotracheal intubation | 1512
ICU | 1512
IRIS | 1512
high dose of IV steroids | 1512
oral prednisolone | 1512
remarkably improved | 1512
returned to the ward | 1512
visual evoked potential tests | 1512
normal baseline visual examination | 1512
bilateral optic neuropathy | 1512
legally blind | 1512
Hepatitis B | 0
HIV | 0
Hepatitis C antibodies | 0
past infection | 0
normal immunoglobulin levels | 0
normal complement levels | 0
discharged | 2016