35 years old | 0
male | 0
common variable immune deficiency (CVID) | 0
monthly maintenance intravenous immunoglobulin (IVIG) infusions | -168
admitted to an outside hospital | 0
fever | -720
headache | -720
progressive shortness of breath | -720
asthma | 0
hypertension | 0
depression | 0
lived in Missouri | 0
never travelled outside of United States | 0
swam in the Tennessee River | -1008
smoked 1.5 packs of cigarettes per day for 20 years | 0
occasionally consumed alcohol | 0
smoked marijuana | 0
son had CVID | 0
no other family members had known immune-deficiencies | 0
construction worker long ago | 0
presently disabled | 0
febrile | 0
tachycardic | 0
left maxillary sinus tenderness | 0
otherwise normal exam | 0
white blood cell count 1.0 × 10−3/μL | 0
neutrophils 36% | 0
lymphocytes 50% | 0
monocytes 14% | 0
hemoglobin 9.4 g/dL | 0
platelets 53 × 10−3/μL | 0
normal serum electrolytes | 0
normal renal function tests | 0
normal liver function tests | 0
chest X-ray chronic blunting of right costo-phrenic angle | 0
clear lung fields | 0
normal cardiac silhouette | 0
CT paranasal sinuses pan sinus mucosal thickening | 0
intravenous vancomycin | 0
ceftazidime | 0
levofloxacin | 0
negative blood cultures | 0
normal urinalysis | 0
negative tick-borne panel | 0
negative Ehrlichia PCR | 0
negative Rocky Mountain spotted fever IgG/IgM | 0
negative tularemia serology | 0
negative Lyme IgG/IgM | 0
negative Babesia serology | 0
negative CMV-PCR | 0
negative monospot | 0
bone marrow biopsy pancytopenia | 0
no blasts | 0
no organisms (acid fast and Giemsa stains) | 0
pancytopenia persisted | 0
fever persisted | 0
micafungin added | 0
transferred to our facility | 0
dyspneic | 0
temperature 39.4 °C | 0
heart rate 118/min | 0
oxygen saturation 93% on nasal oxygen at 11 L/min | 0
firm non-tender massive splenomegaly | 0
bilateral crackles in lower lung fields | 0
no rash | 0
no lymphadenopathy |:
