31 years old | 0
female | 0
pregnant | 0
admitted to the hospital | 0
fever | 0
sinus tachycardia | 0
shortness of breath | 48
cough with sputum | 48
hypoxemia | 48
oxygen therapy | 48
heart failure | 48
pink foaming sputum | 48
cyanosis | 48
emergency cesarean section | 72
cesarean section | 72
fetal heart rate slowed | 72
transferred to ICU | 72
left heart enlargement | 72
left ventricular systolic insufficiency | 72
moderate mitral valve insufficiency | 72
ejection fraction 43% | 72
peripartum cardiomyopathy | 72
bromocriptine | 72
oral heart failure therapies | 72
anticoagulants | 72
vasorelaxant agents | 72
diuretics | 72
cardiac arrest | 78
external cardiac compression | 78
CPR | 78
ECMO team arrival | 330
venoarterial ECMO | 330
right arteriotomy femoral venous cannula | 330
femoral arterial cannula | 330
perfusion distally within the femoral artery | 330
spontaneous circulation | 360
dobutamine | 360
milrinone | 360
intra-aortic balloon pump | 360
continuous renal replacement therapy | 360
activated clotting time | 360
neurological assessments | 360
cardiac function improvement | 360
EF value restored | 360
vital signs stable | 360
lactic acid reduced | 360
bleeding complications | 360
nasal cavity bleeding | 360
gastrointestinal bleeding | 360
incision bleeding | 360
thrombocytopenia | 360
anticoagulant reduction | 360
allogeneic platelet infusion | 360
ECMO assistance stopped | 216
pupils differed in size | 216
cranial computed tomography | 216
intracranial hemorrhage | 216
cranial decompression | 216
intracranial hematoma removal | 216
conscious | 240
recurrent intracerebral hemorrhage | 288
surgery | 288
recovered | 1440
discharged | 1440
follow-up | 8760
good recovery | 8760
returned to work | 8760