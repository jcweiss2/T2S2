60 years old | 0
male | 0
arterial hypertension | -672
fever | -384
chills | -384
malaise | -384
fatigue | -384
anorexia | -384
left flank pain | -384
nausea | -384
vomiting | -384
diarrhea | -384
amoxicillin-clavulanic acid | -336
fever persisted | -336
rash | -336
malaise worsened | -336
fatigue worsened | -336
left flank pain worsened | -336
hematuria | -336
diarrhea reappeared | -336
sepsis | 0
febrile | 0
hypotensive | 0
tachypneic | 0
tachycardic | 0
abdominal ultrasound | 0
enlarged left kidney | 0
leukocytosis | 0
neutrophilia | 0
elevated C-reactive protein | 0
elevated procalcitonin | 0
elevated creatinine | 0
elevated urea | 0
pyelonephritis | 0
parenteral fluids | 0
antimicrobial therapy | 0
cefotaxime | 0
blood culture | 0
urine culture | 0
Salmonella enterica | 0
serovar Enteritidis | 0
resistant to cefuroxime | 0
resistant to ciprofloxacin | 0
resistant to gentamicin | 0
resistant to amikacin | 0
susceptible to ampicillin | 0
susceptible to cefotaxime | 0
susceptible to meropenem | 0
susceptible to trimethoprim/sulfamethoxazole | 0
Clostridioides difficile | 0
positive antigen | 0
positive toxin | 0
trimethoprim/sulfamethoxazole | 0
oral vancomycin | 0
transthoracic echocardiography | 0
native computed tomography | 0
discrete inflammatory changes | 0
fat around the left kidney | 0
discharged | 240
antimicrobial therapy stopped | 264
progressive weakness | 288
night sweating | 288
dull pain | 288
lumbar region | 288
sacral region | 288
elevated CRP | 288
admitted | 288
therapy started | 288
ceftriaxone | 288
oral vancomycin | 288
follow-up blood culture | 288
Salmonella enterica | 288
magnetic resonance imaging | 288
lumbar spine | 288
dilatation of the infrarenal part | 288
abdominal aorta | 288
contrast CT | 288
fusiform aneurysm | 288
abdominal aorta | 288
aneurysm of the left internal iliac artery | 288
saccular shape | 288
compressing the left ureter | 288
dilated left kidney | 288
grade 2 hydronephrosis | 288
vascular surgeons | 288
conservative therapy | 288
ceftriaxone | 288
CT follow-up | 432
progression of the aneurysm diameter | 432
infrarenal aorta recanalized | 432
surgery | 480
ligation of the left internal iliac artery | 480
partial extirpation of the aneurysm | 480
histologic examination | 480
nonspecific inflammation | 480
sterile cultures | 480
parenteral antimicrobial therapy | 480
CT follow-up | 528
complete obliteration | 528
residual aneurysm | 528
discharged | 576
oral therapy | 576
trimethoprim/sulfamethoxazole | 576
CRP level normalized | 624
asymptomatic | 2160
CRP level in reference range | 2160