80 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
non-smoker | 0 | 0 | Factual
hypertension | 0 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
acute dyspnea | -24 | 0 | Factual
fecal incontinence | -6.67 | -6.67 | Factual
left hemiplegia | -6.67 | -6.67 | Factual
dextroversion | -6.67 | -6.67 | Factual
dysarthria | -6.67 | -6.67 | Factual
vomiting | -6.67 | -6.67 | Factual
impaired consciousness | -6.67 | 0 | Factual
Japan coma scale score of Ⅱ-10 | -6.67 | 0 | Factual
right thalamus and putamen bleeding | -6.67 | 0 | Factual
Glasgow coma scale score 12 | 0 | 0 | Factual
systolic blood pressure 91 mmHg | 0 | 0 | Factual
respiratory rate 24/min | 0 | 0 | Factual
oxygen saturation of arterial blood (SpO2) 86% | 0 | 0 | Factual
poor oral hygiene | 0 | 0 | Factual
diminished breath sounds on the left side | 0 | 0 | Factual
coarse crackles in the right lung | 0 | 0 | Factual
decrease in breath sounds in the front of the chest | 0 | 0 | Factual
respiratory condition deteriorated | 0 | 0 | Factual
endotracheal intubation | 0 | 0 | Factual
mechanical ventilation | 0 | 0 | Factual
bilateral infiltration | 0 | 0 | Factual
admitted to the intensive care unit (ICU) | 0 | 0 | Factual
decreased leukocyte count | 0 | 0 | Factual
mildly elevated C-reactive protein (CRP) level | 0 | 0 | Factual
respiratory failure | 0 | 0 | Factual
partial pressure of oxygen in arterial blood (PaO2) 64 mmHg | 0 | 0 | Factual
hepatorenal function normal | 0 | 0 | Factual
extensive infiltration shadows on chest radiography | 0 | 0 | Factual
hematoma extending from the right basal ganglia and putamen to the thalamus | 0 | 0 | Factual
cerebral edema | 0 | 0 | Factual
consolidations admixture with ground-glass opacities on chest CT | 0 | 0 | Factual
A-DROP score corresponded to patient age | 0 | 0 | Factual
increased blood urea nitrogen | 0 | 0 | Factual
decreased SpO2 | 0 | 0 | Factual
impaired consciousness | 0 | 0 | Factual
antigen test for coronavirus disease 2019 negative | 0 | 0 | Factual
Mendelson's syndrome | 0 | 0 | Factual
aspiration bacterial pneumonia | 0 | 0 | Factual
sputum culture showed Streptococcus agalactiae and Klebsiella oxytoca | 0 | 0 | Factual
leukocytopenia | 0 | 0 | Factual
low serum CRP level | 0 | 0 | Factual
respiratory viral pneumonia | 0 | 0 | Possible
management in the ventilator mode | 0 | 288 | Factual
meropenem | 0 | 288 | Factual
levofloxacin | 0 | 288 | Factual
Sivelestat sodium hydrate | 0 | 288 | Factual
lung-protection strategies | 0 | 288 | Factual
prednisolone | 0 | 288 | Factual
partial pressure of oxygen in arterial blood/fraction of inspired oxygen (PaO2/FiO2) 128.75 | 0 | 0 | Factual
P/F ratio improved | 0 | 288 | Factual
infiltration shadows improved | 288 | 288 | Factual
extubated | 288 | 288 | Factual
transferred to the Department of Neurosurgery | 528 | 528 | Factual
transferred to a rehabilitation hospital | 528 | 528 | Factual