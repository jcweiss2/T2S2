79 years old | 0
    female | 0
    admitted to the hospital | 0
    dyspnea | -24
    palpitations | -24
    hypertension | -17520
    type 2 diabetes mellitus | -17520
    atrial fibrillation | -17520
    colonic diverticulosis | -17520
    depressive syndrome | -17520
    osteoporosis | -17520
    mastectomy due to breast cancer | -26208
    ischemic cardiomyopathy | -17520
    acute myocardial infarction | -17520
    percutaneous angioplasty | -17520
    omeprazole 20 mg q.d. | -17520
    metformin 850 mg b.i.d. | -17520
    calcifediol 266 µg q. 1 month | -17520
    calcium 500 mg q.d. | -17520
    alendronate 70 mg q. 1 week | -17520
    acenocumarol 4 mg | -17520
    amiodarone 200 mg q.d. | -1344
    torasemide 5 mg q.d. | -17520
    enalapril 5 mg q.d. | -17520
    letrozole 2.5 mg q.d. | -17520
    citalopram 10 mg q.d. | -17520
    acetaminophen on demand | -17520
    lormetazepam on demand | -17520
    pale | 0
    diaphoretic | 0
    hypothermic (35.6°C) | 0
    tachycardia (146/min) | 0
    aortic murmur II/VI | 0
    chronic venous insufficiency | 0
    no edemas | 0
    hypophonesis | 0
    crackles on the right pulmonary base | 0
    cardiac insufficiency | 0
    atrial fibrillation with fast ventricular response (150/min) | 0
    diuretics | 0
    vasodilators | 0
    digoxin | 0
    echocardiogram apical and mid-segment akinesia | 0
    hypokinesis in basal segments | 0
    elevated cardiac troponin | 0
    slight leucocytosis | 0
    increased inflammatory markers | 0
    thoracic radiography vascular redistribution | 0
    cardiomegaly | 0
    pulmonary edema | 0
    coronary angiography no stenotic or spasmodic changes | 0
    stent stenosis 30% | 0
    ventriculography apical dyskinesia | 0
    Takotsubian apical ballooning | 0
    preserved LVEF | 0
    transdermal nitrates | 0
    digoxin (added) | 0
    decrease in myocardial damage markers | 24
    electrocardiographic stability | 24
    normofrequent atrial fibrillation | 24
    hyperthyroidism (TSH 0.014 µU/mL, FT4 4.48 ng/dL) | 120
    asymptomatic | 120
    no goiter | 120
    no exophthalmos | 120
    no pretibial myxedema | 120
    TSI <0.9 mUI/mL | 120
    anti-thyroperoxidase 6.16 UI/mL | 120
    anti-thyroglobulin 14.88 UI/mL | 120
    amiodarone for past two months | -1344
    type I amiodarone-induced hyperthyroidism | 120
    amiodarone suspended | 120
    methimazole 10 mg q. 8 h | 120
    TSH <0.014 µU/mL | 144
    FT4 7.55 ng/dL | 144
    FT3 4.04 pg/mL | 144
    type II amiodarone-induced hyperthyroidism | 144
    prednisone 45 mg q.d. | 144
    TSH <0.014 µU/mL (after prednisone) | 168
    FT4 3.9 ng/dL | 168
    FT3 1.65 pg/mL | 168
    methimazole stopped | 168
    urgent abdominal surgery (ischemic colitis with perforation) | 168
    right hemicolectomy | 168
    descendant doses of corticoids | 168
    thyroid function normalized | 432
    discharged | 1008
    normal thyroid function | 1008
    complete resolution of TC | 1008
    cardiovascular symptoms back to baseline | 1008
    ischemic colitis with bowel perforation | 4032
    generalized sepsis | 4032
    fatal outcome | 4032
    thyroid function normal | 4032
    