22 years old | 0
female | 0
admitted to the hospital | 0
railway accident | -72
below-knee amputation | -72
interlocking nail in the bilateral femur | -72
open book pelvic bone fracture | -72
Morel-Lavallée lesions | -72
conscious | 0
oriented | 0
stable hemodynamic parameters | 0
heart rate of 90/min | 0
blood pressure of 110/70 mm Hg | 0
respiratory rate of 20/min | 0
iv antibiotics injection meropenem | 0
iv antibiotics injection vancomycin | 0
features of sepsis | 120
surgical debridement of the Morel-Lavallée lesion | 120
hypotension | 120
inotropic support | 120
persistent hypotension | 144
high-grade fever | 144
rising total leukocyte count | 144
black foul smelling necrotic areas | 168
cottony bread mold lesions | 168
surgical debridement | 168
extensive muscle necrosis | 168
breach of peritoneum | 168
bowel exposed | 168
tissue for fungal culture and sensitivity | 168
histopathological examination | 168
nonseptate irregular hyphae of class zygomycetes | 168
provisional diagnosis of mucormycosis | 168
liposomal amphotericin B | 168
fungal culture grew strains of Rhizopus oryzae | 192
invasive mucormycosis | 192
severe septic shock | 216
death | 216