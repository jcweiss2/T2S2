22 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
mild COVID-19 illness | -720 | -720 | Factual
sore throat | -720 | -720 | Factual
loss of sense of smell | -720 | -720 | Factual
positive COVID-19 PCR | -720 | -720 | Factual
full recovery | -336 | -336 | Factual
resolution of symptoms | -336 | -336 | Factual
negative PCR | -336 | -336 | Factual
first dose of inactivated SARS-CoV-2 vaccine | -30 | -30 | Factual
asymptomatic | -30 | 0 | Factual
second dose of inactivated SARS-CoV-2 vaccine | 0 | 0 | Factual
headache | 2 | 2 | Factual
fatigue | 2 | 2 | Factual
fever | 24 | 168 | Factual
sore throat | 24 | 168 | Factual
abdominal pain | 24 | 168 | Factual
high-grade fever | 96 | 96 | Factual
myalgia | 96 | 168 | Factual
nausea | 96 | 168 | Factual
vomiting | 96 | 168 | Factual
diarrhea | 96 | 168 | Factual
faint erythematous non-itchy rash | 96 | 168 | Factual
dry irritant cough | 96 | 168 | Factual
no shortness of breath | 96 | 168 | Negated
no chest discomfort | 96 | 168 | Negated
no urinary symptoms | 96 | 168 | Negated
no pain or swelling of joints | 96 | 168 | Negated
temperature of 39°C | 96 | 96 | Factual
systolic blood pressure of 110 mm Hg | 96 | 96 | Factual
tachycardia | 96 | 168 | Factual
dry mucous membranes | 96 | 96 | Factual
congested throat | 96 | 96 | Factual
bilateral conjunctival injection | 96 | 96 | Factual
left conjunctival hemorrhage | 96 | 96 | Factual
generalised erythematous maculopapular rash | 96 | 168 | Factual
no enlarged peripheral lymph nodes | 96 | 96 | Negated
no audible cardiac murmurs | 96 | 96 | Negated
clear chest | 96 | 96 | Factual
unremarkable abdomen examination | 96 | 96 | Factual
SARS-CoV-2 PCR negative | 96 | 96 | Factual
SARS-CoV-2 IgG positive | 96 | 96 | Factual
throat swab negative for group A streptococcus | 96 | 96 | Factual
sputum culture showed mixed flora | 96 | 96 | Factual
bacterial blood cultures negative | 96 | 96 | Factual
urinalysis showed significant proteinuria | 96 | 96 | Factual
ANA negative | 96 | 96 | Factual
dsDNA negative | 96 | 96 | Factual
c-ANCA negative | 96 | 96 | Factual
p-ANCA negative | 96 | 96 | Factual
C3 reduced | 96 | 96 | Factual
C4 reduced | 96 | 96 | Factual
admitted to ICU | 96 | 96 | Factual
treated with ceftriaxone | 96 | 168 | Factual
treated with levofloxacin | 96 | 168 | Factual
treated with intravenous hydrocortisone | 96 | 120 | Factual
haemodynamic stability | 120 | 120 | Factual
facial puffiness | 120 | 168 | Factual
generalised body oedema | 120 | 168 | Factual
persistent diarrhea | 120 | 168 | Factual
myalgia | 120 | 168 | Factual
anasarca | 120 | 168 | Factual
renal impairment | 120 | 168 | Factual
significant proteinuria | 120 | 168 | Factual
ECG showed sinus tachycardia | 120 | 120 | Factual
non-specific T-wave abnormalities | 120 | 120 | Factual
troponin-I raised | 120 | 120 | Factual
pro-BNP raised | 120 | 120 | Factual
severe tricuspid regurgitation | 120 | 120 | Factual
pulmonary hypertension | 120 | 120 | Factual
right atrium and ventricle moderately dilated | 120 | 120 | Factual
left ventricle cavity size normal | 120 | 120 | Factual
mildly reduced ejection fraction | 120 | 120 | Factual
thin rim of pericardial effusion | 120 | 120 | Factual
bilateral moderate pleural effusion | 120 | 120 | Factual
basal atelectasis | 120 | 120 | Factual
treated with dexamethasone | 168 | 216 | Factual
generalised oedema subsided | 216 | 216 | Factual
skin rash resolved | 216 | 216 | Factual
conjunctivitis resolved | 216 | 216 | Factual
white blood cell count normalised | 216 | 216 | Factual
renal function improved | 216 | 216 | Factual
inflammatory markers normalised | 216 | 216 | Factual
repeat echocardiogram showed trace tricuspid regurgitation | 216 | 216 | Factual
right ventricular systolic function improved | 216 | 216 | Factual
pulmonary artery systolic pressure normalised | 216 | 216 | Factual
discharged home | 240 | 240 | Factual
tapering dose of prednisolone | 240 | 336 | Factual
follow-up | 336 | 336 | Factual
symptoms resolved | 336 | 336 | Factual
general weakness | 336 | 336 | Factual
fatigue | 336 | 336 | Factual
repeat echocardiogram normal | 336 | 336 | Factual