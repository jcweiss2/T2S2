50 years old | 0
Hispanic male | 0
admitted to the hospital | 0
end-stage renal disease | -7200
hypertension | -7200
30-year history of smoking | -26280
bilateral interstitial opacities | -7200
Karnofsky performance status score was 90 | -7200
cytomegalovirus (CMV) IgG was negative | -7200
kidney transplantation | 0
cold ischemic time of 11 hours 59 minutes | 0
warm ischemic time of 63 minutes | 0
immediate graft function | 0
Basiliximab 0.2 mg | 0
Basiliximab 0.2 mg | 96
Valganciclovir 900 mg | 0
sulfamethoxazole/trimethroprim 800/160 mg | 0
Methylprednisolone 250 mg | 0
tacrolimus 2 mg | 0
MMF 1,000 mg | 0
discharged | 120
shortness of breath | 720
cough | 720
respiratory distress | 720
impending respiratory failure | 720
arterial blood gas showed: pH of 7.33, pO2 of 61 mm Hg, pCO2 of 38 mm Hg, and HCO3− of 18.9 mEq/L (FiO2 50%) | 720
intubated | 720
CXR revealed diffuse airspace disease | 720
CT demonstrated patchy ground-glass opacities with interlobular septal thickening, associated with bronchiectasis | 720
bronchoscopy | 720
bronchoalveolar lavage samples were negative | 720
vancomycin 1.5 g | 720
cefepime 1 mg | 720
oseltamivir 150 mg | 720
tacrolimus discontinued | 720
MMF discontinued | 720
prednisone 20 mg changed to methylprednisone 100 mg | 720
aggressive diuresis with furosemide | 720
extubation | 744
arterial blood gas immediately post-extubation showed a pO2 of 89.8 mm Hg, pCO2 of 33.7 mm Hg, pH of 7.44, and a HCO3 of 22.7 mmol/L (FiO2 35%) | 744
MMF resumed | 744
respiratory distress | 768
severe hypoxia | 816
re-intubation | 816
all immunosuppressive drugs discontinued except for methylprednisone | 816
open lung biopsy | 816
extensive areas of interstitial fibrosis | 816
gram negative sepsis | 1008
died | 1008
lung autopsy revealed a picture of extensive intra-alveolar hemorrhages and interstitial fibrosis with thickening of the alveolar septa | 1008