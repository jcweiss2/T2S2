59 years old | 0
male | 0
prostatic cancer | -672
CT guided percutaneous transhepatic core needle liver mass biopsy | -9
angio-embolization of the hepatic mass | -9
admitted to the recovery room | 0
blood pressure 84/55 | 0
heart rate 77 | 0
respiratory rate 26 | 0
acidotic with pH 7.31 | 0
base deficit of 6.5 | 0
INR of 1.6 | 0
PT 17.8 | 0
bladder pressure of 25 mmHg | 0
repeat CT of abdomen and pelvis | 0
perihepatic hematoma expansion | 0
no evidence of blush | 0
admission to the surgical ICU | 0
coagulopathy correction | 0
multiple transfusions of fresh frozen plasma | 0
multiple transfusions of cryoprecipitate | 0
severe intra-abdominal hypertension | 0
compartment syndrome | 0
bladder pressure: 40 mmHg | 0
taken to the operating room | 0
bleeding liver mass located in the dome of segments 7 and 8 | 0
falciform ligament taken down | 0
right upper quadrant packed | 0
patient stabilized | 0
packs were dry at the end of the case | 0
resumed bleeding within twenty-four hours | 24
angiography of the right hepatic artery | 24
no blush | 24
bleeding thought to be venous in origin | 24
fed by a superior right hepatic artery branch | 24
selective right hepatic artery embolization | 24
returned to the OR later that day | 24
hepatic artery branch ligated | 24
laparotomy packing performed in the right upper quadrant | 24
patient stabilized | 24
re-exploration on post-operative day 2 | 48
parenchymal bleeding resumed | 48
Surgicel | 48
Argon beam coagulation | 48
fibrin sealant | 48
more packing | 48
insufficient to create hemostasis | 48
initiated the BOLSA | 48
intraoperative improvements after BOLSA placement | 48
BP at surgery start was 80/45 | 48
BP at end of case was 90/50 | 48
transfusions were described as “massive transfusion protocol ongoing” | 48
total transfusion for case was 3 units packed red blood cells | 48
total transfusion for case was 3 units fresh frozen plasma | 48
estimated blood loss was listed as 2 l | 48
case lasted 19 min | 48
cholecystectomy on POD 4 | 96
ischemic cholecystitis secondary to the right hepatic artery embolization | 96
Wittmann patch placed | 96
serial tightening of the Wittmann patch bedside | 96
pathology report of the liver biopsy returned on POD 7 | 168
hemangioma | 168
BOLSA removed without bleeding | 216
abdomen closed primarily | 216
patient progressed to resumption of activities of daily living | 216
discharged home | 216