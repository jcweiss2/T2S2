15 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
acute myelogenous leukemia | 0 | 0 | Factual
standard induction treatment | -336 | -168 | Factual
chemotherapy | -336 | -168 | Factual
pancytopenia | -168 | 0 | Factual
anti-infective treatment | -168 | 0 | Factual
ciprofloxacin | -168 | 0 | Factual
linezolid | -168 | 0 | Factual
meropenem | -168 | 0 | Factual
tobramycin | -168 | 0 | Factual
liposomal amphotericin | -168 | 0 | Factual
tachycardia | 0 | 0 | Factual
hypotension | 0 | 0 | Factual
lactic acidosis | 0 | 0 | Factual
admitted to pediatric intensive care unit | 0 | 0 | Factual
severely impaired left ventricular ejection fraction | 0 | 0 | Factual
sinus tachycardia | 0 | 0 | Factual
incomplete right bundle branch block | 0 | 0 | Factual
elevated NT-proBNP | 0 | 0 | Factual
elevated high-sensitive troponin T | 0 | 0 | Factual
fluid therapy | 0 | 0 | Factual
noradrenaline | 0 | 0 | Factual
dobutamine | 0 | 0 | Factual
milrinone | 0 | 0 | Factual
deep sedation | 0 | 0 | Factual
mechanical ventilation | 0 | 0 | Factual
lactate acidosis worsened | 0 | 24 | Factual
hypotonic | 0 | 24 | Factual
va-ECMO initiated | 24 | 24 | Factual
cannulation of left femoral artery and vein | 24 | 24 | Factual
Dacron conduit sewed on right femoral artery | 48 | 48 | Factual
second arterial cannula introduced | 48 | 48 | Factual
ECBF enhanced | 48 | 72 | Factual
MAP maintained | 48 | 72 | Factual
PCT levels rose | 48 | 72 | Factual
Hickman catheter explanted | 72 | 72 | Factual
broad-complex tachycardia | 72 | 72 | Factual
esmolol | 72 | 72 | Factual
metoprolol | 72 | 72 | Factual
left ventricular function further decreased | 72 | 96 | Factual
aortic valve ceased to open | 96 | 96 | Factual
second venous cannula placed | 96 | 96 | Factual
left atrium cannulation | 96 | 96 | Factual
ECBF reached 5-6 l/min | 96 | 120 | Factual
lactate levels peaked | 96 | 120 | Factual
MAP rose | 120 | 120 | Factual
cerebral oximetry | 120 | 120 | Factual
left ventricle unloaded | 120 | 120 | Factual
therapeutic anticoagulation | 120 | 168 | Factual
PCT peaked | 120 | 168 | Factual
CRP peaked | 120 | 168 | Factual
leukocytes remained low | 120 | 168 | Factual
high-sensitive troponin T increased | 120 | 168 | Factual
creatine kinase MB increased | 120 | 168 | Factual
cardiac systolic function recovered | 168 | 240 | Factual
ECMO cannulas removed | 240 | 240 | Factual
ECMO completely removed | 288 | 288 | Factual
LVEF recovered | 288 | 288 | Factual
CVVHDF stopped | 288 | 288 | Factual
leucocyte count recovered | 312 | 312 | Factual
respirator weaning | 408 | 408 | Factual
allogenic stem cell transplantation | 1008 | 1008 | Factual
discharged to rehabilitation facility | 1512 | 1512 | Factual
severe critical illness | 1512 | 1512 | Factual
polyneuropathy | 1512 | 1512 | Factual
LVEF recovered | 1512 | 1512 | Factual