47 years old | 0
female | 0
obese | 0
short neck | 0
admitted to the hospital | 0
respiratory distress | 0
asphyxiation | 0
total thyroidectomy | -624
medullary thyroid carcinoma | -624
enlarged fibrotic multinodular goiter | -624
tracheal compression | -624
neck stiffness | -624
throat fullness | -624
hoarseness | -624
orthopnea | -624
difficulty breathing | -624
tracheostomy | -624
tracheomalacia | -624
RLN injury | -624
discharged from the hospital | -48
neck stiffness | -24
throat tightness | -24
dyspnea | -24
pain during swallowing | -24
subfebrile condition | -24
cough | -24
purulent sputum | -24
referred to an otorhinolaryngologist | -24
indirect mirror laryngoscopy | -24
right VCP | -24
decannulation | -18
discharged home | -18
referred to a pulmonologist | -12
bronchodilators | -12
no clinical improvement | -12
admitted to the ED | 0
severe tachy-dyspnea | 0
desaturation | 0
orthodeoxia | 0
biphasic stridor | 0
diaphoresis | 0
impossible swallowing | 0
tachycardia | 0
hypertension | 0
aphonia | 0
fever | 0
post thyroidectomy scar | 0
reddish | 0
previous tracheostomy fully obliterated | 0
large painful submandibular mass | 0
bilateral expiratory rhonchi | 0
purulent sputum | 0
reddish discoloration of the skin | 0
contrast enhanced CT scan | 0
pre-tracheal cavity | 0
gaseous content | 0
closed glottis | 0
immobile glottic musculature | 0
bilateral VCP | 0
intubation | 0
rapid sequence induction | 0
re-tracheostomy | 0
unintentionally retained gauze | 0
gossypiboma | 0
abscess cavity cultures | 0
Streptococcus viridans | 0
antimicrobial course | 0
cured | 720
discharged | 720
decannulated | 744
full recovery | 744
voice rehabilitation | 744
voice fatigue | 960