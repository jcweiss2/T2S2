10 years old | 0
    male | 0
    weight 26 kg | 0
    pain in epigastrium | -72
    dull pain | -72
    mild to moderate pain | -72
    no radiation of pain | -72
    hepatomegaly | -72
    computed tomography scan abdomen | -72
    cystic lesion 12.5 × 8.5 × 11.4 cm in left lobe of liver | -72
    cyst extending to lesser sac and perihepatic area | -72
    small cysts in right kidney | -72
    routine blood investigations | -72
    liver function tests | -72
    anti-Echinococcus IgG antibody positive | -72
    hydatid cyst of liver | -72
    hydatid cyst of kidney | -72
    posted for elective laparoscopic removal of hepatic cysts | 0
    posted for elective laparoscopic removal of renal cysts | 0
    baseline haemodynamic parameters normal | 0
    inhalational induction with sevoflurane | 0
    fentanyl 60 μg administered | 0
    vecuronium 3 mg administered | 0
    trachea intubated | 0
    10% povidone4 iodine injected into hepatic hydatid cyst | 0
    heart rate increased from 110 to 180/min | 1
    hypercarbia | 1
    end-tidal CO2 55 mmHg | 1
    hyperthermia | 1
    temperature increased from 35.1 to 37.4°C | 1
    paracetamol 500 mg administered | 1
    normal saline 0.5 L bolus infused | 1
    arterial blood gas analysis pH 7.14 | 1
    arterial blood gas pCO2 36.5 mmHg | 1
    arterial blood gas pO2 135 mmHg | 1
    arterial blood gas SO2 97.7% | 1
    K+ 7.4 mmol/L | 1
    Na+ 127 mmol/L | 1
    Ca+ 0.81 mmol/L | 1
    Cl− 249 mmol/L | 1
    lactate 4.3 mmol/L | 1
    base deficit -15 mmol/L | 1
    HCO3 12.7 mmol/L | 1
    Hb 16 g/dL | 1
    blood pressure normal | 1
    airway pressures normal | 1
    urine output decreased | 1
    urine output not improved after first fluid bolus | 1
    balanced salt solution 0.5 L bolus infused | 1
    frusemide 15 mg IV administered | 1
    urine output improved | 1
    presumptive diagnosis of anaphylaxis | 1
    hydrocortisone administered | 1
    pheniramine maleate administered | 1
    shifted to ICU | 1
    haemoglobin 17 g/dL | 1
    leukocyte count 49.6 × 103/μL | 1
    serum creatinine 0.9 mg/dL | 1
    serum albumin 1.9 g/dL | 1
    potassium 5.2 mEq/L | 1
    liver function tests normal | 1
    renal function tests normal | 1
    thyroid function tests normal | 1
    severe metabolic acidosis persisted | 1
    plan for haemodialysis made | 1
    tachycardia fluid responsive | 1
    Sterofundin® 100 ml/h started | 1
    albumin 20% 25 ml/h started | 1
    hydrocortisone 6 mg/h started | 1
    echocardiography good cardiac contractility | 1
    under filled heart chambers | 1
    inferior vena cava diameter 0.4 – 0.8 cm | 1
    collapsibility | 1
    haemodialysis initiated | 4
    acidosis corrected | 4
    heart rate settled | 4
    fully awake | 24
    obeying commands | 24
    trachea extubated | 24
    hydrocortisone infusion tapered | 24
    hydrocortisone infusion stopped | 24
    kept in ICU for observation | 24
    shifted to ward | 72
    