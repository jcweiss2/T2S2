49 years old | 0
    female | 0
    presented to a peripheral hospital | 0
    fatigue | 0
    dizziness | 0
    intermittent fever | 0
    minor scratch on left foot | 0
    trauma at left foot | -72
    computed tomography (CT) | 0
    large vegetation at aortic valve cusp | 0
    pericardial effusion | 0
    calculated antibiotic therapy | 0
    referred to department of cardiology | 0
    enormous size of vegetation (~3 cm long) | 0
    increasing pericardial effusion | 0
    referred to center for emergency surgery | 0
    standard sternotomy | 0
    opened pericardium | 0
    hemorrhagic pericardial effusion detected | 0
    placed on cardiopulmonary bypass (CPB) | 0
    aortotomy | 0
    large vegetation identified near left main coronary artery | 0
    thromboembolism prevention during vegetation removal | 0
    two small septic perforations of aortic wall detected | 0
    Prolene 4-0 sutures used for closure | 0
    aortic valve replaced with 21-mm SJM mechanical valve | 0
    uneventful weaning of CPB | 0
    no bleeding in situ | 0
    chest closed | 0
    transferred to ICU | 0
    stable hemodynamic condition | 0
    mild dosages of catecholamines | 0
    arrival in ICU | 0
    sudden large quantities of blood in thoracic drainage (1.5 L) | 1
    hemodynamic instability | 1
    reoperation initiated | 1
    resuscitation on way to operation room | 1
    sternum reopened under resuscitation | 1
    placed on CPB | 1
    preliminary hemodynamic stabilization | 1
    large rupture of left ventricular lateral wall (1.5x1.5 cm) | 1
    attempts for direct closure unsuccessful | 1
    Dor plasty not feasible | 1
    excision of soft phlegmonlike myocardium | 1
    histopathological examination | 1
    myocardial infarction presence | 1
    multiple bacteria in coronary capillary vessels | 1
    bacterial imbibition of myocardial tissue | 1
    myocardial reconstruction with Dacron patch | 1
    larger Dacron patch placed outside myocardium | 1
    additional running suture around second patch | 1
    venous bypass graft using saphenous vein | 1
    BioGlue used on suture | 1
    no bleeding detected after cardiac activity reestablished | 1
    extracorporeal life support (ECLS) via left femoral artery and vein | 1
    CPB weaned | 1
    referred to ICU after chest closure | 1
    mild-to-moderate catecholamine | 1
    ECLS weaned after 5 days | 120
    abscess at left foot lanced | 120
    referred to peripheral hospital after 14 days ICU stay | 336
    antibiotics administered for 6 weeks | 1008
    positive blood cultures for Staphylococcus aureus | 1008
    clindamycin | 1008
    flucloxacillin | 1008
    echocardiography after ECLS weaning | 120
    left ventricular ejection fraction 60% | 120
    mild pericardial effusion | 120
    pseudoaneurysm detected after 1 year | 8760
    reoperation for aneurysm resection | 8760
    7-day postoperative course | 8760
    referred to rehabilitation | 8760
    well at home after half a year | 4392
    