48 years old | 0
male | 0
known diabetic | 0
presented with painful swelling | 0
swelling in the back below the left shoulder | 0
low-grade fever | -756
cough | -756
vaccinated with COVID-19 vaccine | -168
painful swelling on his left arm | -168
spreading to the shoulder and scapular region | -168
decreased limb movements | -168
acute onset of fever | -120
cough with mucoid expectoration | -120
progressive deterioration of his health | -120
receiving anti-tubercular drugs | -120
febrile | 0
left arm swollen and tender | 0
reduced range of movement | 0
unable to raise his arm above the shoulder | 0
ultrasound confirmed an abscess | 0
chest radiographs showed disseminated pulmonary pathology | 0
bilateral lung abscesses | 0
pleural effusions | 0
pus culture yielded pure growth of Burkholderia pseudomallei | 0
treated with intravenous meropenem | 0
improvement | 504
resolution of the abscess | 504
decrease in respiratory symptoms | 504
discharged | 552
advice for oral trimethoprim-sulfamethoxazole | 552 
oral trimethoprim-sulfamethoxazole | 552