23 years old | 0
male | 0
admitted to the ICU | 0
complains of sudden onset of pain abdomen | 0
respiratory distress | 0
intestinal perforation | 0
blood pressure 110/60 mm of Hg | 0
pulse 86 beats/min | 0
respiratory rate 22 breaths/min | 0
SpO2 99% on room air | 0
afebrile on touch | 0
urgent laparotomy | 0
asymptomatic for 2 days after surgery | 48
blood pressure fall up to 84 mmHg | 72
CVC in the right subclavian vein | 72
cannulation of right subclavian vein | 72
CVP catheter placement | 72
USG guidance | 72
lateral approach | 72
guide wire confirmed well in position | 72
guide wire movement free | 72
CVP catheter fixed at 15 cm | 72
dampened CVP waveform | 72
CVP waveform could not be improved | 72
chest radiograph performed | 72
malpositioning of CVC in left subclavian vein | 72
right subclavian CVC removed | 72
reintroduction of CVC under color Doppler guidance | 80
modified Seldinger technique | 80
guide wire confirmed well in position | 80
repeat chest radiograph | 80
correct placement of CVC | 80
normal CVP tracing | 80
discharged | -1 
Note: The time stamp for "discharged" is not explicitly mentioned in the text, so it is assumed to be after the correction of the CVC placement, and the exact time is not known, so it is marked as -1 to indicate that it is not available.