66 years old | 0
male | 0
admitted to the hospital | 0
coronary syndrome | -2640
dual platelet antiaggregant therapy | -2640
chronic kidney failure | -2640
arterial hypertension | -2640
gout arthritis | -2640
obesity | -2640
hyperlipidemia | -2640
necrotizing pancreatitis | -7920
open necrosectomy | -7920
prolonged open abdomen | -7920
incisional hernia | -7920
synthetic mesh | -7920
hypovolemic shock | 0
gastrointestinal bleeding | 0
abdominal wound with mesh exposition | 0
cloudy discharge | 0
high output enterocutaneous fistula diagnosis | 0
oral intake suppressed | 0
subatmospheric pressure device | 0
periodical changes | 0
parenteral nutrition | 0
somatostatin analogous | 0
fistula bleeding | 0
infection | 0
intensive care unit attention | 0
blood transfusions | 0
antibiotics | 0
antifungal management | 0
severe peritoneal adherence syndrome | 0
computed tomography images | 0
laparoscopic access | 0
peritoneal adhesion lysis | 0
paramedian laparotomy | 0
parietectomy | 0
en-bloc resection of the involved small bowel | 0
enteric anastomosis | 0
mechanical sutures | 0
absorbable sutures | 0
open abdomen covered with subatmospheric pressure device | 0
keratinizing and infiltrating giant cell squamous cell carcinoma | 0
moderate and low differentiated | 0
involves all the skin depth | 0
subcutaneous cellular tissue | 0
intestinal wall of all the enterocutaneous fistula | 0
resection margins negative for tumor invasion | 0
keloid scaring | 0
foreign body reactions | 0
clinical deterioration | 48
higher respiratory and hemodynamic support | 48
abdominal drainage turned cloudy | 48
anastomosis dehiscence | 48
anastomosis resection | 48
new enteric anastomosis deferred | 48
severe intestinal edema | 48
new subatmospheric pressure device | 48
septic shock | 96
necrotizing fasciitis of the abdominal wall borders | 96
debridement | 96
subatmospheric pressure device replaced | 96
respiratory and hemodynamic status deterioration | 120
death | 120