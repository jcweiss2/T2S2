3-day-old | 0  
    ex-full term | 0  
    male | 0  
    presented to the emergency department | 0  
    apnea episodes | 0  
    birth weight 3065 g | 0  
    appropriate for gestational age | 0  
    normal spontaneous vaginal delivery | 0  
    maternal polycystic ovarian syndrome | 0  
    maternal metformin treatment during first trimester | 0  
    borderline gestational diabetes concerns | 0  
    elevated glucose tolerance tests | 0  
    normal 3-h glucose test | 0  
    Group B Streptococcal infection | 0  
    antibiotics provided | 0  
    uncomplicated delivery | 0  
    difficulty with breastfeeding | 0  
    poor milk production on day of life 2 | -48  
    formula supplementation | -48  
    discharged home | -48  
    poor feeding at home | -48  
    poor colostrum production | -48  
    continued formula supplementation | -48  
    apnea episodes (ruddy color, limp, eyes rolling back) | -24  
    episodes lasting 10 seconds | -24  
    episodes not associated with feedings | -24  
    return to baseline after stimulation | -24  
    presentation to ED on day of life 3 | 0  
    stable vital signs | 0  
    undetectable glucose | 0  
    Dextrose 10% bolus | 0  
    D 10% infusion | 0  
    glucose 18 mg/dL | 0  
    repeat Dextrose 10% bolus | 0  
    glucose infusion rate 13.85 mg/kg/min | 0  
    sepsis evaluation initiated | 0  
    urinalysis | 0  
    urine culture | 0  
    blood culture | 0  
    empiric ampicillin and gentamicin treatment | 0  
    negative cultures after 48 hours | 48  
    antibiotics discontinued | 48  
    normal chest X-ray | 0  
    negative COVID-19 | 0  
    unremarkable CBC | 0  
    hyperkalemia 5.9 | 0  
    hypocalcemia 7.2 | 0  
    transfer to Cedars-Sinai NICU | 0  
    persistent hypoglycemia requiring high glucose infusion rates | 0  
    normal tone, color, activity level prior to transport | 0  
    blood glucose 44 mg/dL prior to transport | 0  
    arrival to NICU | 0  
    glucose 66 mg/dL | 0  
    D 12.5% infusion at 13.85 mg/kg/min | 0  
    weight 30th percentile | 0  
    length 25th percentile | 0  
    head circumference 55th percentile | 0  
    duplicated earlobes | 0  
    glucose stabilized for 12 hours | 12  
    glucose infusion rate weaned to 12 mg/kg/min | 12  
    pediatric endocrinology consultation | 0  
    persistent hypoglycemia evaluation initiated | 0  
    serum glucose 40 mg/dL | 0  
    normal ammonia 70 µmol/L | 0  
    beta-hydroxybutyrate 0.2 mmol/L | 0  
    cortisol 5.8 µg/dL | 0  
    serum insulin 6.0 µIU/mL | 0  
    hyperinsulinism diagnosis | 0  
    low-dose ACTH stimulation test | 0  
    robust cortisol response | 0  
    adrenal insufficiency excluded | 0  
    diazoxide 8 mg/kg/day initiated | 0  
    chlorothiazide 20 mg/kg/day initiated | 0  
    glucose infusion rate remained elevated at 11.11 mg/kg/min after 36 hours | 36  
    diazoxide increased to 12 mg/kg/day | 36  
    medical genetics consultation | 0  
    chromosomal microarray recommended | 0  
    CH panel recommended | 0  
    intermittent tachypnea | 192  
    oxygen desaturations to 80s | 192  
    chest X-ray concerning for pulmonary edema | 192  
    cardiology consultation | 192  
    echocardiogram showing PDA and PFO | 192  
    left-to-right shunting | 192  
    moderately elevated pulmonary artery pressures | 192  
    chlorothiazide increased to 40 mg/kg/day | 192  
    resolution of pulmonary edema | 192  
    normal repeat echocardiograms | 192  
    CH gene panel negative for ABCC8, KCNJ11, GCK, GLUD1, HADH, HNF1A, HNF4A, SLC16A1, UCP2 | 192  
    chromosome microarray with 17q12 duplication | 192  
    hyperinsulinism improvement | 192  
    diazoxide titrated down to 1.5 mg/kg/day | 192  
    chlorothiazide decreased to 20 mg/kg/day | 192  
    discharged home | 192  
    outpatient follow-up | 192  
    normal cardiac examinations | 192  
    normal echocardiograms | 192  
    weaned off diazoxide and chlorothiazide at 3 months | 2160  

<|eot_id|>
