65 years old | 0
male | 0
non-ischaemic cardiomyopathy | -120
left ventricular ejection fraction (LVEF) 20% | -120
New York Heart Association (NYHA) class II | -120
paroxysmal atrial fibrillation | -120
previous cerebrovascular accident | -120
hypertension | -120
dyslipidaemia | -120
depression | -120
abdominal pain | -120
discharged from community hospital | -120
admitted to hospital | 0
generalized abdominal pain | 0
fatigue | 0
congestive heart failure | 0
transthoracic echocardiography | 0
left ventricular function of 11% | 0
mild right ventricular dysfunction | 0
intravenous furosemide infusion | 0
bisoprolol held | 0
candesartan held | 0
acute kidney injury (AKI) | 8
elevated liver enzymes | 8
lactate normalized | 8
vitals stable | 8
bisoprolol 2.5 mg PO o.d. | 8
sacubitril/valsartan 24/26 mg PO b.i.d. | 8
hypotension | 9
norepinephrine | 9
dobutamine | 9
worsening AKI | 9
transferred to tertiary academic centre | 10
right heart catheterization | 10
vasoplegic shock | 10
sepsis ruled out | 10
adrenal insufficiency ruled out | 10
vasopressor/inotrope | 10
vasoplegic shock resolved | 14
norepinephrine weaned off | 14
creatinine improved | 14
right heart catheterization | 15
resolving vasodilatory shock | 15
cardiogenic shock | 15
dobutamine continued | 15
IV furosemide infusion started | 15
dobutamine weaned off | 17
hydralazine | 17
spironolactone | 17
bisoprolol initiated | 26
ramipril initiated | 32
discharged | 34
net 25 kg lost | 34
oral heart failure therapy | 34
sacubitril/valsartan discontinued | 210
hyperkalaemia | 210