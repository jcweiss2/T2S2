71 years old | 0
male | 0
hypertension | 0
type 2 diabetes | 0
admitted to the hospital | 0
fever | -48
cough | -48
dyspnea | -48
oxygen therapy | -48
noninvasive mechanical ventilation | -48
ceftazidime | -48
corticosteroids | -48
invasive mechanical ventilation | 24
septic shock | 24
renal failure | 24
imipenem/cilastatin | 24
levofloxacin | 24
antithrombotic | 24
estimated GFR with MDRD formulae: 27.5 mL/min/1.73 m2 | 24
oligoanuria | 48
metabolic acidosis | 48
hemodiafiltration | 72
second hemodiafiltration session | 96
urea: 16 | 96
creatinine: 1.9 | 96
improved metabolic acidosis | 96
diuresis | 96
third hemodiafiltration session | 120
leukocytosis | 120
neutrophilia | 120
elevated inflammatory markers | 120
cavitary image in the right upper lobe | 120
hemoculture and urine culture results found no growth | 168
broad-spectrum antibiotics | 168
meropenem | 168
vancomycin | 168
fluconazole | 168
respiratory weaning failure | 288
sedation | 288
relaxation | 288
paralysis | 288
ventilator strategy protection | 288
fiberoptic bronchoscopy | 312
erythematous lesions in the bronchial tree | 312
abundant purulent secretions | 312
cavitary lesion | 312
BAL sample isolated Klebsiella pneumoniae | 336
Pseudomonas aeruginosa carbapenemase Class A | 336
Trichosporon asahii | 336
Ceftazidime/avibactam | 336
colistin | 336
voriconazole | 336
septic shock | 360
multi-organ failure | 360
patient deceased | 384