86 years old | 0
male | 0
admitted to the hospital | 0
abdominal pain | -240
burning sensation while urinating | -240
asthenia | -240
anorexia | -240
weight loss | -360
peripheral arterial disease | -8760
hip replacement surgery | -8760
dehydration | 0
soft abdomen | 0
hypogastric tenderness | 0
palpable mass | 0
full bladder | 0
purulence | 0
hematuria | 0
inflammatory syndrome | 0
CRP at 378 mg/L | 0
leukocytes at 107,000/mm3 | 0
Procalcitonin at 16 ng/mL | 0
acute renal failure | 0
hyperkalemia | 0
creatinine at 1000 μmol/L | 0
emphysematous cystitis | 0
double antibiotic therapy | 0
hydration | 0
hypotension | 0
tachycardia | 0
tachypnea | 0
saturation of 96 % | 0
physiological saline | 0
Urosepsis | 0
Organic acute renal insufficiency | 0
acute pancreatitis | 0
abdomino-pelvic CT scan | 24
parietal enhancement | 24
necrosis | 24
Fresh Frozen Plasma | 24
exploratory laparotomy | 48
cystoscopy | 48
ureteral stent | 48
partial cystectomy | 48
gangrene of the bladder | 48
bladder perforation | 48
total cystectomy | 48
pulmonary embolism | 480
Morganella morganii | 0
radical cystectomy | 48
panparietal necrosis | 48
dense polymorphic suppurative inflammatory infiltrate | 48
favorable postoperative evolution | 720