18 years old | 0
male | 0
primigravida | 0
37 weeks of gestation | 0
referred to our institute | 0
supplemental oxygen | 0
Rapid test diagnosis of Plasmodium falciparum | -1
acute icteric leptospirosis | -1
high grade fever | -1
decreased urine output | -1
yellowish discolouration | -1
altered sensorium | -1
disoriented | -1
febrile | -1
icteric | -1
sub-conjunctival haemorrage | -1
fine basal crepitations | -1
intravenous artesunate | -1
ceftriaxone | -1
doxycycline | -1
anaemia | -1
jaundice | -1
deranged liver function | -1
coagulopathy | -1
thrombocytopenia | -1
increased total leucocyte count | -1
elevated blood urea nitrogen | -1
serum creatinine | -1
abdominal ultrasonography | -1
singleton pregnancy | -1
adequate liquor | -1
umbilical artery systolic-diastolic ratio of 2:1 | -1
mild hepato-splenomegaly | -1
non-reassuring fetal heart rate | -1
aspiration prophylaxis | -1
high-risk consent | -1
emergency caesarean delivery | -1
thiopental | -1
succinylcholine | -1
right internal jugular vein | -1
left radial artery | -1
ultrasonographic guidance | -1
baseline serum glucose level | -1
isoflurane | -1
N2O-O2 mixture | -1
atracurium | -1
delivery of a 2.25 kg baby | -1
fentanyl | -1
oxytocin | -1
Apgar score of 6 | -1
Apgar score of 8 | -1
cord blood pH of 7.28 | -1
base deficit of 5.4 | -1
blood sugar level of 50 mg/dl | -1
hypotension | -1
packed red blood cells | -1
fresh frozen plasma | -1
platelets transfusion | -1
noradrenaline infusion | -1
mild acidosis | -1
normal electrolytes | -1
serum glucose | -1
intensive care unit | -1
intubated state | -1
noradrenaline infusion | -1
ultrasound guided bilateral transverse abdominis plane block | -1
pulmonary haemorrage | -1
blood products | -1
bed side fibre-optic bronchoscopy | -1
erythematous mucosa | -1
blood clots | -1
active oozing | -1
diffuse bleeding from distal airway | -1
Factor VIIa | -1
erythematous mucosa | -1
blood clots | -1
active oozing | -1
diffuse bleeding from distal airway | -1
immediate bleeding cessation | -1
significant reduction of inspired oxygen fraction (FiO2) | -1
chest radiograph | -1
bilateral non-homogeneous opacities | -1
plasmapheresis | -1
dialysis | -1
acute kidney injury | -1
severe hyperbilirubinemia | -1
haemolytic uremic syndrome | -1
high serum lactate dehydrogenase | -1
schistocytes in peripheral blood | -1
computed tomography of the brain | -1
diffuse cerebral oedema | -1
cerebroprotective measures | -1
head elevation | -1
not rotating neck | -1
maintain serum sodium 145-155 Meq/L | -1
keeping blood partial pressure of carbondioxide 32-40 mmHg | -1
blood cultures | -1
urine cultures | -1
Weil-Felix test | -1
typhi dot | -1
dengue | -1
hepatitis viruses serology | -1
stress ulcer prevention | -1
deep vein thrombosis prophylaxis | -1
glycemic control | -1
intensity of fever started reducing | -1
consciousness improved | -1
inotropic support tapered | -1
urine output improved | -1
liver function test with coagulation parameters showed improving trends | -1
Pao2/Fio2 ratio also gradually improved | -1
extubated | -1
wards | -1
safely discharged from the hospital | -1