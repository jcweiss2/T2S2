fever | 0
vomiting | 0
generalized abdominal pain | 0
rash on palms and trunk | 0
severe drowsiness | 0
lethargy | 0
no conjunctivitis | 0
no lymphadenopathy | 0
respiratory rate 25/min | 0
oxygen saturation 93% | 0
tachycardia | 0
hypotension | 0
abdomen tender to palpation | 0
abdominal ultrasound showing enlarged appendix | 0
emergency laparotomy appendectomy | 2
postoperative course toxic | 2
tachycardia | 2
hypotension | 2
fractional shortening | 2
oxygen therapy | 2
bronchopneumonia | 2
treatment with ceftriaxone and amikacin | 2
switched to imipenem | 4
positive history of contact with COVID-19 | 4
positive serology of SARS-CoV-2 | 4
elevated ferritin | 4
elevated IL6 | 4
elevated high-sensitivity troponin | 4
elevated D-dimer | 4
enoxaparin | 4
IV immunoglobulin | 48
aspirin | 48
worsening general condition | 48
febrile | 48
anemic | 48
red blood cell transfusion | 48
pulse dosage of systemic corticosteroids | 72
re-evaluation of emerging shock | 72
aggravation of heart dysfunction | 72
dobutamine | 72
vasoactive drugs discontinued | 120
afebrile | 96
clinical symptoms improved | 96
arterial pressure stable | 96
no pathogenic agents detected | 96
histopathological examination showing catarrhal appendicitis | 96
D-dimer downward trend | 120
troponemia resolved | 120
inflammatory parameters normal | 168
LV function improved | 168
discharge | 288
follow-up outpatient visit | 336
blood tests normalized | 336
COV-2 IgG elevated | 336
abdominal and cardiac ultrasounds normal | 336