23 years old | 0
    multipara | 0
    admitted to the Intensive Care Unit (ICU) | 0
    hemodynamic instability | 0
    spontaneous vaginal delivery | -48
    live full-term male baby | -48
    pregnancy | -48
    no concomitant diseases | 0
    no history of thrombosis | 0
    previous pregnancy | 0
    normal postpartum course | 0
    no uterine instrumentation | 0
    no placental instrumentation | 0
    immediate course of hospitalization | 0
    highly febrile (39.4 °C) | -24
    severe abdominal pain | -24
    hypogastric regions pain | -24
    no nausea | 0
    no vomiting | 0
    lower abdominal quadrant pain | 0
    no uterine pain | 0
    blood pressure 95/65 mm Hg | 0
    pulse rate 107/min | 0
    peripheral oxygen saturation 97% | 0
    abdominal ultrasound | 0
    gynecologic ultrasound | 0
    no useful finding | 0
    cervical swab | 0
    blood culture | 0
    urine culture | 0
    elevated D-dimer (11573 mcg/L) | 0
    elevated C-reactive protein (106.2 mg/L) | 0
    no pyuria | 0
    cefazoline | 0
    low molecular weight heparin (LMWH) prophylactic dose | 0
    analgesics | 0
    hypotensive (64/31 mm Hg) | 24
    pulse rate 110/min | 24
    peripheral oxygen saturation 97% | 24
    aggressive fluid resuscitation | 24
    repeat gynecologic examination | 24
    vaginal ultrasound | 24
    no pathology | 24
    high suspicion of SPT | 24
    contrast-enhanced CT | 24
    thrombus in right pelvic veins | 24
    dilated right ureter | 24
    dilated right renal pelvis | 24
    elevated CRP (401 mg/L) | 24
    elevated procalcitonin (18.75 mg/L) | 24
    elevated urea (8.5 mmol/L) | 24
    elevated creatinine (147 µmol/L) | 24
    decreased D-dimer (5099 mcg/L) | 24
    metronidazole | 24
    transferred to ICU | 24
    hemodynamic instability | 24
    poor response to fluid resuscitation | 24
    vasopressors not needed | 24
    hemodynamic stabilization | 24
    ceftriaxone | 24
    LMWH therapeutic dosage | 24
    episodes of tachypnea | 24
    peaks of body temperature elevation | 24
    falls in peripheral oxygen saturation | 24
    hypoxemia | 24
    hypocapnia | 24
    chest radiography | 24
    pulmonary congestion | 24
    bilateral parenchymal infiltrates | 24
    pleural effusion | 24
    intensive respiratory physiotherapy | 24
    noninvasive ventilation | 24
    no conventional mechanical ventilation | 24
    negative microbiological cultures | 24
    cervical smear Streptococcus pyogenes group A | 24
    transferred to HDU | 72
    peaks of elevated temperature | 72
    tachypnea | 72
    discontinued metronidazole | 168
    LMWH discontinued | 240
    dismissed for home care | 336
    referred to hematologist | 336
    no septic emboli | 0
    no endometritis | 0
    no parametritis | 0
    no pelvic abscess | 0
    no cesarean section wound infection | 0
    no episiotomy infection | 0
    no vaginal lacerations | 0
    no cervical lacerations | 0
    no mastitis | 0
    no drug-induced fever | 0
    no urinary tract infection | 0
    no other infections | 0
    no recurrence | 0
    no other thrombogenic diseases | 0
