60 years old | 0  
    male | 0  
    arterial hypertension | 0  
    visited emergency department | -384  
    fever | -384  
    chills | -384  
    malaise | -384  
    fatigue | -384  
    anorexia | -384  
    left flank pain | -384  
    abrupt onset of chills | -384  
    nausea | -384  
    vomiting | -384  
    diarrhea | -384  
    vomiting subsided | -312  
    diarrhea subsided | -312  
    chills remained | -312  
    malaise remained | -312  
    treated with amoxicillin-clavulanic acid | -312  
    malaise worsened | -312  
    fatigue worsened | -312  
    fever up to 40°C | -312  
    left flank pain developed | -312  
    hematuria | -312  
    diarrhea reappeared | -312  
    sepsis | 0  
    febrile (38.5°Celsius) | 0  
    hypotensive (90/50 mmHg) | 0  
    tachypneic (26 breaths per minute) | 0  
    tachycardic (135 beats per minute) | 0  
    enlarged left kidney | 0  
    leukocytosis (17,280 cells/mL) | 0  
    neutrophilia (15,260 cells/mL) | 0  
    elevated C-reactive protein (388.38 mg/L) | 0  
    elevated procalcitonin (10.61 ng/mL) | 0  
    elevated creatinine (2.68 mg/dL) | 0  
    elevated urea (45.93 mg/dL) | 0  
    diagnosed with pyelonephritis | 0  
    diagnosed with sepsis | 0  
    admitted to intensive care unit | 0  
    parenteral fluids | 0  
    antimicrobial therapy (cefotaxime) | 0  
    blood culture Salmonella enterica | 0  
    urine culture Salmonella enterica | 0  
    resistant to cefuroxime | 0  
    resistant to ciprofloxacin | 0  
    resistant to gentamicin | 0  
    resistant to amikacin | 0  
    susceptible to ampicillin | 0  
    susceptible to cefotaxime | 0  
    susceptible to meropenem | 0  
    susceptible to trimethoprim/sulfamethoxazol | 0  
    Clostridioides difficile antigen positive | 0  
    Clostridioides difficile toxin positive | 0  
    trimethoprim/sulfamethoxazole added | 0  
    oral vancomycin added | 0  
    transthoracic echocardiography | 0  
    native CT abdomen | 0  
    echocardiography unremarkable | 0  
    discrete inflammatory changes of fat around left kidney | 0  
    contrast not used | 0  
    treated with cefotaxime | 0  
    treated with trimethoprim/sulfamethoxazole | 0  
    discharged | 240  
    oral trimethoprim/sulfamethoxazole continued | 240  
    arbitrarily stopped antimicrobial therapy | 288  
    visited emergency department again | 336  
    progressive weakness | 336  
    night sweating | 336  
    dull pain in lumbar and sacral region | 336  
    elevated CRP (66.33 mg/L) | 336  
    physical examination unremarkable | 336  
    abdominal ultrasound unremarkable | 336  
    admitted | 336  
    parenteral ceftriaxone | 336  
    oral vancomycin | 336  
    blood culture Salmonella enterica | 336  
    magnetic resonance imaging of lumbar spine | 336  
    no vertebral affection | 336  
    dilatation of infrarenal part of abdominal aorta | 336  
    contrast CT abdomen | 336  
    fusiform aneurysm of abdominal aorta | 336  
    aneurysm of left internal iliac artery | 336  
    saccular aneurysm | 336  
    compressed left ureter | 336  
    dilated left ureter | 336  
    grade 2 hydronephrosis | 336  
    conservative therapy recommended | 336  
    treated with ceftriaxone | 336  
    CT follow-up progression of aneurysm diameter | 672  
    infrarenal aorta recanalized | 672  
    surgery with ligation of left internal iliac artery | 672  
    partial extirpation of aneurysm | 672  
    tight adhesions between aneurysm and left ureter | 672  
    abdominal aorta aneurysm left intact | 672  
    histologic examination nonspecific inflammation | 672  
    cultures sterile | 672  
    parenteral antimicrobial therapy | 672  
    CT follow-up complete obliteration of residual aneurysm | 840  
    discharged | 840  
    oral trimethoprim/sulfamethoxazole continued | 840  
    asymptomatic at 3-month follow-up | 2160  
    CRP level in reference range | 2160  
    
