32 years old | 0
    female | 0
    Raynaud's phenomenon | 0
    recurrent urinary tract infection | 0
    presented to an outside hospital | -120
    UTI symptoms | -120
    developed shortness of breath | -48
    hypotensive | -48
    altered | -48
    Pressors initiated | -48
    broad spectrum antibiotics initiated | -48
    vancomycin initiated | -48
    cefepime initiated | -48
    metronidazole initiated | -48
    blood cultures obtained | -48
    urine cultures obtained | -48
    E. coli infection | -48
    enterobacter infection | -48
    antibiotic coverage narrowed to cefepime | -48
    anemia | -48
    thrombocytopenia | -48
    coagulopathy | -48
    transfusion of 3 units of platelets | -48
    transfusion of 2 units of red blood cells | -48
    fresh frozen plasma transfusion | -48
    hyponatremic | -48
    sodium 117 mmol/L | -48
    brain MRI obtained | -48
    lumbar puncture obtained | -48
    developed acute respiratory distress | -48
    intubation | -48
    elevated creatinine 6.4 mg/dL | -48
    baseline creatinine 0.6 mg/dL | -48
    urinalysis 3+ blood | -48
    urinalysis 3+ leukocytes | -48
    urinalysis 3+ protein | -48
    urinalysis 4+ bacteria | -48
    continuous renal replacement therapy initiated | -48
    improvement in renal function | -48
    CT abdomen and pelvis obtained | -48
    enlarged kidneys | -48
    hepatosplenomegaly | -48
    developed persistent agitation | -48
    transfer to medical intensive care unit | 0
    anemia | 0
    thrombocytopenia | 0
    hemoglobin 7.6 g/dL | 0
    platelet count 15,000 k/cu mm | 0
    profound leukocytosis | 0
    white blood cell count 30.78k/cu mm | 0
    anion gap metabolic acidosis | 0
    bicarbonate 20 mmol/L | 0
    anion gap 18 | 0
    elevated lactate 5.6 mmol/L | 0
    hyponatremic | 0
    sodium 128 mmol/L | 0
    creatinine 1.8 mg/dL | 0
    differential considerations | 0
    infiltrative diseases | 0
    idiopathic Castleman disease | 0
    malignancy | 0
    IgG4-related disease | 0
    granulomatous disease | 0
    repeat CT abdomen and pelvis with IV contrast obtained | 0
    bilateral nephromegaly | 0
    heterogeneous renal parenchymal enhancement | 0
    loss of corticomedullary differentiation | 0
    focal wedge-shaped hypodensities | 0
    superimposed necrosis | 0
    cinematic rendering CT data | 0
    inflammatory changes in both kidneys | 0
    bilateral renal abscesses | 0
    differential considerations | 0
    infiltrative bilateral renal disease | 0
    glomerulonephritis | 0
    lymphoma | 0
    renal cell carcinoma | 0
    renal biopsy obtained | 0
    recovery of platelet counts | 0
    histiocytic cells infiltration | 0
    focal abscesses | 0
    Gram stain negative | 0
    Gram Weigert stain negative | 0
    Von Kossa stain positive | 0
    Michaelis-Gutman bodies | 0
    CD163 immunostain diffusely positive | 0
    macrophages infiltration | 0
    histiocytes infiltration | 0
    pyelonephritis | 0
    focal micro-abscesses | 0
    malakoplakia | 0
    ultrasound imaging obtained | 0
    left renal biopsy | 0
    right upper quadrant ultrasound | 0
    left nephromegaly | 0
    right nephromegaly | 0
    multiple renal abscesses | 0
    MRI obtained | 0
    bilateral nephromegaly | 0
    intrarenal fluid collections | 0
    perinephric fluid collections | 0
    mild left hydronephrosis | 0
    thickening of left renal pelvis | 0
    thickening of left perinephric fascia | 0
    retroperitoneal soft tissues involvement | 0
    treatment options considered | 0
    antibiotics with intracellular penetration | 0
    tigecycline chosen | 0
    resistance profile considered | 0
    ceftriaxone used | 0
    bethanechol initiated | 0
    vitamin C initiated | 0
    switched to minocycline | 0
    nephrectomy considered | 0
    deferred due to liver involvement | 0
    liver biopsy obtained | 0
    no hepatic malakoplakia | 0
    nephrectomy forgone | 0
    creatinine returned to normal | 0
    leukocytosis | 0
    low-grade fevers | 0
    subsequent MRI showed progression | 0
    extension to left perinephric space | 0
    retroperitoneum involvement | 0
    scheduled for radical left nephrectomy | 0
