52 years old | 0
male | 0
Egyptian | 0
admitted to the hospital | 0
neck pain | -168
dysphagia | -168
difficulty breathing | -168
goiter | -10080
thyroidectomy | -504
post-operative hematoma | -504
evacuation of hematoma | -504
placement of Jackson-Pratt wound drain | -504
bleeding diathesis | -504
anterior neck enlargement | 0
neck tenderness | 0
prothrombin time (PT) | 0
international normalized ratio (INR) | 0
partial thromboplastin time (PTT) | 0
fibrinogen | 0
computerized tomography (CT) scan | 0
neck hematoma | 0
evacuation of neck hematoma | 24
desmopressin (DDAVP) | 24
discharged | 48
severe oral mucosal bleeding | 4320
admitted to the intensive care unit (ICU) | 4320
multiple transfusions | 4320
red blood cells | 4320
platelets | 4320
fresh frozen plasma (FFP) | 4320
DDAVP | 4320
Humate-P | 4320
aminocaproic acid | 4320
surgical packing | 4320
bleeding diathesis workup | 4320
PTT | 4320
Factor II | 4320
Factor V | 4320
Factor VII | 4320
Factor VIII | 4320
Factor IX | 4320
Factor X | 4320
Factor XI | 4320
Factor XII | 4320
Von Willebrand Factor antigen | 4320
Von Willebrand Multimers | 4320
PT/INR | 4320
abdominal pain | 5760
massive hepatosplenomegaly | 5760
coagulopathy workup | 5760
factor VII deficiency | 5760
transjugular biopsy of liver | 5760
prophylactic rFVIIa | 5760
liver biopsy | 5760
AL-amyloidosis-Kappa type | 5760
bleeding at transjugular biopsy site | 5832
retroperitoneal hematoma | 5832
rFactor VIIa infusions | 5832
treatment for AL-amyloidosis-Kappa type | 6312
bortezomib | 6312
dexamethasone | 6312
cyclophosphamide | 6312
colchicine | 7056
prednisone | 7056
GI bleeding | 7056
spontaneous bacterial peritonitis (SBP) | 7056
hepatic encephalopathy | 7056
uncontrolled upper GI hemorrhage | 8760
death | 8760