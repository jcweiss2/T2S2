49 years old | 0
male | 0
obese | 0
BMI-33.9 | 0
ethanol related decompensated liver cirrhosis | -672
recurrent life threatening variceal bleeds | -672
mild ascites | -672
jaundice | -672
CTP score −9 | -672
Child: B | -672
MELD Na: 17 | -672
no previous history of hypertension | 0
no previous history of diabetes | 0
no previous history of asthma | 0
admitted to the hospital | 0
live donor liver transplant | 0
partial MHV right lobe graft | 0
splenic artery ligation | 0
intraoperative course was uneventful | 0
extubated on post-operative day one | 24
post-operative doppler of the recipient showed high portal blood flows | 24
pharmacologically modulated with octreotide infusion | 24
intravenous methylprednisolone 10 mg/kg | 0
tapered to 100 mg | 24
tapered to 80 mg | 48
tapered to 60 mg | 72
tapered to 40 mg | 96
switched over to oral wysolone 20 mg once daily | 120
started on tacrolimus | 48
tacrolimus trough level 8-10 ng/ml | 48
started on mycophenolate mofetil | 192
rising aminotransferases | 120
methylprednisolone pulse therapy | 120
acute cellular rejection | 120
satisfactory hospital course | 480
developed fever | 480
temperature was 101°F | 480
heart rate 110 per minute | 480
respiratory rate 26 per minute | 480
drop in saturation to 88% on ambient air | 480
RT-PCR from nasopharyngeal swab detected the presence of severe acute respiratory syndrome coronavirus-2 | 480
nasopharyngeal aspirate was negative for all other respiratory viruses | 480
immunosuppression was modified | 480
MMF was stopped | 480
oral steroid was changed to intravenous hydrocortisone | 480
tacrolimus in low dose was continued | 480
oxygen saturation was maintained between 94% and 96% with high-flow nasal cannula oxygen therapy | 480
became increasingly tachypnoeic | 504
chest x-ray showed patchy parenchymal bilateral opacities | 504
pre-emptively shifted to intensive care isolation | 504
blood tests for inflammatory markers | 504
started on injection remdesivir | 504
subcutaneous enoxaparin 60 mg | 504
non-invasive ventilation | 504
rapid clinical deterioration of his oxygenation | 528
elevated inflammatory markers | 528
decided against administration of tocilizumab | 528
thrombocytopenia continued to persist | 528
decided to treat him with fresh convalescent plasma | 528
transfused 1st aliquot of 200 ml plasma | 528
transfused 2nd aliquot of 230 ml plasma | 552
transfused 3rd plasma aliquot of 200 ml | 576
showed good recovery | 600
inflammatory markers improved | 600
off oxygen therapy | 960
absolute lymphocyte count increased | 960
radiological resolution of the lung opacities | 960
aminotransferases and total bilirubin continued to show progressive improvement | 960
repeat nasopharyngeal swabs for COVID-19 RT-PCR done thrice | 960
discharged | 1152