47 years old | 0
male | 0
admitted to the hospital | 0
melaena | -168
proximal muscle weakness | -504
weight loss | -504
right hip pain | -336
low energy fall | -336
non-functional pancreatic head neuroendocrine tumour | -5184
pylorus-preserving pancreaticoduodenectomy | -5184
pancreatin | -5184
basal-bolus insulin regime | -5184
insulin glargine | -5184
insulin aspart | -5184
sinus tachycardia | 0
blood pressure 128/63 mm Hg | 0
bilateral pitting oedema | 0
melaena on digital rectal examination | 0
haemoglobin 85 g/L | 0
urea 8.3 mmol/L | 0
creatinine 77 μmol/L | 0
hypokalaemia 2.9 mmol/L | 0
liver function tests | 0
coagulation profile | 0
albumin 41 g/L | 0
2D transthoracic echocardiogram | 0
oesophago-gastro-duodenoscopies | 0
colonoscopy | 0
video capsule endoscopy | 0
CT scan | 0
portal hypertension | 0
variceal dilatation | 0
sub-acute right pubic rami fractures | 0
gallium-68 DOTATATE positron emission tomography | 0
tumour recurrence | 0
invasion of the superior mesenteric vein | 0
porto-mesenteric hypertension | 0
bleeding mesenteric varices | 0
blood transfusions | 24
potassium replacement | 24
lanreotide autogel | 24
discharged | 24
septic shock | 168
Escherichia coli bacteraemia | 168
cytomegalovirus viraemia | 168
discharged to inpatient rehabilitation facility | 336
proximal myopathy | 504
lower back pain | 504
unexplained ecchymosis | 504
hypertension 162/107 mm Hg | 504
oedema | 504
hypokalaemia 2.9 mmol/L | 504
hypernatraemia 148 mmol/L | 504
metabolic alkalosis | 504
osteoporotic vertebral compression fractures | 504
24-h urinary free cortisol collection | 504
low-dose dexamethasone test | 504
Cushing's syndrome | 504
elevated ACTH levels | 504
high-dose dexamethasone suppression test | 504
ectopic ACTH source | 504
pituitary MRI | 504
repeat gallium-68 DOTATATE PET scan | 504
metyrapone | 504
ketoconazole | 504
hydrocortisone replacement | 504
discharged home | 576
lanreotide therapy | 576
reduction in tumour size | 576
community physiotherapy | 576
near pre-morbid performance status | 576
plans to start chemotherapy | 576