50 years old | 0
male | 0
urinary lithiasis | -12000
left renal shockwave lithotripsy | -10920
right pyelotomy | -10560
parathyroidectomy | -10320
left colic pain | 0
mild hyperpyrexia | 0
urinalysis | 0
mixed low burden microbial germs | 0
non-constrast medium CT scan | 0
bilateral lithiasis | 0
left ureteral stenting | 0
antibiotic therapy | 0
Meropenem | 0
Gentamicin | 0
elective left endoscopic combined intrarenal surgery | 0
pre-operative urinalysis | 0
Amoxicillin + clavulanic acid | 0
Valdivia Galdakao position | 0
3-unsuccessful renal puncture | 0
f-URS laser lithotripsy | 0
ureteral access sheath | 0
fever | 24
blood cultures | 24
empirical antibiotic therapy | 24
Tazobactam | 24
Teicoplanin | 24
CT scan | 24
pyelonephritis | 24
antibiotic therapy modified | 48
Meropenem | 48
Linezolid | 48
Pseudomonas Aeruginosa | 48
haemodynamically unstable situation | 72
tachycardia | 72
hypotension | 72
thoracic/abdomen CT scan | 96
pulmonary septic emboli | 96
bilateral pleural effusion | 96
left renal abscess | 96
CT-guided renal drain | 96
ureteral stent replaced | 96
feverish | 240
CT scan | 240
no change from previous control | 240
multidisciplinary counselling | 240
left open nephrectomy | 240
not pyretic | 264
decreasing inflammation indexes | 264
discharged | 336
histological examination | 336
multifocal Xanthogranulomatous pyelonephritis | 336