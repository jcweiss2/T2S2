11 years old | 0
male | 0
admitted to the hospital | 0
acute abdominal pain | -24
abdominal pain started | -24
pushing another boy in a wheelchair | -24
pain worsened | -24
intermittent projectile vomiting | -24
no fever | -24
no chills | -24
no diarrhoea | -24
no bloody stool | -24
otherwise healthy | -24
no medical history | -24
no surgical history | -24
no relevant drug history | -24
no family history | -24
no psychosocial history | -24
no genetic history | -24
septic | 0
lethargic | 0
severely dehydrated | 0
temperature 37.5°C | 0
pulse 157 bpm | 0
blood pressure 97/41 mmHg | 0
moderately distended abdomen | 0
generalised guarding | 0
rebound tenderness | 0
digital rectal examination unremarkable | 0
other systems unremarkable | 0
dehydration | 0
blood urea 10.3 mmol/l | 0
serum creatinine 87 umol | 0
elevated white cell count 14,700/mm3 | 0
haemoglobin 16.8 g/dl | 0
fluid resuscitation | 0
catheterised | 0
nasogastric tube inserted | 0
oxygen administered | 0
taken for surgery | 0
laparotomy | 0
gangrenous small bowel loops | 0
mesenteric cyst | 0
no normal small bowel visible | 0
ischemic loops of bowel | 0
opening in the mesenteric cyst | 0
viable small bowel loops | 0
gangrenous loop of terminal ileum | 0
resection of gangrenous bowel | 0
peritoneal capsule excised | 0
primary jejunum to ascending colon anastomosis | 0
abdomen irrigated | 0
abdomen closed primarily | 0
inotropic support required | 0
post-operative concerns | 0
sepsis | 0
anastomotic leak | 0
short bowel syndrome | 0
inotropic support weaned off | 96
extubated | 96
broad spectrum antibiotics continued | 96
abdominal examination showed no signs of anastomotic leak | 96
discharged | 216
follow-up care | 4320
no clinical evidence of short-bowel syndrome | 4320
no significant morbidity | 4320
peritoneal encapsulation diagnosed | 0
asymptomatic peritoneal encapsulation | -24
acute increase in intra-abdominal pressure | -24
loop of ileum herniated | -24
strangulated | -24
diarrhoea | 216
diarrhoea resolved | 4320
vitamin B12 deficiency considered | 216
fat malabsorption considered | 216
anaemia considered | 216