39 years old | 0
male | 0
arrived at emergency department | 0
endotracheally intubated | 0
medical attention sought five hours after suicidal attempt | -5
suicidal attempt | -5
drain cleaner liquid ingestion | -5
sodium hydroxide | -5
potassium hydroxide | -5
carbonyl diamide | -5
free previous medical history | 0
edematous oral mucosa | 0
chemical injuries to the face | 0
white blood cell count of 12.9 × 103/μL | 0
D-dimer > 5250 ng/mL DDU | 0
chest CT thickening of esophageal and gastric wall | 0
submucosal edema of esophageal and gastric wall | 0
trace para-esophageal stranding | 0
peri-gastric stranding | 0
fluid | 0
no free air | 0
tracheo and broncho esophageal fistulas | 0
massive aspiration | 0
cardiac arrest | 0
proton pump inhibitor | 0
intravenous fluids | 0
prophylactic antibiotics | 0
tracheostomy placement | 312
jejunostomy tube placement | 312
bouts of coughing during sedation-awakening trials | 432
reduction in sedatives | 432
acute hypoxia | 432
oxygen saturation decreased to 50% | 432
pulseless electrical arrest | 432
cardiopulmonary resuscitation | 432
recovery of spontaneous circulation | 432
frothy, yellow-tinted secretions from tracheostomy | 432
no oral secretions during oral cavity suction | 432
nasogastric tube placement | 432
gastric cavity decompression | 432
400-500 mL of fluid suctioned | 432
chest X-ray bibasilar atelectasis | 432
chest X-ray patchy airspace opacities | 432
acute respiratory distress syndrome | 528
recurrent septic shock | 528
aspiration pneumonia | 528
liberated from mechanical ventilation | 960
transition to tracheostomy collar | 960
enteral nutrition through jejunostomy tube | 960
left intensive care unit | 960
discharged home | 2736
endoscopy surveillance progression | 2736
endoscopy surveillance further extend of disease | 2736
bronchoscopy on day 1 | 24
bronchoscopy on day 8 | 192
bronchoscopy after 17 weeks | 2856
new tracheoesophageal fistula | 2856
esophageal lumen opening at mid trachea | 2856
bronchoscopy at 7 weeks | 1176
protrusion of esophageal stent through BEF | 1176
esophagoduodenoscopy at 7 months | 4872
visualization of tracheostomy tube through combined lumen | 4872
double lumen identified | 4872
complete obliteration of stent | 4872
in-growth tissues | 4872
referred for cardiothoracic surgical evaluation | 4872
nutritional optimization | 4872
potential surgical intervention | 4872
admission to hospital/ICU | 0
EGD #1 | 0
bronchoscopy #1 | 24
bronchoscopy #2 | 192
cardiac arrest | 432
esophageal stent placement with EGD #2 | 528
bronchoscopy #3 | 1176
hospital discharge | 2736
bronchoscopy #4 | 2856
EGD #3 | 4872
