59 years old | 0
male | 0
Thai | 0
admitted to the hospital | 0
dry weight 43.6 kg | 0
septic shock | -72
candidemia | -72
vasopressor | -72
norepinephrine | -72
intensive monitoring | -72
hemodynamic instability | -72
acute progressive dyspnea | -72
new-onset ascites | -72
low albumin gradient | -72
high protein | -72
type 2 diabetes | 0
hypertension | 0
old pulmonary tuberculosis | 0
end-stage renal disease | 0
no residual urine output | 0
hemodialysis | 0
triple vessel disease | 0
left ventricular ejection fraction 27% | 0
peripheral artery disease | 0
chronic limb ischemia | 0
dry gangrene | 0
left percutaneous transluminal angioplasty stent | 0
femoral artery endarterectomy | 0
dyspnea | -72
emergency multidetector computed tomography angiography | -72
suspected acute pulmonary embolism | -72
small thrombus in the right atrium | -72
central venous catheter | -72
enoxaparin sodium prefilled syringe | -24
Clexane 4000 IU | -24
40 mg SC once daily | -24
bodyweight 46.8 kg | -24
RA thrombus treatment | -24
anti-Xa level evaluation | -24
4 h after the dose | -24
9 p.m. | -24
non-hemodialysis day | -24
renal impairment | -24
bleeding risk | -24
major bleeding events | -24
retroperitoneal bleeding | -24
intracranial bleeding | -24
anti-Xa level monitoring | -24
peak anti-Xa level | -24
0.5-1 IU/mL | -24
abdominal wall injection | -24
local edema | -24
peripheral edema | -24
ascites | -24
weight gain 6 kg | -24
abdominal paracentesis | -24
TCC removal | -72
enoxaparin hold | -72
4 days | -72
surgery | -72
bleeding | -72
clots in the endotracheal tube | -72
enoxaparin withhold | -72
2 days | -72
airway mucosal injuries | -72
localized inflammation of trachea and bronchi | -72
acquired platelet dysfunction | -72
renal failure | -72
persistent thrombus in the RA | -24
cardiologist examination | -24
repeated echocardiogram | -24
enoxaparin restart | -24
40 mg SC OD | -24
anti-Xa level monitoring | -24
peak anti-Xa level 0.3 IU/mL | -24
subtherapeutic | -24
enoxaparin dose increase | -24
60 mg SC OD | -24
1.17 mg/kg/dose | -24
current bodyweight 55 kg | -24
peak anti-Xa level 0.25 IU/mL | -24
ascites interference | -24
SC enoxaparin absorption | -24
deltoid injection | -24
peak anti-Xa levels 0.45 and 0.51 IU/mL | -24
therapeutic range | -24
enoxaparin dose maintenance | -24
hemodialysis | -24
endotracheal tube bleeding | -24
vasopressor dose | -24
norepinephrine | -24
average norepinephrine doses | -24
abdominal paracentesis | -24
hemodialysis day | -24
TCC removal | -72
enoxaparin hold | -72
surgery | -72
bleeding | -72
clots in the endotracheal tube | -72
enoxaparin withhold | -72
2 days | -72
discharge | 720