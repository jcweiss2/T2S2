17 years old | 0
female | 0
black African | 0
admitted to local clinic | -336
bi-frontal headache | -336
insomnia | -336
subjective fevers | -336
treated for non-specific infection | -336
empiric antibiotics | -336
restlessness | -326
third-person auditory hallucinations | -326
referred to psychiatrist | -326
diagnosed with acute schizoaffective disorder | -326
psychological stressors | -326
death anniversary of mother | -326
final high-school national examinations | -326
admitted to hospital | -321
treated with psychotropic medication | -321
documented fevers | -316
orofacial dyskinesias | -316
tongue-biting | -316
agitation | -316
treated for neuroleptic malignant syndrome | -316
comatose | -316
transferred to tertiary referral hospital | -316
temperature of 39°C | 0
tachycardia | 0
Glasgow Coma Scale 7/15 | 0
grimacing | 0
tongue biting | 0
bruxism | 0
hyper-salivation | 0
abnormal arm movements | 0
intubated | 0
mechanically ventilated | 0
admitted to ICU | 0
investigations for infection | 0
auto-immune disease | 0
toxic causes | 0
polymerase chain reaction for tropical fever pathogens | 0
contrast-enhanced computed tomography scan | 0
cerebrospinal fluid examination | 0
elevated pressures | 0
white cell count of 115/mm3 | 0
lymphocytes | 0
negative PCR for bacterial | 0
tuberculosis | 0
herpes meningo-encephalitis pathogens | 0
contrast-enhanced MRI brain scan | 0
leptomeningeal enhancement | 0
sulcal hyperintensities | 0
electroencephalography | 0
non-specific diffuse slowing | 0
no epileptiform discharges | 0
treated for viral encephalitis | 0
stopped treatment | 24
diagnosed with probable NMDARE | 48
commenced immunosuppression | 48
high-dose intravenous methylprednisolone | 48
intravenous immunoglobulins | 48
orofacial and upper limb movement disorders | 48
controlled with levetiracetam | 48
tetrabenazine | 48
midazolam | 48
propofol infusions | 48
maxillo-mandibular fixation | 48
serum and CSF autoimmune encephalitis panels | 168
positive for antibodies against NMDA receptor | 168
definite diagnosis of NMDARE | 168
MRI pelvis | 168
no ovarian or extra-gonadal teratoma | 168
repeat MRI brain scan | 360
resolution of meningeal enhancement | 360
sulcal hyperintensities | 360
GCS remained low at 8/15 | 360
unrelenting dyskinesias | 360
required higher sedation | 360
repeated IVMP course | 360
concurrent plasma exchange | 360
weekly rituximab | 360
ICU stay complicated by right brachial deep vein thrombosis | 360
treated with low-molecular weight heparin | 360
tongue maceration | 360
required surgical debridement | 360
tracheostomy | 360
percutaneous endoscopic gastrostomy tubes | 360
high-grade fevers | 720
multi-drug resistant Pseudomonas aeruginosa | 720
Klebsiella pneumoniae | 720
isolated from tracheal aspirates | 720
tracheostomy site | 720
septic shock | 720
multi-organ dysfunction | 720
succumbed | 720