28 years old | 0
female | 0
hypothyroidism | 0
hypertension | 0
polycystic ovarian syndrome | 0
admitted to the hospital | 0
fever | -504
myalgias | -504
nausea | -504
vomiting | -504
worked as a paramedic | -504
involved in the care of a SARS-CoV-2-positive patient | -504
initial physical examination | 0
unremarkable physical examination | 0
qualitative BioFire SARS-CoV-2 PCR screen | 0
SARS-CoV-2 virus not detected | 0
febrile | 0
temperature up to 105 °F | 0
upgraded to the intensive care unit | 24
repeat physical examination | 24
palpable liver | 24
no associated rash | 24
no mucosal ulcers | 24
no lymphadenopathy | 24
full septic workup | 24
blood cultures negative | 24
urine cultures negative | 24
acute viral hepatitis panels | 24
hepatitis B virus core immunoglobulin M antibody nonreactive | 24
hepatitis B virus surface antigen nonreactive | 24
hepatitis c virus antibody nonreactive | 24
hepatitis A IgM antibody nonreactive | 24
Monospot testing for EBV infection positive | 24
elevated EBV IgM titers | 24
EBV-PCR positive | 24
computed tomography scan of the chest | 24
unremarkable computed tomography scan of the chest | 24
computed tomography scan of the abdominal | 24
new hepatosplenomegaly | 24
liver measuring 25 cm | 24
repeat qualitative BioFire SARS-CoV-2 PCR screen | 48
SARS-CoV-2 virus detected | 48
transaminitis | 48
developed transaminitis | 48
Hematology/Oncology specialists consulted | 48
concern for early hemophagocytic lymphohistocytosis | 48
ferritin elevated | 48
fibrinogen elevated | 48
triglyceride levels elevated | 48
suspicion of HLH | 48
diagnostic liver biopsy suggested | 48
bone marrow biopsy suggested | 48
biopsies declined by the patient | 48
rituximab started | 72
transferred to a tertiary care center | 96
discharged | 120