78 years old | 0
female | 0
admitted to the emergency department | 0
abdominal pain | 0
hypotension | 0
leukocytosis | 0
pyuria | 0
no increased left hip pain | 0
no edema or erythema surrounding the left hip | 0
initial left total hip arthroplasty | -156
osteoaarthritis | -156
revision of the left total hip arthroplasty | -120
acetabuloplasty with medial acetabular bone grafting | -120
placement of a unipolar hemiarthroplasty | -120
progressive left hip pain | -110
superomedial migration of the unipolar head | -110
placement of an antiprotrusio cage | -30
cervical squamous-cell carcinoma | -216
total hysterectomy | -216
lymphoma | -216
chemotherapy | -216
splenectomy | -216
CT scan of the abdomen and pelvis | 0
small bowel dilatation | 0
severe left hip protrusio | 0
medial migration of the acetabular hardware | 0
hardware penetrating the wall of the sigmoid colon | 0
fluid and gas surrounding the left hip and greater trochanter | 0
sigmoid colon perforation | 0
fistula to the left hip joint and periarticular soft tissues | 0
CT-guided aspiration of the fluid collection | 0
fecal material | 0
Escherichia coli | 0
Streptococcus viridans | 0
Clostridium perfringens | 0
surgery | 24
sigmoidectomy | 24
Hartmann procedure | 24
end-sigmoid colostomy | 24
omental coverage of the hardware | 24
lateral incision over the left hip | 24
brown fluid in the subcutaneous tissues | 24
vastus lateralis muscle involvement | 24
left hip involvement | 24
debridement | 24
cultures from the left hip | 24
Escherichia coli | 24
Streptococcus viridans | 24
Clostridium perfringens | 24
hardware removal | 48
hip disarticulation | 48
femoral hardware removal | 48
partial acetabular hardware removal | 48
femoral-femoral arterial bypass | 48
septicemia | 48
intensive care unit | 48
gastrointestinal bleeding | 336
infected left pelvic hematoma | 336
osteomyelitis of the proximal left femur | 336
decompression of the hematoma | 336
serial irrigation and debridements | 336
removal of remaining acetabulum hardware | 336
congestive heart failure | 336
aspiration | 336
hypotensive | 744
death | 744