5 days old neonate | 0
admitted to neonatal intensive care unit | 0
absence of anal orifice | 0
no meconium passed for 48 hours | -48
meconium passed through urethral orifice | 0
urine passed through urethral orifice | 0
abdominal swelling | 0
no fever | 0
no yellowish discoloration of skin and eyes | 0
no vomiting | 0
no abnormal body movement | 0
female-looking external genitalia | 0
enlarged clitoris | 0
32-year-old para-four mother | 0
amenorrheic for nine months | -6048
antenatal care | -6048
spontaneous vaginal delivery | 0
labor for 14 hours | -14
birth weight 3.2kg | 0
cried immediately after birth | 0
APGAR scores 7 at 1 minute | 0
APGAR scores 10 at 10 minutes | 0
no chronic medical illnesses | 0
prior healthy children | 0
alert general appearance | 0
pulse rate 152 beats per minute | 0
respiratory rate 46 breaths per minute | 0
temperature 36°C | 0
venous oxygen saturation 97% | 0
head circumference 42 cm | 0
anterior fontanel size 2cm | 0
abdomen grossly distended | 0
no anal opening | 0
sacrococcygeal dimple | 0
female external genitalia | 0
labia majora well developed | 0
no fusion of labia majora | 0
labia minora fused to clitoris base | 0
no vaginal opening | 0
phallus 0.8cm | 0
central opening leaking stool | 0
common urethral opening | 0
no palpable gonads | 0
white blood cell 20,000 | 0
neutrophil 53% | 0
lymphocyte 23% | 0
red blood cell 5*10^6 | 0
hemoglobin 15gm/dl | 0
platelet 272*10^3 | 0
blood group A+ | 0
random blood sugar 120gm/dl |8
plain abdominal x-ray | 0
absence of air shadow in distal large bowel | 0
abdominopelvic sonography | 0
left supernumerary kidney | 0
left kidney in renal fossa | 0
left supernumerary kidney on psoas muscle | 0
distinct capsules and blood supply | 0
contralateral single normal kidney | 0
collapsed bladder | 0
diagnosis of cloacal anomaly | 0
diagnosis of ambiguous genitalia | 0
diagnosis of supernumerary kidney | 0
diagnosis of early onset neonatal sepsis | 0
managed with maintenance fluid | 0
intravenous antibiotics | 0
ampicillin 150mg/kg/dose BID | 0
gentamicin 3mg/kg/dose daily | 0
referred to specialized hospital | 48
