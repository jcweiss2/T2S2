10 years old|0
male|0
fever| -168
impetigo| -144
diarrhea| -24
medical history unremarkable|0
family history unremarkable|0
acutely ill|0
uncomfortable|0
irritable|0
unable to stand|0
unable to converse normally|0
heart rate 147 beats/min|0
blood pressure 101/61 mmHg|0
temperature 40.5˚C|0
respiratory rate 42 breaths/min|0
oxygen saturation 100%|0
no nuchal rigidity|0
lung fields clear|0
cheek erythema|0
pharyngeal erythema|0
impetigo on forehead|0
impetigo on jaw|0
abdominal tenderness|0
swelling in left elbow|0
redness in left elbow|0
tenderness in left elbow|0
swelling in left ankle joints|0
redness in left ankle joints|0
tenderness in left ankle joints|0
rapid antigen detection test positive for Group A Streptococcus pharyngitis|0
blood culture positive for Streptococcus pyogenes|0
throat culture positive for Streptococcus pyogenes|0
impetigo pus culture positive for Streptococcus pyogenes|0
minimum inhibitory concentration against ampicillin ≤0.06 µg/ml|0
minimum inhibitory concentration against clindamycin ≤0.12 µg/ml|0
contrast-enhanced CT scan increased fat concentration around cutaneous veins of left lower leg|0
diagnosis of STSS|0
coagulopathy|0
liver involvement|0
generalized erythematous macular rash|0
isolation of Group A Streptococcus|0
DIC score 6 points|0
diagnosis of infectious-type DIC|0
admitted to ICU|0
blood pressure within normal range|0
aggressive intravenous rehydration|0
intravenous amoxicillin-sulbactam|0
intravenous clindamycin|0
intravenous immunoglobulins|0
blood cultures negative on day 3|72
fever persisted until day 10|240
rhTM administration|0
antithrombin-III administration|0
general condition poor on day 2|48
fever persisted on day 2|48
DIC score increased from 5 to 9 points on day 2|48
platelet count ≥30% decrease within 24 h|48
TAT +1 point|48
danaparoid administration on day 2|48
general condition improved after danaparoid + rhTM|48
laboratory findings became less alarming|48
DIC score decreased to 4 points on day 3|72
fibrin degradation products -1 point|72
DIC resolved|72
redness in left lower leg worsening|168
swelling in left lower leg worsening|168
pain in left lower leg worsening|168
redness in left elbow joint worsening|168
swelling in left elbow joint worsening|168
contrast-enhanced CT scan on day 7|168
progressive increase in fat concentration|168
ring-shaped contrast enhancement of left popliteal vein|168
LRINEC score 8|168
skin biopsy performed|168
diagnosis of spongiotic dermatitis|168
diagnosis of suppurative panniculitis|168
soft tissue did not progress to necrosis|168
range of motion of joint not improved|216
MRI performed on day 9|216
MRI showed inflammatory findings in left soleus|216
MRI showed inflammatory findings in left gastrocnemius|216
MRI showed inflammatory findings between the two muscles|216
arthritis not evident|216
osteomyelitis not evident|216
condition improved gradually|216
recovery in legs|216
able to walk|216
discharged on day 20|480
no sequelae|480
no medication-related adverse events|480
no signs of disease during four years of follow-up|480
life returned to regular rhythm|480
