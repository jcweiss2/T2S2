33 years old | 0
female | 0
childhood history of hydronephrosis | -10000
vesicoureteral reflux | -10000
9-year history of erythroderma | -7872
confluent folliculocentric erythematous scaly plaques | -7872
islands of sparing | -7872
orange palmoplantar hyperkeratosis | -7872
eczematous lesions | -7872
differential diagnoses included PRP | -100
differential diagnoses included psoriasis | -100
differential diagnoses included atopic dermatitis | -100
differential diagnoses included epidermotropic cutaneous T-cell lymphoma | -100
search for skin and blood T-cell clone was negative | -100
blood screening did not show Sezary cells | -100
blood screening did not show phenotypically atypical lymphocytes | -100
whole genome sequencing did not find any possible causal mutation | -100
CARD14 sequencing did not find any possible causal mutation | -100
skin biopsy specimens showed epidermal acanthosis | -100
skin biopsy specimens showed alternating orthokeratosis and parakeratosis | -100
skin biopsy specimens showed dermal lymphohistiocytic infiltrate with few neutrophils | -100
type II PRP was diagnosed | 0
intense erythroderma | -100
Staphylococcus aureus septicemia | -100
admitted to the intensive care unit | -100
severe depression | -100
anorexia | -100
loss of 30 kg | -100
previous treatments included topical corticosteroids | -100
previous treatments included acitretin | -100
previous treatments included photochemotherapy | -100
previous treatments included cyclosporine | -100
previous treatments included methotrexate | -100
previous treatments included infliximab | -100
previous treatments included ustekinumab | -100
previous treatments included intravenous immunoglobulin | -100
previous treatments included omalizumab | -100
prednisone was efficient | -100
relapse with less than 0.5 mg/kg/d | -100
cyclosporine was efficient | -100
association with 10 mg prednisone | -100
secukinumab was initiated | 0
informed consent | 0
secukinumab in association with cyclosporine and 10 mg of prednisone | 0
5 subcutaneous 300-mg weekly injections | 0
once-a-month injections | 28
significant and prompt clinical response | 28
quality-of-life improvement | 28
psoriasis area and severity index decreased | 28
dermatologic life quality index score decreased | 28
oral and esophageal candidiasis | 28
treated with fluconazole | 28
fluconazole for 14 days | 28
secukinumab was highly effective | 168
no recurrence of PRP lesions | 168
6-month follow-up | 168