42 years old | 0
female | 0
weight 48.8 kg | 0
height 159 cm | 0
admitted to the hospital | 0
Klatskin tumor | -672
Bismuth type IV | -672
tumor resection | -24
acute hepatic failure | -24
elevated liver function profile | -672
aspartate aminotransferase 170 U/L | -672
alanine aminotransferase 100 U/L | -672
hemoglobin 10.4 g/dl | -24
platelet count 103 × 10^3/µl | -24
prothrombin time (PT) 2.03 | -24
activated partial thrombin time (aPTT) 104.5 seconds | -24
fibrinogen 97 mg/dl | -24
fibrin degradation product >5 µg/ml | -24
D-dimer 3.23 µg/ml | -24
antithrombin III activity 41% | -24
plasminogen activity 30% | -24
protein C activity 43% | -24
metabolic acidosis | -24
pH <7.15 | -24
base deficit >15 mmol/L | -24
hypocalcemia <0.8 mmol/L | -24
hyperglycemia >200 mg/dl | -24
exsanguinating bleeding | -24
transfusion of packed red blood cells | -24
transfusion of fresh frozen plasma | -24
transfusion of platelet concentrates | -24
transfusion of cryoprecipitate | -24
infusion of dopamine | -24
infusion of norepinephrine | -24
total hepatectomy | 0
temporary portocaval shunt | 0
anhepatic state | 0
arterial blood gas analysis | 0
ionic calcium level | 0
dieresis | 0
metabolic acidosis alleviation | 0
pH 7.15-7.25 | 0
base deficit 10-15 mmol/L | 0
hyperchloremia | 0
potassium level 3.5-3.8 mmol/L | 0
magnesium level 1.6-1.7 mg/dl | 0
sodium level 144-146 mmol/L | 0
hypocalcemia <0.8 mmol/L | 0
infusion of calcium gluconate | 0
infusion of sodium bicarbonate | 0
infusion of magnesium | 0
infusion of 5% albumin | 0
infusion of 20% mannitol | 0
infusion of dextrose solution | 0
inotropic support | 0
systolic blood pressure 80-100 mmHg | 0
diastolic blood pressure 60-80 mmHg | 0
urine output <10 ml/hr | 0
elevated creatinine level 1.58 mg/dl | 0
coagulation profile | 0
prolongation of PT (INR) | 0
prolongation of aPTT | 0
fibrinogen <100 mg/dl | 0
living-donor liver transplantation | 15
anesthesia induction | 15
anesthesia maintenance | 15
desflurane | 15
oxygen fraction 0.5 | 15
electrocardiography | 15
SpO2 | 15
radial arterial pressure | 15
femoral arterial pressure | 15
pulmonary arterial pressure | 15
cardiac output | 15
vasoactive support | 15
dopamine | 15
norepinephrine | 15
hemodynamic profile | 15
stable | 15
crystalloid administration | 15
packed red blood cell administration | 15
fresh frozen plasma administration | 15
platelet apheresis | 15
cryoprecipitate administration | 15
postoperative care | 22
cardiovascular support | 22
respiratory support | 22
CCRT | 22
alert | 216
extubation | 384
reintubation | 408
pulmonary effusion | 408
respiratory failure | 408
acute renal insufficiency | 22
peritonitis | 22
bowel anastomosis leakage | 22
sepsis | 22
multiorgan failure | 22
death | 1560