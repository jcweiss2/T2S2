septuagenarian | 0
male | 0
admitted to the hospital | 0
malaise | -72
gait unsteadiness | -72
left arm weakness | -72
fever | -72
vomiting | -72
headache | -72
medication-controlled hypertension | -672
lethargic | 0
opening eyes to voice | 0
pupils were reactive | 0
extraocular movements were full | 0
corneal reflexes were intact | 0
computed tomography of the brain | 0
blood cultures | 0
no oculocephalic movements | 24
cranial nerve functions remained intact | 24
small pupils | 24
intact corneal reflexes | 24
ophthalmology consult was not performed | 24
severe lethargy | 48
left hemiplegia | 48
right gaze preference | 48
poor gag reflex | 48
intubated | 48
admitted to the Intensive Care Unit | 48
computed tomography of the brain | 48
linear band of low attenuation | 48
infarction in the lenticulostriate distribution | 48
analysis of cerebrospinal fluid | 48
moderate neutrophilic pleocytosis | 48
cultures of CSF and blood failed | 48
treated empirically with ceftriaxone | 48
treated empirically with ampicillin | 48
treated empirically with doxycycline | 48
treated empirically with acyclovir | 48
electroencephalography | 48
periodic lateralized epileptiform discharges | 48
empirically loaded with Dilantin | 48
progressive decline in level of consciousness | 72
progressive neurologic impairment | 72
loss of all brainstem reflexes | 72
left-sided pneumothorax | 72
gastrointestinal hemorrhage | 72
bilateral pulmonary edema | 72
recurrent fevers | 72
septic shock | 72
consultants from the Division of Infectious Disease | 72
viral meningoencephalitis | 72
West Nile virus | 72
EEE | 72
Western EE | 72
St. Louis encephalitis | 72
Cache Valley fever | 72
LaCrosse virus infection | 72
rabies | 72
magnetic resonance imaging of the brain | 48
diffuse signal enhancement | 48
meningoencephalitis | 48
CSF obtained | 48
negative India ink examination | 48
fungal culture was negative | 48
serological studies of blood and cerebrospinal fluid | 120
ELISA was positive for serum IgM antibodies to EEE virus | 120
ELISA was negative for serum IgG antibodies | 120
recent infection with EEE virus | 120
ELISA was not positive for IgM antibodies to EEE in the CSF | 120
IgM and IgG antibodies against St. Louis encephalitis virus and LaCrosse virus were not detected | 120
expired secondary to respiratory failure | 168
severe edema | 168
herniation of the cerebellar tonsils | 168
necrosis of the inferior temporal lobe | 168
petechial hemorrhages | 168
perivascular lymphohistiocytic cuffing | 168
meningeal involvement | 168
microglial nodules | 168
acute infarcts | 168
parenchymal edema | 168
hemorrhage | 168
hippocampus demonstrated several areas of microscopic infarction | 168
focal neuronal dropout | 168
cerebellum demonstrated multiple areas of myelin pallor | 168
Purkinje cell dropout | 168
Bergmann's type gliotic reaction | 168
ischemic compromise | 168
punctate hemorrhages | 168
no lesion of the spinal cord | 168
viral inclusions were not identified | 168
retinal hemorrhages | 168
patchy areas that appeared cloudier than usual | 168
decreased number of ganglion cells | 168
microcysts in the ganglion cell and nerve fiber layers | 168
simulating a retinoschisis | 168
T-lymphocytes | 168
macrophages expressing CD68 antigen | 168
coronary artery disease | 168
focally moderate stenosis of the right and left main coronary arteries | 168
acute bronchitis and bronchiolitis | 168
fibrin microthrombi in the kidneys and left adrenal gland | 168
terminal disseminated intravascular coagulation | 168
no generalized lymphohistiocytosis | 168