60 years old | 0
male | 0
Caucasian | 0
merchant ship captain | 0
admitted to the hospital | 0
headache | -24
dizziness | -24
disorientation | -24
ingestion of isopropanol | -24
ingestion of ethanol | -24
consumed most of the liquid in the bottle | -24
empty bottle of rubbing alcohol | -24
labelled as 70% volume per volume isopropyl alcohol | -24
capacity of 473 mL | -24
indication for use as a first aid antiseptic | -24
for rubbing and massaging | -24
disoriented | 0
clinical examination was unremarkable | 0
unenhanced computed tomography scan of the brain | 0
unremarkable | 0
symptomatic treatment was started | 0
collapsed in the hospital | 0.5
deeply comatose | 0.5
Glasgow Coma Scale score of 3/15 | 0.5
hypotension | 0.5
blood pressure of 80/40 mmHg | 0.5
pulse rate of 65 per minute | 0.5
respiratory rate of 8 per minute | 0.5
generalized hypotonia | 0.5
absent tendon reflexes | 0.5
no evidence of trauma to the head or cervical spine | 0.5
administration of intravenous fluids | 0.5
endotracheal intubation | 0.5
admitted to the intensive care department | 0.5
leukocytosis of 26,000 white blood cells per μL | 1
hemoglobin of 15.7 g/dL | 1
mean corpuscular volume of 93 fl | 1
arterial blood gas report | 1
pH of 6.731 | 1
pCO2 level of 28.2 mmHg | 1
pO2 level of 141 mmHg | 1
bicarbonate level of 3.5 mmol/L | 1
oxygen saturation of 95% | 1
blood urea nitrogen of 9.5 mmol/L | 1
serum creatinine of 157 μmol/L | 1
Na+ of 141 mmol/L | 1
K+ of 6 mmol/L | 1
Cl− of 107 mmol/L | 1
HCO3 of 5 mmol/L | 1
capillary blood glucose of 7.2 mmol/L | 1
severe metabolic acidosis | 1
acute renal failure | 1
blood lactic acid level of 8.7 mmol/mL | 1
blood ketones were negative | 1
blood investigations were negative for the presence of ethanol | 1
investigations repeated at 2-hour intervals | 2
increasing renal impairment | 2
hyperglycemia | 2
electrolyte imbalance | 2
low bicarbonate levels | 2
hyperkalemia | 2
follow-up arterial blood gas analysis | 2
severe acidosis | 2
no growth was detected on cultures of urine and blood | 2
no crystals were found in the urine on microscopic examination | 2
serum pseudocholinesterase level of 7,438 U/L | 2
calculated serum osmolarity of 310 mOsmol/L | 2
hemodialysis | 2
norepinephrine | 2
intravenous fluids | 2
fractionated plasma protein | 2
normal saline | 2
unenhanced MRI scans of the brain and spine | 144
bilaterally symmetrical hyperintensities | 144
cerebral and cerebellar cortex and white matter | 144
basal ganglia | 144
thalami | 144
brainstem | 144
swollen and edematous cervical spinal cord | 144
T2-weighted and FLAIR hyperintensities | 144
cerebellar tonsillar herniation | 144
petechial hemorrhages | 144
expired | 240
toxic brain and cervical spinal cord damage | 240