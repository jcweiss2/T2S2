27 years old | 0  
    male | 0  
    transferred to the Emergency Department of Pescara General Hospital | 0  
    car crash | 0  
    awake | 0  
    severe respiratory distress | 0  
    cyanosis | 0  
    hemodynamic instability | 0  
    right pneumothorax | 0  
    thoracic drainage inserted | 0  
    hemodynamic stabilization | 0  
    respiratory stabilization | 0  
    CT scan performed | 0  
    bilateral pneumothorax | 0  
    rib fractures | 0  
    multiple pulmonary contusions | 0  
    sacral wing fracture | 0  
    right tibial plateau fracture | 0  
    no traumatic brain injury | 0  
    ICU admission | 0  
    intubation | 0  
    mechanical ventilation | 0  
    left chest drainage inserted | 0  
    conscious sedation with dexmetomidine | 0  
    conscious sedation with Remifentanil | 0  
    RASS-2 | 0  
    pulmonary contusions managed with bronchial toilet | 0  
    systemic antimicrobial treatment with amikacin | 0  
    systemic antimicrobial treatment with cefazolin | 0  
    plate osteosynthesis for tibial plateau fractures | 0  
    septic episode | 96  
    blood cultures | 96  
    bronchoalveolar lavage | 96  
    empiric antimicrobials modified to piperacillin-tazobactam | 96  
    empiric antimicrobials modified to linezolid | 96  
    Gram-staining | 96  
    Fluorescence in situ hybridization (FISH) of blood culture isolates | 96  
    Pseudomonas spp | 96  
    Staphylococcus spp | 96  
    patient’s conditions unchanged | 168  
    cultural results yielded XDR Pseudomonas aeruginosa (XDR-PA) | 168  
    high-dose meropenem started | 168  
    high-dose colistin started | 168  
    nebulized colistin added | 168  
    XDR-PA isolate from broncho-alveolar lavage | 168  
    pulmonary source for sepsis postulated | 168  
    intense headache | 216  
    neck rigidity | 216  
    lumbar puncture performed | 216  
    cloudy cerebrospinal fluid | 216  
    neutrophils >500/microL | 216  
    glucose 19 mg/dL | 216  
    protein 279 mg/dL | 216  
    Gram-staining of growing colonies | 216  
    Gram-negative bacteria compatible with Pseudomonas spp | 216  
    breakthrough meningitis | 216  
    salvage regimen with high-dose C-T | 216  
    salvage regimen with high-dose Fosfomycin | 216  
    salvage regimen with Rifampicin | 216  
    Dexamethasone added | 216  
    head bone high-resolution CT-scans showed right middle-ear and mastoid suppurative infection | 216  
    no bone fractures | 216  
    meningeal syndrome resolved | 264  
    right mastoidectomy with tympanoplasty postponed | 264  
    extubated | 264  
    transferred to the Infectious Diseases Unit | 264  
    final microbiological characterization of CSF XDR-PA isolates | 264  
    ceftolozane-tazobactam MIC 3 mg/L | 264  
    colistin MIC <0.5 mg/L | 264  
    fosfomycin discontinued | 456  
    ceftolozane-tazobactam discontinued | 336  
    control head bone CT-scans confirmed complete resolution of otomastoiditis | 336  
    discharged | 336  
    no clinically relevant neurological sequelae | 336  
    history of chronic otitis media | -  
    recurring otitis | -  
    treated with quinolones | -  
    treated with cephalosporins | -  
    XDR-PA selection in right mastoid | -  
    severe polytrauma | -  
    multiple chest fractures | -  
    bloodstream infection | -  
    pneumonia | -  
    meningitis | 216  
    CNS escape of XDR-PA | 216  
    otomastoiditis | 216  
    pulmonary contusions | 0  
    sepsis | 168  
    bronchial toilet | 0  
    dexmetomidine sedation | 0  
    Remifentanil sedation | 0  
    amikacin treatment | 0  
    cefazolin treatment | 0  
    piperacillin-tazobactam treatment | 96  
    linezolid treatment | 96  
    meropenem treatment | 168  
    colistin treatment | 168  
    fosfomycin treatment | 216  
    Rifampicin treatment | 216  
    Dexamethasone treatment | 216  
    CSF sampling | 216  
    sterile CSF | 264  
    normalized CSF parameters | 264  
    otomastoiditis resolution | 336  
    Ethical Committee validation | 216  
    off-label prescription | 216  
    synergism between C-T and fosfomycin | 216  
    surgical management of otomastoiditis | 264  
    no competing interests | 336  
    no funding source | 336  
    acknowledgements | 336  
    ethical approval | 336  
    conflict of interest | 336  
    author statement | 336  
    funding source | 336  
