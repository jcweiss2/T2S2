74 years old | 0
female | 0
body mass index 29.3 | 0
chronic AF | 0
VATS-LA maze procedure | 0
sequential one lung ventilation | 0
EZ-Blocker endobronchial blocker | 0
transesophageal echocardiography | 0
bipolar radiofrequency catheter | 0
ablation lesions | 0
persistent fever | -504
altered mental status | -504
left upper extremity weakness | -504
computed tomography of the head | -504
magnetic resonance imaging/angiography of the head | -504
computed tomography of the thorax | -504
air in the posterior LA | -504
suspicion for LA wall abscess or AEF | -504
surgical exploration | -24
median sternotomy | -24
cardiopulmonary bypass | -24
intubation | -24
9F double-lumen central venous catheter | -24
18-G catheter | -24
blood pressure monitoring | -24
blood sampling | -24
esophagogastroduodenoscopy | -24
severe hypotension | -24
phenylephrine | -24
norepinephrine | -24
epinephrine | -24
TEE probe | -24
air in the LA, left ventricle, and aortic root | -24
emergent median sternotomy | -24
institution of CPB | -24
nasogastric tube | -24
aliquots of air | -24
fistula opening into the posterior wall of the LA | -24
patching with bovine pericardium | -24
transfer to surgical intensive care unit | 0
intubated and mechanically ventilated | 0
neurological deterioration | 24
MRI | 24
punctate and confluent hyperintensities | 24
global slowing on EEG | 48
withdrawal of care | 240
death | 240