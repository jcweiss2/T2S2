42-year-old | 0
    gravida 7 para 4 | 0
    presented at 32 weeks of gestation | 0
    reduced fetal movement | 0
    no history of trauma | 0
    mechanical mitral valve replacement | 0
    taking enoxaparin 80 mg twice daily | -672
    switched to warfarin 10 mg/day | -672
    INR of 4.7 | 0
    prothrombin time of 49 s | 0
    activated partial thromboplastin time of 44 s | 0
    fibrinogen 3.4 g/L | 0
    platelets 309,000/mL | 0
    hemoglobin 9 g/dL | 0
    instability of fetal heart rate | 0
    crescent hyperechoic collection suggestive of SDH | 0
    emergency cesarean section | 0
    warfarin stopped 36 h prior to surgery | -36
    born non-vigorous | 0
    no respiratory effort | 0
    pale | 0
    heart rate of 40 BPM | 0
    resuscitation without response | 0
    bagging for 30 s | 0
    heart rate increased to >100 BPM | 0
    no breathing | 0
    intubated at 1 min of age | 0.0167
    oxygen saturation 72–82% | 0.0167
    poor perfusion | 0.0167
    pale color | 0.0167
    umbilical venous catheter inserted | 0.0167
    bolus of normal saline administered | 0.0167
    blood transfusion | 0.0167
    Apgar score 2 at 1 min | 1
    Apgar score 5 at 5 min | 5
    Apgar score 6 at 10 min | 10
    Apgar score 8 at 15 min | 15
    surfactant given | 0.0167
    oxygen saturation improved | 0.0167
    fraction of inspired oxygen 21% | 0.0167
    transferred to NICU | 0.0167
    stable condition | 0.0167
    birthweight 2,010 g | 0
    length 43 cm | 0
    head circumference 31 cm | 0
    bulged anterior fontanelle | 0
    swelling in the right scrotum | 0
    pH 7.11 | 0
    PCO2 58 mm Hg | 0
    base excess −11.6 mmol/L | 0
    bicarbonate 18.4 mmol/L | 0
    hemoglobin 10.4 g/dL | 0
    platelets 119,000/mL | 0
    INR 3.7 | 0
    prothrombin time 38.8 s | 0
    activated partial thromboplastin time 71.9 s | 0
    received 5 mg vitamin K | 0
    higher vitamin K doses for babies with hemorrhage | 0
    brain ultrasound on day 1 | 24
    crescent hypoechoic collection in left frontoparietal region | 24
    echogenic focus in falx | 24
    no midline shift | 24
    no ventricular dilatation | 24
    testes ultrasound on day 1 | 24
    large turbid fluid collection in right scrotal sac | 24
    hemorrhagic fluid | 24
    normal testes appearance | 24
    normal testes perfusion | 24
    head CT on day 2 | 48
    bilateral SDH | 48
    subarachnoid hemorrhage | 48
    diffuse brain edema | 48
    midline shift 6 mm | 48
    brain ultrasound at 20 days | 480
    large subacute/chronic SDH | 480
    midline shift to right | 480
    cystic changes suggestive of severe PVL | 480
    cephalomalacia | 480
    dilated lateral ventricles | 480
    MRI at 24 days | 576
    bilateral acute on subacute SDH | 576
    extensive encephalomalacic changes | 576
    spared basal ganglionic region | 576
    spared frontotemporal area | 576
    spared posterior fossa | 576
    managed conservatively | 0
    no seizure activity | 0
    no hydrocephalus | 0
    right scrotal hemorrhage resolved | 336
    late onset sepsis | 336
    urine culture positive for Klebsiella pneumoniae | 336
    antibiotics for 2 weeks | 336
    discharged at 4 weeks | 672
    tube feeding | 672
    multidisciplinary team follow-up | 672
    spastic quadriplegic cerebral palsy | 87840
    gross motor function classification system level 5 | 87840
    kyphotic posture | 87840
    severe global delays | 87840
    no grasp | 87840
    blindness | 87840
    non-recognized speech | 87840
    