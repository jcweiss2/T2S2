78 years old | 0
male | 0
gastric cancer | 0
type II diabetes mellitus | 0
ischemic heart disease | 0
previous myocardial infarction | -8760
occasional ongoing angina | 0
benign prostatic hypertrophy | 0
open cholecystectomy | -0 (no specific time given, assuming at admission)
adhesions around the cholecystectomy site | 0
dense perisplenic capsular adhesions | 0
fatty liver | 0
bulky left lobe of the liver | 0
Nathanson retractor used | 0
retraction of the left lobe of the liver | 0
laparoscopic mobilization of the stomach and omentum | 0
division of the first part of the duodenum | 0
splenic capsular bleeding | 0
laparoscopic division of the splenic vessels | 0
splenectomy | 0
Roux-en-Y esophagojejunostomy | 0
feeding jejunostomy tube sited | 0
total laparoscopic time of the operation | 3.5
hypotensive | 0
inotropic support | 0
increasing inotropic support | 18
blood pressure stabilized | 24
serum AST levels elevated | 5
serum AST levels came down | 48
serum levels of alkaline phosphatase, gamma-glutamyltransferase, total bilirubin, and C-reactive protein elevated | 24
tachycardia | 48
fever | 48
temperature 38°C | 48
deterioration | 54
ventilatory assistance | 54
suspicion of anastomotic dehiscence | 54
urgent noncontrast abdominal computerized tomogram (CT) | 54
massive destruction in the left lobe of the liver | 54
large loculations of intraparenchymal gas | 54
gas in the portal radicals | 54
exploratory laparotomy | 60
left lobe of the liver necrotic and turgid | 60
left lateral sectionectomy (segments 2,3) | 60
postoperative inotropic support | 60
myocardial infarction | 74
death | 74