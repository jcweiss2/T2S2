74 years old | 0
female | 0
admitted to the emergency department | 0
dizziness | 0
emphysematous chronic obstructive pulmonary disease | -8760
smoking habit | -8760
severe chronic ischemic heart disease | -8760
hypercholesterolemia | -8760
hypoxemic respiratory failure | 0
SpO2 82% | 0
respiratory frequency 24/min | 0
oxygen therapy with a Venturi mask | 0
electrocardiogram negative for ischemia | 0
body temperature 37.6°C | 0
lymphopenia | 0
C-reactive protein increase | 0
centrilobular emphysema | 0
ground glass opacity (GGO) areas | 0
Coronavirus-19 positive | 0
hydroxychloroquine | 0
azithromycin | 0
deteriorated | 168
admitted to the intensive care unit | 168
admitted to the “Covid-19 Sub-ICU” | 168
noninvasive mechanical ventilation (NIMV) | 168
tocilizumab | 168
methylprednisolone | 168
enoxaparin | 168
respiratory failure improved | 216
regression of GGO | 480
arterial blood gasses improved | 480
discontinuation of NIMV | 480
high flow oxygen | 480
clinical conditions deteriorated | 504
increasing respiratory frequency | 504
worsening of hypoxemia | 504
gram-positive sepsis | 504
linezolid | 504
respiratory conditions worsened | 528
NIMV started again | 528
very severe hypoxemic respiratory failure | 1320
radiological progression of pulmonary fibrosis | 1320
death | 1440
severe hypoxemic respiratory failure | 1440