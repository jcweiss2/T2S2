86 years old | 0
    woman | 0
    presented to the emergency department | 0
    nausea | 0
    vomiting | 0
    right upper quadrant abdominal pain | 0
    coronary artery disease | -720
    pulmonary hypertension | -720
    mitral regurgitation | -720
    atrial fibrillation | -720
    chronic kidney disease | -720
    tachycardic | 0
    hypotensive | 0
    right upper quadrant tenderness | 0
    positive Murphy’s sign | 0
    elevated liver enzymes | 0
    alkaline phosphatase 387 U/L | 0
    alanine aminotransferase 89 U/L | 0
    aspartate aminotransferase 78 U/L | 0
    total bilirubin 5.9 mg/dL | 0
    direct fraction of 5.2 mg/dL | 0
    elevated creatinine | 0
    elevated white blood cell count | 0
    normal lipase | 0
    distended gallbladder | 0
    cholelithiasis | 0
    gallbladder wall thickness 3 mm | 0
    14-mm dilated common bile duct | 0
    thickened gallbladder walls | 0
    inflammatory changes within the adjacent fat | 0
    dilated common bile duct | 0
    admitted to the intensive care unit | 0
    sepsis | 0
    acute cholecystitis | 0
    choledocholithiasis | 0
    acute kidney injury | 0
    intravenous hydration | 0
    empiric antibiotics | 0
    endoscopic retrograde cholangiopancreatography | 24
    obstructed cystic duct | 24
    multiple CBD stones | 24
    stone removal after sphincterotomy | 24
    10F x 9 cm plastic stent placed in CBD | 24
    not considered a surgical candidate | 24
    underwent ultrasound-guided PC tube placement | 96
    clinical condition improved | 96
    discharged home | 96
    PC tube in place | 96
    multiple evaluations | 96
    PC tube exchanges | 96
    patent cystic duct | 96
    occluded biliary stent | 96
    some contrast reaching the duodenum | 96
    another ERCP | 2160
    removed biliary stent | 2160
    CBD stones extracted using cholangioscope | 2160
    electrohydraulic lithotripsy | 2160
    CBD completely cleared | 2160
    10F X 7 cm plastic stent placed | 2160
    at risk for recurrent choledocholithiasis | 2160
    hybrid percutaneous–endoscopic technique | 2160
    residual gallstones removed | 2160
    PC tube removed | 2160
    minimized future interventions | 2160
    under sedation and local anesthesia | 2160
    cholecystostomy drain opening dilated | 2160
    28F sheath placed | 2160
    pediatric gastroscope advanced | 2160
    gallbladder visualized | 2160
    multiple stones identified | 2160
    largest stone 14 mm | 2160
    lithotripsy successful | 2160
    gallstones removed | 2160
    Roth net used | 2160
    retrieval basket used | 2160
    20F drainage catheter placed | 2160
    another ERCP performed | 3600
    biliary stent occluded | 3600
    stent removed | 3600
    stone in middle third CBD swept out with 12-mm balloon | 3600
    no other stones remaining | 3600
    percutaneous cholangiogram | 4440
    contrast flow into duodenum | 4440
    no significant obstruction | 4440
    PC tube removed | 4440
    PC site healed | 4440
    no complications | 4440
    asymptomatic at 6-month follow-up | 4320
    asymptomatic at 1-year follow-up | 8760
    