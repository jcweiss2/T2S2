53 years old | 0
male | 0
hypertension | 0
type 2 diabetes mellitus | 0
alcohol abuse | 0
massive bout of alcohol intake | -96
liquid diarrhoea | -96
self-medication by non-steroidal anti-inflammatory drugs (NSAIDs) | -96
febrile respiratory distress | -96
diffuse cutaneous marbling | -96
emergency admission | 0
confused | 0
oligo-anuric | 0
purpuric lesions | 0
acute renal failure | 0
severe inflammation | 0
metabolic acidosis | 0
anaemia | 0
subnormal platelet count | 0
hyperleucocytosis | 0
increased lactate dehydrogenase | 0
free bilirubin | 0
haptoglobinaemia | 0
schizocytosis | 0
prothrombin time | 0
fibrinogen | 0
troponin | 0
pneumonia | 0
global left ventricle hypokinesia | 0
probabilist antibiotherapy | 0
haemodialysis | 0
pneumoccocal infection | 0
cutaneous necrotic lesions | 48
skin biopsy | 48
fibrin thrombi | 48
epidermolysis | 48
haemoglobinaemia | 48
thrombopenia | 48
schizocytes | 48
haptoglobin | 48
plasmatic exchanges | 96
plasma substitution | 96
renal function | 96
haemolysis parameters | 96
anuria | 96
severe thrombopenia | 96
schizocytosis | 96
skin lesions | 96
necrosis | 96
confusion | 96
obnubilation | 96
cardiac parameters | 96
troponin | 96
left ventricular function | 96
ECZ treatment | 120
mental confusion | 120
platelet count | 120
haptoglobin | 120
platelets | 144
diuresis | 240
renal function | 240
dialysis withdrawal | 336
renal function | 600
ECZ therapy | 720
skin lesions | 720
trans-tibial amputation | 2160
investigations | 0
ADAMTS13 activity | 0
monoclonal gammapathy | 0
human immunodeficiency virus (HIV) | 0
hepatitis C | 0
Parvovirus B19 | 0
cytomegalovirus | 0
stool culture | 0
shigatoxin genes | 0
direct Coombs’ test | 0
indirect Coombs’ test | 0
plasma levels of complement factors | 0
C3 | 0
C4 | 0
CH50 | 0
complement alternative pathway (CAP) regulators | 0
factor I (CFI) | 0
factor H (CFH) | 0
CD46 leucocyte expression | 0
plasmatic C5b9 | 0
anti-CFH antibodies | 0
genetic screening | 0
complement genes | 0
complement factor H (CFH) | 0
complement factor I (CFI) | 0
C3 | 0
factor B | 0
membrane cofactor protein (MCP or CD46) | 0
thrombomodulin (THBD) | 0
ECZ discontinuation | 4320
biological parameters | 8760
renal function | 8760
serum creatinine | 8760