41 years old | 0
female | 0
menorrhagia | -2520
dysmenorrhea | -2520
tranexamic acid | -2520
mefenamic acid | -2520
iron supplements | -2520
regular ultrasound pelvis | -2520
normal endometrial thickness | -2520
normal ovaries | -2520
stable adenomyoma | -2520
levonorgestrel-releasing intra uterine device (IUD) inserted | -720
levonorgestrel-releasing intra uterine device (IUD) expelled | -720
norethisterone | -720
palpitations | -720
total hysterectomy bilateral salpingectomy | 0
adenomyotic uterus | 0
normal tubes and ovaries | 0
estimated blood loss of 200 mL | 0
mild chronic endocervicitis | 0
leiomyoma | 0
adenomyosis | 0
recovery | 24
ambulating independently | 24
soft diet | 24
fever | 48
epigastric discomfort | 48
nausea | 48
diarrhoea | 48
CT of abdomen and pelvis | 72
fluid collection superior to the bladder | 72
intravenous clindamycin | 72
intravenous meropenem | 120
intra-abdominal drain inserted | 168
green-debris-laden fluid drained | 168
Candida on cultures | 168
investigations to screen for an immunocompromised state | 168
investigations to screen for bowel injury | 168
intravenous fluconazole | 168
symptoms resolved | 240
drain removed | 240
discharged home | 288
oral antibiotics | 288
oral fluconazole | 288
repeat scans | 672
marked reduction in collection | 672
HIV screen | 0
non-reactive HIV screen | 0
diabetes mellitus (DM) screen | 0
haemoglobin A1c (HbA1c) 4.9% | 0
blood culture | 0
no bacterial growth | 0
urine culture | 0
no bacterial growth | 0
stool culture | 0
no Salmonella | 0
no Shigella | 0
no Campylobacter | 0
no Vibrio species | 0
no Clostridium difficile | 0
stool microscopy | 0
no ova | 0
no cysts | 0
no trophozoites | 0
no parasites | 0
fluid culture | 168
Candida albicans | 168
Gram stain smear | 168
blastoconidia with pseudohyphae | 168 
vaginal swab | 192
negative vaginal swab | 192
recurrent inflammatory smears | -2520
vaginal candidiasis | -2520
PAP smears | -2520
lower genital swabs | -2520 
CT abdomen and pelvis | 72
CT abdomen and pelvis image | 672 
white cell count | 168
C reactive protein | 168 
intra-abdominal candidiasis | 168 
antifungal treatment | 168 
source control interventions | 168 
multidisciplinary team management | 168 
percutaneous catheter drainage | 168 
echinocandin | 168 
fluconazole | 168 
abscess formation | 168 
bloodstream invasion | 168 
sepsis | 168 
mortality | 0 
immunocompromised state | 0 
gastrointestinal tract injuries | 0 
vaginal infections | 0 
vaginal discharge | 0 
lower genital tract infection | 0 
screening test | 0 
surgery | 0 
intraoperative findings | 0 
specimen retrieval | 0 
transvaginal retrieval | 0 
ascending infection | 0 
intra-abdominal fluid | 168 
high clinical suspicion | 168 
intra-abdominal candidiasis (IAC) | 168 
gastrointestinal tract injuries | 72 
bowel injury | 72 
peritoneal dialysis | 0 
immunocompromised state | 0 
diabetes mellitus | 0 
multiple antibiotics | 0 
candidaemia | 0 
candida peritonitis | 0 
caesarean section | 0 
candida chorioamnionitis | 0 
vaginal swab | 192 
DNA probe test | 192 
sensitivity | 192 
specificity | 192 
inflammatory markers | 168 
white cell count | 168 
C reactive protein | 168 
antifungal therapy | 168 
echinocandin | 168 
fluconazole | 168 
abscess | 168 
peritonitis | 168 
sepsis | 168 
bloodstream invasion | 168 
mortality | 0 
intra-abdominal candidiasis | 0 
healthy woman | 0 
uncomplicated routine hysterectomy | 0 
risk factors | 0 
intra-abdominal candidiasis (IAC) | 168 
candida species | 0 
fungal peritonitis | 0 
candida albicans | 168 
intra-abdominal fluid | 168 
CT scan | 72 
collection | 72 
drainage | 168 
antifungal treatment | 168 
fluconazole | 168 
recovery | 240 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 0 
healthy woman | 0 
uncomplicated routine hysterectomy | 0 
risk factors | 0 
candida species | 0 
fungal peritonitis | 0 
candida albicans | 168 
intra-abdominal fluid | 168 
CT scan | 72 
collection | 72 
drainage | 168 
antifungal treatment | 168 
fluconazole | 168 
recovery | 240 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 672 
follow-up | 672 
CT scan | 672 
collection | 672 
reduction | 672 
intra-abdominal candidiasis | 168 
diagnosis | 168 
treatment | 168 
management | 168 
outcomes | 