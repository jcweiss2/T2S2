58 years old|0
woman|0
presented to the emergency department|0
altered mental status|0
difficulty breathing|0
intermittent weakness|-720
fever|-720
rash|-720
history of multiple tick exposures|-720
hypotensive|0
hypoxic|0
intubated|0
vasopressors initiated|0
creatinine of 203.32 μmol/L|0
albumin of 17 g/L|0
aspartate aminotransferase of 110 unit/L|0
white blood cell count of 3.4 × 109/L|0
hemoglobin level of 80 g/L|0
hematocrit level of 26%|0
platelet count of 36 × 109/L|0
admitted to the intensive care unit|0
lumbar puncture performed|0
urinalysis|0
urine culture|0
blood culture|0
blood test for tick-borne infections|0
septic shock|0
acute respiratory distress syndrome|0
vancomycin administered|0
cefepime administered|0
doxycycline added|0
chest x-ray showed bilateral diffuse infiltrates|0
hypoxia worsened|0
acute respiratory distress syndrome management protocol started|0
troponin level of 10 ng/mL|0
electrocardiogram (ECG) revealed no acute abnormality|0
transthoracic echocardiogram revealed no acute abnormality|0
left ventricular ejection fraction (LVEF) of 55% to 60%|0
left ventricular end-systolic volume index of 26 mL/m2|0
left ventricular end-diastolic volume index 67 mL/m2|0
normal wall motion|0
elevated troponin thought to be type 2 myocardial infarction|0
troponin I level increased to > 40 ng/mL|24
telemetry showed episodes of nonsustained ventricular tachycardia (NSVT)|24
repeat ECG revealed low-voltage QRS with ST-segment elevation|24
ST-segment elevation of 2 mm in leads I and AVL|24
Q waves in leads V1 and V2|24
taken emergently to the cardiac catheterization laboratory|24
coronary angiography showed normal coronary arteries|24
blood cultures negative for 5 days|-120
urine cultures negative for 5 days|-120
urinalysis elevated myoglobin levels|0
polymerase chain reaction (PCR) negative for herpes simplex virus|0
polymerase chain reaction (PCR) negative for cytomegalovirus|0
Ehrlichia chaffeensis PCR positive|0
hepatitis panel showed no immunity or prior exposure to hepatitis A, B, or C|0
Rocky Mountain Spotted Fever titers showed elevated immunoglobulin-G antibody (Ab)|0
anti-nuclear Ab negative|0
anti–double-stranded DNA negative|0
anti-smith negative|0
anti-ribonuclear protein negative|0
anti-Sjögren syndrome type A and B negative|0
rheumatoid factor negative|0
serum protein electrophoresis negative|0
cytoplasmic antineutrophil cytoplasmic Ab negative|0
perinuclear antineutrophil cytoplasmic Ab negative|0
vancomycin stopped|0
cefepime stopped|0
doxycycline continued|0
respiratory status improved|192
extubated|192
frequent premature ventricular contractions|192
multiple episodes of NSVT|192
high suspicion for myocarditis|192
cardiac magnetic resonance imaging revealed global hypokinesis|192
LVEF of 32%|192
left ventricular mass of 45 g/m2|192
delayed enhancement in myocardium and pericardium|192
myopericarditis|192
carvedilol administered|192
lisinopril administered|192
discharged to inpatient rehabilitation|384
cardiomyopathy persisted|2400
repeat transthoracic echocardiogram revealed LVEF of 25%|2400
repeat ECG revealed improvement in QRS voltages|2400
intermittent episodes of NSVT|2400
amiodarone administered|2400
cardioverter-defibrillator implanted|2400
two admissions for acute heart failure exacerbation|8760
human monocytic ehrlichiosis|0
acute febrile tick-borne illness caused by E. chaffeensis|0
vector ticks found in Southeastern to South Central United States|0
cardiac complications rarely reported with ehrlichiosis|0
ehrlichiosis-induced myocarditis|0
cardiac enzyme elevation|0
new cardiomyopathy|0
dysregulated inflammatory response|0
early doxycycline therapy|0
favorable outcome|0
survived|0
