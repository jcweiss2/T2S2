69 years old | 0
male | 0
admitted to the emergency department | 0
abdominal pain | -168
nausea | -168
vomiting | -168
fever | -24
mental status change | -24
chronic renal disease | 0
primary hypertension |* 0
diabetes mellitus | 0
history of coronary bypass surgery | 0
elevated fever (37.6°C) | 0
tachycardia (110 beats per minute) | 0
normal blood pressure (105/65 mmHg) | 0
Glasgow coma scale score 11 | 0
tenderness in all four quadrants | 0
right lower quadrant tenderness | 0
abdominal distension | 0
no signs of acute abdomen | 0
obstipation | -72
decreased bowel sounds | 0
empty rectum | 0
leukocytosis (12.9 103/uL) | 0
increased serum C-reactive protein (27.1 mg/dL) | 0
increased procalcitonin (11.5 ng/mL) | 0
increased creatinine (5.3 mg/dL) | 0
increased glucose (388 mg/dL) | 0
increased lactate (2.3 mmol/L) | 0
abdominal ultrasound minimal free fluid | 0
abdominal tomography 13 × 7 cm fluid collection | 0
diffuse free air within fluid collection | 0
extension to bilateral pararenal fascia | 0
extension to perirenal space | 0
interpreted as duodenal perforation | 0
retroperitoneal abscess | 0
received prophylactic broad-spectrum antibiotics | 0
underwent emergency surgery | 0
retrocecally appendicitis | 0
perforated appendicitis | 0
purulent contents spreading to retroperitoneal area | 0
appendectomy | 0
drained abscess | 0
inserted multiple drains | 0
no perforation in upper gastrointestinal tract | 0
abscess cultures negative | 0
followed in intensive care unit for 4 days | 0
septicemia | 0
septicemia subsided | 0
discharged on 15th postoperative day | 360
painful swelling in left scrotum | 720
fluctuation in left scrotum | 720
purulent discharge from left scrotum | 720
no signs of peritonitis | 720
fistula orifice in left scrotum | 720
purulent discharge | 720
abdominal tomography 17 × 7 cm abscess cavity | 720
normal leukocyte (7.09 103/uL) | 720
increased C-reactive protein (7.27 mg/dL) | 720
increased procalcitonin (0.58 ng/mL) | 720
increased lactate (2.7 mmol/L) | 720
percutaneous drainage | 720
broad-spectrum antibiotics | 720
abscess culture negative | 720
control tomography abscess regressed | 720
drainage from fistula orifice | 720
discharged after 17 days | 1128
