47 years old | 0
female | 0
diabetes mellitus | -7920
nausea | -48
vomiting | -48
decreased oral intake | -48
back pain | -48
headache | -24
levothyroxine | -336
subcutaneous long-acting insulin | -336
topiramate | -336
canagliflozin | -336
post-thyroidectomy Graves’ disease | -6336
cholecystectomy | -6336
depression | -6336
fibromyalgia | -6336
hyperlipidemia | -6336
spinal fusion surgery | -6336
volume depleted | 0
dry mucosal membranes | 0
absence of axillary sweat | 0
mild epigastric tenderness | 0
glucose 152 mg/dL | 0
sodium 138 mEq/L | 0
potassium 4.4 mEq/L | 0
chloride 105 mEq/L | 0
total carbon dioxide 16 mEq/L | 0
anion gap 17 | 0
serum blood urea nitrogen 16 mg/dL | 0
creatinine 0.76 mg/dL | 0
mixed acid-base disorder | 0
primary respiratory acidosis | 0
pH 7.18 | 0
PCO2 47.6 mmHg | 0
bicarbonate 17 mEq/L | 0
urinalysis pH 5 | 0
2+ ketones | 0
3+ glucose | 0
thyroid function tests unremarkable | 0
liver function tests unremarkable | 0
serum lactic acid 1 mEq/L | 0
withholding insulin | 0
discontinuing canagliflozin | 0
intravenous volume expansion | 0
cultures unremarkable | 12
spine MRI unremarkable | 12
lumbar puncture unremarkable | 12
nausea partially responded to ondansetron | 12
vomiting partially responded to ondansetron | 12
serum glucose <200 mg/dL | 12
insulin not administered | 12
serum bicarbonate 10 mEq/L | 12
transferred to medical intensive care unit | 12
repeat arterial blood gas | 12
pH 7.05 | 12
PCO2 26.9 mmHg | 12
bicarbonate 7 mEq/L | 12
total serum carbon dioxide 5 mEq/L | 12
isotonic bicarbonate started | 12
ingested soft diet | 24
blood glucose increased | 24
renal and endocrine consultants diagnosis of atypical diabetic ketoacidosis | 24
IV infusion of regular insulin | 24
serum bicarbonate normalized | 36
anion gap normalized | 36
regular diet resumed | 48
C-peptide level undetectable | 48
discharged | 72