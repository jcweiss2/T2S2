56 years old | 0
    female | 0
    referred to surgical unit with left-sided liver mass | 0
    denied previous history of chronic hepatitis | 0
    denied alcohol abuse | 0
    denied blood transfusion | 0
    transabdominal subtotal hysterectomy | prior to 2014
    unilateral oophorectomy | prior to 2014
    uterine leiomyoma | prior to 2014
    benign ovarian cyst | prior to 2014
    normal physical examination | 0
    normal routine laboratory tests | 0
    serum alpha-fetoprotein level 3.2 ng/mL | 0
    CA19-9 level 488.43 U/mL | 0
    contrast-enhanced abdominal ultrasonography revealed multiple liver tumors | 0
    maximum tumor dimensions 12.1 cm ×7.1 cm | 0
    magnetic resonance cholangiopancreatography performed | 0
    diagnosis of left-sided liver cancer | 0
    Child-Pugh class A | 0
    laparotomic left-sided hepatectomy | 0
    hilar lymphadenectomy | 0
    cholecystectomy | 0
    moderately differentiated ICC | 0
    chronic cholecystitis | 0
    uneventful postoperative course | 0
    follow-up ultrasonography on eighth postoperative week | 168
    three recurrent tumors in right lobe | 168
    sizes 1.5 cm ×1.3 cm, 1.2 cm ×1.0 cm, 0.9 cm ×1.0 cm | 168
    liver function remains Child-Pugh class A | 168
    serum alpha-fetoprotein 2.9 ng/mL | 168
    Doppler ultrasound-guided RFA performed | 168
    three sessions of RFA at 78 W for 16 minutes | 168
    follow-up ultrasound post-RFA day 3 | 192
    filling defect in ablated area | 192
    residual mass 1.0 cm ×0.8 cm in segment VIII | 192
    no significant liver/coagulation abnormalities | 192
    second RFA performed | 192
    initial power 50 W for 7 minutes | 192
    febrile (39.2°C) on second day after second RFA | 216
    hemoglobin 80 g/L | 216
    white cell count 10.4×109/L | 216
    alanine transferase 5,304 IU/L | 216
    aspartate transferase 7,906 IU/L | 216
    albumin 30.7 g/L | 216
    total bilirubin 38.9 μmol/L | 216
    prothrombin time 22.4 seconds | 216
    international normalized ratio 1.91 | 216
    emergency MRI showed extensive liver necrosis | 216
    diagnosis of RFA-associated ALF | 216
    prophylactic antimicrobial therapy | 216
    blood transfusion | 216
    nutritional liver support | 216
    lactose enemas | 216
    intravenous aspartic acid, ornithine, arginine | 216
    hyperammonemia (102 μmol/L) | 216
    respiratory distress | 216
    agitated | 216
    confused | 216
    increased heart rate | 216
    deteriorating pulse oxygen saturation | 216
    arterial blood gas PO2 71 mmHg | 216
    PCO2 50 mmHg | 216
    pH 7.32 | 216
    chest X-ray bilateral pulmonary inflammation | 216
    pleural effusion | 216
    contrast echocardiogram diagnosed HPS | 216
    diagnosis of HPS | 216
    ALF | 216
    ARF | 216
    excluded acute respiratory distress syndrome | 216
    excluded systemic inflammatory response syndrome | 216
    transnasal intubation | 216
    transferred to respiratory care unit | 216
    mechanical ventilation | 216
    tracheostomy | 216
    repeated chest X-ray showing improving pulmonary sepsis | 216
    improving pleural effusion | 216
    weaned from ventilator after 2 weeks | 360
    liver function improvement from fifth week | 840
    discharged at eleventh week after RFA | 1848
    followed up at outpatient clinic | 1848
    survived free of recurrence at 1 year | 8760
    <|eot_id|>