injury to the cervical esophagus during spinal surgery | -168
emergency esophageal diversion | -168
gastric pull-up procedure | -132
postoperative anastomotic leakage | -132
endoscopy and esophageal stent placement | -132
discharge with fully covered esophageal stent | -115
local cervical infection and sepsis | -99
transfer to tertiary university hospital | -99
admission | 0
clear signs of malnutrition and systemic inflammation | 0
jugular and cervical phlegmon | 0
hemoglobin level of 6.7 g/dL | 0
white blood cell count of 6400 cells/μL | 0
platelet count of 210 × 10^3/μL | 0
creatinine level of 0.76 mg/dL | 0
unremarkable liver and cholestasis parameters | 0
albumin level of 2.8 g/dL | 0
chest computed tomography scan | 0
endoscopy | 0
dislodged esophageal stent | 0
esophageal perforation 2 cm distal to the pharynx | 0
infected cavity | 0
5 cm-long stenosis of the esophagus | 0
stent removal | 0
endoscopic vacuum therapy | 12
EsoSponge system placement | 12
jugular and cervical phlegmon resolution | 24
repeated endoscopic balloon dilatation | 24
subtotal esophageal resection and reconstruction | 168
free-jejunal graft interposition | 168
CT angiography | 168
partial sternotomy | 168
laparotomy | 168
jejunal segment harvest | 168
graft implantation | 168
cervical anastomosis | 168
upper mediastinal gastro-jejunostomy | 168
sternocleidomastoid muscle flap | 168
abdominal reconstruction | 168
end-to-end jejunojejunostomy | 168
postoperative course uneventful | 192
oral alimentation reestablished | 192
daily speech therapy | 192
anastomotic healing confirmed | 216
transfer to rehabilitation clinic | 216
discharge in good clinical condition | 240