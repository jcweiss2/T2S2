42 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
granular dystrophy | 0 | 0 | Factual
DALK | 0 | 0 | Factual
big bubble technique | 0 | 0 | Factual
8 mm recipient stromal flap | 0 | 0 | Factual
air injected into stroma | 0 | 0 | Factual
donor button cut 8.25 mm | 0 | 0 | Factual
DM peeled off | 0 | 0 | Factual
donor button sutured | 0 | 0 | Factual
age of donor cornea 36 years | 0 | 0 | Factual
in situ cornea excision | 0 | 0 | Factual
surgery went well | 0 | 0 | Factual
whitish infiltrates | 24 | 24 | Factual
severe anterior chamber reaction | 24 | 24 | Factual
postoperative keratitis | 24 | 24 | Factual
graft removed | 24 | 24 | Factual
graft replaced | 24 | 24 | Factual
corneal scrapings sent for microbiology | 24 | 24 | Factual
host DM clear and intact | 24 | 24 | Factual
topical vancomycin started | 27 | 0 | Factual
topical ceftazidime started | 27 | 0 | Factual
Gram-stain showed Gram-negative Bacilli | 48 | 48 | Factual
infiltrates along entire graft host junction | 48 | 48 | Factual
hypopyon | 48 | 48 | Factual
topical antibiotics increased | 48 | 48 | Factual
corneal scrapings report | 72 | 72 | Factual
Klebsiella pneumoniae | 72 | 72 | Factual
resistant to multiple antibiotics | 72 | 72 | Factual
sensitive to imipenem | 72 | 72 | Factual
imipenem drops started | 72 | 0 | Factual
infiltration extended | 96 | 96 | Factual
hypopyon persisted | 96 | 96 | Factual
therapeutic penetrating keratoplasty | 120 | 120 | Factual
infiltrates in host DM | 120 | 120 | Factual
graft clear | 144 | 144 | Factual
no infiltrates or hypopyon | 144 | 144 | Factual
gatifloxacin drops added | 144 | 0 | Factual
prednisolone drops added | 168 | 0 | Factual
unaided vision 6/60 | 432 | 432 | Factual
vision improved to 6/18 with pin hole | 432 | 432 | Factual
graft clear | 432 | 432 | Factual
anterior segment quiet | 432 | 432 | Factual
intraocular pressure normal | 432 | 432 | Factual
pathogen eradicated | 432 | 432 | Factual