44 years old | 0
female | 0
South East Asian | 0
admitted to the Otolaryngology outpatient clinic | 0
hoarseness | -1314
loss of voice | -1314
reduction in effort tolerance | -1314
short of breath | -1314
unintentional weight loss | -1314
loss of appetite | -1314
laryngeal irritation | -1314
globus sensation in the throat | -1314
recurrent non-productive cough | -1314
choking and coughing on swallowing liquids | -1314
denies dysphagia | -1314
denies odynophagia | -1314
no significant past medical history | 0
no significant past surgical history | 0
breathing difficulties | -672
noisy breathing | -672
admitted to a district hospital | -672
treated for bronchial asthma | -672
readmitted to the district hospital | -504
nursed in the intensive care unit | -504
otolaryngology consult | -504
referred to UKM Medical Centre | -504
apyrexial | 0
haemodynamically stable | 0
audible biphasic stridor at rest | 0
able to count up to 10 in a single breath | 0
no respiratory distress | 0
cardiopulmonary assessment unremarkable | 0
bulky right false cord | 0
limited mobility of the right vocal cord | 0
severe bilateral subcordal edema | 0
narrowing the airway | 0
nasal and oral cavities normal | 0
abnormal Voice Handicap Index-10 score | 0
abnormal Eating Assessment Tool-10 score | 0
microcytic hypochromic anaemia | 0
haemoglobin of 9.0 g/dl | 0
immunological screening negative | 0
unremarkable chest x-ray findings | 0
thickening of the right false cord | 0
thickening of the true cord | 0
thickening of the aryepiglottic fold | 0
edema of the subglottis | 0
endolaryngeal microsurgery | 0
firm mass arising from the right ventricle | 0
mass extending into the right paraglottic space | 0
right subcordal mass ablated | 0
dilated up to 30 French Bougie | 0
worsening inspiratory stridor | 6
tachypnoea | 6
emergency tracheostomy | 6
sheets of small to medium-sized neoplastic cells | 6
neoplastic cells infiltrating the muscle fibres | 6
round to oval nuclei | 6
finely-dispersed chromatin | 6
inconspicuous nucleoli | 6
scanty cytoplasm | 6
immunoreactive for LCA | 6
immunoreactive for MPO | 6
immunoreactive for CD117 | 6
negative for CKAE1/AE3 | 6
negative for CD20 | 6
negative for Cd79a | 6
negative for CD3 | 6
negative for CD34 | 6
negative for TdT | 6
investigated for myeloproliferative disease | 6
bone marrow biopsy and trephine confirmed primary AML | 6
received chemotherapy with HiDAC protocol | 6
mass on the right false cord not visualised | 168
bilateral severe subcordal edema not visualised | 168
developed neutropenic sepsis | 168
developed invasive pulmonary aspergilosis | 168
repeat bone marrow biopsy showed refractory AML | 168
passed away | 720