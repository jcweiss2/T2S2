83 years old | 0
    male | 0
    type 2 diabetes | 0
    hypertension | 0
    atrial fibrillation | 0
    myocardial infarction | 0
    rectum carcinoma | -48
    low anterior resection | -48
    gas leakage at resection site | -48
    fecal leakage at resection site | -48
    perforations in colon transversus | -48
    sacral abscess | -48
    aspiration during intubation | 0
    ICU admission | 0
    sedation | 0
    hemodynamically stable | 0
    respiratory stable | 0
    baseline sublingual microcirculatory measurement | 0
    deterioration | 24
    shock | 24
    cardiopulmonary resuscitation | 24
    cardiac arrest | 24
    hypoxia | 24
    atelectasis of right lung | 24
    administration of nor-adrenaline | 24
    administration of adrenaline | 24
    vasoactive-inotropic score 99 | 24
    rising serum lactate up to 9.2 mmol/L | 24
    declining renal function | 24
    urine output 17 mL/24 h | 24
    sepsis diagnosis | 24
    CRRT with CytoSorb hemoadsorber | 24
    microcirculatory measurement at 24 h | 24
    microcirculatory measurement at 36 h | 36
    microcirculatory measurement at 48 h | 48
    microcirculatory measurement at 120 h | 120
    hemoadsorber replacement every 24 h | 24
    decreased lactate levels to 2.2 mmol/L | 24
    decreased VIS by 43% | 24
    76% decrease in lactate levels | 48
    VIS decreased by 87% | 48
    reduced TVD | 0
    reduced perfused vessel density | 0
    reduced microcirculatory flow index | 0
    heterogeneous plugged capillaries | 0
    high lactate levels | 0
    improved microcirculatory parameters within 12 h of CytoSorb | 12
    normalized microcirculatory flow index | 12
    increased TVD | 12
    reduced lactate levels | 12
    brisk flow at 36 h | 36
    no plugged vessels | 36
    improved clinical condition | 36
    fluid ultrafiltration initiated at 48 h | 48
    restoration of fluid balance | 48
    aggressive fluid resuscitation | 24
    progressive decline in TVD | 24
    blood transfusion | 48
    increased TVD during de-escalation | 120
    stable condition | 120
    regained consciousness | 120
    return to surgery ward on day 19 | 456
    total hospital stay 59 days | 1416
    discharge to nursing facility | 1416
    normalized renal function | 1416
    