41 years old | 0
female | 0
history of untreated hypertension | -672
history of morbid obesity | -672
history of chronic back pain | -672
history of IVDU | -672
low back pain | -336
diffuse abdominal pain | -336
lower extremity weakness | -336
anorexia | -336
fever | -336
chills | -336
shortness of breath | -336
dizziness | -336
constipation | -336
recent use of acetaminophen | -336
recent use of gabapentin | -336
recent use of hydrocodone | -336
recent use of methamphetamines | -336
recent use of marijuana | -336
admitted to the hospital | 0
blood pressure of 79/53 mmHg | 0
heart rate of 149 bpm | 0
lactic acid of 4.2 mg dl-1 | 0
white blood cell count (WBC) 37 500 u l-1 | 0
erythrocyte sedimentation rate 75 mm h-1 | 0
urine toxicology was positive for cannabis | 0
urine toxicology was positive for amphetamines | 0
midline tenderness of the lumbar spine | 0
3/5 strength in bilateral lower extremities | 0
bilateral shoulder warmth | 0
bilateral shoulder erythema | 0
bilateral shoulder tenderness | 0
limited range of motion | 0
multiple needle puncture sites on the antecubital fossas | 0
puncture wounds on the right foot | 0
blood cultures were collected | 0
started on vancomycin | 0
started on metronidazole | 0
started on aztreonam | 0
started on IV fluids | 0
MRSA bacteraemia | 0
sensitivities to vancomycin | 0
sensitivities to rifampin | 0
sensitivities to levofloxacin | 0
sensitivities to clindamycin | 0
sensitivities to daptomycin | 0
sensitivities to linezolid | 0
bilateral shoulder plain radiographs | 0
arthrocentesis of the acromioclavicular (AC) joints | 0
WBC of 93 137 u l-1 in one shoulder | 0
WBC of 32 043 u l-1 in the other shoulder | 0
aspirates were cultured | 0
grew MRSA | 0
emergent surgical debridement of the shoulders | 24
intubated | 24
MRI of the lumbar spine | 24
L3-L5 osteomyelitis | 24
facet septic arthritis | 24
dorsal paraspinous myositis | 24
L2-L5 epidural abscess | 24
bilateral psoas myositis | 24
bilateral psoas abscesses | 24
MRI of the bilateral shoulders | 48
septic arthritis of the AC joints | 48
right distal trapezius abscess | 48
left supraclavicular abscess | 48
MRI of the brain | 48
no acute intracranial processes | 48
transthoracic echocardiogram (TTE) | 48
no valvular vegetations | 48
cardiology deferred acquiring a transoesophageal echocardiogram | 48
repeat surgical debridement of the shoulders | 72
neurosurgery evaluated the patient | 72
leukocytosis continued to rise | 72
peaked at 52 100 u l-1 | 96
trough levels of vancomycin were being monitored | 96
repeat blood cultures continued to be positive for MRSA | 96
antibiotics were escalated to daptomycin | 240
antibiotics were escalated to ceftaroline | 240
blood cultures became negative | 336
rifampin was added | 336
infectious disease physician | 336
management of the patient’s concurrent osteomyelitis | 336
management of the patient’s concurrent facet septic arthritis | 336
management of the patient’s concurrent bilateral psoas abscesses | 336
management of the patient’s concurrent left supraclavicular abscess | 336
management of the patient’s concurrent right distal trapezius abscess | 336
required critical care | 336
extubation | 336
repeat MRI of the lumbar spine | 432
worsening epidural abscess | 432
neurosurgery took the patient for surgical drainage | 432
drain placement | 432
intraoperative wound cultures were positive for MRSA | 432
intraoperative wound cultures were positive for Proteus mirabilis | 432
improved clinically | 504
all drains were removed | 504
discharged | 504
prescribed oral levofloxacin | 504
prescribed oral rifampin | 504
lost to follow-up | 504