61 years old | 0
    male | 0
    undifferentiated schizophrenia | 0
    admitted to the intensive care unit | 0
    syncopal episode | 0
    agitation | -840
    aggressive behavior | -840
    hypothyroidism | -336
    levothyroxine | -336
    free thyroid-stimulating hormone of 1.20 | -336
    seizure disorder | -840
    divalproex sodium extended release 1000 mg daily | -840
    levetiracetam 750 mg twice daily | -840
    clozapine treatment started | -840
    clozapine 150 mg every morning | -840
    clozapine 150 mg every evening | -840
    clozapine evening dose increased to 175 mg | -120
    glaucoma | -840
    dorzolamide/timolol eye drops | -840
    regular diet | -840
    encouraged to take plenty of fluids and fibers | -840
    walk around the nursing station | 0
    syncopal episode | 0
    temperature 98°F | 0
    blood pressure 86/54 mmHg | 0
    pulse 127 beats/min | 0
    respiratory rate 16 breaths/min | 0
    oxygen saturation 100% | 0
    intravenous access obtained | 0
    normal saline 500 mL bolus administered | 0
    responsive within few minutes | 0
    tried to get up | 0
    moving all limbs | 0
    no focal motor deficits | 0
    no seizure activity | 0
    confused | 0
    agitated | 0
    unable to provide history | 0
    transferred to intensive care unit | 0
    abdominal distension | 0
    hypoactive bowel sounds | 0
    rectal examination revealed hard impacted stool | 0
    stool guaiac test negative | 0
    leukocyte count 17300/mm3 | 0
    neutrophil differential 52% | 0
    absolute neutrophil count 9000/mm3 | 0
    band neutrophils 12% | 0
    leukocyte count 7100/mm3 (Week 1) | -168
    neutrophil differential 45% (Week 1) | -168
    absolute neutrophil count 3195/mm3 (Week 1) | -168
    leukocyte count 6600/mm3 (Week 2) | -336
    neutrophil differential 61% (Week 2) | -336
    absolute neutrophil count 4026/mm3 (Week 2) | -336
    leukocyte count 5400/mm3 (Week 3) | -504
    neutrophil differential 65% (Week 3) | -504
    absolute neutrophil count 3510/mm3 (Week 3) | -504
    leukocyte count 5200/mm3 (Week 4) | -672
    neutrophil differential 60% (Week 4) | -672
    absolute neutrophil count 3120/mm3 (Week 4) | -672
    leukocyte count 6500/mm3 (Week 5) | -840
    neutrophil differential 67% (Week 5) | -840
    absolute neutrophil count 4355/mm3 (Week 5) | -840
    hemoglobin 18.6 g/dL | 0
    elevated BUN/creatinine 34/1.4 | 0
    low serum bicarbonate 18 mmol/L | 0
    low serum chloride 100 mmol/L | 0
    elevated anion gap 17 | 0
    serum lactic acid elevated 115.4 mg/dL | 0
    serum valproic level 60 µg/mL | 0
    sinus tachycardia | 0
    no acute ST-T segment changes | 0
    serum troponin I normal | 0
    urine specific gravity high | 0
    no bacteria in urine | 0
    no elevated nitrate in urine | 0
    urine toxicology negative | 0
    chest X-ray elevated hemidiaphragm | 0
    chest X-ray low lung volumes | 0
    chest X-ray clear lung fields | 0
    abdominal X-ray fecal content in colon | 0
    abdominal X-ray dilated small bowel | 0
    started on broad spectrum antibiotics | 0
    intravenous fluids administered | 0
    worsening hypotension | 0
    surgical evaluation requested | 0
    deemed too unstable for surgery | 0
    managed per surviving sepsis guidelines | 0
    cardiac arrest | 12
    expired | 12
    blood culture Escherichia coli | 24
    urine culture no growth | 24
    no history of constipation | 0
    no fecal impaction | 0
    minimally communicative | 0
    mumbling incoherent words | 0
    disorganized | 0
    aggressive at times | 0
    intra-abdominal sepsis | 0
    bowel obstruction | 0
    fecal impaction | 0
    hypotension | 0
    sepsis | 0
    septic shock | 0

<|eot_id|>