80 years old | 0
male | 0
admitted to the hospital | 0
urinary tract infection | -120
fever | -120
dysuria | -120
cephalexin | -120
urine analysis | -120
large leukocyte esterase | -120
bacteria | -120
Escherichia coli | -120
resistance to ampicillin | -120
resistance to levofloxacin | -120
resistance to trimethoprim | -120
resistance to sulfamethoxazole | -120
intermediate sensitivity to ampicillin/sulbactam | -120
sensitivity to cefazolin | -120
sensitivity to gentamicin | -120
sensitivity to nitrofurantoin | -120
cephalexin 500 mg three times daily | -48
erythematous rash | -48
sloughing of the skin | -48
discontinued cephalexin | -24
transferred to a local burn intensive care unit | -24
chronic obstructive pulmonary disease | 0
type 2 diabetes mellitus | 0
coronary artery disease | 0
hypertension | 0
hypothyroidism | 0
depression | 0
end-stage renal disease | 0
hemodialysis | 0
multiple myocardial infarctions | 0
ischemic cardiomyopathy | 0
atrial fibrillation | 0
hydrocodone/acetaminophen | 0
levothyroxine | 0
escitalopram | 0
carvedilol | 0
guaifenesin | 0
docusate | 0
calcitriol | 0
albuterol | 0
amiodarone | 0
pulmonary infiltrates | 24
respiratory failure | 24
intubated | 24
difficulty swallowing | 24
endotracheal tube | 24
toxic epidermal necrolysis syndrome | 24
56% of the total body surface area | 24
skin detachment | 24
blood pressure 81/45 mm Hg | 24
respiratory rate 12 breaths/min | 24
temperature 36.8 °C | 24
white blood cell count 1.5 × 103/mm3 | 24
neutrophils 73% | 24
platelet count 77,000/µL | 24
serum creatinine 2.12 mg/dL | 24
venous serum lactate 3.1 mmol/L | 24
oxygen saturation 99% | 24
norepinephrine | 24
vasopressin | 24
albumin 25% | 24
lactated Ringer’s | 24
tetanus–diphtheria toxoids vaccine | 24
gentamicin 120 mg | 24
fluconazole 100 mg | 24
WBC 5.4 × 103/mm3 | 48
SCr 1.98 mg/dL | 48
venous serum lactate 1.8 mmol/L | 48
random serum gentamicin level 2.4 mg/dL | 48
gentamicin 120 mg | 48
fluconazole 200 mg | 48
Candida species | 48
Gram-negative rods | 48
Gram-positive rods | 48
wide complex tachycardia | 96
amiodarone | 96
gentamicin held | 96
random serum gentamicin level 2.2 mg/dL | 96
gentamicin 120 mg | 96
Pseudomonas aeruginosa | 96
expired | 144