81 years old | 0
male | 0
hypertension | 0
hyperlipidemia | 0
remote smoking | 0
chronic obstructive pulmonary disease (COPD) | 0
peptic ulcer disease (PUD) | 0
maroon stools | -72
bright red blood per rectum | -72
lightheadedness | -72
daily intake of baby aspirin | -672
previous melena episode | -1344
no recent melena | 0
no abdominal pain | 0
no nausea | 0
no vomiting | 0
no fevers | 0
no chills | 0
orthostatic | 0
unsuccessfully managed with intravenous (IV) fluids | 0
emergency colonoscopy | 0
3 colonic polyps removed | 0
diverticuli | 0
re-hospitalized for COPD | 720
massive painless hematochezia episode | 720
received IV steroids | 720
hypovolemic shock | 720
intubation | 720
ICU care | 720
extubation | 720
another massive painless hematochezia episode | 720
initial bleeding scan negative | 720
large transfusion requirement | 720
stabilized | 720
another episode of massive hematochezia | 720
2nd bleeding scan positive | 720
splenic flexure | 720
sigmoid colon | 720
increased uptake in the distal abdominal aorta | 720
right common iliac | 720
angiography did not reveal a specific bleeding site | 720
active hematochezia | 720
hypotension | 720
9 units of blood | 720
differential diagnoses of diverticular bleed | 720
PUD | 720
arteriovenous malformations | 720
severe hemorrhoids | 720
repeat urgent colonoscopy | 720
transverse and descending colon diverticular disease | 720
left hemicolectomy | 720
previous abdominal aortic aneurysm (AAA) | 720
aortoenteric (AE) fistula | 720
exploratory laparotomy | 720
total abdominal colectomy | 720
excision of the AE fistula | 720
massive lower GI bleed | 720
right iliac artery aneurysm | 720
good health at a one-year follow-up | 8760