41 years old | 0
female | 0
history of untreated hypertension | -672
morbid obesity | -672
chronic back pain | -672
IVDU | -672
low back pain | -336
diffuse abdominal pain | -336
lower extremity weakness | -336
anorexia | -336
fever | -336
chills | -336
shortness of breath | -336
dizziness | -336
constipation | -336
acetaminophen | -336
gabapentin | -336
hydrocodone | -336
methamphetamines | -336
marijuana | -336
admitted to the hospital | 0
blood pressure of 79/53 mmHg | 0
heart rate of 149 bpm | 0
lactic acid of 4.2 mg dl-1 | 0
WBC 37 500 u l-1 | 0
erythrocyte sedimentation rate 75 mm h-1 | 0
urine toxicology positive for cannabis | 0
urine toxicology positive for amphetamines | 0
midline tenderness of the lumbar spine | 0
3/5 strength in bilateral lower extremities | 0
bilateral shoulder warmth | 0
bilateral shoulder erythema | 0
bilateral shoulder tenderness | 0
limited range of motion | 0
multiple needle puncture sites on the antecubital fossas | 0
puncture wounds on the right foot | 0
vancomycin | 0
metronidazole | 0
aztreonam | 0
IV fluids | 0
MRSA bacteraemia | 0
sensitivities to vancomycin | 0
sensitivities to rifampin | 0
sensitivities to levofloxacin | 0
sensitivities to clindamycin | 0
sensitivities to daptomycin | 0
sensitivities to linezolid | 0
bilateral shoulder plain radiographs | 0
arthrocentesis of the AC joints | 0
WBC of 93 137 u l-1 in one shoulder | 0
WBC of 32 043 u l-1 in the other shoulder | 0
MRSA in aspirates | 0
emergent surgical debridement of the shoulders | 0
intubation | 0
MRI of the lumbar spine | 0
L3-L5 osteomyelitis | 0
facet septic arthritis | 0
dorsal paraspinous myositis | 0
L2-L5 epidural abscess | 0
bilateral psoas myositis | 0
bilateral psoas abscesses | 0
MRI of the bilateral shoulders | 0
septic arthritis of the AC joints | 0
right distal trapezius abscess | 0
left supraclavicular abscess | 0
MRI of the brain | 0
TTE | 0
no valvular vegetations | 0
cardiology deferred transoesophageal echocardiogram | 0
repeat surgical debridement of the shoulders | 24
neurosurgery evaluation | 24
leukocytosis | 24
peak WBC of 52 100 u l-1 | 48
trough levels of vancomycin | 48
repeat blood cultures positive for MRSA | 48
antibiotics escalated to daptomycin | 240
antibiotics escalated to ceftaroline | 240
blood cultures became negative | 336
rifampin added | 336
repeat MRI of the lumbar spine | 336
worsening epidural abscess | 336
surgical drainage with drain placement | 432
intraoperative wound cultures positive for MRSA | 432
intraoperative wound cultures positive for Proteus mirabilis | 432
improved clinically | 480
all drains removed | 480
discharged | 672
oral levofloxacin | 672
oral rifampin | 672
lost to follow-up | 672