59 years old | 0
male | 0
admitted to the hospital | 0
intermittent diarrhea | -120
diarrhea with water-like stools | -120
abdominal pain | -120
nausea | -120
vomiting | -120
decreased production of dark-colored urine | -72
fatigue | -72
limb weakness | -72
Klebsiella pneumoniae bacteraemia | 0
sepsis | 0
septic shock | 0
septic AKI | 0
Acute Physiology and Chronic Health Evaluation score 18 | 0
Sequential Organ Failure Assessment score 10 | 0
temperature 38.5 °C | 0
pulse 128 beats/min | 0
respiration 22 breaths/min | 0
blood pressure 70/40 mmHg | 0
abdomen slightly puffy and soft | 0
upper abdominal pressure | 0
back pain | 0
bowel “chirping” 5-6 times/min | 0
hemoglobin level 18.3 g/dL | 0
total white blood cell count 21.4 × 10^9/L | 0
neutral granulocytes 71.9% | 0
platelet count 169 × 10^9/L | 0
metabolic acidosis | 0
blood gas pH 7.35 | 0
PCO2 30 mmHg | 0
PO2 66 mmHg | 0
PO2/FiO2 110 mmHg | 0
bicarbonate 16.6 mmol/L | 0
base excess -9.0 mmol/L | 0
lactate 3.5 mmol/L | 0
aspartate aminotransferase 573.1 U/L | 0
alanine aminotransferase 47 U/L | 0
total bilirubin 7.58 µmol/L | 0
serum creatinine 708.8 µmol/L | 0
urea 20.48 mmol/L | 0
albumin 26.9 g/L | 0
prothrombin time 12.5 s | 0
activated partial thromboplastin time 31.3 s | 0
international normalized ratio 1.08 | 0
procalcitonin 32.60 ng/mL | 0
empirical treatment with meropenem | 0
blood cultures | 0
Klebsiella pneumoniae | 0
meropenem sensitive | 0
intravenous crystalloid fluid | 0
invasive dynamic hemodynamic monitoring | 0
noradrenaline | 0
CRRT with oXiris hemofilter | 0
CVVHDF | 0
regional citrate anticoagulation | 0
mild hypocalcemia | 12
intravenous calcium supplementation | 12
noradrenaline infusion reduced | 65
noradrenaline infusion stopped | 65
lactate level 2.1 mmol/L | 6
lactate clearance rate 40% | 6
endotoxin level decreased | 6
interleukin-6 decreased | 6
interleukin-10 decreased | 6
procalcitonin level decreased | 72
urine volume increased | 240
SCr decreased | 72
SOFA score decreased | 72
APACHE II score decreased | 72
CRRT discontinued | 480
kidney function recovered | 480
discharged | 600