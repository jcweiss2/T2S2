63 years old | 0
farm worker | 0
admitted to infection ward | 0
weakness | 0
headache | 0
fever | 0
working in farm | -168
generalized myalgia | -168
malaise | -168
vomiting | -168
no abdominal pain | 0
no jaundice | 0
denied contact with animals | 0
positive surgical history | 0
no consumption of dairy products | 0
no travel to endemic areas | 0
alert | 0
oriented | 0
pyrexial (39.5°C) | 0
conjunctival suffusion | 0
no scleral jaundice | 0
normal skin | 0
normal heart | 0
normal lung | 0
bladder not felt | 0
liver not felt | 0
normal rectal examination |6 0
cranial nerves unremarkable | 0
kerning sign negative | 0
brudzinski sign negative | 0
headache increased permanently | 48
hiccup | 120
photophobia | 120
diplopic vision | 120
ptosis | 120
right preorbital edema | 120
normal eye movement | 120
eye deviation to medial site | 144
brainstem involvement | 168
unable to sit without support | 168
ataxic | 168
dysarthric | 168
uvula deviated to left | 168
lack of gag reflex | 168
right facial paresis | 168
transported to ICU | 168
decreased consciousness | 168
hemoptysis | 168
gastrointestinal bleeding | 168
normal abdominal sonography | 168
leptospirosis suspicion | 168
serum sample sent for testing | 168
L. serjoe hardjo 1/1600 | 168
neurological consultation | 168
MRI/MRV prescribed | 168
CST syndrome | 168
axial CT scan showed increased intensity | 168
no focal lesions | 168
normal cranial ventricles | 168
normal cisterns | 168
MRV loss of flow cavernous sinus | 168
right cavernous sinus expansion | 168
longitudinal filling defect | 168
parietal irregularities | 168
superior sagittal sinus normal | 168
transverse sinus normal | 168
sigmoid sinus normal | 168
internal jugular vein normal | 168
leptospirosis diagnosis | 168
