57 years old|0
female|0
hospitalized for acute respiratory failure from cardiogenic shock|0
chronic congestive heart failure|-4320
postpartum cardiomyopathy|-4320
type 2 diabetes|-4320
hypothyroidism|-4320
acute respiratory failure|-24
cardiogenic shock|-24
new-onset nonischemic cardiomyopathy|0
left ventricular ejection fraction drop from 57% to 5%|0
prolonged hospitalization|0
worsening preexisting hypokalemia|0
loop diuretics|0
spironolactone|0
losartan|0
serum morning cortisol elevated to 122.4 μg/dL|0
ACTH elevated to 181 pg/mL|0
serum morning cortisol repeated 75.7 μg/dL|0
ACTH repeated 170 pg/mL|0
low aldosterone/renin ratio|0
aldosterone <1.0 ng/dL|0
renin 0.92 ng/mL/h|0
24-hour free urine cortisol elevated to 6100 μg/24h|0
DHEA sulfate levels 62.3 μg/dL|0
Metanephrine plasma levels <10 pg/mL|0
CT abdomen showed symmetrical enlargement of both adrenal glands|0
right adrenal maximum diameter 7 cm|0
left adrenal maximum diameter 9 cm|0
pre-contrast Hounsfield units 40–45|0
postcontrast washout about 40%|0
denied recent weight gain|0
denied headaches|0
denied vision change|0
denied abdominal striae|0
denied proximal muscle weakness|0
denied hirsutism|0
denied acne|0
denied history of kidney stones|0
denied steroid use|0
blood pressure within normal range|0
no evidence of cushingoid features|0
pituitary MRI revealed normal pituitary gland|0
transthoracic echocardiogram showed LVEF 5%|0
improved cardiac condition with medical management|72
vasopressors|72
diuretics|72
3-week follow-up CT abdomen near resolution of adrenal enlargement|504
morning cortisol normalized 9.55 µg/dL|504
ACTH normalized 8.3 pg/mL|504
24-h free urine cortisol normalized 2 μg/24h|504
potassium levels normalized|504
minimal need for potassium replacement|504
LVEF improved from 5% to 10%|504
discharged from the hospital|504
cortisol and ACTH checks within normal limits at 6 weeks post-discharge|-504
readmitted 5 months later for septic shock due to pneumonia|3624
worsening cardiac failure|3624
subsequent liver failure|3624
gastrointestinal bleeding|3624
died|3624
morning cortisol level normal 9.11 µg/dL|3624
no autopsy completed|3624
admitted to intensive care unit|0
dobutamine 5 µg/kg/min|0
milrinone|0
diuresis with IV bumetamide|0
diuresis achieved|72
cardiovascular stability achieved|72
milrinone weaned off|72
transitioned to oral bumetamide|72
adrenal enlargement significantly improved|504
normalization of morning cortisol|504
normalization of ACTH|504
normalization of 24-h free urine cortisol|504
readmitted 5 months later|3624
septic shock due to pneumonia|3624
liver failure|3624
death|3624
cortisol normal during readmission|3624
no autopsy|3624
