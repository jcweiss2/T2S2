40 years old | 0
male | 0
admitted to ICU | 0
height 175 cm | 0
weight 90 kg | 0
type 1 diabetes mellitus | -8760
kidney transplant | -8760
diabetic kidney disease | -8760
mechanical ventilation | 0
agitation | 0
percutaneous thrombectomy | 0
acute ischemic stroke | 0
aspiration pneumonia | 24
septic shock | 24
increasing vasopressors requirements | 24
respiratory support | 24
transthoracic echocardiography | 24
new onset heart systolic murmur | 24
hypertrophic left ventricle | -120
no other pathological conditions | -120
dynamic left ventricular outflow tract obstruction | 24
severe mitral regurgitation | 24
systolic anterior motion of the mitral valve | 24
mean arterial pressure 65 mmHg | 24
norepinephrine 1.8 μg/kg/min | 24
non-fluid responsive | 24
control assisted ventilation | 24
FiO2 100% | 24
PEEP 15 mm Hg | 24
transesophageal echocardiography | 24
hypertrophic septum | 24
dynamic LVOTO | 24
maximum intraventricular gradient 165 mm Hg | 24
severe eccentric MR | 24
esmolol bolus | 24
hemodynamic improvement | 24
increase in MAP | 24
reduction in norepinephrine dose | 24
esmolol perfusion | 24
titrate esmolol dose | 24
norepinephrine reduction | 48
FiO2 reduction | 48
venous oxygen saturation augmentation | 48
lactate levels decrease | 48
hemorrhagic transformation of stroke | 288
neurological deterioration | 288
death | 288