high-grade fever | -48
influenza B virus infection | -48
wife diagnosed with influenza B virus infection | -72
daughters diagnosed with influenza B virus infection | -72
rapid test positive for influenza B antigens | -48
oseltamivir administered | -48
persistent fever | -24
dyspnea at rest | -24
admitted to hospital | 0
temperature 38.7°C | 0
blood pressure 117/80 mmHg | 0
heart rate 76 beats/min | 0
oxygen saturation level 88% | 0
fine crackles in lung fields | 0
white blood cell count 7400/mm3 | 0
C-reactive protein 18.1 mg/dL | 0
aspartate transaminase 91 IU/L | 0
L-lactate dehydrogenase 362 IU/L | 0
creatine kinase 793 IU/L | 0
Krebs von den Lungen-6 1772 U/mL | 0
arterial blood gas analysis showed hypoxemia | 0
high-flow nasal oxygen support started | 0
intravenous peramivir administered | 0
antibiotics administered | 0
Gram staining did not show bacterial infection | 0
Ziehl-Neelsen staining did not show bacterial infection | 0
periodic acid-Schiff stain did not show fungal infection | 0
sputum culture did not show bacterial or fungal infection | 0
blood cultures did not show bacterial infection | 0
reticular shadow on chest CT worsened | 72
PaO2/FiO2 ratio deteriorated to 83 | 72
diagnosed with severe ARDS | 72
mechanical ventilation proposed | 72
high levels of positive end-expiratory pressure proposed | 72
patient and family refused intubation | 72
polymyxin B-immobilized fiber column hemoperfusion performed | 72
intravenous methylprednisolone administered | 144
noninvasive positive pressure ventilation support started | 144
immunosuppressant therapy administered | 144
patient's condition worsened | 240
patient died | 3120
autopsy performed | 3120
pathological findings showed diffuse alveolar damage | 3120
no specific abnormality in other organs | 3120