18 years old male | 0
underwent orthotopic heart transplant for familial hypertrophic cardiomyopathy | -216
closely monitored in the cardiothoracic Intensive Care Unit postoperatively | 0
immunosuppressant regimen included prednisone | 0
immunosuppressant regimen included mycophenolate mofetil | 0
immunosuppressant regimen included tacrolimus | 0
extubated successfully | 48
developed sudden onset of shortness of breath | 72
hypoxic respiratory failure | 72
endotracheal intubation | 72
mechanical ventilation | 72
hemodynamically unstable | 72
requiring vasopressor support | 72
total white blood cell count of 48,000 cells/mm3 | 72
80% neutrophils | 72
14% bands | 72
3% lymphocytes | 72
3% monocytes | 72
renal function tests within normal range | 72
liver function tests within normal range | 72
blood cultures obtained | 72
broad-spectrum antibiotics initiated | 72
intravenous vancomycin | 72
cefepime | 72
azithromycin | 72
computed tomography of the chest revealed bilateral pulmonary consolidations | 72
computed tomography of the chest revealed air bronchograms | 72
computed tomography of the chest revealed bilateral pneumothoraces | 72
bronchoscopy performed | 96
bronchial washings performed | 96
bronchoalveolar lavage cultures revealed normal respiratory flora | 96
bronchoalveolar lavage cultures revealed Candida albicans | 96
blood cultures showed no microbial growth after 5 days of incubation | 168
marked leukocytosis persisted | 168
blood cultures repeated | 168
repeat CT chest demonstrated worsening diffuse pulmonary consolidations | 168
bronchoscopy performed | 216
BAL cultures of mycobacteria showed no growth | 216
BAL cultures of Mycoplasma pneumoniae showed no growth | 216
BAL cultures of Legionella showed no growth | 216
BAL viral cultures of adenovirus negative | 216
BAL viral cultures of Cytomegalovirus negative | 216
BAL viral cultures of influenza negative | 216
BAL viral cultures of parainfluenza negative | 216
BAL viral cultures of respiratory syncytial virus negative | 216
blood CMV viral load by PCR undetectable | 216
HIV serology nonreactive | 216
serum cryptococcal antigen sent | 216
serum Aspergillus galactomannan assay sent | 216
serum (1→3)-β-D-glucan assay sent | 216
urine for Histoplasma antigen sent | 216
BAL cytology demonstrated acute inflammatory cells | 216
Gomori's methenamine silver stain of BAL cytology negative for Pneumocystis jirovecii | 216
Gomori's methenamine silver stain identified acute angle septated hyphae suggestive of Aspergillus species | 216
BAL cultures isolated Aspergillus flavus | 216
minimal inhibitory concentration of voriconazole to A. flavus susceptible | 216
empiric therapy with intravenous voriconazole initiated | 216
empiric therapy with micafungin initiated | 216
serum Aspergillus galactomannan elevated at 4.8 OD | 216
serum (1→3)-β-D-glucan high at 263 pg/mL | 216
serum cryptococcal antigen negative | 216
urine Histoplasma antigen negative | 216
diagnosis of invasive pulmonary aspergillosis | 216
responded dramatically to combined antifungal therapy | 240
vasopressor support discontinued | 240
micafungin discontinued | 240
voriconazole transitioned to oral route | 240
review of day 4 BAL fungal cultures confirmed only Candida colonies | 216
patient's family denied gardening or spreading mulch prior to admission | 216
other organ recipients from same donor not diagnosed with invasive aspergillosis | 216
no hospital construction or renovation | 216
air sampling cultures conducted in patient's room | 216
air sampling cultures conducted in adjacent rooms | 216
mold spore concentrations in patient's room 78 S/m3 | 216
mold spore concentrations in adjacent rooms 26 S/m3 | 216
basidiospore variety detected | 216
no Aspergillus spore identified | 216
immunosuppression decreased | 216
bilateral chest tubes placed | 216
persistent air leak | 216
patient discharged on the 43rd posttransplant day | 1032
voriconazole maintenance monotherapy | 1032
repeat serum Aspergillus galactomannan assay 0.61 OD | 2016
voriconazole therapy for 6 months | 4320
complete pulmonary recovery achieved | 4320
off antifungal therapy for 1½ years | 13176
no clinical signs of relapse of Aspergillus infection | 13176
