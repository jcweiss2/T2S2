69 years old | 0
female | 0
breast cancer | -168
surgery for breast cancer | -168
zoledronic acid | -140
diabetes | 0
atrial fibrillation | 0
osteonecrosis | -84
necrosis involving the upper and lower jaw | -84
histological examination | -84
mechanical debridement | -84
washing with hydrogen peroxide | -84
iodopovidone | -84
1% chlorhexidine gel | -84
disinfected the oral cavity | -84
H2O2 | -84
0.2% chlorhexidine | -84
mandibular pain | -28
slight temperature | -28
signs of local inflammation | -28
spontaneous emission of pus | -28
amoxicillin and clavulanic acid | -28
metronidazol | -28
facial computed tomography scan | -28
multiple radiotransparent areas | -28
bilateral reactive laterocervical lymphadenopathy | -28
worsened local and general symptoms | -14
temperature of 39.1℃ | -14
tachycardia | -14
dysphagia | -14
dyspnea | -14
tachypnea | -14
extensive swelling of the face and neck | -14
bright red extended skin | -14
positive foveal sign | -14
incipient trismus | -14
mandible deviated to the right | -14
major discharge of pus | -14
panoramic radiograph | -14
full-thickness mandibular fracture | -14
CT scan of the face, neck, and chest | -14
thickening of the soft tissue | -14
multiple bilateral abscesses | -14
normal thoracic-mediastinal district | -14
right mandibular fracture | -14
white blood cell count of 42,100/mm3 | -14
C-reactive protein 31.7 mg/dL | -14
glycemia 183 mg/dL | -14
metronidazole | 0
ceftriaxone | 0
surgically drained | 0
necrosis of the superficial cervical fascia | 0
thrombosis in the anterior jugular veins | 0
necrotizing fasciitis | 0
empyema | 0
Staphylococcus epidermidis | 0
Pseudomonas aeruginosa | 0
Candida albicans | 0
ciprofloxacin | 4
imipenem | 4
hydrogen peroxide | 4
ceftazidime | 4
impaired cardiovascular function | 4
calcium antagonists | 4
beta blockers | 4
antiplatelet agents | 4
diuretics | 4
electrolytes | 4
albumin | 4
absence of empyema | 8
diffuse signs of pneumonia | 8
massive involvement on the left side | 8
septic shock | 10
kidney failure | 10
liver failure | 10
death | 10