76 years old | 0
female | 0
hypertension | -26280
type II diabetes mellitus | -21840
coronary heart disease | -13140
myocardial infarction | -13140
senile dementia | -13140
open cholecystectomy | -31920
abdominal wall hernia repairs | -6720
morbid obesity | 0
body mass index (BMI) 37.8 kg/m2 | 0
progressive abdominal pain | -120
admitted to the hospital | 0
septico-toxic shock | 0
acute abdomen | 0
recurrent, incarcerated and eventrated abdominal wall hernia | 0
eventrated hernia | 0
local defense musculaire | 0
abdominal ultrasonography | 0
laboratory tests | 0
chest X-ray | 0
native abdominal X-ray | 0
securing central venous access | 0
epidural cannulation | 0
intravesical catheter insertion | 0
urgent right upper transverse laparotomy | 0
local feculent peritonitis | 0
incarcerated and perforated ascending colon | 0
perforated terminal ileum | 0
extended right hemicolectomy | 0
resection of terminal ileum | 0
side-to-side ileo-transversostomy | 0
necrectomy | 0
abdominal gap | 0
biological graft unavailable | 0
synthetic mesh implantation not considered | 0
dermal-subcutaneous pannicule removed | 0
epidermis removed | 0
subcutaneous adipose tissue removed | 0
defect completed with dermal flaps | 0
first dermal graft inserted | 0
dermal graft fixed to abdominal wall | 0
external dermal graft fixed | 0
external dermal graft perforated | 0
greater omentum spared | 0
direct abdominal sutures not applied | 0
surgery took 250 min | 0
preparation of dermal grafts took 50 min | 0
intraoperative blood loss 740 mL | 0
intensive care | 0
empiric imipenem/cilastatin i.v. antibiotic therapy started | 0
thrombosis prophylaxis with enoxaparine s.c. started | 6
fever ceased | 96
bowel movement restarted | 120
red blood cell transfusions administered | 120
nasogastric tube left in place | 0
nasogastric tube removed | 72
oral nourishment started | 120
mobilisation started | 120
elastic abdominal belt put on | 120
intra-abdominal drain removed | 144
left subcutaneous drain removed | 168
right subcutaneous drain removed | 240
skin sutures removed | 360
discharged | 432
thrombosis prophylaxis prescribed | 432
wound healed per primam intentionem | 432
follow-up physical examinations | 720
follow-up blood tests | 720
follow-up abdominal wall ultrasonographies | 720
abdominal computed tomography | 1440
no hernia recurrency | 1440
no subcutaneous fistula or seroma formation | 1440