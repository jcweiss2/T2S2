42 years old | 0
male | 0
generalized weakness | -2160
fever | -2160
cough | -2160
12 kg weight loss | -2160
living in Guatemala | -2160
serum HIV-antibody test positive (ELISA) | -2160
sputum AFB smear positive | -2160
HIV-1 Western blot test positive | 0
CD4 cell count 10/µL | 0
HIV RNA titer 18,000 copies/mL | 0
anti-tuberculosis medications (isoniazid, rifampin, ethambutol, pyrazinamide) | 0
fluconazole | 0
trimethoprim/sulfamethoxazole | 0
generalized weakness persisted | 0
fever persisted | 0
admitted to KU hospital | 0
body temperature 37.6℃ | 0
oral thrush | 0
hepatosplenomegaly | 0
ascites | 0
hemoglobin 10.6 g/dL | 0
white blood cell 2,700/µL | 0
platelet 58,000/µL | 0
total bilirubin 2.4 mg/dL | 0
AST/ALT 131/48 IU/L | 0
ALP 114 IU/L | 0
GGT 133 IU/L | 0
chest X-ray costophrenic angle blunting | 0
chest X-ray fluid shifting in right hemithorax | 0
chest X-ray mild pneumonic infiltration in left lung | 0
disseminated tuberculosis suspected | 0
Mycobacterium tuberculosis identified from sputum culture | 0
anti-tuberculosis medication continued | 0
sputum AFB smear negative | 0
anti-retroviral agents (zidovudine, lamivudine, efavirenz) | 0
pancytopenia progressed rapidly | 0
hemoglobin 7.4 g/dL | 0
white blood cell count 1,070/µL | 0
platelet count 13,000/µL | 0
rifampin discontinued | 0
zidovudine discontinued | 0
trimethoprim/sulfamethoxazole discontinued | 0
pancytopenia persisted | 0
new pulmonary infiltrates | 120
septic shock | 120
empirical antibiotic therapy (piperacillin/tazobactam) | 120
transferred to intensive care unit | 144
mechanical ventilator support | 144
gram stain from sputum negative | 144
ordinary culture from sputum negative | 144
gram stain from blood negative | 144
ordinary culture from blood negative | 144
pancytopenia not improved | 144
pneumonia not improved | 144
hepatosplenomegaly not improved | 144
bone marrow aspiration | 216
bone marrow biopsy | 216
died | 240
Histoplasma capsulatum identified | 216
disseminated histoplasmosis confirmed | 216
