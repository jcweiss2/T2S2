67 years old | 0
male | 0
Indian | 0
admitted to the hospital | 0
type 2 diabetes mellitus | -8760
primary hypothyroidism | -8760
depression | -8760
gliclazide | -8760
thyroxine | -8760
venlafaxine | -8760
fever | -24
stupor | -24
generalized rigidity | -24
agitation | -72
visual hallucinations | -72
auditory hallucinations | -72
olanzapine | -24
clonazepam | -24
conscious | 0
irrelevant talk | 0
febrile | 0
tachycardia | 0
hypertension | 0
symmetric rigidity | 0
preserved deep tendon reflexes | 0
absent clonus | 0
flexor plantar reflex | 0
pupils equal and reacting to light | 0
intravenous fluids | 0
intravenous paracetamol | 0
physical cooling | 0
labetalol | 0
blood cultures | 0
routine haematology | 0
biochemistry | 0
creatinine phosphokinase levels | 0
NCCT head | 0
cerebro-spinal fluid analysis | 0
intubated | 12
mechanical ventilatory support | 12
dantrolene | 12
bromocriptine | 12
broad spectrum antibiotics | 12
supportive treatment | 12
neurological deterioration | 12
right extensor plantar response | 12
right hemiparesis | 12
acute haemorrhage | 12
left frontal deep and peri-ventricular white matter | 12
mild surrounding edema | 12
poly-microbial sepsis | 48
hospital-acquired pneumonia | 48
escalation of antibiotics | 48
anti-fungal drugs | 48
CPK values declined | 192
tracheostomised | 192
prolonged intubation | 192
gradual weaning trial | 192
uneventful recovery | 240
discharged | 240
mild residual weakness | 240
right upper limb | 240
right lower limb | 240