73 years old | 0 | 0 
female | 0 | 0 
hypertension | 0 | 0 
syphilis | 0 | 0 
type 2 diabetes mellitus | 0 | 0 
admitted to the hospital | 0 | 0 
altered mental status | 0 | 0 
mechanical fall | -720 | -720 
pruritic scalp | -720 | 0 
purulent drainage from sinuses on the scalp | -720 | 0 
temperature of 97.9°F | 0 | 0 
heart rate of 127 bpm | 0 | 0 
respiratory rate of 22 breaths/min | 0 | 0 
blood pressure of 144/80 mmHg | 0 | 0 
oxygen saturation of 98% on room air | 0 | 0 
oriented to person | 0 | 0 
oriented to place | 0 | 0 
not oriented to time | 0 | 0 
face, scalp and right ear were erythematous and edematous | 0 | 0 
large fluctuant mass with purulent drainage over the occipital and parietal portions of the scalp | 0 | 0 
posterior auricular mass without signs of active drainage | 0 | 0 
hyperglycemia to 700 | 0 | 0 
anion gap metabolic acidosis with serum bicarbonate of 20 | 0 | 0 
ketonuria | 0 | 0 
non-contrast head computed tomography (CT) | 0 | 0 
extensive multifocal scalp swelling along the right temporal, right posterior parietal and left frontal regions | 0 | 0 
no acute intracranial abnormalities | 0 | 0 
diabetic ketoacidosis | 0 | 0 
cellulitis of the scalp | 0 | 0 
concern for underlying abscesses | 0 | 0 
continuous infusion of insulin | 0 | 192 
intravenous Vancomycin | 0 | 192 
intravenous Cefepime | 0 | 192 
incision and drainage of scalp lesion | 48 | 48 
10-cm subgaleal abscess with large amounts of purulence evacuated | 48 | 48 
initial admission blood cultures grew MRSA | 72 | 72 
paranasal sinus CT with intravenous contrast | 72 | 72 
no involvement | 72 | 72 
transesophageal echocardiogram | 72 | 72 
no evidence for endocarditis | 72 | 72 
pulse irrigation of the wounds | 96 | 96 
sharp debridement | 96 | 96 
involvement of plastic surgery | 96 | 96 
serial bedside debridements | 96 | 192 
scalp wound measured 20 cm in length, 10 cm in width and 2 cm depth | 192 | 192 
right posterior auricular wound measured 7 × 7 × 2 cm | 192 | 192 
split-thickness skin grafts harvested from the right thigh | 192 | 192 
100% take of the grafts | 192 | 192 
discharged | 768 | 768 
intravenous Vancomycin to complete a full 7-week course | 768 | 1008 
skin graft healed well | 1008 | 1008 
some surrounding areas of hyperpigmentation | 1008 | 1008 
no areas of the graft were rejected | 1008 | 1008