57 years old | 0
male | 0
admitted to the hospital | 0
industrial accident | -744
C2 vertebral body fracture | -744
high cervical SCI at the C3 level | -744
no key muscle activity in all extremities | -744
last intact sensory level was the C3 dermatome | -744
deep anal pressure | -744
no voluntary anal contraction | -744
C3 AIS B | -744
pulmonary function test | -304
severely decreased pulmonary function | -304
tidal volume 220 mL | -304
vital capacity 800 mL | -304
peak cough flow 130 L/min | -304
continuous hypercapnia | -304
PaCO2 over 45 mmHg | -304
diaphragm fluoroscopy | -304
average length of the diaphragm apex decreased | -304
portable ventilator with volume controlled assisted ventilation mode | -304
active pulmonary rehabilitation techniques | -304
air stacking exercise with an Ambu bag | -304
sputum expectoration by mechanical insufflation-exsufflation | -304
accessory respiratory muscle training | -304
readmitted to the intensive care unit | -168
septic shock | -168
urinary tract infection | -168
tracheostomy | -168
step-by-step pulmonary rehabilitation program | -168
tracheostomy tube removed | -24
total weaning | -24
respiratory insufficiency | -24
concomitant sleep apnea | -24
aging | -24
intermittent NIV with pressure support ventilation mode | 0
nasal mask | 0
oral air leak | 0
full face mask | 0
anxiety | 0
limited communication | 0
novel alarm system | 0
microcontroller board | 0
sound generator | 0
pressure transducer | 0
endotracheal tube | 0
neck rotation | 0
sensor | 0
intended motion | 0
pressure exceeded 10 cm H2O | 0
single beep sound | 0
loud alarm sound | 0
discharged home | 24
no complications | 24