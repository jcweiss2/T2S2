67 years old | 0
male | 0
coronary artery disease | 0
type II diabetes | 0
hypertension | 0
peripheral vascular disease | 0
normal renal function | 0
admitted with septic arthritis of the right knee | 0
coronary artery bypass | -2904
Staphylococcus aureus infection at the site of the saphenectomy | -2904
numerous septicemias | -2904
disseminated Staphylococcus aureus infections involving the lungs | -2904
disseminated Staphylococcus aureus infections involving the right knee | -2904
disseminated Staphylococcus aureus infections involving the sternal wound | -2904
disseminated Staphylococcus aureus infections involving the surgical wound at the right femur | -2904
five surgical revisions | -2904
mechanically ventilated | -2904
ARDS | -2904
haemodynamically unstable | -2904
vasopressors required | -2904
broad-spectrum antibiotics | -2904
renal function deteriorated | 360
oliguric acute renal failure | 360
sepsis | 360
nephrotoxic medication | 360
COX-2 inhibitor | 360
gentamycin | 360
ACEI | 360
continuous venovenous haemofiltration | 912
uraemia | 912
metabolic acidosis | 912
encephalopathy | 912
serum creatinine stabilized | 1056
anuric ARF | 1344
no response to hydration | 1344
no response to diuretics | 1344
10% pentastarch received | 264
intermittent haemodialysis | 1608
normal sized kidneys | 1608
no hydronephrosis | 1608
dirty brown casts | 1608
no eosinophilia | 1608
fractional excretion of sodium 1.2% | 1608
furosemide | 1608
marked bilateral hypoperfusion | 1608
renal blood flow 255 ml/min | 1608
severe hydropic changes of the cytoplasm of tubular cells | 1608
discharged after a 6-month stay | 4320
chronic haemodialysis | 4320
By systematically parsing the timeline and converting all mentioned days into hours relative to admission, I constructed the comprehensive event table.</s>|
