79 years old | 0
male | 0
admitted to the hospital | 0
acute abdominal pain | -2
HPVG detected | -2
abdominal CT | -2
transferred to hospital | -2
stable vital signs | 0
body temperature: 37.2°C | 0
blood pressure: 112/74 mmHg | 0
pulse rate: 68 beats/min | 0
abdominal distention | 0
rebound tenderness | 0
abdominal guarding | 0
peritoneal irritation | 0
acute inflammation | 0
white blood cell count of 18 400/μL | 0
C-reactive protein concentration of 17.7 mg/dL | 0
dehydration | 0
metabolic acidosis | 0
base excess of −7.0 mmol/L | 0
elevated creatine kinase | 0
plain abdominal radiographs | 0
distention of the small intestine | 0
subileus | 0
contrast-enhanced abdominal CT | 0
HPVG | 0
contrast defect in a region of the small intestine | 0
small amount of ascites around the intestine | 0
no thrombus in any artery | 0
thickened appendix wall | 0
urgent laparotomy | 2
generalized peritonitis | 2
intestinal necrosis | 2
turbid ascites | 2
dilated small intestine | 2
discoloration of the appendix | 2
wall thickening of the appendix | 2
gangrenous appendicitis | 2
appendectomy | 2
abdominal drainage | 2
pathological findings | 4
no evidence of malignancy | 4
Escherichia coli positive in ascitic culture | 4
intravenous antibiotic treatment | 4
meropenem | 4
septic shock | 12
disseminated intravascular coagulation | 12
blood purification therapy | 12
admitted to ICU | 12
CT images on Day 7 | 168
HPVG disappeared | 168
left ICU | 168
discharged from hospital | 240