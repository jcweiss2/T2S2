37 years old|0
male|0
close contact with COVID-19 patient|-96
high-grade fever|-72
myalgia|-72
dry cough|-72
tested positive for COVID-19|-48
advised to self-isolate|-48
worsening shortness of breath|-24
bibasal crackles|0
gallop rhythm|0
resting tachycardia|0
no pedal oedema|0
lymphopaenia|0
raised CRP (74 mg/L)|0
lactate dehydrogenase (303 U/L)|0
BNP (247 pg/mL)|0
mildly deranged liver function tests|0
sinus tachycardia on ECG|0
bibasal infiltrates on chest X-ray|0
TTE showing LVEF 10%-15%|0
dilated left ventricle|0
ordered serial cardiac monitoring|0
high-grade temperature spikes (39°C–40°C)|0
CRP <100 mg/L|0
prescribed ceftriaxone|0
negative blood and urine cultures|0
CRP creeping up|72
changed to piperacillin/tazobactam|72
vancomycin added|72
renal functions deteriorating|120
creatinine clearance worsening|120
vancomycin levels normal|120
creatinine clearance <10 mL/min/1.73 m2|168
creatinine 657 μmol/L|168
oliguria|168
started haemodialysis|168
renal biopsy showing acute tubular injury|168
vancomycin stopped|168
intermittent haemodialysis for 8 days|168
improvement in ejection fraction|336
ejection fraction 25%-30%|336
renal function improving|336
no longer oliguric|336
stopped dialysis|336
follow-up cardiac MRI EF 46%|2064
renal function within normal range|2064
advised to self-isolate|2064
booked heart failure clinic follow-up|2064
booked renal clinic follow-up|2064
outcome symptom free|336
outcome ejection fraction improved|336
outcome renal function recovered|336
low-dose beta blocker|0
ACE inhibitor started|0
ACE inhibitor held|120
intravenous antibiotics|0
monitoring heart function|0
intensive care unit admission|168
discharged|336
learning points multisystemic COVID-19|0
learning points breathlessness non-respiratory|0
learning points atypical cardiorenal complications|0
learning points need for further research|0
