64 years old | 0
woman | 0
admitted for elective radical total gastrectomy | 0
feeding jejunostomy | 0
poorly differentiated T1 gastric carcinoma | 0
hypertension | -infinity (background history)
anemia | -infinity (background history)
no significant family history | 0
no significant psychosocial history | 0
no previous surgical history | 0
antihypertensive medication | -infinity (ongoing before admission)
progressed as expected postoperatively | 0
no immediate intraoperative complications | 0
jejunostomy feeds commenced | 24 (following day after admission)
routine postoperative contrast CT scan | 48 (day 2)
no anastomotic leak | 48
bilateral pleural effusions | 48
multiple vomits | 96 (day 4)
no bowel opening since procedure | 96
tachycardic (HR 140 bpm) | 96
febrile (39.4°C) | 96
dyspnoeic (RR 27, SpO2 96% on 6L O2) | 96
mildly tender abdomen | 96
cool peripheries | 96
pH 7.45 | 96
lactate 4.2 mmol/L | 96
white cell count 1.9 × 10^9/L | 96
CRP 456 mg/L | 96
septic workup | 96
repeat CT chest abdomen pelvis | 96
broad-spectrum antibiotics commenced | 96
suspected aspiration pneumonia | 96
markedly dilated Roux loop (obstruction) | 96
distended caecum and ascending colon (caecal volvulus) | 96
bilateral pleural effusions | 96
urgent exploratory laparotomy | 96
grossly distended caecal volvulus compressing jejunostomy | 96
obstruction of small bowel at jejunostomy sutures | 96
right hemicolectomy performed | 96
jejunostomy un-kinked | 96
small bowel viability confirmed | 96
feeding tube removed | 96
small bowel defect repaired | 96
bacteraemia developed | 96
intravenous antibiotics | 96
prolonged ICU admission | 96
tracheostomy | 96
ARDS | 96
pericardial effusion | 96
pleural effusions | 96
full recovery | 96
histology confirmed ischemic changes | 96
