22 years old | 0
female | 0
referred to trauma center | -96
railway accident | -96
below-knee amputation | -96
interlocking nail in bilateral femur | -96
open book pelvic bone fracture | -96
extensive Morel-Lavallée lesions over left flank | -96
conscious | 0
oriented | 0
stable hemodynamic parameters | 0
heart rate 90/min | 0
blood pressure 110/70 mm Hg | 0
respiratory rate 20/min | 0
regular dressing | 0
use of iv antibiotics meropenem | 0
use of iv antibiotics vancomycin | 0
sepsis | 0
surgical debridement of Morel-Lavallée lesion | 120
general anesthesia | 120
extensive necrotic area from left 12th rib to left thigh | 120
pelvic bone exposed | 120
hypotension | 120
inotropic support | 120
shifted to ICU | 120
persistent hypotension | 120
higher inotropic support | 120
high-grade fever 41°C | 120
rising total leukocyte count 30000/ml | 120
postoperative day 3 | 168
black foul smelling necrotic areas on wound | 168
cottony bread mold lesions on edges | 168
immediate surgical debridement | 168
extensive muscle necrosis | 168
peritoneum breached | 168
bowel exposed | 168
tissue for fungal culture | 168
histopathological examination | 168
nonseptate irregular hyphae of class zygomycetes | 168
provisional diagnosis of mucormycosis | 168
liposomal amphotericin B started | 168
fungal culture grew Rhizopus oryzae | 168
invasive mucormycosis | 168
died | 216
severe septic shock | 216
