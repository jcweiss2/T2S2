60 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
PAN | -8760 | 0 | Factual
paroxysmal atrial fibrillation | -8760 | 0 | Factual
hypertension | -8760 | 0 | Factual
dyslipidemia | -8760 | 0 | Factual
non-insulin dependent diabetes mellitus | -8760 | 0 | Factual
septic shock | -17520 | -17520 | Factual
scrotal pain | 0 | 0 | Factual
fever | 0 | 0 | Factual
fatigue | 0 | 0 | Factual
tachycardia | 0 | 0 | Factual
hypotension | 0 | 0 | Factual
vancomycin | 0 | 24 | Factual
Zosyn | 0 | 24 | Factual
broad-spectrum antibiotics | 0 | 24 | Factual
kidney function worsened | 24 | 48 | Factual
meropenem | 48 | 120 | Factual
creatinine level continued to rise | 48 | 120 | Factual
macular rash | 120 | 168 | Factual
axillary area rash | 168 | 192 | Factual
chest rash | 168 | 192 | Factual
head rash | 168 | 192 | Factual
neck rash | 168 | 192 | Factual
abdomen rash | 168 | 192 | Factual
mental status decline | 168 | 192 | Factual
bullae | 192 | 216 | Factual
vesicles | 192 | 216 | Factual
dermatology team involved | 192 | 216 | Factual
biopsy obtained | 216 | 216 | Factual
local steroid cream | 216 | 216 | Factual
AGEP diagnosis | 216 | 216 | Factual
kidney injury | 216 | 216 | Factual
neutrophilia | 216 | 216 | Factual
cyclic fevers | 216 | 216 | Factual
rash became pustular | 216 | 216 | Factual
high grade fever | 216 | 216 | Factual
transfer to ICU | 216 | 216 | Factual
pulse steroids | 216 | 240 | Factual
fever subsided | 240 | 240 | Factual
rash improvement | 240 | 240 | Factual
sloughing decreased | 240 | 240 | Factual
acute kidney injury resolution | 240 | 240 | Factual
steroid taper | 240 | 240 | Factual
skin biopsy | 0 | 0 | Factual
urine analysis | 0 | 0 | Factual
CT chest/abdomen/pelvis | 0 | 0 | Factual
CBC/BMP/coagulation | 0 | 0 | Factual
DRESS | 0 | 0 | Negated
GPP | 0 | 0 | Negated
PAN typical rash | 0 | 0 | Negated
Steven Johnson syndrome | 0 | 0 | Negated
leukocytoclastic vasculitis | 0 | 0 | Negated
subcorneal pustular dermatosis | 0 | 0 | Negated
cutaneous candidiasis | 0 | 0 | Negated
T cell-mediated neutrophilic inflammation | 0 | 0 | Factual
CD4+ T cells | 0 | 0 | Factual
cytotoxic CD8+ T cells | 0 | 0 | Factual
inflammatory cytokines | 0 | 0 | Factual
chemokines | 0 | 0 | Factual
CXCL8 | 0 | 0 | Factual
GM-CSF | 0 | 0 | Factual
neutrophil apoptosis | 0 | 0 | Factual
superficial infiltrate | 0 | 0 | Factual
interstitial infiltrate | 0 | 0 | Factual
mid-dermal infiltrate | 0 | 0 | Factual
dermal edema | 0 | 0 | Factual
intra- and subcorneal spongiform | 0 | 0 | Factual
PAN mechanism | 0 | 0 | Factual
immune complex-mediated disease | 0 | 0 | Factual
medium-sized arterial inflammation | 0 | 0 | Factual
arterioles | 0 | 0 | Negated
capillaries | 0 | 0 | Negated
venules | 0 | 0 | Negated
tender erythematous nodules | 0 | 0 | Negated
purpura | 0 | 0 | Negated
livedo reticularis | 0 | 0 | Negated
ulcers | 0 | 0 | Negated
bullous eruption | 0 | 0 | Negated
vesicular eruption | 0 | 0 | Negated
subcorneal accumulation of neutrophils | 0 | 0 | Negated
perivascular infiltrate of neutrophils | 0 | 0 | Negated
keratinocyte damage | 0 | 0 | Negated
systemic corticosteroids | 240 | 240 | Factual
immunosuppression | 240 | 240 | Factual
negative cultures | 0 | 0 | Factual
penicillin antibiotics | 0 | 0 | Negated