77 years old | 0
male | 0
Iraqi | 0
admitted to the hospital | 0
hypertension | -672
diabetes | -672
ischemic heart disease | -672
captopril | -672
metformin | -672
aspirin | -672
atorvastatin | -672
progressive weakness in lower limbs | -72
retention of urine | -72
loss of sensations in lower limbs | -72
febrile illness | -96
no shortness of breath | -96
no cough | -96
low-grade fever | 0
fine crackles | 0
normal S1 and S2 heart sounds | 0
distended bladder | 0
full consciousness | 0
normal vital signs | 0
normal higher cerebral function | 0
intact cranial nerves | 0
normal strength in upper limbs | 0
normal sensory examination in upper limbs | 0
flaccid paralysis in lower limbs | 0
hypotonia in lower limbs | 0
sensory level at T10 | 0
loss of sensations below T10 | 0
retention of urine | 0
elevated WBC count | 0
lymphopenia | 0
elevated renal indices | 0
typical feature of COVID-19 on chest CT | 0
normal degenerative change on cervical dorsal area MRI | 0
normal degenerative change on lumbosacral spine MRI | 0
negative PCR screening for other viruses | 0
negative serology tests for other infections | 0
negative interferon gamma release assays test | 0
methylprednisolone treatment | 0
insulin therapy | 0
ceftriaxone treatment | 0
azithromycin treatment | 0
positive RT-PCR test result | 24
shortness of breath | 48
admitted to intensive care unit | 48
mechanical ventilation | 48
multiorgan failure | 72
septicemia | 72
death | 72