44 years old | 0
male | 0
admitted to the hospital | 0
unknown history of diabetes mellitus | 0
10 days history of progressive left facial necrosis | -240
blurred vision of the left eye | -240
left periorbital pain | -240
swelling | -240
fever | -240
general malaise | -240
self-extracted left upper second decayed molar | -336
decayed tooth | -672
intermittent sharp pain | -672
poor oral hygiene | -672
loss of appetite | -672
hyperglycemic | 0
plasma glucose 576 mg/dL | 0
crepitus | 0
fluctuation | 0
local heat | 0
computed tomography | 0
diffuse subcutaneous emphysematous changes | 0
leukocytosis | 0
high CRP level | 0
metabolic acidosis | 0
high procalcitonin level | 0
septic status | 0
urgent operation | 0
tracheostomy | 0
naso-gastric tube | 0
surgical drainage | 0
debridement | 0
intensive care unit | 0
oxacillin | 0
ceftazidime | 0
blood cultures | 0
oxacillin-sensitive staphylococcus bacteremia | 0
staged and targeted surgeries | 24
extensive fasciotomy | 216
fasciectomy | 216
bicoronal incision | 216
upper blepharoplasty incision | 216
anterior facial flap | 216
occipital flap | 216
wound culture | 216
Pseudomonas aeruginosa | 216
Klebsiella pneumoniae | 216
vancomycin | 216
imipenem/cilastatin | 216
left medial thigh meshed split thickness skin graft | 432
discharged | 888
visual acuity of left eye preserved | 888