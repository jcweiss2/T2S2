74 years old | 0
female | 0
admitted to the hospital | 0
dyspnea on exertion | -48
dry cough | -48
chest pain | -48
myalgias | -720
malaise | -720
anorexia | -720
diagnosed with polymyalgia rheumatica | -720
treated with prednisolone | -720
tachypneic | 0
central cyanosis | 0
use of inspiratory accessory muscles | 0
bilateral inspiratory crackles | 0
severe hypoxemia | 0
pH 7.48 | 0
partial pressure of oxygen 49 mmHg | 0
partial pressure of carbon dioxide 31 mmHg | 0
oxygen saturation 83% | 0
anemia | 0
hemoglobin level 10.9 g/dL | 0
leukocytosis | 0
white blood cell count 11.5x10^9/L | 0
neutrophils 82% | 0
normal platelet count | 0
platelet count 213x10^9/L | 0
elevated inflammatory marker levels | 0
erythrocyte sedimentation rate 80 mm/h | 0
C-reactive protein 3710 mg/dL | 0
impaired kidney function | 0
serum creatinine 1.73 mg/dL | 0
diffuse bilateral patchy opacities on chest x-ray | 0
normal sinus radiographs | 0
treated with ceftriaxone | 0
treated with azithromycin | 0
noninvasive ventilation | 0
high-resolution computed tomography | 0
extensive ground-glass opacities | 0
consolidation in right upper lobe | 0
relative subpleural sparing | 0
abdomen computed tomography | 0
no pathological findings on abdomen computed tomography | 0
transferred to ICU | 96
rapidly worsening respiratory distress | 96
commencing circulatory failure | 96
intubated | 96
mechanical ventilation | 96
cardiovascular support | 96
fluids | 96
vasopressors | 96
decline of hemoglobin concentration | 96
hemoglobin level 7.9 g/dL | 96
marked leukocytosis | 96
white blood cell count 18.5x10^9/L | 96
neutrophils 92% | 96
worsening renal function | 96
creatinine 2.06 mg/dL | 96
active urine sediment | 96
dysmorphic red blood cells | 96
red blood casts | 96
negative transthoracic echocardiogram | 96
left ventricular systolic function normal | 96
fiberoptic bronchoscopy | 120
no endobronchial lesions | 120
hemorrhagic bronchoalveolar lavage fluid | 120
negative bacterial cultures | 120
negative mycobacterial cultures | 120
no cytological evidence of malignancy | 120
blood in stool | 120
colonoscopy | 120
mild edema on gut biopsy | 120
histopathologic changes of chronic colitis | 120
positive ANCA | 120
PR3-cANCA titer 1/80 | 120
negative antiglomerular basement membrane | 120
negative antinuclear antibodies | 120
negative extractable nuclear antigens | 120
negative serology for hepatitis B and C virus | 120
rheumatoid factor 10 IU/mL | 120
normal complement levels | 120
diagnosed with ANCA-associated vasculitis | 120
treated with high-dose steroids | 120
treated with cyclophosphamide | 120
treated with plasmapheresis | 120
clinical stabilization | 240
improvement of arterial blood gases | 240
resolution of ARDS on chest x-ray | 240
weaned from mechanical ventilation | 960
referred to rehabilitation unit | 960
died of sepsis | 1920
nosocomial pneumonia | 1920