58 years old | 0
male | 0
admitted to the hospital | 0
headache | -4320
progressive right hemiparesis | -4320
hyperreflexia | 0
positive right Babinski reflex | 0
left thalamic lesion | 0
ring-enhancement pattern | 0
leukocytosis | 0
anti-HIV antibodies negative | 0
N. beijingensis infection | 0
triple antibiotic therapy | 0
closed ventriculostomy system | 0
extensive swelling | 0
Ommaya reservoir insertion | 0
blood culture negative | 0
cerebrospinal fluid culture negative | 0
thoracoabdominal CT scan negative | 0
transthoracic echocardiogram negative | 0
transesophageal echocardiogram negative | 0
clinical improvement | 168
seizure episode | 168
anisocoria | 168
emergency CT scan | 168
orotracheal intubation | 168
severe swelling | 168
increased abscess size | 168
supratentorial ventriculomegaly | 168
cisternal obstruction | 168
emergency Ommaya puncture | 168
turbid-yellow liquid retrieved | 168
surgical intervention | 168
abscess drained | 168
capsule partially resected | 168
contralateral ventriculostomy system attached | 168
SIRS | 168
Pseudomonas aeruginosa tracheitis | 168
Klebsiella pneumoniae tracheitis | 168
vancomycin administration | 168
fever | 168
tachycardia | 168
chest X-ray multilobed opacities | 168
gram-positive bacilli presence | 168
septic shock suspected | 168
multiple antibiotic regimen | 168
vasoactive support required | 336
anticonvulsive management | 336
myoclonic movements | 336
CT scans without new development | 336
SIRS suggestive of multisystem infection | 504
increased blood urea nitrogen | 504
increased creatinine | 504
anuria | 504
increased ventilation requirements | 504
death | 504
no history of concomitant disease | 0
no immunosenescence | 0
no HIV co-infection | 0
no cancer chemotherapy | 0
no long-term immunomodulatory therapy | 0
no endocarditis | 0
no hydrocephalus | 336
no new development at abscess | 336
no mass or solid organ lesion | 0
no chest pain | 0
no shortness of breath | 0
no septic shock with pulmonary foci confirmed | 168
