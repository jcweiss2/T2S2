72 years old | 0
female | 0
admitted to the hospital | 0
decreased consciousness level | 0
stupor status | 0
history of elective left internal carotid artery stenting | -72
transient ischemic attack | -72
history of diabetes mellitus | 0
hypertension | 0
ischemic heart disease | 0
aspirin | -72
clopidogrel | -72
statins | -72
amlodipine | -72
valsartan | -72
antidiabetics | -72
sudden fall in consciousness level | -48
right hemiplegia | 0
brain computed tomography scan | 0
Doppler sonography | 0
totally occluded LICA | 0
unfractionated heparin | 0
carotid artery wired | 0
thrombosuction | 0
alteplase | 0
carotid stent thrombosis | 0
second carotid stenting procedure | 0
iatrogenic edge dissection | 0
LICA stenting | 0
postdilation | 0
patency of the LICA flow | 0
M1 and M3 branches of the middle cerebral artery normal | 0
M2 branch occluded | 0
transferred to intensive care unit | 0
intravenous nitroglycerin | 0
systolic blood pressure maintained | 0
control brain CT scan | 48
massive infarction in the MCA area | 48
expired | 96
sepsis | 96
ventilator-associated pneumonia | 96
disseminated intravascular coagulation | 96