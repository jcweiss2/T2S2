76 years old | 0
    woman | 0
    metastatic lung adenocarcinoma | -2160
    palliative chemoimmunotherapy | -2160
    fevers | 0
    dyspnea | 0
    cough | 0
    invasive ductal carcinoma of the right breast | -5520
    lumpectomy | -5520
    aromatase inhibitor | -5520
    20 pack-year tobacco use history | -306240
    ceased smoking 35 years ago | -306240
    recently traveled to the Southwest United States | -720
    no history of chest radiation | 0
    hypoxemia on exertion | -2160
    right upper lobe mass | -2160
    lung metastases | -2160
    liver metastases | -2160
    biopsy of the lung | -2160
    biopsy of the liver | -2160
    metastatic adenocarcinoma consistent with lung origin | -2160
    no actionable mutations on standard tumor molecular profiling | -2160
    carboplatin | -2160
    pemetrexed | -2160
    pembrolizumab | -2160
    administered intravenously every 21 days | -2160
    stable disease | -1080
    fevers (midway through the fourth cycle) | -1080
    dyspnea on exertion (midway through the fourth cycle) | -1080
    cough (midway through the fourth cycle) | -1080
    CT angiogram of the chest | 0
    no pulmonary embolism | 0
    confluent regions of consolidation in the lungs bilaterally | 0
    significantly worse on the left | 0
    small left pleural effusion | 0
    bilateral cavitary lung lesions | 0
    admitted to the intensive care unit | 0
    severe hypoxemic respiratory failure | 0
    PaO2/FiO2 ratio of 87 | 0
    broad-spectrum antibiotics | 0
    worsening hypoxemia on day three | 72
    endotracheal intubation | 72
    mechanical ventilation | 72
    positive end-expiratory pressure titrated | 72
    lung protective ventilation utilizing a low tidal volume strategy | 72
    bronchoscopy on day three | 72
    thin secretions in the left lower lobe | 72
    bronchoalveolar lavage studies | 72
    neutrophilic predominance (70%) | 72
    neutrophilic predominance (54%) | 72
    negative gram stain | 72
    negative bacterial culture | 72
    negative viral culture | 72
    negative legionella culture | 72
    negative fungal culture | 72
    negative nocardia culture | 72
    negative acid-fast bacteria culture | 72
    negative Aspergillus galactomannan antigen | 72
    negative blood markers of infection | 72
    negative urine markers of infection | 72
    transthoracic echocardiogram | 72
    mild symmetric left ventricular hypertrophy | 72
    normal right ventricular size | 72
    normal right ventricular systolic function | 72
    no significant valvular disease | 72
    no signs of increased filling pressures | 72
    no atrial septal defect | 72
    deferred lung biopsy | 72
    immune checkpoint inhibitor pneumonitis suspected | 72
    intravenous methylprednisolone (2 mg/kg/day) | 72
    significant desaturations on day nine | 216
    FiO2 of 0.8 | 216
    positive end-expiratory pressure of 10 cmH2O | 216
    negative total body fluid balance | 216
    steroid-refractory pembrolizumab-induced pneumonitis | 216
    intravenous immunoglobulin (IVIg) | 216
    IVIg administered on days 9–13 | 216
    rapid and significant clinical improvement | 216
    radiographic improvement | 216
    successful extubation on day 12 | 288
    repeat chest CT imaging on day 12 | 288
    marked improvement in severe interstitial abnormality | 288
    organizing phase of acute lung injury | 288
    clinical response to immunomodulatory therapy | 288
    transitioned to prednisone (1 mg/kg/day) | 336
    supplemental oxygen requirement decreased | 336
    weaned to an oxymizer device | 336
    discharged on day 23 | 552
    oxygen needs decreased to 1.5 L per minute | 1344
    improved exercise tolerance | 1344
    prednisone decreased to 0.5 mg/kg/day | 1344
    slow taper over 2 months | 1344
    re-staging CT of the torso performed six weeks after admission | 1008
    continued improvement of the left-sided infiltrate | 1008
    remaining bilateral subpleural interstitial fibrotic abnormality | 1008
    stable malignant disease burden | 1008
    <|eot_id|>
    