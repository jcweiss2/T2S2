42 years old|0
    male|0
    admitted to the hospital|0
    severe abdominal pain|0
    fever|0
    body temperature of 39°C|0
    jaundice|0
    severe weakness|0
    sick for at least 3 weeks|-504
    rise in body temperature to subfebrile ranges|-504
    pain in the right hypochondrium|-504
    radiating to the lower back|-504
    chills|-504
    body temperature rose to 38.5°C|-504
    went to the doctor| -240
    absence of instrumental confirmation|-240
    acute pyelonephritis diagnosed|-240
    antibiotic therapy prescribed|-240
    oral ciprofloxacin|-240
    analgesics|-240
    ketoprophen|-240
    nimesulide|-240
    treatment had no effect|-240
    abdominal pain sharply increased|0
    spread to the entire right half of the abdomen|0
    yellowness of the skin|0
    sclera|0
    darkening of the urine|0
    severe jaundice|-175200
    viral hepatitis excluded|-175200
    cholecystostomy performed|-175200
    transferred to university surgical clinic|-175200
    tumor of the pancreatic head suspected|-175200
    operated upon|-175200
    surgical revision|-175200
    study of biopsy specimens|-175200
    pancreatic cancer not excluded|-175200
    pancreatoduodenectomy performed|-175200
    cholecystectomy performed|-175200
    external drainage of pancreatic remnant duct|-175200
    postoperative period|-175200
    pancreatic drainage spontaneously migrated|-175200
    no further complications|-175200
    spontaneous internal fistula suspected|-175200
    discharged|-175200
    histological examination|-175200
    chronic pancreatitis confirmed|-175200
    final diagnosis|-175200
    chronic pancreatitis with pancreatic head fibrosis|-175200
    multiple small pancreatic abscesses|-175200
    compression of the common bile duct|-175200
    obstructive jaundice|-175200
    felt relatively good|0
    diagnosed with diabetes mellitus|-17520
    insulin therapy prescribed|-17520
    worked as a driver|0
    smoked for about 20 years|0
    consumed alcohol very rarely|0
    followed medical recommendations|0
    severe general condition|0
    ill|0
    adynamic|0
    moderate yellowness of the skin|0
    sclera|0
    hot skin|0
    body temperature 38.9°C|0
    heart rate 100 beats per minute|0
    blood pressure 110/70 mm Hg|0
    abdomen painful|0
    moderately tender|0
    rebound tenderness present|0
    hemoglobin 113 g/l|0
    erythrocytes 4.0×10^12/l|0
    leukocytes 13.9×10^9/l|0
    neutrophils 90%|0
    platelets 279×10^9/l|0
    ALT 810 U/l|0
    AST greater than 913 U/l|0
    amylase 5 U/l|0
    total bilirubin 277 μmol/l|0
    glucose 28.0 mmol/l|0
    creatinine 49 μmol/l|0
    prothrombin index 65%|0
    INR 1.28|0
    free gas under right hemidiaphragm|0
    heterogeneity of liver shadow|0
    gas-fluid levels in liver tissue|0
    signs of bowel paresis|0
    dissimilarity of liver tissue|0
    hyperechoic lesions|0
    thick fluid|0
    gas in right subdiaphragmatic space|0
    signs of portal hypertension|0
    portal vein diameter 14 mm|0
    chronic pancreatitis in pancreatic remnant|0
    no free fluid in abdominal cavity|0
    rupture of liver abscess suspected|0
    peritonitis suspected|0
    perforation of ulcer not excluded|0
    emergency surgery scheduled|0
    midline laparotomy|0
    brownish muddy fluid in right paracolic gutter|0
    iliac fossa|0
    organs forming conglomerate|0
    purulent8hemorrhagic fluid outflow|0
    liver tissue debris|0
    abscess cavity 12x10x8 cm|0
    intraoperative endoscopy|0
    no ulcer in gastric stump|0
    jejunal loop freed from adhesions|0
    abscess cavity flushed|0
    abdominal cavity flushed|0
    postoperative period|0
    prolonged mechanical ventilation|36
    inotropic support with epinephrine|36
    sepsis diagnosed|36
    procalcitonin 5.1 ng/ml|36
    Staphylococcus haemolyticus in blood|36
    Klebsiella pneumoniae in urine|36
    Escherichia coli in urine|36
    E. coli in pus|36
    S. haemolyticus in pus|36
    Klebsiella in peritoneal exudate|36
    Acinetobacter in peritoneal exudate|36
    vancomycin|36
    meropenem|36
    amikacin|36
    right8sided pneumonia|36
    bilateral pleural effusions|36
    pleural cavities drained|240
    transferred to surgical ward|336
    gradual improvement|336
    reduction of liver lesion|336
    discharged|960
    subphrenic drains|960
    serous8purulent fluid|960
    bile staining|960
    drains removed|2736
    satisfactory condition|1344
    works as driver|1344
    receives insulin|1344
    enzyme replacement therapy|1344
    liver tissue healed|1344
    no biliary hypertension|1344
    non8dilated bile ducts|1344
    atrophic pancreatic remnant|1344
    non8dilated Wirsung duct|1344
    mild hyperglycemia|1344
    low serum amylase|1344
    normal blood test parameters|1344
    normal biochemistry|1344
    normal coagulograms|1344