66 years old | 0\
    male | 0\
    coronary artery bypass surgery | -17520 (assuming medical antecedent from 66 years old, approximate 20 years ago)\
    percutaneous coronary intervention | -17520\
    chronic obstructive pulmonary disease | -17520\
    diabetes | -17520\
    myelo-dysplastic syndrome | -17520\
    75-pack years of smoking | -17520\
    ongoing pain during defecation | -1344 (2 months before admission)\
    hematochezia observed during bowel preparation | -1344\
    colonoscopy | 0\
    unstable bleeding in the sigmoid colon | 0\
    admitted to the hospital | 0\
    alert | 0\
    hypotensive | 0\
    normal heart rate | 0\
    fever of 38.9 °C | 0\
    tenderness in the lower left quadrant | 0\
    anaemic (haemoglobin 6.0 mmol/L) | 0\
    intravenous fluid stabilization | 0\
    blood cultures made | 0\
    intravenous antibiotics given | 0\
    contrast-enhanced CT revealed retroperitoneal bleeding from left external iliac artery | 0\
    emergency damage control endo-grafting | 0\
    temperature fluctuating between 37−39 °C | 72 (3 days after admission)\
    intermittent left-sided abdominal pain | 72\
    septic | 72\
    CT-scan showed hematoma with air near covered stent and sigmoidal colon | 72\
    Clostridium tertium found in blood cultures | 72\
    white blood count decreasing | 72\
    C-reactive-protein concentration decreasing | 72\
    control CT-scan after nine days revealed regression of infected hematoma | 216 (9 days after admission)\
    thickening of the sigmoid colon | 216\
    informed about surgical options | 216\
    exploratory laparotomy | 216\
    confirmed fistula | 216\
    Hartmann’s procedure performed | 216\
    infected stent removed | 216\
    femoro-femoral bypass operation performed | 216\
    intensive care unit stay for 5 days | 216\
    hypotension during ICU stay | 216\
    pain during ICU stay | 216\
    slow recovery | 216\
    good recovery | 216\
    histological examination revealed diverticulitis with abscess, inflammation, perforation | 504 (3 weeks post-operatively)\
    signs of infection in left groin | 504\
    CT-scan confirmed infection | 504\
    treated with intravenous antibiotics | 504\
    re-incision with drainage | 504\
    rinsing of abscess cavity | 504\
    discharged | 672 (3 weeks + discharge after 2 weeks treatment, total 5 weeks)\
    oral antibiotics for 2 weeks | 672\
    control appointment after 2 weeks | 840 (2 weeks post-discharge)\
    no signs of vascular prosthesis infection | 840\
    antibiotics discontinued | 840\
    no further follow-up | 840\
    patient experienced stress regarding colostomy | 840\
    expressed gratefulness about recovery | 840\
    