41 years old | 0
woman | 0
followed up in the outpatient clinic for menorrhagia | 0
no significant medical history | 0
no significant surgical history | 0
no significant social history | 0
no significant family history | 0
drug allergy to amoxicillin | 0
presented to the outpatient clinic for menorrhagia | -103248
presented to the outpatient clinic for dysmenorrhea | -103248
managed with tranexamic acid | -103248
managed with mefenamic acid | -103248
managed with iron supplements | -103248
regular ultrasound pelvis done every 6 months | -103248
normal endometrial thickness | -103248
normal ovaries | -103248
stable adenomyoma (4.5 cm) | -103248
on regular follow-up | -103248
symptom of heavy menstrual flow worsened | -103248
requiring multiple hospital admissions for blood transfusions | -103248
requiring multiple hospital admissions for intravenous iron infusion | -103248
levonorgestrel-releasing IUD (Mirena) inserted on three occasions | -103248
expelled soon after insertion | -103248
trial of norethisterone | -103248
developed palpitations | -103248
offered definite surgical treatment with total hysterectomy bilateral salpingectomy | -103248
decided to proceed with the operation | 0
total laparoscopic hysterectomy bilateral salpingectomy (TLHBS) | 0
adenomyotic, 12-week size uterus | 0
normal tubes | 0
normal ovaries | 0
specimen retrieved vaginally | 0
estimated blood loss of 200 mL | 0
TLHBS completed uneventfully | 0
retrieval of the specimen difficult due to bulky and globular uterus | 0
adenomyotic uterus 'cored' with tissue scissors | 0
manipulated forward and backward into the abdominal cavity and vagina | 0
mild chronic endocervicitis in the cervix | 0
benign findings (leiomyoma and adenomyosis) | 0
recovering well | 24
ambulating independently | 24
on soft diet | 24
developed fever | 48
developed epigastric discomfort | 48
developed nausea | 48
developed diarrhea | 48
CT abdomen and pelvis performed | 72
fluid collection superior to the bladder | 72
symptoms not improving despite escalating antibiotic regimen | 120
symptoms worsened | 120
became unwell with high-grade temperatures | 120
developed abdominal bloating | 120
developed epigastric pain | 120
developed vomiting | 120
developed watery green stools | 120
intra-abdominal drain inserted under ultrasound guidance | 168
fluid collection superior to the bladder drained | 168
green-debris-laden fluid drained | 168
fluid culture grew Candida | 168
immunocompromised state screen negative | 168
bowel injury screen negative | 168
symptoms resolved after intravenous fluconazole | 240
drain removed | 240
discharged home | 288
oral antibiotics (ciprofloxacin and metronidazole) | 288
fluconazole to complete for 2 weeks | 288
repeat scans in 4 weeks showed marked reduction in collection | 672
CT abdomen and pelvis revealing the collection (predrainage) | 72
CT abdomen and pelvis image at 4-week follow-up | 672
HIV screen non-reactive | 168
DM screen HbA1c 4.9% | 168
blood culture no bacterial growth | 168
urine culture no bacterial growth | 168
stool culture no Salmonella | 168
stool culture no Shigella | 168
stool culture no Campylobacter | 168
stool culture no Vibrio species isolated | 168
stool culture no Clostridium difficile isolated | 168
stool microscopy no ova | 168
stool microscopy no cysts | 168
stool microscopy no trophozoites | 168
stool microscopy no parasites seen | 168
fluid culture Candida albicans | 168
Gram stain smear blastoconidia with pseudohyphae | 168
intravenous fluconazole commenced | 168
marked improvement in clinical state | 168
symptoms resolved | 240
asymptomatic at 4-week follow-up | 672
repeat CT abdomen and pelvis showed marked reduction in collection | 672
vaginal swab performed on POD 8 | 192
vaginal swab negative | 192
recurrent inflammatory smears | 0
vaginal candidiasis on PAP smears | 0
lower genital swabs | 0
DNA probe test for Candida | 192
white cell count normal | 168
C reactive protein elevated | 168
Candida peritonitis post caesarean section | 0
Candida chorioamnionitis | 0
screening test for lower genital tract infection | 0
