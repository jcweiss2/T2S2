64 years old| 0
male | 0
penetrating abdominal trauma | -22*24
emergency surgery | -22*24
intra-abdominal exsanguinating bleeding | -22*24
duodenal disruption | -22*24
multiple small bowel perforation | -22*24
duodenojejunostomy | -22*24
resection of about 150 cm of small bowel | -22*24
anastomosis | -22*24
bleeding control | -22*24
sepsis | -22*24+delta
multiorgan failure | -22*24+delta
referred to our institution | -22*24
surgical reexploration | -22*24+22*24
enteroenteric anastomosis failure | -22*24+22*24
large amount of bilestained fluid in the abdomen | -22*24+22*24
remaining small bowel less than 1 m | -22*24+22*24
pyloric exclusion not considered | -22*24+22*24
pancreaticoduodenectomy not considered | -22*24+22*24
enteroenterostomy | -22*24+22*24
duodenal primary repair | -22*24+22*24
feeding tube placement distal to perforated duodenum | -22*24+22*24
massive irrigation | -22*24+22*24
multiple drain tube placement | -22*24+22*24
intensive care | -22*24+22*24
ventilator weaning | -22*24+22*24
transfer to general ward | -22*24+22*24
enteral feeding through jejunal feeding tube | -22*24+22*24
severe retraction of duodenum | -22*24+22*24
duodenal disruption gap approximately 5 cm | -22*24+22*24
abdominal wall defect | -22*24+22*24
impossible to close duodenum primarily | -22*24+22*24
impossible to close wall defect primarily | -22*24+22*24
decision to use free flap for abdominal wall defect repair | -22*24+22*24
persistent leakage of gastric, bile, and pancreatic juice | -22*24+22*24
diversion of bile and pancreatic juices via endoscopic retrograde cholangiopancreaticography | -22*24+22*24
placement of pancreatic duct drainage tube | -22*24+22*24
placement of bile duct drainage tube | -22*24+22*24
placement of first covered expandable metallic stent (16mm diameter, 90mm long) | -22*24+22*24
reestablished duodenal continuity | -22*24+22*24
diversion through endoscopic nasobiliary drainage | -22*24+22*24
diversion through endoscopic nasopancreatic drainage | -22*24+22*24
first stent migration downward 5 days after placement | (-22*24+22*24) +5*24
removal of first stent through abdominal defect | (-22*24+22*24) +5*24
placement of second covered expandable metallic stent (16mm diameter, 130mm long) | (-22*24+22*24) +5*24
stent sutured tightly to duodenum | (-22*24+22*24) +5*24
debridement | (-22*24+22*24) +5*24 +7*24
closure of abdominal wall defect with free flap | (-22*24+22*24) +5*24 +7*24
duodenostomy with drainage tube placement | (-22*24+22*24) +5*24 +7*24
decompression of duodenum | (-22*24+22*24) +5*24 +7*24
prevention of infection | (-22*24+22*24) +5*24 +7*24
endoscopic images at 3 months post-stent placement | ((-22*24+22*24) +5*24 +7*24) + (112-7)*24
stent electively removed 112 days after placement | ((-22*24+22*24) +5*24 +7*24) + (112-7)*24
removal of pancreatic duct drainage tube | ( ((-22*24+22*24) +5*24 +7*24) + (112-7)*24 ) +13*24
removal of bile duct drainage tube | ( ((-22*24+22*24) +5*24 +7*24) + (112-7)*24 ) +13*24
oral food intake after stent removal | ( ((-22*24+22*24) +5*24 +7*24) + (112-7)*24 ) +13*24
complete healing of abdominal wall defect | ( ((-22*24+22*24) +5*24 +7*24) + (112-7)*24 ) +13*24
small enterocutaneous fistula observed | ( ((-22*24+22*24) +5*24 +7*24) + (112-7)*24 ) +13*24
upper gastrointestinal water-soluble contrast study on 234th postoperative day | 234*24
good passage of contrast | 234*24
small enterocutaneous fistula | 234*24
no significant obstruction | 234*24
