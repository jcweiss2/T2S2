54 years old|0
male|0
decompensated nonalcoholic steatohepatitis cirrhosis|0
orthotopic liver transplant (OLT)|0
side-to-side cavoplasty|0
duct-to-duct biliary anastomosis|0
end-to-end portal vein anastomosis|0
end-to-end common hepatic artery (HA) anastomosis|0
discharged home|168
physical therapy|168
19 months post-OLT|-1314
syncope|-1314
trimalleolar left ankle fracture|-1314
ibuprofen 800 mg 3 times per day|-1314
arthralgias|-1314
advised to discontinue ibuprofen|-1314
not taking proton pump inhibitors|-1314
dark stools|0
vomiting fresh blood with clots|0
hemoglobin drop (5 g)|0
intubated|0
urgent upper endoscopy|0
hemorrhagic shock|0
resuscitated with blood products|0
duodenal ulcer (2-3 cm)|0
large visible vessel in ulcer|0
endoscopic epinephrine injection|0
endoclips|0
bipolar electrocautery|0
unsuccessful hemostasis|0
no antral biopsies|0
stool Helicobacter pylori testing recommended|0
mesenteric angiogram|0
no active extravasation|0
proper HA luminal narrowing and irregularity|0
nonfilling of gastroduodenal artery (GDA)|0
aspartate aminotransferase 2,686 U/L|0
alanine aminotransferase 3,406 U/L|0
ischemic hepatitis|0
computed tomography angiogram|0
severe proper HA stenosis|0
moderate common HA stenosis|0
GDA occlusion|0
multifocal hepatic infarcts|0
duodenal thickening|0
surgical intervention|0
exploratory laparotomy|0
duodenum adherent to donor HA|0
full-thickness ulceration of duodenum|0
HA folded at anastomosis|0
HA pseudoaneurysm|0
resection of aneurysmal segment|0
new end-to-end HA anastomosis|0
ultrasound demonstrating excellent flow|0
Graham patch sutured on duodenum|0
right upper quadrant drain|0
intubated in ICU|0
perioperative antibiotics|0
Streptococcus mitis group infection|0
Haemophilus influenzae infection|0
extubated|48
open reduction and internal fixation of left ankle|96
liver functions normalized|96
normal HA flow on ultrasound|96
discharged|312
subacute rehab facility|312
medically stable|312
