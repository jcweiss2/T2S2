64 years old | 0
female | 0
Hepatitis C-induced liver cirrhosis | 0
end-stage renal disease | 0
chronic anemia | 0
hypothyroidism | 0
admitted to the emergency department | 0
fatigue | 0
weakness | 0
blurry vision | 0
shortness of breath |#0
fell | -72
abrasion on left forearm | -72
developed blisters on left forearm | 0
hyperpigmentation | 0
edema | 0
hemorrhagic bullae | 0
diminished breath sounds | 0
bibasilar crackles | 0
white blood cell count 19,550 | 0
lactic acid 10.7 | 0
chest CT scan bibasilar atelectasis | 0
chest CT scan consolidation | 0
abdominal CT scan hepatosplenomegaly | 0
abdominal CT scan cirrhosis | 0
abdominal CT scan portal venous hypertension | 0
abdominal CT scan ascites | 0
diagnosed septic shock | 0
cellulitis | 0
pneumonia | 0
placed on pressors | 0
admitted to intensive care unit | 0
infectious disease consultation | 0
Aeromonas infection suspected | 0
gentamicin | 0
Levaquin | 0
vancomycin | 0
Zosyn | 0
orthopedic surgery consultation | 0
blisters aspirated | 0
no excisional debridement | 0
white blood cell count 12,350 | 24
blood cultures released | 72
Aeromonas veronii complex | 72
isolate resisted ampicillin-sulbactam | 72
isolate resisted piperacillin-tazobactam | 72
antibiotics narrowed to ceftazidime | 72
antibiotics narrowed to gentamicin | 72
received post-dialysis vancomycin | 72
remained stable | 0
discharged | 240
