38 years old | 0
male | 0
rectal mucous discharge | -1728
no rectal bleeding | -1728
no altered bowel habits | -1728
family history of pancreatic cancer | 0
colonoscopy | -48
nodular-mixed type lateral spreading tumor | -48
tumor in the lower rectum | -48
tumor measuring 40 mm | -48
histopathology | -48
tubular-villous adenoma | -48
high-grade dysplasia | -48
endorectal ultrasound | -24
mixed echogenicity image | -24
uTisN0 | -24
tumor on the posterior wall of the rectum | -24
tumor located 4.0 cm from the anal verge | -24
endoscopic transanal resection | 0
no complications | 0
no rectal perforation | 0
wound closed by running suture | 0
transanal endoscopic operation system | 0
colon mechanical preparation | -12
surgical antibiotic prophylaxis | -12
ciprofloxacin | -12
metronidazole | -12
resected lesion histologically analyzed | 12
tubular-villous adenoma | 12
high-grade dysplasia | 12
intramucosal carcinoma | 12
surgical margins negative | 12
no abdominal discomfort | 24
no nausea | 24
no fever | 24
solid food tolerated | 24
diffuse abdominal pain | 48
asthenia | 48
heart rate 122 beats/min | 48
respiratory rate 25 breaths/min | 48
painful abdomen | 48
white blood cell count 10,270/mm3 | 48
immature forms 14% | 48
serum C-reactive protein level 25 mg/dL | 48
metabolic acidosis | 48
elevated lactic acid | 48
diagnosis of abdominal focus of sepsis | 48
volume expansion initiated | 48
antibiotics changed | 48
piperacillin-tazobactam | 48
admitted to intensive care unit | 48
abdominal radiography | 72
pneumoretroperitoneum | 72
computed tomography of abdomen | 72
retroperitoneal air | 72
laparotomy | 96
diffuse retroperitoneal gas infiltration | 96
loop colostomy | 96
opening of rectal wound | 96
hospitalized in intensive care unit | 96
discharged | 264
stoma closed | 4320