55 years old| 0
    male | 0
    presented to the emergency department | 0
    malaise | -336
    fever | -336
    weakness | -336
    weight loss | -336
    sore throat | -336
    dry cough | -336
    stab wounds | -672
    splenectomy | -672
    denied tick bites | -672
    febrile (38.2 C) | 0
    tachypneic | 0
    tachycardic | 0
    jaundice | 0
    acute renal injury | 0
    creatinine 5.2 mg/dl | 0
    creatinine increased to 10 mg/dl | 24
    mild liver injury | 0
    elevated INR (1.47) | 0
    mixed hyperbilirubinemia (10.7 mg/dl) | 0
    direct bilirubin 7.4 mg/dl | 0
    elevated lactate dehydrogenase (975 U/L) | 0
    undetectable haptoglobin | 0
    peripheral blood smear intracellular parasites | 0
    parasitemia 11.8% | 0
    B. microti detected by PCR | 0
    fulminant babesiosis infection | 0
    multi-organ systemic failure | 0
    atovaquone | 0
    azithromycin | 0
    transferred to medical intensive care unit | 0
    deteriorating kidney function | 24
    positive c-ANCA | 24
    positive ANA | 24
    low complement levels | 24
    exchange transfusions | 24
    parasitemia dropped to 2% | 24
    parasitemia dropped to 0.1% | 24
    clinical status improved | 24
    laboratory parameters improved | 24
    resolution of parasitemia | 1440
    creatinine 0.9 mg/dl | 1440
    negative c5-ANCA | 1440
    