92 years old | 0
female | 0
admitted to the hospital | 0
hypertension | -672
atrial fibrillation | -672
dementia with Lewy bodies | -672
sick sinus syndrome | -672
orthostatic hypotension | -672
falls at home | -672
rabeprazole | -672
mianserin | -672
clean 2 cm wound on the right leg | -672
fever | -648
erythema | -648
edema of the right leg | -648
lymphangitis | -648
dermohypodermitis | -648
antimicrobial treatment with amoxicillin | -648
venous Doppler | -648
no thrombosis | -648
injury extended to the entire lower limb | -645
purplish discoloration of the skin | -645
bullae | -645
necrosis | -645
severe pain | -645
morphine administration | -645
limited leg movements | -645
necrotizing fasciitis | -645
blood cultures | -645
broad-spectrum antibiotic therapy | -645
piperacillin | -645
tazobactam | -645
gentamicin | -645
deteriorated condition | -645
low blood pressure | -645
high heart rate | -645
low body temperature | -645
high respiratory rate | -645
low oxygen saturation | -645
reduced consciousness | -645
distended abdomen | -645
dyspnea | -645
computed tomography scan | -645
no pneumonia | -645
no abdominal or pelvic infection | -645
low white cell count | -645
low hemoglobin | -645
low platelet count | -645
high C-reactive protein | -645
low blood glucose | -645
high procalcitonin | -645
high troponin | -645
low pH | -645
low HCO3 | -645
high blood lactate | -645
no urine infection | -645
septic shock | -645
fluid challenge | -645
transfer to intensive care unit | -645
mechanical ventilation | -645
inotropic support | -645
antibiotic administration | -645
death | 0
Klebsiella pneumoniae | -648
hyper mucoviscous colonies | -648
positive string test | -648
resistance to amoxicillin | -648
resistance to piperacillin | -648
resistance to ticarcillin | -648
capsular serotype K2 | -648
RmpA | -648
aerobactin | -648
yersiniabactin | -648
sequence type ST86 | -648