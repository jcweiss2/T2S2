31 years old | 0
female | 0
admitted to the hospital | 0
chronic hypertension | -672
SLE | -672
hydroxychloroquine | -672
deep venous thrombosis | -672
enoxaparin | -672
postpartum | -96
heavy vaginal bleeding | 0
tachycardia | 0
hypotension | 0
fever | 0
anemia | 0
thrombocytopenia | 0
liver function tests normal | 0
fibrinogen normal | 0
renal function normal | 0
intravenous fluid resuscitation | 0
red blood cells transfusion | 0
platelet transfusion | 0
broad-spectrum antibiotics | 0
enoxaparin discontinued | 0
hydroxychloroquine discontinued | 0
intrauterine balloon tamponade | 0
vaginal bleeding ceased | 0
hemodynamics improved | 0
platelet count decreased | 24
anemia | 24
schistocytes | 48
haptoglobin normal | 48
bilirubin normal | 48
reticulocyte count normal | 48
autoimmune panel evaluation | 72
complement levels | 72
cardiolipin antibodies | 72
antinuclear antibody | 72
anti-Smith | 72
dsDNA | 72
SSA/SSB | 72
ADAMTS-13 activity | 72
antibodies against hydroxychloroquine | 72
heparin-induced thrombocytopenia panel | 72
persistent-elevated blood pressure | 72
epigastric pain | 72
acute kidney injury | 72
magnesium sulfate | 72
granular casts | 72
proteinuria | 72
absent dysmorphic red blood cells | 72
acute aphasia | 120
altered mental status | 120
PLEX | 144
rituximab | 216
vincristine | 264
methylprednisolone | 168
discharged | 432