65 years old | 0
male | 0
Caucasian | 0
admitted to the hospital | 0
hypertension | -8760
persistent AF | -8760
irritative cough | 336
respiratory origin | 336
severe headache | 504
persistent cough | 504
fever | 504
unremarkable vital signs | 504
excessive coughing | 504
anticoagulant therapy | 504
leukocytosis | 504
brain computed tomography | 504
subarachnoid hemorrhage | 504
warfarin withheld | 504
broad-spectrum antibiotics | 504
shortness of breath | 504
transthoracic echocardiography | 504
bubbles in left ventricle | 504
bubbles in left atrium | 504
communication with esophagus | 504
communication with bronchial tree | 504
mechanical ventilation | 504
endotracheal tube | 504
right main bronchus | 504
upper endoscopy | 504
large clot | 504
distal esophageal wall | 504
covered stent | 504
cardiac arrest | 504
resuscitation attempts | 504
futile | 504
pronounced dead | 504
autopsy | 504
fistula | 504
esophagus | 504
left atrium | 504
radiofrequency pulmonary vein isolation procedure | -336
catheter-based procedure | -336
DRESS syndrome | -10080
minocycline | -10080
acne | -10080
fever and rash | -10080 
diffuse erythematous or maculopapular eruption | 0
pruritus | 0
increased WBC count | 0
eosinophilia | 0
systemic involvement | 0
discharged | 24