35 years old | 0
male | 0
admitted to the hospital | 0
right-sided upper back and flank pain | 0
cupping procedure | -24
intermittent fevers | -504
cough | -504
anorexia | -504
general malaise | -504
seen multiple naturopathic physicians | -504
urgent care visit | -168
started on azithromycin | -168
started on doxycycline | -168
presumptive diagnosis of pneumonia | -168
improvement in febrile symptoms | -168
improvement in overall well-being | -168
blood pressure of 116/75 mmHg | 0
heart rate of 119 beats per minute | 0
respiratory rate of 20 breaths per minute | 0
temperature of 36.2°C | 0
O2 saturation of 97% | 0
alert | 0
appropriate | 0
no signs of respiratory distress | 0
cupping marks on his back | 0
absence of breath sounds on the right side of the chest | 0
abdomen was soft | 0
abdomen was non-tender | 0
chest radiograph | 0
80% opacification of the right hemithorax | 0
pneumonia | 0
parapneumonic effusion | 0
bedside ultrasound | 0
hepatic abscess | 0
CT of the chest, abdomen and pelvis | 0
10.2 × 8.9 × 12.6 cm abscess in the right lobe of the liver | 0
white blood cell count of 25×10^9/L | 0
creatinine of 92 mmol/L | 0
lactate of 3.5 mmol/L | 0
liver transaminases were within normal limits | 0
international normalized ratio was within normal limits | 0
O2 requirements increased to 4L | 0
blood pressure started to trend down | 0
blood pressure dropped to 90/60 | 0
heart rate of 108 | 0
treated with 2 liters of normal saline | 0
started on levofloxacin | 0
started on vancomycin | 0
started on piperacillin/tazobactam | 0
thoracocentesis | 0
33,688 u/L white blood cells | 0
93% neutrophils | 0
initial gram stain was negative | 0
antibiotics switched to ceftriaxone | 0
antibiotics switched to metronidazole | 0
admitted to the surgical intensive care unit | 0
central line placement | 0
interventional radiology guided liver abscess drainage | 0
percutaneous drain placement | 0
tube thoracostomy | 0
VATS decortication procedure | 0
diaphragmatic defect was found | 0
continuous with the hepatic abscess cavity | 0
no microorganisms found on gram stain | 0
no microorganisms found on subsequent cultures | 0
discharged from hospital | 720
spent 1 month on intravenous ceftriaxone | 720
spent 1 month on intravenous metronidazole | 720
antibiotics discontinued | 720