43 years old | 0
female | 0
sickle cell disease | 0
admitted to the hospital | 0
headache | -1440
dizziness | -1440
personality changes | -1440
behavioral changes | -1440
recurrent vomiting | -1440
axillary temperature 37.4°C | 0
heart rate 156 bpm | 0
respiratory rate 22 cpm | 0
blood pressure 112/84 mmHg | 0
SpO2 99% | 0
endoscopic evaluation of the sinuses | 0
sinus infection | 0
functional endoscopic sinus surgery | 0
debridement of the slough and dead tissue | 0
local intranasal ceftriaxone | 0
local intranasal caspofungin | 0
brain CT scan | 0
left frontal intra-axial thick-walled ring-enhancing lesion | 0
extensive surrounding edema | 0
craniotomy | 24
excisional biopsy of the frontal lobe lesion | 24
intraoperative diagnosis | 24
left granulomatous invasive fungal sinusitis | 24
erosion of the sella turcica and lateral sphenoid bone | 24
cavernous sinus | 24
Aspergillus flavus | 48
resistant to amphotericin B | 48
susceptible to voriconazole | 48
susceptible to itraconazole | 48
susceptible to posaconazole | 48
Aspergillus antigen test negative | 48
invasive sinus aspergillosis | 48
intracerebral aspergilloma | 48
voriconazole treatment | 48
caspofungin treatment | 48
seizures | 168
sepsis | 168
renal impairment | 168
malnutrition | 168
pancytopenia | 168
high risk of aspiration pneumonia | 168
intubated | 168
drowsy | 168
Glasgow coma scale 11/15 | 168
convulsive movements | 168
Salmonella sepsis | 168
ventriculitis | 168
renal function tests abnormal | 168
high creatinine | 168
blood urea nitrogen levels high | 168
second craniotomy | 192
subgaleal abscess | 192
left epidural abscess | 192
subdural abscess | 192
intraventricular abscess | 192
external ventricular drain | 192
cerebrospinal fluid analysis | 192
red blood cell count 50/mm3 | 192
WBC 700×106/L | 192
polymorphs 90% | 192
mononuclear cells 10% | 192
ampicillin-resistant Salmonella | 192
ciprofloxacin-resistant Salmonella | 192
ceftriaxone treatment | 192
brain CT scan | 192
purulent fluid | 192
edema | 192
mass effect on the frontal horn of the lateral ventricles | 192
communication with the left frontal horn | 192
abscess collection in the left lateral ventricle | 192
ventriculitis | 192
died | 240