14 years old | 0
    female | 0
    admitted to the hospital | 0
    fatigue | -672
    nose bleeding | -672
    generalized ecchymosis over the body | -672
    arthralgia | -672
    pallor | 0
    tachycardia | 0
    dermal/mucosal petechiae | 0
    ecchymosis | 0
    liver palpable 6 cm below mid-costal line | 0
    spleen palpable 4 cm below mid-costal line | 0
    leukocyte count of 333,000/mm3 | 0
    hemoglobin level of 4 g/dl | 0
    platelet count of 29,000/mm3 | 0
    peripheral blood smear with 97% L1-type blasts | 0
    myeloperoxidase negative blastic cells | 0
    pre-B-cell ALL detected by immunophenotyping | 0
    normal transaminases | 0
    normal blood urine nitrogen | 0
    normal creatinine | 0
    normal uric acid | 0
    normal phosphor | 0
    high lactate dehydrogenase (2,970 IU/ml) | 0
    leukopheresis performed two times | 0
    lumbar puncture done on 4th day | 96
    no cells in cerebrospinal fluid | 96
    benign cerebrospinal fluid cytology | 96
    modified BFM protocol (Turk ALL 2000) given | 0
    PBS smear on 8th day showing 1,395/mm3 blast count | 192
    no hematologic remission in bone marrow aspiration on 15th day | 360
    blast rate 27% on 15th day | 360
    no hematologic remission in bone marrow aspiration on 33rd day | 792
    blast rate 12% on 33rd day | 792
    high-risk group inclusion | 792
    BCR)ABL fusion gene positive | 0
    t(9;22) in 11 out of 20 metaphases | 0
    first course of HR1 block therapy given | 0
    imatinib started (400 mg/m2/day) | 0
    severe mucositis developed | 0
    total parenteral nutrition initiated | 0
    severe intractable gastrointestinal hemorrhage | 0
    erythrocyte transfusion | 0
    platelet transfusion | 0
    severe neutropenia | 0
    fever reached 39°C | 0
    CRP positive (26 mg/dl) | 0
    HR2 block treatment not started | 0
    imatinib continued regularly | 0
    bone marrow aspiration 37 days after HR1 completion | 888
    remission seen in bone marrow | 888
    depressive mood | 888
    no verbal cooperation | 888
    decreased muscle strength | 888
    increased muscle tonus | 888
    deep tendon reflex increased | 888
    Babinski test positive | 888
    normal cranial MRI | 888
    severe mucositis ongoing after 43 days | 1032
    hemorrhagic diarrhea | 1032
    typhlitis | 1032
    hyperemesis | 1032
    TPN continued | 1032
    sudden unconsciousness | 1032
    Glasgow coma score 7 | 1032
    cardiac pulse 34/min | 1032
    arterial blood pressure 70/30 mm Hg | 1032
    capillary perfusion time 3 s | 1032
    hypothermia | 1032
    WBC 2,030/mm3 | 1032
    absolute neutrophil count 1,640/mm3 | 1032
    hemoglobin 5.09 g/dl | 1032
    platelets 44,000/mm3 | 1032
    CRP 6.8 mg/dl | 1032
    urea 113 mg/dl | 1032
    creatinine 0.9 mg/dl | 1032
    glucose 136 mg/dl | 1032
    AST 77 IU/l | 1032
    ALT 91 IU/l | 1032
    bilirubin 0.3 mg/dl | 1032
    GGT 88 IU/l | 1032
    prothrombin time 17.6 s | 1032
    INR 1.4 | 1032
    activated partial thromboplastin time 43 s | 1032
    D-dimer 1,211 ng/ml | 1032
    fibrinogen 190 mg/dl | 1032
    normal blood electrolytes | 1032
    metabolic acidosis (lactic acid 12.6 mmol/l) | 1032
    transfer to Pediatric Intensive Care Unit | 1032
    intensive fluid replacement | 1032
    positive inotropic support | 1032
    erythrocyte suspension | 1032
    thrombocyte suspension | 1032
    left ventricular ejection fraction 64% | 1032
    broad-spectrum antibiotics for sepsis and septic shock | 1032
    encephalopathy progression | 1032
    generalized tonic-clonic convulsions | 1032
    intubation | 1032
    mechanical ventilation | 1032
    cranial CT showing 9-mm bleeding region | 1032
    peripheral edema in left basal ganglion | 1032
    supportive treatment with NaHCO3 for 12 h | 1032
    lactic acidosis progression (lactic acid 20 mmol/l) | 1032
    hemodiafiltration performed | 1032
    thiamine deficiency suspected | 1032
    intravenous thiamine 4 × 25 mg/day started | 1032
    lactic acidosis regression | 1032
    thiamine continued for 3 months | 1032
    transfusion-dependent anemia | 0
    transfusion-dependent thrombocytopenia | 0
    prolonged febrile neutropenia | 0
    persistent severe mucositis | 0
    gastrointestinal hemorrhage | 0
    encephalopathy | 0
    convulsions | 0
    chemotherapy discontinuation | 0
    bone marrow examination two months after HR1 completion | 1488
    bone marrow remission | 1488
    BCR-ABL gene fusion negative | 1488
    mechanical ventilation for 1 month | 0
    extubation | 720
    PEG performed | 2880
    swallowing dysfunction | 2880
    54 days in intensive care unit | 1296
    cognitive functions returned to normal after 6 months | 4320
    mucositis slow regression | 4320
    physiotherapy for spastic tetraparesis | 4320
    discharge home after 9 months | 6480
    imatinib continued | 6480
    no convulsions recurrence | 6480
    started walking with support at 9 months post-discharge | 9720
    walked independently at 12 months post-discharge | 13104
    PEG closed after 5 months | 3600
    oral feeding resumed | 3600
    no transfusion needed after 6 months post-HR1 | 4320
    bone marrow examinations every 3 months | 4320
    morphological remission observed | 4320
    molecular remission observed | 4320
    no matched donor found | 4320
    morphological remission at 30 months post-diagnosis | 21600
    molecular remission at 30 months post-diagnosis | 21600
    <|eot_id|>
    