56 years old | 0
female | 0
admitted to the hospital | 0
weakness | -744
numbness | -744
lower extremities | -744
hands | -744
neck | -744
type 2 diabetes mellitus | -8760
hypertension | -8760
necrotizing pancreatitis | -8760
gallstones | -8760
total parenteral nutrition (TPN) | -4380
albuminocytologic dissociation | 0
cerebrospinal fluid (CSF) | 0
Guillain-Barré syndrome (GBS) | 0
intravenous immunoglobulin (IVIG) | 0
encephalopathy | 120
pancytopenia | 120
hypotensive | 168
blood pressure of 64/48 mmHg | 168
unresponsive to verbal stimuli | 168
minimally responsive to painful stimuli | 168
Glasgow Coma Scale (GCS) score of 6 | 168
anasarcic | 168
flaccid paralysis | 168
calcium of 6.7 mg/dL | 168
hemoglobin of 9.4 g/dL | 168
white cell count of 2.1×10^9/L | 168
phosphorus of 1.1 mg/dL | 168
creatinine <0.2 mg/dL | 168
albumin <1.5 gm/dL | 168
lactate of 4 mmol/L | 168
malnutrition | 168
sepsis | 168
meropenem | 168
vancomycin | 168
anidulafungin | 168
intravenous fluids | 168
norepinephrine | 168
high-dose intravenous thiamine | 168
electroencephalogram (EEG) | 168
diffuse slow waves | 168
severe metabolic encephalopathy | 168
brain magnetic resonance imaging (MRI) | 168
hyperintensity of the bilateral medial thalamus | 168
Wernicke’s encephalopathy | 168
serum thiamine level of 104 nmol/L | 168
improved mental status | 336
able to understand simple commands | 336
discontinued norepinephrine | 336
discontinued antimicrobial treatment | 336
extubated | 360
electromyography (EMG) | 504
severe sensorimotor polyneuropathy | 504
transferred out of the intensive care unit (ICU) | 1008