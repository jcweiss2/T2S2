66 years old | 0
woman | 0
presented with fever | -192
fever | -192
close contact with confirmed COVID-19 case | -192
SARS-CoV-2 RNA detected | -192
initial supportive treatment | -192
headache | 0
fatigue | 0
muscle aches | 0
mild abdominal pain | 0
diarrhoea | 0
vomiting | 0
presented to hospital | 0
hypertension | 0
osteopenia | 0
Perindopril/Amlodipine | 0
Cholecalciferol | 0
ex-smoker | 0
20 pack years | 0
no history of immunosuppression | 0
no chronic organ dysfunction | 0
no history of fungal colonization | 0
independent in activities of daily living | 0
fever (40°C) | 0
respiratory rate 26/min | 0
pulse 80/min | 0
blood pressure 120/70 mmHg | 0
oxygen saturation 89% on room air | 0
increase in work of breathing | 0
bibasal coarse crepitations | 0
arterial blood gas | 0
pH 7.44 | 0
PaO2 70 mmHg | 0
PaCO2 34 mmHg | 0
lactate 0.9 mmol/L | 0
white blood cell count 5.3 ×109/L | 0
neutrophil differential count 3.9 ×109/L | 0
lymphocyte count 1.2 ×109/L | 0
AST 52U/L | 0
ALT 32 U/L | 0
GGT 61U/L | 0
LDH 429 U/L | 0
normal renal function | 0
blood cultures isolated Facklamia hominis | 0
urine culture isolated Escherichia coli | 0
susceptible to Ceftriaxone | 0
chest radiology demonstrated pulmonary opacities | 0
admitted to COVID-19 respiratory ward | 0
Ceftriaxone 1g daily | 0
Azithromycin 500mg daily | 0
supplemental oxygen | 0
subcutaneous enoxaparin sodium | 0
no specific COVID-19 therapy | 0
condition deteriorated | 24
progressive dyspnoea | 24
increasing oxygen requirement | 24
admitted to ICU | 24
temperature 39.5°C | 24
respiratory rate 40/min | 24
oxygen saturation 91% on HFNP | 24
FiO2 40% | 24
airflow 40 L/m | 24
no heart failure signs | 24
echocardiogram demonstrated normal biventricular function | 24
mild right ventricular dilatation | 24
arterial blood gas on FiO2 40% | 24
pH 7.46 | 24
PaO2 59 mmHg | 24
PaCO2 31 mmHg | 24
awake prone positioning | 24
no improvement in oxygenation | 24
endotracheal intubation | 24
mechanical ventilation | 24
lung-protective ventilation | 24
deterioration in ventilatory parameters | 24
severe ARDS criteria | 24
worsening respiratory function | 192
hypercapnoea | 192
fever absent | 192
CRP 351mg/L | 192
ALT 125 U/L | 192
AST 154 U/L | 192
GGT 611 U/L | 192
ALP 229 U/L | 192
ferritin 1295 μg/L | 192
D-dimer 0.99mg/L | 192
fibrinogen 5.8g/L | 192
chest radiology progression | 192
ETT sample obtained | 192
SARS-CoV-2 RNA persistent | 192
7-day Piperacillin/Tazobactam | 192
prone ventilation | 192
improvement in ventilatory parameters | 192
fungal elements on Gram stain | 192
Aspergillus fumigatus complex isolated | 192
three subsequent ETT cultures isolated Aspergillus | 192
new onset fever | 240
bilateral consolidation | 240
intravenous Voriconazole initiated | 240
fever settled | 264
inflammatory markers improved | 264
liver function normalized | 264
Voriconazole trough levels 2.72mg/L | 264
extubated | 288
oral Voriconazole 300mg twice daily | 288
two negative SARS-CoV-2 RT-PCR | 360
discharged home | 360
CECT chest | 432
bilateral organising pneumonia | 432
fibrosis | 432
segmental pulmonary embolism | 432
Voriconazole ceased | 432
Apixaban | 432
liver function testing | 432
Voriconazole trough level 3.6mg/L | 432
mild dry cough | 432
improved effort tolerance | 432
no systemic features | 432
