50 years old | 0
Japanese man | 0
idiopathic pulmonary fibrosis | -192
hypoxia | -192
acute exacerbation of idiopathic pulmonary fibrosis | -192
broad-spectrum antibiotics | -192
prednisolone | -192
deteriorated clinical condition | -192
intubated | -192
mechanically ventilated | -192
aggressive mechanical ventilation | -192
PaCO2 88 mmHg | -192
PaO2 48 mmHg | -192
FIO2 1.0 | -192
V-V ECMO | -192
21-Fr drainage cannula in left femoral vein | -192
19-Fr return cannula in right femoral vein | -192
condition stabilized | -192
tracheostomy | -192
no improvement | -192
legal issues preventing LTx in Singapore | -192
transported to ICU in Japan | 0
sedated | 0
mechanically ventilated | 0
ECMO blood flow 4 L/min | 0
SpO2 over 85% | 0
sweep gas flow 100% oxygen | 0
PaCO2 30-35 mmHg | 0
mechanical ventilation lung rest settings | 0
driving pressure 5 cmH2O | 0
PEEP 10 cmH2O | 0
FIO2 0.4 | 0
heart rate 50 beats/min | 0
blood pressure 156/104 mmHg | 0
no inotropes | 0
echocardiography ejection fraction 60.7% | 0
TR-PG 10 mmHg | 0
normal renal function | 0
heparin anticoagulant | 0
activated partial thromboplastin time 50D80 seconds | 0
vancomycin prophylaxis | 0
other antibiotics as required | 0
gradual improvement | 24
mechanical ventilation discontinued | 912
awake | 1008
tracheostomy tube removed | 1008
speech cannula inserted | 1008
speech cannula removed | 1008
low-flow oxygen therapy | 1008
high-flow oxygen therapy | 1008
nasal cannula | 1008
Venturi mask | 1008
SpO2 over 85% | 1008
oral intake | 1128
severe respiratory failure | 1128
no other organ failure | 1128
target SpO2 achieved | 1128
target PaCO2 achieved | 1128
fine adjustment of ECMO blood flow | 1128
fine adjustment of sweep gas flow | 1128
supplemental oxygen through native lung | 1128
analgesia with morphine | 1128
fully awake | 1128
oriented | 1128
communicative | 1128
physiotherapist daily | 1128
exercise | 1128
respiratory training | 1128
clinical decision for irreversible respiratory failure | 1128
listed on LTx registry | 1128
LTx evaluation consultation | 1416
changed membrane oxygenator 23 times | 1416
changed cannula 10 times | 1416
membrane oxygenator changes due to gas exchange failure | 1416
membrane oxygenator changes due to thrombus | 1416
membrane oxygenator changes due to acute platelet reduction | 1416
average oxygenator lifespan 16 days | 1416
cannula changes due to sepsis | 1416
cannula changes due to blood stream infection | 1416
two-site cannulation mode | 1416
right internal jugular vein drainage four times | 1416
right femoral vein drainage four times | 1416
left femoral vein drainage three times | 1416
left internal jugular vein return three times | 1416
right femoral vein return three times | 1416
left femoral vein return one time | 1416
25 or 23-Fr cannula for drainage | 1416
23 or 21-Fr cannula for return | 1416
no technical complications | 1416
dyspnea | 5352
SpO2 90% | 5352
ECMO flow 5 L/min | 5352
echocardiography D shape | 5352
TR-PG 56 mmHg | 5352
TR-PG 27 mmHg on day 201 | 4824
bosentan | 5352
sildenafil | 5352
worsening right failure | 5424
TR-PG 78 mmHg | 5424
ECMO conversion to VV-A | 5424
condition improved | 5424
TR-PG decreased to 43 mmHg | 5424
ECMO conversion back to V-V | 6768
listed on LTx registry | 6816
attempted cannula change | 7320
occluded veins due to thrombosis | 7320
unable to access veins | 7320
used same cannula from day 276 | 7320
septic shock | 8904
attempted cannula change again | 8904
no flow in veins by echocardiography | 8904
relatively stable | 8904
able to talk | 8904
maintained oral intake | 8904
decided to disconnect ECMO | 8904
ECMO disconnected | 9672
patient died | 9672
no autopsy | 9672
