63 years old|0
    male|0
    employed as a dentist|0
    outpatient dental clinics|0
    experienced systemic reaction|0
    acute and diffuse urticaria|0
    recurrent loss of consciousness|0
    treated with steroids|0
    treated with epinephrine|0
    anaphylactic shock suspected|0
    transitory loss of consciousness|-8760
    laryngeal hyper-reactivity|-8760
    Skin Prick Tests for common inhalant allergens negative|0
    Skin Prick Tests for latex allergens negative|0
    Immuno-CAP for chlorhexidine-specific IgE 0.04 kU/L|0
    total IgE 46.7 kU/L|0
    BAT performed for phenol|0
    BAT performed for ortho-phthalaldehyde|0
    BAT performed for chlorhexidine|0
    CD63 expression 14.5%|0
    stimulation index SI 6.0|0
    mouthwash containing chlorhexidine CD63 9.6%|0
    mouthwash containing chlorhexidine SI 4.0|0
    other disinfectants tested negative|0
    2.0% solution chlorhexidine digluconate|0
    mixed with tetradecyltrimethylammonium bromide|0
    mixed with dodecyltrimethylammonium bromide|0
    mixed with isopropanol|0
    itching|0
    redness|0
    urticaria|0
    occupational asthma|0
    mild dyspnea|0
    facial erythematous|0
    pruritic eruption|0
    localized edema|0
    papular eruption|0
    recurrent episodes of dermatitis|0
    chest tightness|0
    dyspnea|0
    rhinorrhea|0
    paroxysmal sneezing|0
    non-productive cough|0
    wheezing|0
    secondary infection|0
    hand dermatitis|0
    urticaria of forearms|0
    rhinitis|0
    contact dermatitis|0
    allergy to aspirin|0
    anaphylactic reaction during specific inhalation challenge test|0

<|eot_id|>