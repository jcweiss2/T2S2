67 years old | 0
male | 0
admitted to the hospital | 0
hypertension | -6720
degenerative joint disease | -6720
bilateral knee replacement | -6720
substance abuse | -6720
trauma to face and chest wall | -24
lightheadedness | 0
fatigue | 0
leukocytosis | 0
hemoglobin of 10.2 g | 0
venous lactic acid of 2.4 mol/l | 0
intramuscular and subpectoral hematoma | 0
extrapleural extension into the chest | 0
acute right second through fifth anterior rib fractures | 0
bilateral lower lobe bronchopneumonia | 0
blood cultures obtained | 0
started on empiric antibiotics with intravenous piperacillin–tazobactam | 0
afebrile | 0
hypotensive | 0
admitted to intensive care unit | 0
suspected septic shock | 0
initiation of vasopressors | 0
antibiotics broadened to intravenous vancomycin, cefepime and metronidazole | 48
repeat blood, urine and sputum cultures obtained | 48
sputum cultures grew methicillin-resistant Staphylococcus aureus | 96
antibiotics narrowed to intravenous vancomycin | 96
left knee pain | 120
notable swelling on physical exam | 120
concern for infection of prosthetic knee joint | 120
sterile left knee aspiration | 120
synovial fluid cloudy, amber colored | 120
white blood cells of 9.28 × 10^3/mcL | 120
calcium pyrophosphate crystals | 120
complete washout and debridement of the joint | 144
retention of prosthesis | 144
infected knee with purulence | 144
antibiotic regimen transitioned to intravenous cefazolin | 168
cultures from infected area obtained | 168
joint specimen, tissue specimen and fluid specimen cultured | 168
C. bifermentans grew in two sets of cultures | 264
antibiotic regimen transitioned to intravenous ampicillin–sulbactam | 264
contrast computerized tomography scan of abdomen | 264
human immunodeficiency virus screening | 264
discharged to rehabilitation facility | 384
referral to gastroenterology for outpatient colonoscopy | 384
follow-up with internal medicine | 744
recovered full range of motion of left knee | 744
no signs of lingering joint or systemic infection | 744
taking Augmentin | 744
reported medication adherence | 744
had not yet opted to undergo colonoscopy | 744