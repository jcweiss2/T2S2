17 years old | 0
    female | 0
    admitted to a tertiary medical pediatric gastroenterology unit | 0
    abdominal pain | 0
    fever | 0
    severe sideropenic anemia | 0
    hemoglobin level of 70 g/L | 0
    ferritin value of 9 µg/L | 0
    diarrhea | 0
    diagnosed with ulcerative colitis (pancolitis, E4 localization, Mayo score 2) | 0
    treated with mesalamine | 0
    symptoms improved | 0
    laboratory results improved | 0
    discharged home | 168
    well for the first 9 days | -216
    developed fever (up to 38.7℃) | -216
    sore throat | -216
    right neck swelling | -216
    tenderness | -216
    Group A streptococcal rapid antigen test (negative) | -216
    diagnosed with viral pharyngitis | -216
    symptoms worsened | -240
    neck swelling enlarged | -240
    pain became severe (could not move head) | -240
    came to emergency department | -264
    physical examination revealed right sided supraclavicular very painful edema | -264
    reduced neck movement | -264
    no skin changes | -264
    red tonsils without exudate | -264
    spleen palpable 1 cm below left costal margin | -264
    normal clinical examination (rest) | -264
    unremarkable family history for chronic illness | -264
    elevated leukocytes | -264
    elevated platelets count | -264
    elevated inflammatory markers | -264
    coagulation test results slightly out of reference range | -264
    neck ultrasound revealed complete thrombosis of right external and IJVs (5 cm) | -264
    thrombus within right subclavian vein | -264
    neck MRI | -264
    MRI venography performed | -264
    thrombosis of right subclavian vein | -264
    thrombosis of right jugular veins | -264
    thrombosis of truncus brachiocephalicus | -264
    partial thrombosis of right sigmoid | -264
    partial thrombosis of transverse sinus | -264
    chest ultrasound revealed bilateral pleural effusion | -264
    heart ultrasound revealed apical pericardial effusion | -264
    normal heart contractility | -264
    diagnosed with Lemierre syndrome | -264
    transported to intensive care unit | -264
    treated with intravenous antibiotics (ceftriaxone and clindamycin for first 5 days) | -264
    treated with clindamycin for following 9 days | -264
    received subcutaneous low-molecular-weight heparin | -264
    heparin titrated based on anti-Xa activity | -264
    paired blood cultures taken | -264
    throat swabs taken | -264
    no pathogen isolated | -264
    afebrile after 72 hours of antibiotic treatment | -192
    comprehensive thrombophilia testing | -192
    factor V Leiden normal | -192
    protein C normal | -192
    protein S normal | -192
    factor VIII normal | -192
    antithrombin III normal | -192
    antinuclear antibodies negative | -192
    anticardiolipin antibodies negative | -192
    homocysteine levels normal | -192
    F2 gene mutation G20210A c. *97G>A not found | -192
    FV Leiden c.1691G>A, p. Arg534GIn mutation not found | -192
    discharged from hospital | -96
    continue anticoagulation therapy at home | -96
    low-molecular-weight heparin replaced by apixaban after 9 months | 2160
    subsequent follow-ups showed amelioration of neck edema | 2160
    neck ultrasound confirmed regression of thrombosis | 2160
    color Doppler confirmed recanalization of jugular vein | 2160
    UC in clinical remission | 2160
    Paediatric Ulcerative Colitis Activity Index was 0 | 2160
    normal calprotectin levels | 2160
    no signs of anemia | 2160
    <|eot_id|>
    