18 year old male | 0
admitted to hospital | 0
fever | -72
shortness of breath | -72
chest X-ray bilateral interstitial infiltrates | 0
empirical therapy for community-acquired pneumonia | 0
weight loss | -2160
lethargy | -2160
swallowing difficulties | -2160
hypoxic respiratory failure | 0
intubated | 0
CT scan widespread nodular infiltrates | 24
mediastinal abscess | 24
septic | 0
high-dose vasopressors | 0
hemodynamic instability resolved | 72
lung-protective mechanical ventilation | 0
intermittent prone positioning | 0
negative bronchoalveolar lavage cultures | 0
negative viral PCR assays | 0
negative Ziehl-Neelsen staining | 0
indeterminable IGRA for tuberculosis | 0
negative infectious work-up | 0
negative malignant work-up | 0
negative immunological work-up | 0
expanded antibiotic therapy | 0
empirical corticosteroids | 0
empirical immunoglobulins | 0
transbronchial biopsies | 432
bilateral tension pneumothoraces | 432
pneumopericardium | 432
subcutaneous emphysema | 432
pleural drainage | 432
critical oxygenation | 432
veno-venous ECMO therapy | 432
acid-fast bacilli in transbronchial biopsies | 432
tuberculosis treatment initiation | 432
rifampicin | 432
isoniazid | 432
ethambutol | 432
pyrazinamide | 432
confirmed miliary tuberculosis | 624
Mycobacterium tuberculosis growth in admission samples | 624
bacteria in tracheal aspirate | 624
bacteria in urine | 624
bacteria in cerebrospinal fluid | 624
granulomas in bone marrow | 624
granulomas in liver | 624
granulomas in lung | 624
susceptible to first-line agents | 624
dysphagia related to mediastinal tuberculosis | 624
mediastinal abscess related to tuberculosis | 624
multiple lung bullae | 432
persistent pneumothoraces | 432
subtherapeutic isoniazid levels | 432
subtherapeutic rifampicin levels | 432
escalated doses | 432
intravenous administration | 432
acid-fast bacilli in tracheal aspirates | 672
multi-resistant Pseudomonas aeruginosa | 672
Stenotrophomonas maltophilia | 672
eradicated with inhaled colistin | 672
eradicated with inhaled tobramycin | 672
eradicated with intravenous amikacin | 672
eradicated with meropenem | 672
eradicated with ceftazidime/avibactam | 672
low amikacin levels | 672
signs of recovery | 1080
increasing lung compliance | 1080
lung re-expansion | 1080
weaned from ECMO | 1200
thrombocytopenia | 1200
minor bleedings | 1200
sensory symptoms in lower limbs | 1200
stayed in ICU for 76 days | 1824
rehabilitation | 2160
resumed activities | 2160
resumed sports | 2160
