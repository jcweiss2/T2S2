56 years old | 0
male | 0
diagnosed with nodular sclerosing cluster of differentiation (CD) 30+, CD15+ HL | -8760
stage IV disease | -8760
diffuse involvement of the lymph nodes | -8760
diffuse involvement of the bone marrow | -8760
diffuse involvement of the liver | -8760
power-injectable port inserted | -8400
six cycles of ABVD chemotherapy | -8400
partial response | -6720
two other lines of chemotherapy | -6720
poor clinical response | -6720
evaluated for autologous hematopoietic stem cell transplant (HSCT) | 0
pretransplant transthoracic echocardiogram (TTE) | 0
2.2 × 1.8 cm RA mass | 0
normal cardiac function | 0
sent to the emergency room | 0
hemodynamically stable | 0
asymptomatic | 0
physical examination unremarkable | 0
leukocytosis of 15,000 cells/mm3 | 0
hemoglobin of 7.5 mg/dL | 0
normal platelet count | 0
computed tomography (CT) imaging | 24
RA mass with unclear etiology | 24
extra-cardiac findings consistent with diffuse HL | 24
transesophageal echocardiogram (TEE) | 48
RA mass attached to the posterior atrial wall | 48
RA mass attached to the central venous catheter (CVC) | 48
cardiac magnetic resonance imaging (CMR) | 72
no enhancement of the RA mass with gadolinium contrast injection | 72
diagnosis of CRAT | 72
heparin for anticoagulation | 72
cardiac thoracic surgery consulted | 72
possible thrombectomy | 72
fever | 96
hypotension | 96
pancytopenia | 96
managed in the intensive care unit | 96
broad spectrum antibiotics | 96
vasopressors | 96
rapidly deteriorated | 120
succumbed to the disease | 120