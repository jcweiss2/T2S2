60 years old | 0
male | 0
alcoholic | 0
admitted to medical casualty | 0
self-induced vomiting | -72
cough with expectoration | -72
hiccups | -72
altered behavior | -72
dizziness | -72
fall in washroom | -24
past history of admission for symptomatic hyponatremia | -216
serum sodium: 123 mEq L−1 | -216
serum potassium: 4.9 mEq L−1 | -216
managed with 3% hypertonic saline | -216
serum sodium: 129 mEq L−1 | -204
discharged home | -144
presented to neurology department | -120
complain of imbalance | -120
slurred speech | -120
drowsiness | -120
fever | -120
cough | -120
Glasgow Coma Scale (GCS) E4V1M1 | -120
hypertonic bilateral upper and lower limbs | -120
hyperreflexia | -120
bilateral extensor plantar | -120
nystagmus | -120
restricted extraocular muscle movements | -120
shifted to intensive care unit (ICU) | -120
intubated | -120
antibiotics | -120
antimalarials | -120
stress ulcer prophylaxis | -120
deep venous thrombosis prophylaxis | -120
injection thiamine | -120
intravenous fluids | -120
differential diagnosis of CPM | -120
extrapontine myelinolysis | -120
subdural hemorrhage | -120
associated sepsis with delirium | -120
hepatic encephalopathy | -120
Wernicke–Korsakoff syndrome | -120
autoimmune encephalitis | -120
routine blood, urine and radiological investigations | -120
Magnetic resonance imaging (MRI) brain | -120
hyperintensities in the central part of pons | -120
relative sparing of peripheral pons | -120
bilateral corticospinal tracts | -120
transverse pontine fibers | -120
trident pattern in the upper pons | -120
involvement of tegmentum of midbrain | -120
bilateral thalamic | -120
globus pallidus | -120
tracheostomy | -112
weaned from ventilator | -105
put on T-piece | -105
multidisciplinary approach | -105
neurology | -105
ophthalmology | -105
psychiatry | -105
physical medicine rehabilitation | -105
medicine | -105
conscious oriented (GCS – E4VTM6) | -60
vitals stable | -60
rigidity and hyperreflexia | -60
shifted from ICU | -30
followed up until discharge | 0
physical rehabilitation | 0
able to walk with support | 60