69 years old | 0
male | 0
admitted to the hospital | 0
fever | -20
altered consciousness | -20
prostate cancer | -2520
chemotherapy | -2520
prednisolone | -2520
proton pump inhibitor | -2520
Cabazitaxel Acetonate | -2520
Glasgow Coma Scale E3V3M5 | 0
temperature 40.6°C | 0
blood pressure 142/80 mmHg | 0
pulse rate 126/min | 0
respiratory rate 30/min | 0
percutaneous oxygen saturation 98% | 0
conjunctive pale | 0
no icterus | 0
no abnormal findings in chest | 0
median surgical scar | 0
mildly edematous lower extremities | 0
no palpable surface lymph nodes | 0
no rash | 0
no neck stiffness | 0
highly elevated white blood cell count | 0
anemia | 0
cytoplasmic vacuolation of white blood cells | 0
anisocytosis | 0
spherocytes | 0
high lactate dehydrogenase | 0
high creatine kinase | 0
severe hemolysis | 0
piperacillin/tazobactam | 0
blood pressure dropped | 2
cardiopulmonary arrest | 2
cardiopulmonary resuscitation | 2
circulation recovered | 2
blood cell transfusion | 2
vasopressors | 2
hypothermia treatment | 2
hemolysis worsened | 2
difficulty maintaining blood pressure | 2
death | 30
Clostridium perfringens detected | 30
Gram-positive bacilli identified | 30
bacilli phagocytized by white blood cells | 30
Clostridium perfringens isolate serotype TW62 | 30
non-enterotoxin producing | 30
α toxin-producing type A | 30
susceptible to penicillins | 30
susceptible to β-lactams | 30