73 years old | 0
male | 0
medical history of multiple thromboses | 0
deep vein thrombosis in 1995 | -172440
deep vein thrombosis in 2011 | -172440
pulmonary embolism in 1995 | -172440
pulmonary embolism in 2004 | -172440
presented in 2013 | 0
two consecutive acute coronary syndromes within 1-month interval | -720
continuous anticoagulation with vitamin K antagonists (fluindione) | 0
admitted to cardiology department | -720
acute thoracic pain | -720
electrocardiogram evidenced inferior Q waves with ST elevation | -720
echography revealed antero-inferior akinesia | -720
serum troponins not quantified | -720
transferred for coronarography | -720
coronary catheterization revealed intraluminal thrombus in right coronary artery | -720
balloon angioplasty performed | -720
no stent inserted due to unexplained fever | -720
antiplatelet therapy with acetylsalicylic acid and clopidogrel added | -720
presented again with typical acute chest pain | -672
electrocardiogram evidenced inferior Q waves | -672
echography found antero-inferior akinesia | -672
ultrasensitive troponins elevated (560 ng/L) | -672
new coronary catheterization performed | -672
evidenced thrombosis in right coronary artery | -672
asymptomatic incomplete intraluminal obstruction of circumflex artery | -672
angioplasty performed without vascular stenting | -672
persistent fever since 2 months | -1440
marked inflammatory syndrome | 0
additional investigations performed | 0
fatigue | 0
signs of anemia | 0
hemoglobin level 90 g/L | 0
reticulocytes 52 × 10^9/L | 0
white blood cells 6.6 × 10^9/L | 0
normal differential | 0
platelet count 52 × 10^9/L | 0
C-reactive protein (CRP) level 147 mg/L | 0
tests for infectious diseases negative | 0
tests for systemic inflammatory diseases negative | 0
tests for vasculitis negative | 0
serum haptoglobin decreased | 0
lactate dehydrogenase (LDH) markedly elevated | 0
direct antiglobulin test negative | 0
computerized tomography (CT) scan showed thrombosis of hepatic vein | 0
multiple thromboses despite anticoagulation | 0
signs of hemolysis | 0
flow cytometry test disclosed big-sized PNH clone | 0
neutrophils lacking CD66b, CD16, CD24 antigens | 0
monocytes lacking CD24 antigen | 0
BM smears normocellular | 0
mild signs of dysmegacaryocytopoiesis | 0
no excess blasts (2%) | 0
karyotype normal | 0
diagnosis of classical PNH | 0
presence of fever | 0
inflammatory syndrome | 0
increased risk of severe infections | 0
decision to start eculizumab postponed | 0
acute abdomen | 0
hypotension | 0
functional renal insufficiency | 0
admitted to intensive care unit | 0
CT scan not helpful | 0
surgical exploration of abdomen performed | 0
no major abnormality found | 0
acute abdomen linked to multiple thromboses of small abdominal vessels | 0
treatment with eculizumab started | 0
prophylaxis including vaccination against meningococcal and pneumococcal infection | 0
penicillin V therapy | 0
anticoagulation maintained | 0
antiplatelet treatments maintained | 0
fever resolved | 0
abdominal pain resolved | 0
inflammatory syndrome resolved | 0
LDH level returned to normal | 0
required repeated transfusions of red blood cell packs | 0
severe thrombocytopenia occurred | 672
no signs of hemolysis | 672
BM examination showed normocellular BM | 672
dysplasia of 3 myeloid lineages | 672
11% blasts | 672
diagnosis of refractory anemia with excess blast-2 | 672
BM karyotype normal | 672
vitamin K antagonists stopped | 672
antiplatelet treatment maintained | 672
platelet transfusions performed | 672
red blood cell transfusions performed | 672
only transient improvement | 672
not eligible for BM transplantation | 672
hypomethylating treatment with 53-azacytidine (AZA) added | 672
cytopenias remained unchanged after 2 cycles | 672
admitted to intensive care unit | 1344
septic shock due to Aeromonas veronii infection | 1344
implantable chamber infection | 1344
multiorgan failure | 1344
death despite broad-spectrum antibiotics and vasopressor medication | 1344
