55 years old | 0
male | 0
African American | 0
chronic pulmonary obstructive disease | -175200
alcohol dependence | -175200
alcohol withdrawal symptoms | 0
headache | 0
tremors | 0
sweating | 0
denied liver disease | 0
denied sleep disturbances | 0
denied memory changes | 0
denied seizures | 0
anxious | 0
tremulous | 0
slow and delayed response to questions | 0
unsteady gait | 0
scleral icterus | 0
skin icterus | 0
gynecomastia | 0
bibasilar crackles | 0
liver edge palpable 3cm below costal margin | 0
asterixis | 0
nail clubbing | 0
non-pitting edema of the legs | 0
macrocytic anemia | 0
hemoglobin 11.3 g/dl | 0
Mean Corpuscular Volume 101.8 fL | 0
platelet count 83,000/μL | 0
total protein 8.2 g/dL | 0
albumin 2.8 g/dL | 0
total Bilirubin 3.9 mg/dL | 0
AST 69 U/L | 0
ALT 36 U/L | 0
ammonia level 124 mcg/dl | 0
INR 1.6 | 0
computed tomography of the abdomen showing early cirrhosis | 0
admitted to the hospital | 0
diagnosis of alcohol withdrawal | 0
possible hepatic encephalopathy | 0
chlordiazepoxide-based alcohol withdrawal protocol started | 0
tapering doses | 0
lactulose for hepatic encephalopathy | 0
300 mg chlordiazepoxide over 9 days | 0
good control of withdrawal symptoms | 0
mental status deteriorated | 216
upgraded to intensive care unit | 216
urine drug screen positive for benzodiazepines | 216
repeat ammonia level 121 mcg/dl | 216
septic work-up unremarkable | 216
diagnosis of benzodiazepine-induced hepatic encephalopathy | 216
flumazenil 1mg IV given | 216
significant improvement of mental status | 216
effect short-lived (20 minutes) | 216
mental status deteriorated again | 216
repeated single doses of flumazenil failed | 216
flumazenil drip started at 0.25 mg/hour | 216
persistent nausea | 216
treated with ondansetron | 216
flumazenil well tolerated | 216
attempts to decrease infusion rate resulted in deterioration | 216
repeated urine benzodiazepine testing positive three times | 216
flumazenil maintained for 28 days | 216
flumazenil tapered off successfully | 672
mental status returned to normal | 672
repeat urine benzodiazepine test negative | 672
discharged home | 672
