38 years old | 0 | 0 
female | 0 | 0 
13th week of pregnancy | 0 | 0 
admitted to the emergency room | 0 | 0 
abdominal discomfort | -24 | 0 
nausea | -24 | 0 
vomiting | -24 | 0 
no fever | -24 | 0 
no vaginal discharge | -24 | 0 
evaluated in the Obstetric Emergency Department | 0 | 0 
discharged home | 0 | 0 
persistent abdominal pain | 144 | 144 
nausea | 144 | 144 
vomiting | 144 | 144 
tachycardic | 144 | 144 
diffuse abdominal pain | 144 | 144 
guarding on the right quadrants | 144 | 144 
neutrophilia | 144 | 144 
low prothrombinemia | 144 | 144 
acute renal failure | 144 | 144 
high procalcitonin | 144 | 144 
high c-reactive protein | 144 | 144 
abdominal ultrasound | 144 | 144 
moderate fluid in all quadrants | 144 | 144 
good foetal vitality | 144 | 144 
surgical consultation | 144 | 144 
hypotension | 144 | 144 
general abdominal guarding | 144 | 144 
hyperlacticaemia | 144 | 144 
hypokalaemia | 144 | 144 
hyperglycaemia | 144 | 144 
septic shock with an abdominal source | 144 | 144 
emergency exploratory laparotomy | 144 | 144 
generalised purulent peritonitis | 144 | 144 
perforated acute appendicitis | 144 | 144 
appendicectomy | 144 | 144 
abdominal washing | 144 | 144 
laparostomy | 144 | 144 
admitted to the Intensive Care Unit | 144 | 144 
septic shock | 144 | 144 
need for vasopressor therapy | 144 | 144 
dialysis | 144 | 144 
intravenous piperacillin-tazobactam antibiotherapy | 144 | 192 
laparostomy revision | 192 | 192 
marked bowel oedema | 192 | 192 
bowel distention | 192 | 192 
mild intraabdominal soiling | 192 | 192 
peritoneal lavage | 192 | 192 
new laparostomy with progressive closure technique | 192 | 192 
recovered progressively | 192 | 336 
surgical revision | 336 | 336 
abdominal cavity primary closed | 336 | 336 
antibiotherapy adjusted | 336 | 336 
piperacillin-tazobactam suspended | 336 | 336 
amoxicillin with clavulanic acid started | 336 | 336 
transferred to the obstetrics ward | 432 | 432 
discharged home | 504 | 504 
elective caesarean section | 1008 | 1008 
gave birth to a healthy child | 1008 | 1008 
ventral hernia | 1344 | 1344 
incisional hernia correction | 1344 | 1344 
child thriving without neurological or other impairments | 1344 | 1344