27 years old | 0
Gravida 4 | 0
Para 3 | 0
17 weeks’ gestation | 0
fever | -72
dry cough | -72
shortness of breath | -72
COVID-19 diagnosis | 0
SARS-CoV-2 positive | 0
first COVID-19 vaccine dose | -264
admission | 0
3-day history of fever | -72
3-day history of shortness of breath | -72
3-day history of dry cough | -72
conscious | 0
stable hemodynamic parameters | 0
body temperature 39.0°C | 0
SpO2 84% | 0
FiO2 60% |4 0
respiratory rate 30 breaths/minute | 0
blood pressure 130/80 mmHg | 0
pulse 125 beats per minute | 0
transferred to ICU | 0
severe ARDS | 0
increased AST | 0
increased ALT | 0
increased CRP | 0
increased LDH | 0
increased ferritin | 0
severe hypoxia | 0
moderate hypercapnia | 0
normal renal function | 0
normal coagulation tests | 0
bilateral alveolar infiltration | 0
live fetus | 0
sinus tachycardia | 0
HFNC | 0
HFNC FiO2 100% | 0
HFNC flow 60 l/min | 0
BiPAP | 24
BiPAP EPAP 8 cmH2O | 24
BiPAP IPAP 13 cm | 24
BiPAP FiO2 100% | 24
intubation | 96
IMV | 96
IMV VC mode | 96
IMV RR 20/min | 96
IMV PEEP 10 cmH2O | 96
IMV Vt 300 ml | 96
IMV I/E ratio 1/2 | 96
IMV FiO2 100% | 96
dexamethasone 6 mg/day | 0
enoxaparin 60 mg twice daily | 0
clopidogrel 75 mg daily | 0
ceftriaxone 2 g/day | 0
multivitamin | 0
magnesium | 0
zinc | 0
enteral feeding | 0
parenteral nutrition | 0
TPE | 144
fever 39°C | 288
antibiotic change to meropenem | 288
antibiotic change to linezolid | 288
extubation | 312
CPAP | 312
CPAP FiO2 60% | 312
HFNC | 360
HFNC flow reduced | 360
FiO2 reduced | 360
oxygen support discontinued | 504
discharged | 648
healthy 20-week gestational fetus | 648
