75 years old | 0
    male | 0
    acute ischemic stroke due to thrombotic occlusion of the M1 segment of the left A. cerebri media | 0
    coronary angiography | -384
    intervention for non-ST-elevation myocardial infarction | -384
    right-sided hemiplegia | 0
    mechanical thrombectomy | 0
    aspiration pneumonia | 0
    piperacillin/tazobactam | -168
    recurrent sinus bradycardia | 0
    intermittent ventricular escape rhythm | 0
    third-degree sinoatrial block | 0
    2-chamber pacemaker implantation | -96
    povidone-iodine solution | -96
    discharge to neurological rehabilitation facility | -72
    readmitted | 168
    fever | 168
    hyperthermic, reddened pacemaker incision site | 168
    leucocytosis | 168
    elevated C-reactive protein | 168
    blood cultures collected | 168
    ampicillin/sulbactam | 168
    pacemaker pocket infection suspected | 168
    system extraction | 168
    intraprocedural inspection of pacemaker pocket | 168
    no pus | 168
    old hematoma | 168
    swab samples of pacemaker and pocket | 168
    explanted leads retained for microbiological diagnostic | 168
    transferred to intensive care unit | 168
    persisting sinoatrial block | 168
    transesophageal echocardiography | 168
    mobile vegetation from the right atrium to the superior vena cava | 168
    presence of ghosts | 168
    device-associated endocarditis | 168
    blood cultures positive for C. difficile | 168
    pacemaker samples positive for C. difficile | 168
    stool sample obtained | 168
    toxigenic C. difficile strains | 168
    nontoxigenic isolate | 168
    antimicrobial testing | 168
    ribotyping | 168
    minimum inhibitory concentration testing | 168
    genotyping detected RT014 | 168
    clonality confirmed by whole-genome sequencing | 168
    RT020 detected in stool | 168
    unclassified nontoxigenic isolate | 168
    no signs of previous C. difficile infection | 168
    no history of infectious diarrhea | 168
    no contact with infectious diarrhea | 168
    abdominal ultrasound revealed no pathologies | 168
    intravenous vancomycin | 168
    oral metronidazole | 168
    normalization of leukocytes | 168
    normalization of C-reactive protein | 168
    liver enzymes increased | 168
    oral antibiotic therapy switched to vancomycin | 168
    repeated blood cultures negative | 168
    stool samples during therapy negative | 168
    transferred back to rehabilitation facility | 168
    intravenous vancomycin continued | 168
    oral vancomycin for decolonization | 168
    tapering regime | 168
    readmitted for pacemaker reimplantation | 168
    TEE revealed elimination of vegetations | 168
    blood cultures negative | 168
    skin swabs negative | 168
    colonoscopy showed noninflamed sigmoid diverticula | 168
    toxigenic C. difficile isolated from stool | 168
    RT005 detected | 168
    intravenous vancomycin treatment | 168
    reimplantation of pacemaker | 168
    oral vancomycin tapering regime | 168
    follow-up visit | 168
    normal pacemaker function | 168
    no sign of infection | 168
    