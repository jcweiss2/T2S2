40 years old | 0
male | 0
admitted to the Haematology Clinic | 0
recurrent ALL | 0
allogeneic bone marrow transplantation | 0
extensive maculopapular skin rash | -84
GVHD | -84
systemic corticosteroids | -84
treatment with systemic steroids | -84
gradually reducing regime | -84
monitored as an outpatient | -84
unexplained fever | -360
admitted to the Haematology Clinic | -360
treatment with intravenous antibiotics | -360
apyrexial | -360
non-specific abdominal disturbance | -24
acute onset of depressive effect | -24
low mood | -24
stopped eating | -24
severely disturbed night sleep | -24
stopped communicating | -24
reluctant to see his wife and children | -24
reduced motivation | -24
reduced energy | -24
fear of death | -24
abdominal CT scans | -24
no specific cause for abdominal disturbance | -24
ALL in remission | -24
deteriorating mood | -24
consultation by the Liaison Psychiatric team | -24
profoundly low mood | -14
anhedonia | -14
reduced energy | -14
severely disturbed sleep | -14
reduced appetite | -14
weight loss | -14
hopelessness | -14
helplessness | -14
passive death wishes | -14
suicidal thoughts | -14
well-orientated | -14
MMSE score 30/30 | -14
severe depressive episode | -14
HAM-D score 25 | -14
treatment with duloxetine | -14
duloxetine titrated up to 60 mg daily | -7
partial response | -7
death wishes subsided | -7
low mood | -7
biological symptoms of depression | -7
HAM-D score 17 | -7
vague abdominal disturbance | -7
localized abdominal pain | 0
intestinal leakage | 0
explorative laparotomy | 0
sepsis | 2
death | 2