23 years old | 0
    male | 0
    methicillin-resistant Staphylococcus aureus (MRSA) impetigo at the forearm | -8760
    right tibia fracture | -8760
    intramedullary fixation (IMN) | -8760
    interlocking screws removed due to skin irritation and pain | -672
    redness at the surgical site | -552
    swelling at the surgical site | -552
    stitch abscess | -552
    MRSA positive cultures from the surgical site | -552
    oral antibiotic treatment | -552
    fever | -216
    right groin pain | -216
    viral infection | -216
    systemic fever (39 °C) | -168
    myalgia | -168
    difficult and painful ambulation | -168
    right forearm cellulitis | -168
    right sudden onset uveitis | -168
    systemic rash | -168
    right hip lymphadenopathy | -168
    increased CRP (30 mg/dL) | 0
    increased WBC (14,000) | 0
    elevated hepatic enzymes | 0
    elevated lactic dehydrogenase (LDH) | 0
    elevated creatine phosphokinase (CPK) | 0
    unremarkable radiograph of both hips | 0
    IV antibiotics against MRSA | 0
    hemodynamic deterioration | 0
    fulminant MRSA sepsis | 0
    admitted to the intensive care unit (ICU) | 0
    ultrasound-guided drainage | 0
    enlargement of the abscesses diameter | 72
    persistent fever | 72
    CRP level of 36 mg/dL | 72
    WBC count of 20,000 | 72
    surgical intervention | 72
    combined approach of Smith-Peterson and modified Stoppa | 72
    general condition improving after surgery | 72
    less frequent fever spikes | 72
    decrease in CRP | 504
    decrease in WBC | 504
    almost complete recovery | 1344
    ambulate normally without pain | 1344
    no functional limitations | 1344
    returned to daily activities | 1344