50 years old | 0
male | 0
admitted to the hospital | 0
urinary lithiasis history | 0
left colic pain | 0
mild hyperpyrexia (37.5°C) | 0
left renal shockwave lithotripsy (SWL) in 1990 | -175200
right pyelotomy for phosphatic/oxalate stones in 1998 | -175200
parathyroidectomy in 2000 | -175200
urinalysis revealing mixed low burden microbial germs | 0
non-contrast medium CT scan (NCCT) finding bilateral lithiasis | 0
left kidney lithiasis (1.2×2.7 cm, 1400 HU) | 0
right lower pole lithiasis (1.5×1.4 cm, 1350 HU) | 0
treated with left ureteral stenting | 0
antibiotic therapy (Meropenem and Gentamicin) | 0
referred for elective left endoscopic combined intrarenal surgery (ECIRS) | 0
pre-operative urinalysis negative | 0
Amoxicillin + clavulanic acid administered | 0
Valdivia Galdakao position during procedure | 0
3 unsuccessful renal puncture attempts | 0
converted to f;URS laser lithotripsy | 0
100WATT Holmium Quanta System used | 0
ureteral access sheath 10/12FR | 0
1 hour operative time | 0
procedure stopped | 0
deferred to second look | 0
fever (>38°C) on first day | 24
blood cultures performed | 24
empirical antibiotic therapy with Tazobactam and Teicoplanin administered | 24
CT scan showing pyelonephritis with no abscesses or perirenal haematoma | 24
antibiotic therapy modified based on Pseudomonas Aeruginosa in blood cultures | 24
Meropenem and Linezolid administered | 24
admitted to Intensive Care Unit due to haemodynamically unstable situation | 24
tachycardia | 24
hypotension | 24
thoracic/abdomen CT scan performed at 4 days post-surgery | 96
pulmonary septic emboli | 96
bilateral pleural effusion | 96
left renal abscess | 96
CT-guided renal drain placed | 96
ureteral stent replaced | 96
continued fever on tenth day | 240
CT scan showing no change from previous control | 240
multidisciplinary counselling with anesthesiologists, radiologists, and infectivologists | 240
counselled for left open nephrectomy | 240
left open nephrectomy performed | 240
not pyretic on first day post-nephrectomy | 264
decreasing inflammation indexes | 264
discharged on 7 days post-OP | 336
histological examination showing multifocal Xanthogranulomatous pyelonephritis | 336
- 50 years old | 0
7 male | 0
left renal shockwave lithotripsy (SWL) in 1990 | -262800
right pyelotomy for phosphatic/oxalate stones in 1998 | -192720
converted to f-URS laser lithotripsy | 0
no abscesses | 24
no perirenal haematoma | 24
discharged on 7 days post-OP | 408
histological examination showing multifocal Xanthogranulomatous pyelonephritis | 408
