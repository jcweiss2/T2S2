breast cancer | 0
chemotherapy | 0
radiation to the chest | 0
severe aortic stenosis | 0
concomitant coronary artery disease | 0
90% occlusion of the left anterior descending artery | 0
tissue aortic valve replacement | 0
saphenous vein graft bypass to the left anterior descending artery | 0
induction of anesthesia | 0
intubation | 0
dissection of the left internal mammary artery | 0
use of the greater saphenous vein | 0
discontinuation of cardiopulmonary bypass | 0
decline in cerebral head saturations | -0.5
use of vasopressors | -0.5
extubation | 2
persistent lactic acidosis | 2
high-dose vasopressor support | 2
mixed cardiogenic and vasoplegic shock | 2
lethargy | 15
leftward gaze | 15
right upper extremity weakness | 15
resolution of symptoms | 15.25
progressive bilateral tongue ecchymoses | 15
tongue numbness | 15
dysgeusia | 15
CT scan of the head | 15
CT angiogram of the brain and neck | 15
mild calcification at the bifurcation of the right common carotid artery | 15
50% focal stenosis of the distal left common carotid artery | 15
complete occlusion of the right lingual artery | 15
mild distal collateral flow | 15
multifocal irregularities of the left lingual artery | 15
normal postoperative platelet count | 15
normal prothrombin time | 15
normal international normalized ratio | 15
normal fibrinogen | 15
no prior history of known vasculitic disease | 15
normal ADAMTS13 inhibitor screen | 15
volume resuscitation with crystalloid and colloid | 15
low-dose epinephrine | 15
high-dose norepinephrine | 15
high-dose vasopressin | 15
improvement of systemic vascular resistance | 17
otolaryngology service consultation | 17
serial examinations of the patient’s tongue | 17
evaluation with multiple flexible bronchoscopes | 17
persistent tongue numbness | 17
persistent dysgeusia | 17
supportive therapy | 17
improvement of examination and symptoms | 48
return of tongue sensation and taste to baseline | 72
transient ischemic attack | 15 
no shortness of breath | 0
denies chest pain | 0