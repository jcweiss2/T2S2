26 years old | 0
male | 0
admitted to the hospital | 0
febrile illness | -168
involuntary, hyperkinetic movements | -168
weakness of both upper and lower limbs | -168
excessive sweating | -168
insomnia | -168
autonomic dysfunction | -168
behavioral abnormalities | -168
auditory hallucinations | -168
resting pulse rate above 110 beats/min | 0
elevated blood pressure above 160/100 mm of Hg | 0
wasting of muscles of all four limbs | 0
hypokalemia | 0
hypoproteinemia | 0
low total protein | 0
low albumin | 0
low globulin | 0
positive serum anti-CASPR2 antibody | 0
treatment with high-dose steroids | 0
treatment with intravenous immune globulin (IVIG) | 0
no improvement with high-dose steroids and IVIG | 336
decision to carry out therapeutic plasma exchange (TPE) | 336
placement of double-lumen femoral line | 336
establishment of peripheral venous access | 336
correction of potassium levels | 336
start of TPE | 336
use of FFP and saline as replacement fluid | 336
calculation of total plasma volume | 336
exchange of 100% of total plasma volume | 336
persistent hyperkinetic movements | 336
obstruction of femoral line and tubing | 336
restraint of limbs | 336
administration of tablet methyl prednisolone | 336
administration of tablet clonazepam | 336
allergic reaction to FFP | 336
treatment with antihistamines | 336
premedication with antihistamines | 432
elevated blood pressure above 160/100 mm of Hg | 432
tachycardia above 110 bpm | 432
transfusion of four units of FFP | 432
enhancement of FFP support | 432
rectification of total serum proteins | 432
clinical signs of improvement | 528
ability to sit with support | 528
ability to eat and walk with support | 720
mild, occasional hyperkinetic movements | 720
improvement of autonomic dysfunction | 720
normalization of pulse rate | 720
normalization of blood pressure | 720
subsidence of excessive sweating | 720
subsidence of restlessness | 720
subsidence of insomnia | 720
absence of behavioral abnormalities | 720
decline of anti-CASPR2 antibodies | 720
treatment with oral prednisolone | 720
remission | 2160