36 years old | 0
male | 0
butcher | 0
history of smoking | 0
cannabinoid consumption | 0
admitted to the hospital | 0
severe headache | 0
fever | 0
dysarthria | 0
confusion | 0
psychomotor agitation | 0
Glasgow Coma Scale of 13 | 0
nuchal rigidity | 0
respiratory distress | 0
desaturation | 0
diminished breath sounds bilaterally | 0
Brudzinski's sign absent | 0
Kernig's sign absent | 0
Lasegue's sign absent | 0
leukocytosis | 0
neutrophilia | 0
elevated C-reactive protein | 0
thrombocytopenia | 0
renal function unremarkable | 0
hepatic function unremarkable | 0
ionogram unremarkable | 0
serology tests unremarkable | 0
urine toxicology tests negative | 0
cerebral computerized tomography | 0
hydrocephalus in the third ventricle | 0
cerebrospinal fluid analysis | 0
glucose levels of 1mg/dL | 0
protein concentration of 671 mg/dL | 0
white blood cell count of 104cells/mm3 | 0
cerebrospinal fluid Gram stain with Gram-positive diplococci | 0
acute bacterial meningitis diagnosed | 0
ceftriaxone started | 0
vancomycin started | 0
acyclovir started | 0
dexamethasone started | 0
thiamine supplementation started | 0
SARS-CoV-2 infection positive | 0
sedated | 0
mechanically ventilated | 0
vasopressor support started | 0
intracranial pressure monitored | 0
intracranial hypertension | 0
cerebrospinal fluid drainage through a lumbar drain | 0
seizures | 0
anticonvulsant therapy started | 0
levetiracetam started | 0
cerebrospinal fluid culture positive for Streptococcus suis II | 0
antibiotic therapy administered for 14 days | 0
dexamethasone discontinued after 5 days | 0
improvement in oxygenation | 0
hemodynamic stability | 0
sedation stopped | 0
mechanically ventilated weaned | 0
discharged to a district hospital | 0
complete resolution of symptoms | 0
Streptococcus suis meningitis diagnosed | 0 
working as a butcher without adequate work protection | -672 
frequent contact with the nasal and oral cavity | -672 
no hearing loss | 0 
no focal neurological deficits | 0 
no recurrence of seizures | 0 
no shortness of breath | 0 
no chest pain | 0 
no other risk factors | 0 
no asplenia | 0 
no diabetes mellitus | 0 
no alcoholism | 0 
no malignancy | 0 
no structural heart disease | 0 
no COVID-19 symptoms | 0 
no alterations in other diagnostic exams that suggested COVID-19 disease | 0 
COVID-19 pandemic | -10000 
Streptococcus suis reported in pigs in Portugal | -10000 
limited case reports of infection in humans in Portugal | -10000 
patient consent obtained | 0 
patient consent for publication | 0 
patient understands anonymity cannot be guaranteed | 0 
no conflicts of interest | 0 
no financial support and sponsorship | 0