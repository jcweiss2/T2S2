70 years old | 0
male | 0
type 2 diabetes mellitus | -6720
previous kidney transplantation | -5040
previous kidney transplantation | -336
end-stage renal disease | -6720
focal segmental glomerulosclerosis | -6720
chronic antibody-mediated rejected | -336
admitted to the intensive care unit | 0
distributive shock | 0
vasopressor support | 0
piperacillin-tazobactam | 0
blood cultures bottles grew a non-lactose fermenting gram-negative bacillus | 19
cystoscopy | -96
microscopic hematuria | -96
bilobar prostatic hypertrophy | -96
Pseudomonas aeruginosa | 19
piperacillin-tazobactam dosing | 19
defervesced | 19
normalized hemodynamic parameters | 19
transferred to the ward | 19
oral ciprofloxacin | 19
persistent P. aeruginosa bacteremia | 19
high-dose ceftazidime | 19
persistently bacteremic | 168
no indwelling catheters | 168
no perinephric abscess | 168
no hydronephrosis | 168
no clinical or radiographic evidence of pneumonia | 168
no known cardiac valvulopathy | 168
no arterial aneurysms | 168
delirium | 168
rectal pain | 168
digital rectal examination | 168
enlarged and tender prostate | 168
endorectal ultrasound | 168
prostatomegaly | 168
increased vascularity | 168
multiple prostatic abscesses | 168
ultrasound-guided transrectal needle aspirate | 168
purulent fluid | 168
cultures grew the same phenotypic strain of P. aeruginosa | 168
transurethral resection of the prostate gland | 192
unroofing of prostatic abscess | 192
surgical pathology specimen | 192
sheets of foamy histiocytes | 192
abundant necrotic debris | 192
rare hemosiderin deposition | 192
Auramine-rhodamine and Grocott-Gomori’s methamine silver stains | 192
negative for acid-fast bacilli | 192
negative for fungi | 192
histicocytes did not express cytokeratin AE1/AE3 | 192
immunohistochemistry | 192
excluding the possibility of an epithelial neoplasm | 192
pathologic findings | 192
diagnostic of XG prostatitis | 192
completed 10 days of oral ciprofloxacin | 240
surveillance urine cultures grew Pseudomonas aeruginosa | 240
new lower urinary tract symptoms | 240
6 additional weeks of ciprofloxacin | 240
no significant adverse events | 480
follow-up assessment | 720
clinically doing very well | 720
no infectious or urinary tract symptoms | 720