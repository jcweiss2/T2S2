59 years old | 0
    male | 0
    hypertensive | 0
    non-diabetic | 0
    admitted for stapled hemorrhoidopexy | 0
    rectal bleeding | -2592
    prolapsing piles | -2592
    tablet metoprolol 50 mg | -17520
    tablet amlodipine 5 mg | -17520
    4th degree piles | 0
    large external component | 0
    pre-operative investigations within normal limits | 0
    prophylactic antibiotics | -0.5
    ceftriaxone | -0.5
    gentamycin | -0.5
    standard SH performed | 0
    spinal anesthesia | 0
    difficulty in closure | 0
    hemorrhoids excised | 0
    intraoperative uneasiness | 0
    intraoperative discomfort | 0
    sedated with midazolam 1mg | 0
    MAP fell below 65 mm Hg | 0
    hypotensive for 10-12 min | 0
    Ringer lactate 500 ml | 0
    tetrastarch 500 ml | 0
    MAP stabilisation above 70 mm Hg | 0
    total fluid administered 1300 ml | 0
    shifted to post-operative ward | 0
    pain at operative site | 120
    intranasal butorphanol nasal spray 1 mg | 120
    uneventful post-operative period | 120
    did not pass urine | 720
    generalized weakness | 720
    breathlessness | 720
    BP falling to MAP below 60 mm Hg | 960
    1L 0.9% normal saline | 960
    shifted to ICU | 960
    did not pass urine until 4 pm | 1080
    BP 70 mm Hg systolic | 1080
    central line inserted | 1080
    CVP guided fluid therapy | 1080
    targeted CVP around 10 mm Hg | 1080
    ABG analysis | 1080
    oxygen administered through venturi mask | 1080
    monitoring of non-invasive BP | 1080
    pulse rate monitoring | 1080
    heart rate monitoring | 1080
    SpO2 monitoring | 1080
    temperature monitoring | 1080
    continuous CVP monitoring | 1080
    urine output monitoring | 1080
    abdominal girth monitoring | 1080
    temperature 102°F | 1080
    BP 74 mm Hg systolic | 1080
    pulse rate 134 bpm | 1080
    respiratory rate 32/min | 1080
    SpO2 78% | 1080
    decreased air entry in both lungs | 1080
    fine crepts present | 1080
    abdominal distension | 1080
    no abdominal tenderness | 1080
    absent bowel sounds | 1080
    urinary catheterization | 1080
    electrocardiogram sinus tachycardia | 1080
    cardiac markers within normal limits | 1080
    noradrenaline infusion | 1080
    dopamine infusion | 1080
    routine investigations | 1080
    coagulation profile | 1080
    serum procalcitonin levels | 1080
    ABG metabolic acidosis | 1080
    pO2 51.9 mm Hg | 1080
    pCO2 37.8 mm Hg | 1080
    pH 7.27 | 1080
    HCO3- 17.5 mmol/L | 1080
    BE –8.7 mmol/L | 1080
    biphasic positive airway pressure ventilation | 1080
    blood cultures | 1080
    fungal staining | 1080
    meropenem 2 g IV | 1080
    meropenem 1 g in 100 ml NS twice daily | 1080
    teicoplanin 400 mg IV stat | 1080
    teicoplanin 400 mg once daily on alternate days | 1080
    blood urea 69 mg/dl | 1080
    serum creatinine 3.7 mg/dl | 1080
    metronidazole 500 mg IV three times daily | 1080
    vasopressors started | 1080
    MAP maintained 60'70 mm Hg | 1080
    urine output 50 ml in 1 h | 1080
    sequential organ failure assessment score 14 | 1080
    deranged coagulation profile | 1080
    6 units fresh frozen plasma transfused | 1080
    chest physiotherapy | 1080
    nebulization | 1080
    general nursing care | 1080
    hemodynamic parameters improved | 1080
    urine output improved | 1080
    ABG improved | 1080
    noradrenaline tapered | 1080
    dopamine tapered | 1080
    intermittent oxygen through Hudson mask | 1080
    improved after 4 days | 4320
    shifted to room care | 4320
    discharged after nine days | 216
    
    