83 years old | 0 | 0 
male | 0 | 0 
admitted to the hospital | 0 | 0 
leg ecchymosis | 0 | 0 
anuric | 0 | 0 
rhabdomyolysis-induced AKI | 0 | 0 
sepsis | 0 | 0 
acute prostatitis | 0 | 0 
syncope | -12 | -12 
fell to the ground | -12 | -12 
lying on the floor | -12 | 0 
increased urea | 0 | 0 
increased creatinine | 0 | 0 
increased myoglobin | 0 | 0 
increased CPK | 0 | 0 
increased LDH | 0 | 0 
increased CRP | 0 | 0 
increased PCT | 0 | 0 
increased total bilirubin | 0 | 0 
increased direct bilirubin | 0 | 0 
increased AST | 0 | 0 
increased ALT | 0 | 0 
increased PSA | 0 | 0 
increased white blood cell count | 0 | 0 
volume expansion | 0 | 504 
diuretic treatment | 0 | 504 
antibiotic treatment | 0 | 504 
furosemide | 0 | 192 
femoral central venous catheter placement | 0 | 0 
HFR-Supra | 0 | 120 
extracorporeal treatment | 0 | 120 
myoglobin removal | 0 | 120 
inflammatory status reduction | 0 | 120 
fluid balance maintenance | 0 | 120 
low molecular weight heparin administration | 0 | 0 
urea reduction | 96 | 96 
creatinine reduction | 96 | 96 
myoglobin reduction | 96 | 96 
CPK reduction | 96 | 96 
LDH reduction | 96 | 96 
CRP reduction | 96 | 96 
PCT reduction | 96 | 96 
urine output increase | 96 | 504 
furosemide tapering | 192 | 192 
oral furosemide administration | 192 | 504 
antibiotic therapy switch | 48 | 48 
piperacillin/tazobactam | 0 | 48 
meropenem | 48 | 504 
HFR-Supra sessions | 0 | 120 
blood flow | 0 | 120 
endogenous ultrafiltrate flow | 0 | 120 
ultrafiltration rate adjustment | 0 | 120 
femoral hemodialysis catheter removal | 120 | 120 
right jugular central venous catheter placement | 120 | 120 
on-line hemodiafiltration | 120 | 168 
high-flux hemodialysis | 168 | 192 
dialysis therapy prolongation | 120 | 192 
renal failure | 0 | 504 
chronic kidney disease | 504 | 504 
discharge | 504 | 504 
urea level at discharge | 504 | 504 
creatinine level at discharge | 504 | 504 
CRP level at discharge | 504 | 504 
total bilirubin level at discharge | 504 | 504 
ASL level at discharge | 504 | 504 
ALT level at discharge | 504 | 504 
PSA level at discharge | 504 | 504 
white blood cell count at discharge | 504 | 504 
urea level 6 months after discharge | 1512 | 1512 
creatinine level 6 months after discharge | 1512 | 1512 
GFR 6 months after discharge | 1512 | 1512