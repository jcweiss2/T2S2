70 years old | 0
male | 0
T3V1N0M0 rectal tumor | -8760
laparoscopic APR | -8760
adjuvant chemotherapy | -8760
oxaliplatin | -8760
fluorouracil | -8760
calcium folinate | -8760
perineal hernia | -408
reconstruction of the pelvic floor | -408
biological mesh | -408
Permacol | -408
transperineal approach | -408
postoperative course uneventful | -408
pelvic-abdominal CT scan | -136
no signs of locoregional recurrence | -136
no reherniation | -136
weight loss | -72
thoracic-abdominal CT scan | -72
multiple metastases to the liver | -72
multiple metastases to the lungs | -72
chemotherapy | -72
bevacizumab | -72
irinotecan | -72
calcium folinate | -72
fluorouracil | -72
signs of sepsis | 0
high temperature | 0
tachycardia | 0
hypotension | 0
pain in the right buttock | 0
infection at the area | 0
acute US examination | 0
abscess | 0
US-guided drainage | 0
intravenous fluids | 0
broad-spectrum antibiotics | 0
CT scan with contrast | 24
subcutaneous abscess cavity | 24
communication to the small bowel | 24
laparotomy | 48
perineal fistula from the distal ileum | 48
resection of the small bowel | 48
primary anastomosis | 48
fluid and electrolyte disturbances | 48
intensive care unit | 48
pressors | 48
parenteral nutrition | 48
perineal wound | 48
vacuum-assisted closure | 48
hospice for terminal care | 672
discharged | 672