9 years old | 0
female | 0
rhabdomyosarcoma | -504
fever | -168
jaundice | -168
right upper quadrant abdominal pain | -168
VAC chemotherapy | -504
vincristine | -504
actinomycin-D | -504
cyclophosphamide | -504
wide excision of the tumor | -252
postoperative VAC chemotherapy | -252
mild abdominal pain | -192
neutropenic fever | -192
white blood cell 0.78×10^3/μL | -192
hemoglobin 6.9 g/dL | -192
platelets 4×10^3/μL | -192
intravenous broad-spectrum antibiotics | -192
piperacillin | -192
tazobactam | -192
transfusion | -192
red blood cells | -192
platelets | -192
granulocyte colony stimulating factor | -192
mild elevation of liver enzymes | -192
aspartate transaminase 103 U/L | -192
alanine transaminase 77 U/L | -192
total bilirubin 1.5 mg/dL | -192
abdominal pain aggravated | -168
persistent fever | -168
pancytopenia | -168
white blood cell 0.42×10^3/μL | -168
hemoglobin 8.1 g/dL | -168
platelet 6×10^3/μL | -168
marked increase in liver enzymes | -168
aspartate transaminase 519 U/L | -168
alanine transaminase 370 U/L | -168
hyperbilirubinemia | -168
total bilirubin 4.8 mg/dL | -168
prothrombin time 1.17 international normalized ratio | -168
active partial thromboplastin time 55.2 seconds | -168
hepatomegaly | -168
icteric sclerae | -168
abdominal distension | -168
body weight increased by 6.1% | -168
severe abdominal pain | -144
fever peaked to 38.9°C | -144
reversed blood flow of the right portal vein | -144
defibrotide treatment | -144
transfer to intensive care unit | -144
condition became unstable | -144
diffuse pleural effusion | -144
irritable | -144
did not recognize mother and medical personnel | -144
liver enzyme levels peaked | -144
aspartate transaminase 2,110 U/L | -144
alanine transaminase 1,908 U/L | -144
total bilirubin 15.1 mg/dL | -144
direct bilirubin 8.6 mg/dL | -144
ammonia level increased | -144
hepatic encephalopathy | -144
vasopressor infusion | -144
paracentesis of the ascites | -144
glycerin enema | -144
rifaximin | -144
lactulose | -144
mechanical ventilation | -120
condition gradually improved | -96
recovery from myelosuppression | -96
defibrotide treatment continued for 10 days | -96
body weight began to decrease | -72
fever gradually subsided | -72
laboratory results showed improvement | -72
weaned from mechanical ventilator | 0
abdominal US showed normalized blood flow of the right portal vein | 120
discharged | 216
bilirubin level normalized | 432
parents refused further chemotherapy | 432
surveillance imaging studies showed no evidence of recurrence of cancer or any sequelae to the liver | 528