35 years old | 0
female | 0
brought in by emergency medical services | 0
level 1 trauma code | 0
struck by motor vehicle | 0
loss of consciousness | 0
Glasgow Coma Scale 15 | 0
severe respiratory distress | 0
complaints of shortness of breath | 0
pulse rate 125 beats per minute | 0
BP 67/20 | 0
respiratory rate 45 breaths per minute | 0
ecchymoses around left eye | 0
facial laceration | 0
decreased breath sounds on right side | 0
no other obvious external signs of trauma | 0
FAST performed | 0
FAST negative | 0
one liter of isotonic fluid administered | 0
blood pressure normalized | 0
chest X-ray obtained | 0
large right pneumothorax | 0
chest tube placed | 0
lung re-expansion successful | 0
vitals normalized | 0
intubated for agitation | 0
CT scan workup | 0
non-contrast CT head/C-spine | 0
CT Chest/Abdomen/Pelvis with IV contrast | 0
grade 5 liver laceration | 0
grade 5 right kidney laceration | 0
grade 1 splenic laceration | 0
left clavicle fracture | 0
bilateral small pneumothoraces | 0
hypotensive after CT scan | 0
decision for operating room | 0
entered abdomen | 0
large amount of blood encountered | 0
blood evacuated | 0
four-quadrant packing | 0
right medial visceral rotation performed | 0
large hematoma in retroperitoneum | 0
exploration of hematoma | 0
shattered inferior portion of kidney | 0
superior portion of kidney bleeding significantly | 0
renal vessels ligated with 2–0 silk suture | 0
nephrectomy performed | 0
right ureter unable to be located | 0
hemostasis of spleen and liver | 0
removal of packs | 0
no other abdominal injuries | 0
repacked | 0
Barker vac placed | 0
brought to ICU | 0
received 7 units packed red blood cells | 0
received 3 units fresh frozen plasma | 0
received 4 liters crystalloid | 0
taken to Interventional Radiology | 24
no active extravasation from hepatic or splenic artery | 24
returned to OR on POD#2 | 48
active bleeding over dome of liver | 48
packs removed | 48
repacked | 48
hemostasis achieved | 48
monitored in ICU | 48
returned to OR on POD#5 | 120
third laparotomy | 120
packs removed | 120
no bleeding noted | 120
right ureterectomy performed | 120
abdomen closed primarily | 120
brought back to ICU | 120
extubated on POD#7 | 168
persistently elevated WBC | 312
CT abdomen/pelvis with IV contrast on POD#13 | 312
right kidney remnant isolated | 312
large rim-enhancing collection | 312
urinoma | 312
ultrasound-guided drainage on POD#16 | 384
8 French drainage catheter placed | 384
cultures without growth | 384
persistent drainage | 384
options discussed | 384
IR angioembolization vs completion nephrectomy | 384
decision for angioembolization | 384
embolization performed on POD#19 | 456
two traumatic pseudoaneurysms found | 456
embolized with 300–500 micron embospheres | 456
lower renal artery occluded with tornado microcoil | 456
completion arteriogram successful occlusion | 456
post-embolization febrile | 456
complaints of severe flank pain | 456
antibiotics continued for 24 hours | 456
afebrile | 480
pain resolved | 480
drain removed on POD#25 | 600
stable for discharge on POD#26 | 624
no residual functional deficits | 624
follow-up BUN/Cr 17/1.16 | 624
