32 weeks | 0
preterm | 0
baby boy | 0
vaginal delivery | 0
28 years old | 0
primigravida mother | 0
antenatal steroids | -24
premature rupture of membranes | -24
spontaneous labour | -24
Apgar 9-10 | 0
normal examination at birth | 0
birth weight 1800 g | 0
head circumference 30.5 cm | 0
admitted to neonatal intensive care unit | 0
orally fed | 0
antibiotics | 0
elevated procalcitonin 0.45 ng/ml | 0
fever 38.5°C | 24
screeches | 24
CRP 77 mg/L | 24
WBC 4.81 x 10^9/L | 24
normal lumbar puncture | 24
haemoculture positive for Gram-negative bacillus | 24
intubated | 48
severe apnoea | 48
altered hemodynamic status | 48
painful abdomen | 48
distended abdomen | 48
contractured abdomen | 48
large gastric residual volume | 48
clear appearance of gastric residual | 48
regular stools | 48
normal stools | 48
abdominal X-ray | 48
ultrasound | 48
non-abnormal signs on imaging | 48
CRP 155 mg/L | 48
normal WBC | 48
thrombocytopenia | 48
exploratory laparotomy | 48
perforated appendicitis | 48
peritonitis | 48
appendectomy | 48
peritoneal lavage with warm saline | 48
favourable outcome | 48
histopathology confirmed appendicitis | 48
no Hirschprung's disease | 48
follow-up at 5 months | 3600
