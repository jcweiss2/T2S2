17 years old|0
    African American|0
    male|0
    depression|0
    transferred from an outside hospital|0
    3-day history of nonbilious, nonbloody vomiting|0
    new-onset erythematous blanching macular rash on trunk, arms, legs|0
    tachycardic (134 beats per minute)|0
    hypertensive (142/98 mm Hg)|0
    febrile with temperature of 38.5°C|0
    hypotensive (90/60 mm Hg)|4
    remained tachycardic|4
    concerns of septic shock|4
    blood cultures drawn|4
    empiric antibiotic treatment|4
    admitted to the hospital|4
    hyponatremia (135 mMol/L)|4
    direct hyperbilirubinemia (6.18 mg/dL)|4
    low lactate dehydrogenase (111 units/L)|4
    polymorphic neutrophil dominant leukocytosis (12 800/mm3)|4
    elevated C-reactive protein (99.3 mg/L)|4
    sterile pyuria|4
    direct hyperbilirubinemia continued to rise|192
    peaked at 14.12 mg/dL 8 days after admission|192
    γ-glutamyl transferase within normal limits|192
    lipase within normal limits|192
    amylase within normal limits|192
    transaminases within normal limits|192
    alanine aminotransferase at 51 Units/L|192
    further laboratory investigations for causes of direct hyperbilirubinemia negative|192
    ultrasound showed over distended gallbladder|192
    computed tomography negative for obstruction|192
    magnetic resonance cholangiopancreatography negative for obstruction|192
    extensive infectious disease workup negative|192
    cytomegalovirus negative|192
    Epstein-Barr virus negative|192
    group A Streptococcus negative|192
    human immunodeficiency virus negative|192
    hepatitis panel negative|192
    blood cultures negative|192
    urine cultures negative|192
    remained hypotensive|192
    remained tachycardic|192
    several fluid boluses|192
    developed S3 gallop|192
    orthopnea|192
    elevated brain natriuretic peptide (2749 pg/mL)|192
    respiratory distress|192
    heart failure|192
    chest X-ray demonstrated bilateral lower lobe pleural effusions|192
    echocardiogram demonstrated mild decrease in left ventricular function|192
    mild mitral valve regurgitation|192
    tricuspid valve regurgitation|192
    small posterior pericardial effusion|192
    coronary arteries did not demonstrate pathology|192
    transferred to pediatric intensive care unit|192
    concerns of new-onset heart failure|192
    worsening leukocytosis|192
    heart failure stabilized|192
    respiratory distress stabilized|192
    new-onset microcytic anemia|192
    thrombocytosis|192
    elevated ferritin|192
    low albumin|192
    significant systemic inflammation|192
    diagnosed with incomplete Kawasaki disease|192
    clinical features (2 or 3)|192
    fever ≥5 days|192
    peripheral extremity changes|192
    polymorphous rash|192
    elevated CRP|192
    echocardiogram changes|192
    thrombocytosis after seventh day of fever|192
    albumin ≤3.0 g/dL|192
    elevated ALT level|192
    WBC count ≥15 000/mm|192
    ≥10 WBC/hpf on urinalysis|192
    hyperbilirubinemia likely from acalculous cholecystitis|192
    treated with ursodiol|192
    intravenous immunoglobulin (IVIG)|192
    moderate dose of 30 mg/kg/day divided every 6 hours|192
    supportive treatment for shock|192
    improved|360
    discharged from hospital|360
    feeling back at baseline|360
    scleral icterus|360
    direct bilirubin remained elevated at 4.24 mg/dL|360
    low-dose aspirin (5 mg/kg/day)|360
    ursodiol 300 mg QID|360
    scheduled follow-up 10 days after discharge|360
    minimal residual peeling of palms and soles|360
    bilirubin normalized|360
    echocardiogram demonstrated grossly normal coronary arteries|360
    previous abnormalities no longer appreciated|360
    final diagnosis incomplete KD with atypical features|360
    Kawasaki disease shock syndrome (KDSS)|360
    <|eot_id|>