12 years old | -9360
male | -9360
admitted to the hospital | 0
abdominal lymphoma | -9360
infection with methicillin-resistant Staphylococcus aureus (MRSA) | 0
isolation | 0
chemotherapy scheduled | 0
chemotherapy could not commence | 0
treated with local antiseptic (octenidin) | 0
treatment with octenidin for 12 days | 12
no improvement | 12
treated with Australian medical honey (Medihoney) | 12
wound free of bacteria | 14
chemotherapy started | 14
discharged | 14 
leukemia | -9360
chemotherapy | -9360
wound healing problems | -9360
wound infections | -9360
bloodstream infections | -9360
immunocompromized patients | -9360
nosocomial spread | 0
diffuse erythematous or maculopapular eruption | 0
pruritus | 0
DRESS syndrome | 0
fever persisted | 0
rash persisted | 0 
infection cleared | 14
medical honey effective | 0
hygroscopic | 0
glucose oxidase | 0
gluconic acid | 0
hydrogen peroxide | 0
antibacterial properties | 0
pH level of honey | 0
bacterial colonization | 0
infection | 0
recalcitrant wound healing | 0
acidification of wounds | 0
speeds healing | 0
anti-inflammatory effects | 0
debriding action | 0
malodour | 0
medical honey irradiated | 0
Clostridium botulinum spores | 0
gamma irradiation | 0
Medihoney | 0
mixture of two honeys | 0
antibacterial activity | 0
licensed for wound care | 0
practical advances | 0
easy to change | 0
no pain | 0
no harm | 0
regenerating tissue | 0
malodour abandoned | 0
anti-inflammatory | 0
debriding effects | 0
diabetes | 0
well accepted | 0
drawbacks | 0
pain | 0
atopic reactions | 0
systemic atopic reaction | 0
cost | 0
dressing changes | 0
scientific evidence | 0
prospectively randomized controlled study | 0
in vitro studies | 0
animal studies | 0
clinical experiences | 0
observational studies | 0
what makes medical honey effective | 0
mechanism of action | 0
antibacterial properties | 0
anti-inflammatory effects | 0
debriding action | 0
pH level | 0
why is the final product irradiated | 0
Clostridium botulinum | 0
spores | 0
anaerobic environment | 0
botulinum toxin | 0
systemic effects | 0
paralysis | 0
cardiac arrhythmia | 0
gamma irradiation | 0
safety measure | 0
Medihoney not an antiseptic | 0
antiseptic criteria | 0
fast onset of activity | 0
broad spectrum effect | 0
enhancement of wound healing | 0
no adverse effects | 0
moderate cost | 0
conventional wound care products | 0
paediatric oncology | 0
silver dressings | 0
povidone iodine | 0
iodine products | 0
systemic absorption | 0
thyroid function | 0
alcohol-containing antiseptics | 0
systemic antibiotics | 0
neutropenia | 0
fever | 0
local sign | 0
soft tissue infection | 0
bacterial resistance | 0
frequency of dressing changes | 0
exudate | 0
stable wound care | 0
prospective studies | 0
compliance issues | 0
pain relief | 0
odour control | 0
patient satisfaction | 0
leg ulcers | 0
compression therapy | 0
Medihoney dressings | 0
ulcer pain | 0
size decreased | 0
odorous wounds | 0
deodorized | 0
patient acceptance | 0
concordance | 0
adverse effects | 0
stinging pain | 0
local atopic reactions | 0
systemic atopic reaction | 0
cost issues | 0
randomized controlled trial | 0
natural honey | 0
IntraSite Gel | 0
healing time | 0
adverse events | 0
satisfaction with treatment | 0
cost of treatment | 0
WoundViewer database | 0
prospective collection | 0
datasets | 0
clinical use | 0
medical honey products | 0
wound care | 0
clinical evidence | 0
comparative studies | 0
conclusion | 0
prospective randomized studies | 0
safety | 0
efficacy | 0
medical honey | 0
wound care | 0
CE-certified honey dressings | 0
Medihoney products | 0
alternative treatment | 0
wounds | 0
acknowledgements | 0
Humboldt Foundation | 0
German Chancellor Scholarship | 0
WoundViewer database | 0
Medihoney Inc | 0