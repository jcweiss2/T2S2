75 years old | 0
    female | 0
    recurrent urinary tract infections | 0
    hypothyroidism | 0
    chronic pain | 0
    depression | 0
    opioid dependence | 0
    presented to the emergency department | 0
    altered mental status | 0
    poor historian | 0
    family not present | 0
    temperature 100 °F | 0
    heart rate 130 bpm | 0
    blood pressure 114/60 mmHg | 0
    pulse oximetry 86% on room air | 0
    using accessory muscles | 0
    diminished air entry | 0
    scattered rhonchi | 0
    wheezes bilaterally | 0
    bilateral lower extremity edema | 0
    alert | 0
    awake | 0
    oriented only to self | 0
    WBC count 19,000 | 0
    neutrophilic predominance | 0
    BUN 43 mg/dl | 0
    creatinine 2.1 mg/dl | 0
    albumin 3 g/dl | 0
    lactic acid 2.2 mg/dL | 0
    ABG pH 7.37 | 0
    ABG PaCO2 29.9 mmHg | 0
    ABG PaO2 45.5 mmHg | 0
    acute hypoxic respiratory failure | 0
    admission CXR bilateral infiltrates | 0
    placed on BiPAP | 0
    improvement within 24-48 hours | 24
    respiratory status worsened | 72
    unable to maintain oxygen saturation | 72
    repeat CXR stable bilateral infiltrates | 72
    worsening hypoxia | 72
    sinus tachycardia | 72
    new onset paroxysmal atrial fibrillation | 72
    EKG S1QIIITIII pattern | 72
    received ceftriaxone | 0
    received azithromycin | 0
    prophylactic low molecular weight heparin | 0
    chest CTA revealed saddle PE | 72
    lethargic | 72
    hypoxia not improving | 72
    upgraded to ICU | 72
    intubated | 72
    Mycoplasma IgM > 950 U/mL | 72
    Mycoplasma IgG > 320 U/mL | 72
    WBC count improved | 72
    lactic acid normalized | 72
    sputum culture negative | 72
    blood culture negative | 72
    anticardiolipin antibody | 72
    lupus anticoagulant | 72
    protein C | 72
    protein S | 72
    prothrombin gene mutation | 72
    factor V Leiden mutation | 72
    decreased protein C activity | 72
    increased cold agglutinin titers | 72
    started on tPA | 72
    started on heparin drip | 72
    intubated for three days | 72
    weaned off mechanical ventilation | 96
    antibiotics discontinued | 96
    maintaining oxygen saturation on 6 L nasal cannula | 96
    severely hypoxic | 144
    on 100% high flow nasal cannula | 144
    unable to maintain oxygen saturation | 144
    reintubated | 144
    concern for intraalveolar hemorrhage | 144
    bronchoscopy serosanguinous secretions | 144
    no overt bleeding | 144
    placed on cefepime | 144
    placed on vancomycin | 144
    placed on fluconazole | 144
    repeat cultures negative | 144
    antibiotics discontinued | 144
    extubated again | 144
    downgraded to medical telemetry | 144
    physical deconditioning | 144
    required rehabilitation | 144
    discharged to rehabilitation facility | 144
    PE | 72
    Mycoplasma pneumonia | 72
    saddle PE | 72
    anemia | 72
    cold agglutinins | 72
    hemolysis | 72
    increased indirect bilirubin | 72
    low haptoglobin levels | 72
    catheter directed thrombolysis | 72
    anticoagulation with heparin | 72
    full recovery | 144
    focal infiltrate | 72
    multiple areas of atelectasis | 72
    S1QIIITIII pattern | 72
    empiric treatment | 72
    thrombolysis | 72
    acute saddle PE | 72
    prothrombotic state | 72
    venous thromboembolism | 72
    early treatment initiation | 144
    