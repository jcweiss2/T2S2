33 years old | 0
male | 0
minor superficial injury on lower left leg | -240
ski vacation | -240
deterioration of wound conditions | -240 to -168
outpatient visit to general medicine center | -168
initiation of oral Cefuroxime | -168
progressive clinical deterioration | -168 to -144
aching hematoma | -144
admitted to hospital | -144
surgical treatment of hematoma | -144
two further wound debridements | -144 to -96
application of vacuum-assisted closure | -144 to -96
antibiotic therapy escalated to Clindamycin and Tazobactam | -144
transferred to university hospital | 0
awake | 0
oriented | 0
stable respiratory condition | 0
stable circulatory condition | 0
temperature 37.2°C | 0
blood pressure 171/85 mmHg | 0
pulse 140 beats per minute | 0
rhythmic pulse | 0
oxygen saturation 95% | 0
somnolent | 0
easily aroused | 0
severe pain in both axillae | 0
severe pain in both groins | 0
swellings in both axillae | 0
swellings in both groins | 0
increased WBC count (23.1×10³/μL) | 0
increased CRP (298.8 mg/dL) | 0
surgical wound excisions | 0
large debridement in left lower leg | 0
antibiotic therapy changed to Meropenem, Penicillin G, and Clindamycin | 0
tissue samples taken | 0
swabs taken | 0
blood cultures taken | 0
no causative pathogen identified | 0
increased inflammation markers | 24
clinical deterioration | 24
Levofloxacin added | 24
Daptomycin added | 24
Caspofungin added | 24
hole-body computed tomography scan | 72
fasciitis of left upper and lower leg | 72
symmetrical bilateral pulmonary edema | 72
bilateral pleural effusions | 72
basal atelectasis | 72
generalized barrier disruption | 72
progredient lung edema | 72
respiratory dysfunction | 72
mechanical ventilation | 72
operational inspection of axillae | 96
large debridement of both axillae | 96
left thigh surgically explored | 96
fasciotomy performed | 96
increase of necrotic area | 96
positive serological evidence of Herpes simplex virus-I | 96
Acyclovir initiated | 96
Corynebacterium tuberculostearicum detected | 96
Acinetobacter baumanii detected | 96
direct pathogen detection unsuccessful | 96
Hydrocortisone initiated | 120
IVIg (Pentaglobin) initiated | 120
hyperinflammation diminished | 120
general condition improved | 120
weaning from respirator | 168
CRP decreased | 168
WBC decreased | 168
procalcitonin decreased | 168
hemodynamic support reduced | 168
vacuum-assisted wound closure | 240
moved to primary care station | 768
wound closure with split-skin graft | 936
discharged | 1152
healthy at follow-up | 4320
