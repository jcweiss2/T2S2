39 years old | 0
    male | 0
    admitted to the hospital | 0
    hematemesis | 0
    hemorrhagic shock | 0
    arterial hypertension | 0
    autoimmune thyroiditis | 0
    type 2 diabetes mellitus | 0
    diabetic neuropathy | 0
    retinopathy | 0
    nephropathy | 0
    stage 3 chronic renal failure | 0
    no history of liver disease | 0
    no alcohol abuse | 0
    no exposure to hepatotoxic substances | 0
    assumption of non-steroidal anti-inflammatory drugs | -168
    neuropathic lower limbs pain | -168
    emergency esophagogastroduodenoscopy | 0
    huge clot in the stomach | 0
    active bleeding | 0
    source of hemorrhage not identified | 0
    cardiac arrest | 0
    cardiopulmonary resuscitation | 0
    hemodynamic stability achieved | 0
    transferred to intensive care unit | 0
    administration of high-dose proton pump inhibitors | 0
    abdominal Doppler ultrasonography | 0
    no sign of liver disease | 0
    normal flow into vena porta | 0
    pancreas poorly assessed | 0
    spleen region poorly assessed | 0
    important abdominal meteorism | 0
    further esophagogastroduodenoscopy | 24
    source of bleeding not identified | 24
    celio-mesenteric arteriography | 24
    no arterial blush | 24
    two episodes of gastrointestinal hemorrhage | 48
    transfused with packed red blood cells | 48
    transfused with plasma | 48
    abdominal contrast-enhanced computed tomography | 72
    severe atrophy of pancreas | 72
    chronic pancreatitis | 72
    thrombosis of splenic vein | 72
    splenomegaly | 72
    cavernomatous transformation of splenic hilum | 72
    third esophagogastroduodenoscopy | 96
    remission of bleeding | 96
    large isolated varices of gastric fundus | 96
    signs of recent bleeding | 96
    left-sided portal hypertension | 96
    gastrointestinal hemorrhage from gastric varices | 96
    scheduled for splenectomy | 96
    splenomegaly (17 cm) | 96
    laparoscopic approach deemed feasible | 96
    splenic artery embolization | 96
    two vascular plugs | 96
    coil | 96
    spleen ischemic | 120
    reticulum of varices at splenic hilum | 120
    laparoscopic dissection | 120
    splenic artery divided | 120
    gastroepiploic vein divided | 120
    splenic vein divided | 120
    short gastric vessels divided | 120
    minimal blood losses | 120
    no intraoperative complications | 120
    spleen extracted | 120
    postoperative course uneventful | 124
    discharged on postoperative day 4 | 124
    no further episodes of gastric bleeding | 8760
    <|eot_id|>
    