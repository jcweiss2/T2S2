29 years old | 0
    male | 0
    hepatic transplantation in 2009 | -105192
    autoimmune hepatitis | -105192
    hepatic rejection | -168
    hepatic transplantation considered again | 0
    minimal shortness of breath | 0
    orthopnea | 0
    vital signs within normal limits | 0
    loud, superficial, systodiastolic murmur | 0
    palpable thrill along right and left lower parasternal border | 0
    hepatic failure findings | 0
    edema | 0
    ascites | 0
    hypoalbuminemia | 0
    albumin 2.6 g/dL | 0
    thrombocytopenia | 0
    platelets 56,000/mm3 | 0
    hyperbilirubinemia | 0
    total bilirubin 15.6 mg/dL | 0
    direct bilirubin 11.2 mg/dL | 0
    transthoracic echocardiography (TTE) | 0
    transesophageal echocardiography (TEE) | 0
    ruptured aneurysm from noncoronary sinus of valsalva | 0
    turbulent flow from aortic aneurysm toward left atrium | 0
    mild aortic regurgitation | 0
    moderate mitral regurgitation | 0
    continuous high-velocity jet 4.0 m/s | 0
    evaluated at cardiology and cardiovascular surgeon's council | 0
    surgical operation recommended | 0
    refused surgery | 0
    hepatic transplant preparations delayed | 0
    discharged | 168
    admitted to gastroenterology clinic after 3 months | 2160
    elevated hepatic enzymes | 2160
    peak alanine aminotransferase 1895 U/L | 2160
    peak aspartate aminotransferase 2356 U/L | 2160
    ascites | 2160
    diffuse edema | 2160
    fever 39°C | 2160
    increased infection parameters | 2160
    peak C-reactive protein 89 mg/dL | 2160
    peak white blood cell 33,000/mm3 | 2160
    decreased complement values | 2160
    C3 6.6 mg/dL | 2160
    C4 18 mg/dL | 2160
    four blood cultures taken | 2160
    viridans group streptococcus | 2160
    bedside portable echocardiography | 2160
    two gross vegetations on atrial surface of anterior mitral leaflet | 2160
    posterior mitral leaflet | 2160
    ampicillin initiated | 2160
    gentamicin initiated | 2160
    infective endocarditis | 2160
    septic shock | 2160
    died due to multiple organ dysfunction syndrome | 2160