72 years old | 0  
    woman | 0  
    primary biliary cholangitis | 0  
    admitted to the hospital | 0  
    general fatigue | 0  
    dyspnea on effort | 0  
    lumbar vertebral compression fracture | -113880  
    osteoporosis | -113880  
    heart failure | -113880  
    tachycardia-induced cardiomyopathy | -113880  
    persistent atrial fibrillation | -113880  
    rapid ventricular response | -113880  
    radiofrequency catheter ablation | -113880  
    paroxysmal atrial flutter | -113880  
    sinus bradycardia | -113880  
    bisoprolol fumarate | -113880  
    enalapril maleate | -113880  
    rivaroxaban | -113880  
    ursodeoxycholic acid | -113880  
    CelestamineⓇ | -113880  
    marked sarcopenia | 0  
    blood pressure 90/42 mmHg | 0  
    regular pulse rate 60 beats/min | 0  
    no cardiac murmur | 0  
    no respiratory crackles | 0  
    normocytic anemia | 0  
    elevated serum brain natriuretic peptide | 0  
    elevated anti-mitochondrial antibody M2 | 0  
    chest radiography no cardiomegaly | 0  
    no congestion | 0  
    no pleural effusion | 0  
    electrocardiogram normal sinus rhythm | 0  
    P-waves extremely low voltage | 0  
    T-wave inversion in precordial leads | 0  
    transthoracic echocardiography mild generalized hypokinesis | 0  
    ejection fraction 52% | 0  
    bilateral atrial dilatation | 0  
    no left ventricular dilatation | 0  
    no hypertrophy | 0  
    no pericardial effusion | 0  
    transmitral Doppler inflow pseudo-normalization | 0  
    E/A ratio 1.02 | 0  
    mitral annulus velocity impaired left ventricular relaxation | 0  
    e' 5.3 cm/s | 0  
    coronary angiography intact coronary arteries | 0  
    right heart catheterization | 0  
    mean pulmonary capillary wedge pressure 6 mmHg | 0  
    pulmonary artery pressure 22/8 mmHg | 0  
    mean right atrial pressure 6 mmHg | 0  
    cardiac index 1.73 L/min/m2 | 0  
    anti-mitochondrial M2 antibody-associated cardiomyopathy | 0  
    endomyocardial biopsy | 0  
    right ventricular perforation | 24  
    cardiogenic shock | 24  
    pericardiocentesis | 24  
    surgical closure | 24  
    percutaneous cardiopulmonary support | 24  
    hemodynamic instability | 24  
    transfer to cardiac care unit | 24  
    dobutamine 5 μg/kg/min | 24  
    intubated | 24  
    medications discontinued | 24  
    biventricular Takotsubo cardiomyopathy | 24  
    progressive reduction in blood pressure | 24  
    reduced daily urine output | 24  
    no deterioration in echocardiographic assessment | 24  
    rapid improvement in biventricular Takotsubo cardiomyopathy | 24  
    central venous pressure >12 mmHg | 24  
    inferior caval vein diameter >18 mm | 24  
    serum electrolyte levels stable | 24  
    no hypovolemic shock | 24  
    no septic shock | 24  
    serial monitoring cardiac output | 24  
    systemic vascular resistance reduction | 24  
    serum glucose 77 mg/dL | 72  
    intravenous hyperalimentation | 72  
    systemic vascular resistance 740 dynes・sec・cm-5 | 72  
    acute adrenal insufficiency | 72  
    discontinuation of CelestamineⓇ | 72  
    long-term CelestamineⓇ use | -113880  
    hydrocortisone 150 mg/day | 72  
    hemodynamic stabilization | 72  
    systemic vascular resistance normalization | 72  
    serum adrenocorticotropic hormone 167.9 pg/mL | 72  
    serum cortisol 32.6 μg/dL | 72  
    uneventful clinical course | 72  
    hydrocortisone tapered | 72  
    oral hydrocortisone 10 mg/day | 72  
    discharged | 72  
    
