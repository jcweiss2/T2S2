62 years old | 0 | 0 
male | 0 | 0 
admitted to the hospital | 0 | 0 
bilateral otalgia | -120 | 0 
use of olive oil ear drops | -120 | 0 
Glasgow Coma Scale score 8 | -1 | -1 
bilateral otalgia not improved | -120 | 0 
past medical history of CRS with nasal polyposis | 0 | 0 
past medical history of chronic obstructive pulmonary disease | 0 | 0 
past medical history of hypertension | 0 | 0 
past medical history of glaucoma | 0 | 0 
past medical history of right sided keratoconus | 0 | 0 
past medical history of hypercholesterolaemia | 0 | 0 
beclomethasone/formoterol inhaler | 0 | 0 
salbutamol inhaler | 0 | 0 
amlodipine | 0 | 0 
simvastatin | 0 | 0 
beclometasone dipropionate nasal spray | 0 | 0 
tachypnoeic | 0 | 0 
tachycardic | 0 | 0 
pyrexial | 0 | 0 
Glasgow Coma Scale score 11 | 0 | 0 
bilateral green purulent rhinorrhea | 0 | 0 
bilateral proptosis | 0 | 0 
right sided chemosis | 0 | 0 
flexible nasendoscopy | 0 | 0 
thick green secretions | 0 | 0 
raised CRP | 0 | 0 
raised white cell count | 0 | 0 
raised neutrophil count | 0 | 0 
low lymphocyte count | 0 | 0 
raised lactate | 0 | 0 
pus aspirates collected | 0 | 0 
Streptococcus pneumoniae isolated | 0 | 0 
no evidence of fungal infection | 0 | 0 
contrast-enhanced computed tomography | 0 | 1 
opacification of the paranasal sinuses | 0 | 1 
bony erosion of the lateral walls of both ethmoid sinuses | 0 | 1 
soft tissue bulging into the right orbit | 0 | 1 
bilateral proptosis | 0 | 1 
no intracranial abnormality | 0 | 1 
increasingly combative | 1 | 24 
confused | 1 | 24 
aversion to light | 1 | 24 
lumbar puncture | 1 | 24 
pale cloudy fluid | 1 | 24 
extremely cellular specimen | 1 | 24 
high protein | 1 | 24 
low glucose | 1 | 24 
Streptococcus pneumoniae isolated | 1 | 24 
no evidence of fungal infection | 1 | 24 
treatment for sepsis and presumed meningitis initiated | 0 | 0 
intravenous ceftriaxone | 0 | 240 
fluticasone nasal spray | 0 | 240 
xylometazoline hydrochloride nasal spray | 0 | 240 
regular saline nasal irrigation | 0 | 240 
admitted to the critical care unit | 0 | 0 
intubated and ventilated | 12 | 12 
successfully extubated | 192 | 192 
completed a 10-day course of intravenous antibiotics | 240 | 240 
discharged home | 312 | 312 
ongoing input from the physiotherapy and occupational therapy teams | 312 | 312 
outpatient follow-up with the critical care and ENT teams | 312 | 312 
prescribed a 2-week course of betamethasone nasal drops | 312 | 336 
prescribed a 6-week course of fluticasone nasal spray | 336 | 504 
regular saline nasal irrigation | 312 | 504 
recovering well at 3-month follow-up | 744 | 744 
returned to work full time | 744 | 744 
some vivid memories of his stay on CCU | 744 | 744 
no signs of post-traumatic stress disorder | 744 | 744 
managed medically as an outpatient by the ENT team | 744 | 744 
ongoing CRS with nasal polyposis | 744 | 744 
did not wish for further sinus surgery | 744 | 744 
6-month follow-up contrast-enhanced magnetic resonance imaging | 1512 | 1512 
extensive bilateral ethmoid polyposis | 1512 | 1512 
hypertrophied inferior turbinates | 1512 | 1512 
left sided smooth dural enhancement | 1512 | 1512 
Aspergillus and Alternaria specific IgE levels within normal range | 1512 | 1512