59 years old | 0
male | 0
decreased general well-being | 0
somnolent | 0
cachexia | 0
arterial hypotension | 0
heart rate 90 bpm | 0
respiratory frequency 25 per minute | 0
urinary incontinence | 0
severe necrosis of the scrotum | 0
severe necrosis of the perineum | 0
spontaneously perforated necrosis | 0
smell suggesting moist gangrene | 0
inflammatory syndrome | 0
hemoglobin 6.7 mmd/L | 0
hemoglobin 5.3 mmd/L | 0
hemoglobin 5.5 mmd/L | 0
hemoglobin 4.8 mmd/L | 0
hemoglobin 5.1 mmd/L | 0
leukocytes 9.8 Gpt/L | 0
leukocytes 9.5 Gpt/L | 0
leukocytes 22.5 Gpt/L | 0
leukocytes 11 Gpt/L | 0
leukocytes 10.6 Gpt/L | 0
fibrinogen 8.7 g/L | 0
fibrinogen >9 g/L | 0
fibrinogen 7.7 g/L | 0
fibrinogen 6.3 g/L | 0
fibrinogen 4.5 g/L | 0
fibrinogen 6 g/L | 0
C-reactive protein 327 mg/L | 0
C-reactive protein 298 mg/L | 0
C-reactive protein 87 mg/L | 0
procalcitonin 7.24 μg/L | 0
procalcitonin 4.62 μg/L | 0
procalcitonin 2.2 μg/L | 0
procalcitonin 0.51 μg/L | 0
procalcitonin 0.34 μg/L | 0
partial thromboplastin time 42.3 seconds | 0
colonization of Bacteroides pyogenes | 0
colonization of Staphylococcus haemolyticus | 0
colonization of Escherichia coli | 0
colonization of Clostridium innocuum | 0
colonization of Enterococcus faecium | 0
colonization of Enterococcus faecalis | 0
colonization of Candida albicans | 0
colonization of non-albicans Candida | 0
Enterococcus faecium sensitive to macrolide-lincosamide-streptogramin | 0
Enterococcus faecium sensitive to glycylcycline | 0
Enterococcus faecium sensitive to glycopeptide class antibiotics | 0
Enterococcus faecium resistant to beta-lactam antibiotic | 0
Enterococcus faecium resistant to aminoglycoside antibiotic | 0
Enterococcus faecium resistant to fluoroquinolone drug class | 0
injury of the right lumbar plexus | 0
calcified chronic pancreatitis | 0
pancreatic pseudocyst | 0
applied two stents | -43200
stent dislocation | -43200
eliminated stent | -43200
replaced stent with inflatable balloon | -43200
X-ray CT examination | -43200
foreign structure ~10 cm in sigmoid colon | -43200
double perforation | -43200
air in peritoneal cavity | -43200
massive inflammation of perivisceral structures | -43200
stent extraction | 0
sigmoidoscopy | 0
colostomy | 0
sigmoidal anus praeter | 0
debridement of scrotum | 0
debridement of peritoneum | 0
distal colon rinsed with saline | 0
sigmoid colon rinsed with saline | 0
no evidence of perforation | 0
surgical necrosis removal | 0
repeated debridement | 0
antimicrobiotic protection | 0
transferred to urologic ward | 24
debridement in urologic ward | 24
suprapubic catheter change | 24
subcutaneous testicle relocation | 24
released with no sign of local infection | 168
recommendation for plastic surgery | 168
scrotal area covered by skin transplantation | 168
periscrotal area covered by skin transplantation | 168
right testicle repositioned into inguinal area | 168
vacuum therapy applied | 168
rejection of transplanted skin | 240
necrosis of transplanted skin | 240
necrotic areas removed | 240
vacuum therapy continued | 240
released from hospital | 240
wound showed granular phenotype | 240
patches changed daily | 240
ileus induced by adhesion pathology | 480
laparotomy with adhesiolysis | 480
released in good mental health | 480
spatial and time oriented | 480
cooperative | 480
stable blood pressure | 480
sustained spontaneous breathing frequency | 480
no visible necrotic tissue | 480
control examination in January 2014 | 2160
operated areas no indications of inflammation | 2160
edges smooth and easily movable | 2160
wounds dry and well covered on right side | 2160
left side smooth pink shiny area with clean edges | 2160
both testicles slightly smaller | 2160
right testicle located in upper femur area | 2160
left testicle located in palpable inguinal area | 2160
scrotal skin slightly raised below penoscrotal angle | 2160
preputium tight | 2160
balanitis developed | 2160
investigation described as painful | 2160
no arbitrary anal sphincter contractions | 2160
recommended stationary intervention | 2160
vacuum patch therapy | 2160
digital cleaning of ampulla recti | 2160
check up on micturition features | 2160
balanitis therapy | 2160
circumcision if required | 2160
ambulant therapy preferred | 2160
suprapubic catheter closed off | 2160
spontaneous micturition via urethra | 2160
Fournier necrotizing fasciitis diagnosis | 0
peripheral necrosis considered septic embolism | 0
septic embolisms lead to acral necrosis | 0
lower extremity amputation | 0
clinical tableau different from Fournier fasciitis | 0
pale marbled skin | 0
patient in shock | 0
acral necrosis | 0
no rotten odor | 0
myositis caused by β#hemolytic group A streptococcus considered | 0
Fournier fasciitis marked by localized pain | 0
streptococcal myositis marked by widespread pain | 0
myalgia misinterpretation | 0
muscle edema later for myalgia | 0
cold skin without obvious erythema | 0
therapeutic approach streptococcal myositis early antibiotics | 0
radical debridement | 0
leg amputation | 0
broad spectrum antibiotics FG | 0
infection resistance occurred | 0
dislocated stent triggering factor | 0
no bowel wall perforation | 0
bacterial colonization favored by immunodeficiency | 0
FG age range 53-58 years | 0
FG increasingly older patients | 0
LRINEC score >8 | 0
increased risk NSTI | 0
high mortality FG | 0
urgent diagnosis required | 0
debridement under antibiotic protection | 0
maggot utilization considered | 0
higher cost maggot treatment | 0
limited compliance maggot treatment | 0
defect not covered with muscle flap | 0
vacuum-assisted closure used | 0
hyperbaric oxygen therapy with VAC considered | 0
HBO inhibits anaerobic bacteria | 0
reduces tissue necrosis extension | 0
HBO favors neutrophilic phagocytic function | 0
HBO angiogenesis | 0
HBO fibroblast proliferation | 0
HBO intracellular antibiotic transport | 0
Grabe et al questionable HBO effect | 0
HBO efficiency not demonstrated | 0
comorbidities treatment important | 0
alcoholism | -43200
malnutrition | -43200
cachexia | -43200
hepatic involvement | -43200
renal involvement | -43200
chronic pancreatitis | -43200
FG cause dislocated stent | 0
immunodeficiency favored by alcoholism | -43200
bacterial multiplication | -43200
necrosis of overlying skin | 0
radiologists did not detect stent on CT | -43200
no bowel perforation confirmed during surgery | 0
laparotomy required | 480
colostomy required | 480
rectal incontinence | -43200
defects not properly cleaned | 0
continuous contamination | 0
sigmoidal anus praeter decision | 0
severe clinical history | -43200
chronic hepatitis | -43200
calcified chronic pancreatitis | -43200
decreased metabolism | -43200
immunodeficiency | -43200
negative nitrogen balance | -43200
Korsakoff’s syndrome | -43200
sensory dysfunction lumbar plexus | -43200
motor dysfunction lumbar plexus | -43200
incontinence | -43200
FG spread to male genital organs | 0
therapeutic challenges | 0
multidisciplinary collaboration required | 0
optimal wound management | 0
lower risk retractile scarring | 0
