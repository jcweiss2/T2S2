63 years old | 0
female | 0
admitted to the hospital | 0
RA | -972
Steinbrocker radiographic stage IV | -756
no history of IM | 0
no hypersensitivity to mosquito bites | 0
cervical and axillary lymphadenopathy | -144
treatment with methotrexate | -144
treatment with infliximab | -144
biopsy of a lymph node | -144
LPD | -144
discontinuation of MTX and IFX | -144
leukocytoclastic vasculitis | -96
antineutrophil cytoplasmic antibody-negative pauci-immune crescentic glomerulonephritis | -96
treatment with etanercept | -96
EBV DNA level 940 copies/106 WBC | -96
anti-EBV VCA IgG 1:320 | -96
anti-EBV VCA IgM negative | -96
anti-EBV EBNA antibody negative | -96
spleen enlargement | -96
lymphadenopathy | -96
CAEBV | -96
initiation of ABT treatment | -540
mild hepatocellular injury | -540
recurrent fever | -240
liver injury | -240
final dose of ABT | -144
persistent liver injury | -120
pancytopenia | 0
admission to the hospital | 0
pulse 101 beats/min | 0
blood pressure 103/52 mmHg | 0
body temperature 37°C | 0
respiratory rate 22 breaths/min | 0
oxygen saturation 99% | 0
Eastern Cooperative Oncology Group Performance Status Grade 4 | 0
tenderness in the right upper quadrant | 0
pancytopenia | 0
liver injury | 0
hyperbilirubinemia | 0
inflammatory response | 0
high levels of ferritin | 0
high levels of soluble interleukin-2 receptor | 0
low levels of IgG | 0
low levels of albumin | 0
normal prothrombin time international normalized ratio | 0
CMV pp65 antigen positive | 0
Aspergillus antigen positive | 0
anti-VCA IgG positive | 0
elevated EBV DNA level | 0
diagnosis of HLH | 0
systemic inflammatory response syndrome | 0
sepsis | 0
treatment with meropenem | 0
treatment with micafungin | 0
treatment with ganciclovir | 0
death | 648
hepatic failure | 648
autopsy | 648
liver atrophy | 648
bridging fibrosis | 648
zonal necrosis of hepatocytes | 648
infiltration of medium-sized to large atypical lymphocytes | 648
infiltration of EBV-infected CTLs | 648
hemophagocytosis | 648
infiltration of atypical lymphocytes in the spleen, lymph nodes, and bone marrow | 648
invasive pulmonary aspergillosis | 648
CMV antigenemia | 648