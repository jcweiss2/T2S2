74 years old|0
    male|0
    admitted to the emergency department|0
    altered mental status|0
    fever|-48
    cough with mucopurulent sputum|-48
    abdominal pain|-48
    hypertension|0
    gastroesophageal reflux|0
    moderate alcohol consumption|0
    lansoprazole|-48
    perindopril|-48
    amlodipine|-48
    disoriented|0
    uncooperative|0
    blood pressure 135/85 mmHg|0
    heart rate 103 beats/min|0
    respiratory frequency 18 breaths/min|0
    peripheral oxygen saturation 85%|0
    tympanic temperature 39.6 °C|0
    livedo reticularis|0
    increased capillary refill time|0
    bilateral rhonchi|0
    intense epigastric pain|0
    right hypochondrium pain|0
    muscle guarding|0
    hypoxic respiratory failure|0
    leukocytosis|0
    neutrophilia|0
    aspartate aminotransferase 1896 U/L|0
    alanine aminotransferase 640 U/L|0
    lactate dehydrogenase 2499 U/L|0
    alkaline phosphatase 230 U/L|0
    total bilirubin 4.78 mg/dL|0
    blood lactate level increased|0
    C-reactive protein increased|0
    procalcitonin 83.86 ng/mL|0
    blood cultures sent|0
    empiric broad-spectrum antibiotics started|0
    piperacillin/tazobactam|0
    abdominal computed tomography scan with contrast|0
    diffuse heterogeneous structure|0
    hypodensity within the right lobe of the liver|0
    two relatively extensive areas with gas|0
    no evidence of abscess formation|0
    no significant changes|0
    emphysematous hepatitis|0
    acute liver failure|0
    severe metabolic acidosis|0
    distributive shock|0
    vasopressor support|0
    admitted to intensive care unit|0
    supportive therapy instituted|0
    clinical state deteriorated|24
    blood analysis deteriorated|24
    antimicrobial spectrum extended|24
    vancomycin|24
    metronidazole|24
    fluconazole|24
    multiorgan failure|48
    death|72
    multi-sensitive Escherichia coli|72

