59 years old | 0
white | 0
female | 0
shortness of breath | -720
exertional dyspnea | -720
cough | -720
weakness in legs | -720
atrial fibrillation | -720
rapid ventricular rate | -720
amiodarone | -720
anticoagulant | -720
hospitalizations for worsening dyspnea | -720
respiratory rate of 27 | 0
SpO2 of 83% on room air | 0
microscopic hematuria | 0
diffuse alveolar hemorrhage (DAH) | 0
positive cytoplasmic anti-neutrophil cytoplasmic antibodies (C-ANCA) | 0
high proteinase 3 IgG | 0
Granulomatosis with Polyangiitis (GPA) suspicion | 0
infectious disease workup | 0
positive qualitative CMV PCR | 0
low viral load in bronchoscopy | 0
concern for active CMV infection was low | 0
rituximab for induction of remission for GPA | 0
high-dose steroids | 0
prophylaxis for Pneumocystis jirovecii pneumonia (PJP) | 0
1 gm of rituximab | 0
ganciclovir | 0
nausea | 0
chills | 0
rigors | 0
IV hydrocortisone | 0
second dose of rituximab (1 gm) | 720
IgG and IgM levels below normal | 744
IgG of 308 mg/dL | 744
IgM 27 mg/dL | 744
no fevers or concern for infection | 744
plan to monitor closely | 744
acute respiratory failure | 1440
septic shock | 1440
E. coli bacteremia | 1440
intubated and sedated | 1440
death | 1440