61 years old | 0
male | 0
admitted to the hospital | 0
systemic erythema | -720
oedema of the lower limbs | -540
allopurinol tablets | -720
systemic rash | -720
gout | -720
elevated white blood cell count | -720
high C-reactive protein | -720
high ALT | -720
drug-induced dermatitis | -720
glucocorticoid | -720
loratadine | -720
cetirizine | -720
rash disappeared | -540
discharged | -540
hypertension | -4380
diabetes mellitus | -120
secondary diabetes | -120
blood pressure 129/86 mmHg | 0
heart rate 124 beats/min | 0
temperature 38.7 °C | 0
respiration 17 breaths/min | 0
saturation 95% | 0
localized red-purplish discoloration | 0
white blood cell count 13.2 × 10^9/L | 0
neutrophilia 93% | 0
hemoglobin 79 g/L | 0
elevated CRP 302 mg/L | 0
procalcitonin 2.84 ng/mL | 0
degraded albumin 24 g/L | 0
high serum creatinine 4.95 mg/dL | 0
elevated B-type natriuretic peptide 1791.6 pg/mL | 0
glycosylated haemoglobin 9.2% | 0
metabolic acidosis | 0
ultrasonography scan | 0
oedema of the dorsum of the feet | 0
intermuscular abscess | 0
magnetic resonance imaging | 24
multiple muscle and subcutaneous soft tissue swelling | 24
intermuscular abscesses | 24
broad-spectrum intravenous antibiotics | 0
cefoperazone sodium/sulbactam sodium | 0
caspofungin | 0
serum albumin | 0
fluids | 0
immunoglobulins | 0
blood glucose monitoring | 0
insulin | 0
ultrasound-guided abscess puncture and drainage | 24
bloody purulent fluid | 24
Gram-positive cocci | 48
Staphylococcus aureus | 48
surgical debridement | 48
necrotic tissue | 48
vacuum sealing drainage | 72
negative pressure | 72
saline | 72
continuous irrigation | 72
second debridement | 168
unhealed right leg | 168
coughed up bloody sputum | 216
short of breath | 216
saturation 93% | 216
oxygen concentration 33% | 216
remarkable wheezes | 216
echocardiography | 216
slight enlargement of the left ventricular cavity | 216
ejection fraction 57% | 216
pericardial effusions | 216
moderate anaemia | 216
elevated brain natriuretic peptide | 216
lactate dehydrogenase | 216
computed tomography scan | 216
acute bilateral pulmonary oedema | 216
pleural effusions | 216
non-invasive positive pressure ventilation | 216
glucocorticoids | 216
diuretics | 216
immunoglobulin | 216
thymosin | 216
red blood cells | 216
erythropoietin | 216
repeated debridement | 336
skin grafting | 2880
discharged | 2880
follow-ups | 4320
well-controlled diabetes | 4320