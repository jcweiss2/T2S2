54 years old | 0
male | 0
presented to the hospital | 0
melena | 0
hemoglobin of 6.7 g/dL | 0
history of transhiatal esophagectomy | -7776
esophageal adenocarcinoma | -7776
esophagogastroduodenoscopy | 0
5-cm clean-based ulcer | 0
ulcer on the anterior surface of the gastric conduit | 0
ischemic etiology | 0
biopsies of the ulcer edge | 0
reactive foveolar mucosa | 0
intraepithelial lymphocytosis | 0
fibrinopurulent exudate | 0
no dysplasia | 0
outpatient surgical referral | 0
discharged | 0
proton pump inhibitors | 0
hematemesis | 720
hemoglobin nadir of 4.8 g/dL | 720
esophagogastroduodenoscopy in the intensive care unit | 720
deeper, hematin-stained ulcer base | 720
rhythmic pulsations | 720
corresponding to cardiac contractions | 720
chest computed tomography | 720
suspicion of ulcer erosion to the heart | 720
urgent thoracic surgery consult | 720
gastrocardiac fistula | 720
intraoperative visualization | 720
large defect in the ventricular wall | 720
bovine pericardial patch | 720
repair of gastrocardiac fistula | 720
failure to wean from mechanical ventilation | -7776
pneumonia | -7776
reintubation | -7776
sepsis | -7776
pulmonary edema | -7776
deep wound infection | -7776
recurrent malignancy | -7776
Candida albicans infection | -7776
severe peptic ulcer disease | -7776
trauma | -7776
sepsis | 720
gastrointestinal bleeding | 720
intermittent bleeding | 720
exsanguination | 720
surgical repair | 720
closing the defect | 720
pericardial patches | 720
surgical management | 720
good outcomes | 720
informed consent | 0