55 years old | 0
male | 0
nonalcoholic steatohepatitis | -672
alpha 1 antitrypsin deficiency | -672
orthotopic liver transplant | 0
incarcerated inguinal hernia | 24
hernia repair | 24
cytomegalovirus viremia | 24
valganciclovir | 24
discharged | 336
mycophenolate mofetil | 0
tacrolimus | 0
prednisone | 0
encephalopathy | 336
increasing home oxygen requirements | 336
sparse speech | 336
disorientation | 336
nonfocal neurologic examination | 336
white blood cell count 9.3 × 10^9/L | 336
creatinine 2.12 mg/dL | 336
blood urea nitrogen 53 mg/dL | 336
arterial ammonia 204 µmol/L | 336
induction dosing of intravenous ganciclovir | 336
empiric antibiotic coverage with vancomycin, meropenem, micafungin | 336
intravenous micronutrient supplementation for B1, B6, and levocarnitine | 336
lumbar puncture | 336
encapsulated yeast suspicious for Cryptococcus | 336
liposomal amphotericin B | 336
flucytosine | 336
continuous renal replacement therapy (CRRT) | 336
rifaximin | 336
zinc | 336
lactulose | 336
ammonia 692 µmol/L | 360
neurological deterioration | 360
mechanical ventilation | 360
empiric intravenous doxycycline | 360
urine and bronchial aspirate for Mycoplasma and Ureaplasma polymerase chain reaction (PCR) | 360
ammonia <100 µmol/L | 432
Cryptococcal serum and cerebrospinal fluid (CSF) antigen titers >1:2560 | 432
cultures from bronchoalveolar lavage, CSF, and blood revealed cryptococcal growth | 432
repeat lumbar punctures | 480
opening pressures greater than 45 cmH2O | 480
large volume drainage | 480
thrombocytopenia | 480
mental status improvement | 528
tracheostomy | 528
persistent hydrocephalus | 576
oliguric renal failure | 576
progressive splenic infarcts with necrosis | 576
splenectomy | 576
sepsis | 624
duodenal leak | 624
renal failure | 624
failure to thrive | 624
comfort care in hospice | 720
urea cycle disorder screening studies | 720
low urine orotic level | 720
normal serum citrulline and arginine level | 720