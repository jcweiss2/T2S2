43 years old | 0
female | 0
presented with continuing fever | -336
lower abdominal pain | -336
foul-smelling discharge from left perianal region | -336
duration of 2 weeks | -336
no previous medical illness | 0
physical examination of the perineum | 0
necrotic tissue | 0
foul-smelling thin pus | 0
surgery | 0
left perianal region debrided | 0
deep pockets of abscess | 0
second postoperative day | 48
lower abdominal pain worsened | 48
ultrasound showed fluid collection | 48
laparotomy | 48
thick abscess in entire anterior abdominal wall | 48
necrotic rectus muscle | 48
superiorly extending to subcostal region | 48
inferiorly extending to retro-pubic space | 48
abscess in peritoneal cavity | 48
laterally extending to para-renal retroperitoneal region | 48
abscess drainage | 48
debridement | 48
abdomen left open with Bogota bag | 48
pockets packed | 48
drainage tubes in situ | 48
transferred to intensive care unit | 48
antibiotics changed to wider spectrum | 48
relaparotomy done 48 hours later | 96
no disease progression | 96
stayed in ICU | 96
continued antibiotics for 2 weeks | 336
on 35th day following initial debridement | 840
15 × 30 cm sub@-umbilical fascia defect | 840
reconstructed with non-vascularized bilateral tensor fascia-lata graft | 840
abdomen closed | 840
secondary closure of perianal wound | 840
3-month follow-up | 2160
6-month follow-up | 4320
9-month follow-up | 6480
computed tomography scan shows normal anterior abdominal fascia | 6480
