29 years old | 0
male | 0
ingested metformin | -5.5
ingested ethanol | -5.5
vomiting | -5.5
diarrhea | -5.5
thirst | -5.5
abdominal pain | -5.5
bilateral leg pain | -5.5
agitated | -5.5
fingerstick glucose level of 180 mg/dL | -5.5
history of psychosis | 0
history of depression | 0
prior suicide attempts | 0
discontinued olanzapine | 0
discontinued sertraline | 0
family history of type II diabetes | 0
daily ethanol use | 0
daily tobacco use | 0
admitted to the Emergency Department | 0
temperature of 35.2°C | 0
pulse of 113 beats/min | 0
blood pressure of 129/59 mmHg | 0
respirations at 28 breaths/min | 0
100% saturation via pulse oximetry on room air | 0
awake and oriented x4 | 0
agitated and slightly confused | 0
GCS=14 | 0
pupils were equal and reactive at 4mm | 0
oral mucous membranes were dry | 0
tachycardia | 0
heart and lung exams were unremarkable | 0
abdomen was mildly tender to palpation diffusely | 0
incontinent of feces | 0
stool was guaiac-negative | 0
normal rectal tone | 0
narrow-complex sinus tachycardia | 0
repeat fingerstick glucose of 364 mg/dL | 0
combative | 0
intravenous lorazepam 2 mg | 0.75
intravenous dolasetron 12.5 mg | 0.75
intravenous morphine sulfate 4 mg | 0.75
hydration with 0.9% saline | 0.75
physical restraints removed | 1
laboratory evaluation | 0.5
serum glucose level of 707 mg/dL | 0.5
elevated anion-gap metabolic acidosis | 0.5
arterial blood gas analysis | 0.5
pH 7.10 | 0.5
pCO2 18.8 mmHg | 0.5
pO2 133.1 mmHg | 0.5
serum lactate level >11.1 mmol/L | 0.5
osmolal gap >20 mOsm/kg | 0.5
urinalysis | 0.5
glycosuria | 0.5
moderate hemoglobin | 0.5
no calcium oxalate crystalluria | 0.5
no blood cells | 0.5
no signs of infection | 0.5
urine drug screen | 0.5
admitted to the medical intensive care unit | 1
nephrology service consulted | 1
repeat laboratory analysis | 4
decreasing bicarbonate | 4
severe hyperglycemia | 4
unresponsive | 5
vomit | 5
aspirate | 5
pulseless electrical activity | 5
heart rate of 29/min | 5
resuscitated | 5
chest compressions | 5
endotracheal intubation | 5
intravenous epinephrine 2 mg | 5
intravenous atropine 1 mg | 5
intravenous sodium bicarbonate 176 mEq | 5
heart rate of 110/min | 5
blood pressure 121/88 mmHg | 5
intra-resuscitative ABG | 5
pH 6.95 | 5
pCO2 55.7 mmHg | 5
pO2 88.1 mmHg | 5
bicarbonate 12.4 mEq/L | 5
bicarbonate drip | 5
transferred to the ICU | 5
non-sustained episodes of ventricular tachycardia | 6
blood pressure fell to 72/44 mmHg | 6
dopamine drip | 6
coagulopathic | 6
INR 3.08 | 6
fibrinogen 113 mg/dL | 6
d-dimer >8.0 mcg/mL | 6
platelet count 390 k/mm3 | 6
hematocrit 47.7% | 6
echocardiogram | 6
mildly decreased left ventricular function | 6
serial cardiac enzymes | 6
elevated CK-MB fraction | 6
elevated troponin I | 6
hemodialysis | 12
PEA recurred | 15
expired | 19
last set of laboratory results | 14
serum lactate level >11.1 mEq/L | 14
bicarbonate 12 mEq/L | 14
glucose 327 mg/dL | 14