60 years old | 0
woman | 0
DM | 0
chronic renal failure | 0
admitted to the hospital | 0
severe pain in upper lip | -96
bullous lesion in upper lip | -96
suspected cellulitis in upper lip | -96
denied special trauma history | 0
suspected zoster infection | 0
antiviral treatment | 0
not regularly adhering to DM medication | 0
serum glucose level of 346 mg/dL | 0
hemoglobin A1c of 7.8% | 0
white blood cell count of 12,000/μL | 0
C-reactive protein level of 93.7 mg/L | 0
sudden chest pain | 12
NSTEMI | 12
moved to intensive care unit | 12
transferred to department of internal medicine | 12
sudden high fever exceeding 38°C | 18
hypotension | 18
mental status deteriorated to stupor | 18
worsened general condition | 18
swelling of upper lip increased | 18
inflammation of upper lip increased | 18
ulcerative lesion on oral mucosa of upper lip | 18
intra-oral wound with foul odor | 18
purulent discharge | 18
white blood cell count of 23,000/μL | 18
C-reactive protein level of 385.8 mg/L | 18
septic shock | 18
blood culture tests | 18
pus culture tests | 18
coronary angiography | 18
3-vessel disease | 18
severe stenosis | 18
intravenous broad-spectrum antibiotics | 18
boosters | 18
adjunctive treatment measures | 18
upper lip gangrene | 48
upper lip necrosis | 48
diffuse gaseous necrosis on facial CT | 48
cutaneous fistula of upper lip | 48
chest CT | 48
persistent dyspnea | 48
abscess-like lung nodule in right upper lobe | 48
septic emboli from upper lip infection | 48
Laboratory Risk Indicator for Necrotizing Fasciitis score of 10 | 48
immediate surgical intervention | 48
debridement under general anesthesia | 48
full-layer necrosis of upper lip | 48
orbicularis oris muscle necrosis | 48
K. pneumoniae confirmed in blood culture | 120
K. pneumoniae confirmed in pus culture | 120
antibiotic regimen with ceftriaxone | 120
antibiotic regimen with metronidazole | 120
serial debridement | 120
purulent discharge ceased | 312
follow-up pus culture confirmed K. pneumoniae | 312
follow-up pus culture confirmed MRSA | 312
full-layer skin defect | 840
soft tissue defect | 840
scar contracture | 840
discharged | 1200
scar release | 4320
Abbe flap coverage | 4320
flap detachment | 5280
flap division | 6240
favorable correction of upper lip drooling | 6240
patient satisfied with results | 6240
