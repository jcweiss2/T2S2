44 years old | 0
female | 0
admitted to the hospital | 0
intermittent headache | -672
progressive memory loss | -672
hypothyroidism | -672
electroconvulsive therapy | -672
major depressive disorder | -672
craniotomy | 0
gross total resection of the right temporal mass | 0
anaplastic astrocytoma | 0
radiation | 0
temozolomide | 0
grade-1 toxicity of the skin | 24
gastritis | 24
lymphopenia | 168
thrombocytopenia | 168
adjuvant temozolomide | 168
Atovaquone | 168
neutropenia | 216
dyspnea | 336
rash | 336
paronychia | 336
severe pancytopenia | 336
platelet transfusion | 336
red blood cell transfusion | 336
cefuroxime | 336
fluconazole | 336
cellulitis | 336
bone marrow biopsy | 336
hypocellular bone marrow | 336
HIV negative | 336
HBV negative | 336
HCV negative | 336
EBV negative | 336
CMV negative | 336
parvovirus negative | 336
B12 supplementation | 336
neutropenic fever | 504
septic shock | 504
Bartholin gland abscess | 504
rectovaginal fistula | 504
broad-spectrum antibiotics | 504
Enterococcus VRE bacteremia | 504
repeat bone marrow biopsy | 504
pan-hypoplasia | 504
granulocyte monocyte-colony stimulating factor | 504
eltrombopag | 504
cord blood stem cell transplantation | 504
fludarabine | 504
melphalan | 504
lung abscesses | 504
pyelonephritis | 504
acute hypoxic respiratory failure | 504
septic shock | 504
multiple organ failure | 504
death | 504