27 years old | 0
    pregnant | 0
    G4P2 | 0
    28th GW | 0
    born in Western Africa | 0
    living in Italy since 2012 | 0
    presented to the emergency department | 0
    headache | 0
    vomiting | 0
    diarrhea | 0
    pelvic pain | 0
    low back pain | 0
    contracted malaria in 2007 | -87600
    slight increase in LDH | 0
    mild anemia | 0
    hemoglobin 9.9 g/dl | 0
    no morphological abnormalities on renal echography | 0
    discharged | 0
    returned due to persistent symptoms | 48
    hyperpyrexia | 48
    admitted to the obstetric ward | 48
    prophylactic ceftriaxone | 48
    peak hyperthermia 39.4℃ | 72
    loss of consciousness | 72
    recovered in 15 minutes | 72
    residual aphasia | 72
    evident cognitive impairment | 72
    improved slowly over a few hours | 72
    no rigor nucalis | 72
    no signs of focal deficit | 72
    no pathological abnormalities of the central nervous system | 72
    respiratory parameters stable | 72
    hemodynamic parameters stable | 72
    SpO2 99% in room air | 72
    BP 135/70 mmHg | 72
    HR 95 bpm | 72
    increased CRP | 72
    increased bilirubin | 72
    increased LDH | 72
    hemoglobin decreased to 7.8 g/dl | 72
    malaria parasites found on peripheral blood smear | 72
    blood parasites 7% | 72
    quinine prescribed | 72
    clindamycin prescribed | 72
    tight control of glycemia | 72
    tight control of BP | 72
    tight control of electrocardiography | 72
    fetal parasitemia suspected | 72
    hemolysis suspected | 72
    cesarean delivery planned | 72
    general condition stable | 72
    no coagulation abnormalities | 72
    platelet count slightly lower than normal | 72
    PLT 98.000 /ml | 72
    lactated Ringer's solution administered | 72
    ranitidine administered | 72
    spinal anesthesia | 72
    hyperbaric bupivacaine 0.5% injected | 72
    sufentanil injected | 72
    anesthetic block reached T4 level | 72
    BP decreased slightly | 72
    BP remained stable throughout surgery | 72
    baby had slight respiratory depression | 72
    Apgar score 8 at 1 and 5 min | 72
    bloodless umbilical cord | 72
    baby weight 1.77 kg | 72
    required immediate oxygen support | 72
    hypoxemia | 72
    SpO2 decreased to <80% | 72
    oxytocin started | 72
    postoperative analgesia | 72
    patient-controlled analgesia pump | 72
    morphine 1 mg/h for 24 h | 72
    acetaminophen prescribed | 72
    surgery uncomplicated | 72
    blood loss estimated 500 ml | 72
    Plasmodium falciparum identified | 168
    blood parasites decreased to 1% | 240
    antibiotic therapy continued | 72
    symptoms resolved two days after childbirth | 96
    oxygen therapy discontinued for baby | 96
    no parasites in baby's blood | 120
    no signs of fetal hemolysis | 120
    