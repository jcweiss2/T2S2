47 years old | 0
    man | 0
    hepatitis C | 0
    hemophilia A | 0
    Factor VIII | 0
    ulcerative colitis | 0
    prednisone | -240
    admitted to MICU | 0
    temperature 34.4°C | 0
    heart rate 96 bpm | 0
    blood pressure 107/51 | 0
    respiratory rate 14 | 0
    oxygen saturation 97% | 0
    cachectic | 0
    abdomen distended | 0
    diffusely tender | 0
    no rebound tenderness | 0
    no guarding | 0
    rectal examination positive for gross blood | 0
    non-contrast abdomen and pelvis CT scan | 0
    pancolitis | 0
    started on antibiotics | 0
    transferred to SICU | 0
    hypotension | 0
    vasopressors | 0
    respiratory failure | 0
    mechanical ventilation | 0
    leukocytosis | -48
    lactic acidosis | -48
    normalized leukocytosis | -24
    normalized lactic acidosis | -24
    weaned off vasopressors | -24
    extubated | -24
    Clostridium difficile antigen negative | -24
    antibiotics narrowed | -24
    sudden onset sharp abdominal pain | -168
    peritoneal signs | -168
    non-contrast abdominal CT scan | -168
    pneumoperitoneum | -168
    colitis | -168
    ascites | -168
    deemed too high a surgical risk | -168
    loop ileostomy | -168
    small bowel normal | -168
    ascites clear | -168
    extubated postoperatively | -168
    initially improved | -168
    supraventricular tachycardia | -240
    respiratory failure requiring mechanical ventilation | -240
    hypotension requiring vasopressors | -240
    large-volume serosanguinous ascites drainage | -240
    ascites cultures grew Candida | -240
    ascites cultures grew Methicillin-resistant Staphylococcus aureus | -240
    ascites cultures grew E. coli | -240
    appropriate antibiotic therapy initiated | -240
    sputum cultures grew 1+ Aspergillus fumigatus | -240
    repeat ET aspirate culture negative for fungus | -240
    non-contrast chest CT scan | -240
    no fungal pneumonia | -240
    intubated | -240
    weaned off vasopressors | -240
    abdominal examination improved | -240
    peritoneal signs | -336
    acute hypotension | -336
    vasopressors | -336
    black ileostomy output | -336
    bleeding from intra-abdominal drain | -336
    bright red blood per rectum | -336
    exploratory laparotomy | -336
    small bowel necrotic | -336
    distal jejunum necrosis | -336
    distal ileum necrosis | -336
    73 centimeters resected | -336
    primary anastomosis | -336
    profuse intra-abdominal bleeding | -360
    hemodynamically unstable | -360
    massive transfusion | -360
    aggressive attempts to correct coagulopathy | -360
    deteriorated | -360
    goals of care changed | -360
    died | -384
    third ET aspirate culture positive for A. fumigatus | -384
    hemorrhagic bowel | 0
    gangrenous bowel | 0
    granular friable mucosa | 0
    ulcerated mucosa | 0
    transmural bowel necrosis | 0
    fungi within bowel wall | 0
    fungi within artery wall | 0
    fungi within lumen | 0
    Gomori Methenamine Silver stain positive | 0