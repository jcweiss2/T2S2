64 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
severe headache | -24 | 0 | Factual
right periorbital and mid-facial swelling | -24 | 0 | Factual
fever | -336 | -168 | Factual
headache | -336 | -168 | Factual
light pain in the right ear | -336 | -168 | Factual
purulent secretion from the ear | -336 | -168 | Factual
swelling and redness of the skin behind the right ear | -336 | -168 | Factual
tinnitus | -336 | -168 | Factual
hearing disorder | -336 | -168 | Factual
right acute mastoiditis | -336 | -168 | Factual
Amoxicillin | -336 | -168 | Factual
painkillers | -336 | -168 | Factual
anti-inflammatory drugs | -336 | -168 | Factual
arterial hypertension | 0 | 0 | Factual
angiotensin-converting enzyme inhibitors | 0 | 0 | Factual
right facial and periorbital swelling | 0 | 0 | Factual
right blepharoptosis | 0 | 0 | Factual
chemosis | 0 | 0 | Factual
proptosis | 0 | 0 | Factual
visual acuity of 7/12 on her right eye | 0 | 0 | Factual
no visual fields abnormalities | 0 | 0 | Factual
normal intraocular pressures | 0 | 0 | Factual
no relative afferent pupillary defect | 0 | 0 | Factual
normal color vision | 0 | 0 | Factual
no signs of optic disc swelling | 0 | 0 | Factual
febrile | 0 | 0 | Factual
conscious | 0 | 0 | Factual
somnolent | 0 | 0 | Factual
no neurological deficits | 0 | 0 | Factual
normal cardiovascular examination | 0 | 0 | Factual
normal respiratory examination | 0 | 0 | Factual
elevated white blood cells count | 0 | 0 | Factual
elevated erythrocyte sedimentation rate | 0 | 0 | Factual
elevated C-reactive protein | 0 | 0 | Factual
normal renal and liver functions | 0 | 0 | Factual
negative tests for vasculitis | 0 | 0 | Factual
negative tests for human immunodeficiency virus | 0 | 0 | Factual
negative tests for diabetes | 0 | 0 | Factual
prothrombin G20210A mutation | 0 | 0 | Factual
normal coagulation profile | 0 | 0 | Factual
normal urinalysis | 0 | 0 | Factual
non-opacification of the right cavernous sinus | 0 | 0 | Factual
Ceftriaxone | 0 | 48 | Factual
Enoxaparin | 0 | 48 | Factual
no corticosteroids | 0 | 0 | Factual
shortness of breath | 96 | 96 | Factual
reduced oxygen saturation | 96 | 96 | Factual
unilateral homogeneous opacification on right lobar lung | 96 | 96 | Factual
air bronchograms | 96 | 96 | Factual
right lobar pneumonia | 96 | 96 | Factual
Amikacin | 96 | 168 | Factual
Piperacillin–Tazobactam | 96 | 168 | Factual
improvement | 168 | 168 | Factual
transfer back to the Service | 168 | 168 | Factual
control contrast-enhanced magnetic resonance angiography | 168 | 168 | Factual
persistence of the lacunar image in the right cavernous sinus | 168 | 168 | Factual
improved ophthalmological symptoms | 168 | 168 | Factual
diminished periorbital swelling | 168 | 168 | Factual
discharged | 336 | 336 | Factual
oral anticoagulant – Acenocoumarol | 336 | 0 | Factual
follow-up CT venogram | 720 | 720 | Factual
full recovery | 720 | 720 | Factual