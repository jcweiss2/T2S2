69 years old | 0
    female | 0
    admitted to the emergency department | -2
    oral ingestion of ∼300 ml Roundup | -2
    vomiting | -2
    lethargy | -2
    conscious | -2
    disoriented | -2
    Glasgow coma scale of 12 | -2
    blood pressure of 91/56 mm Hg | -2
    SpO2 of 91% in room air | -2
    abdominal tenderness | -2
    unremarkable systemic examination | -2
    gastric lavage | -2
    transferred to emergency ICU | 0
    hydration with normal saline | 0
    correction of acidosis with sodium bicarbonate | 0
    arterial blood gas analysis | 0
    serum lactate level of 19.1 mmol/l | 0
    hemoperfusion | 0
    decreased consciousness level | 6
    required ventilatory support | 6
    vasoactive support needed | 6
    BP drop | 6
    total leukocyte count high | 0
    creatinine 122 μmol/l | 0
    glutamic oxalacetic transaminase 212 IU/l | 0
    alanine aminotransferase 307 IU/l | 0
    alkaline phosphatase 1131 IU/l | 0
    creatine kinase 246 U/l | 0
    uncontrolled seizures | 8
    elevated lactate levels | 8
    worsening metabolic acidosis | 8
    norepinephrine 16 µg/kg/min | 8
    metaraminol bitartrate 3 µg/kg/min | 8
    structured fat emulsion injection 50 g/day | 8
    large amount of fluid | 8
    BP remained low | 8
    hemoglobin 185 g/l | 8
    hematocrit 0.55 l/l | 8
    serum creatinine 164 mg/dl | 8
    total protein 59.6 g/l | 8
    albumin 31.6 g/l | 8
    glutamic oxalacetic transaminase 1012 IU/l | 8
    alanine aminotransferase 570 IU/l | 8
    alkaline phosphatase 2152 IU/l | 8
    C-reactive protein 134.7 mg/l | 8
    creatine kinase 7201 U/l | 8
    myoglobin >3769 ng/ml | 8
    IL-6 7411 pg/ml | 8
    IL-10 37.4 pg/ml | 8
    pulmonary effusion | 8
    fluid accumulation in intestinal wall and lumen | 8
    edema in interstitial spaces | 8
    capillary leak syndrome | 8
    CRRT initiation | 8
    plasma infusion 1000 ml | 8
    albumin infusion | 8
    small doses of glucocorticoids | 8
    ulinastatin 0.4 million every 8 h | 8
    increased urine output | 8
    BP stabilization | 8
    CRRT discontinued | 72
    extubated | 168
    transferred out of ICU | 240
    discharged | 480
    no abnormal signs at 3 months | 2160
   