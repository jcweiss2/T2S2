64 years old | 0
female | 0
Han nationality | 0
admitted to the hospital | 0
cough | -360
fever | -120
chest tightness | -120
shortness of breath | -120
stayed in Wuhan | -600
came back to Shenzhen | -120
temperature 37.5 ºC | 0
blood pressure 124/74 mmHg | 0
SpO2 91% | 0
pulse 85 times/min | 0
respiration rate 22 times/min | 0
thick respiratory sounds | 0
no obvious dry or wet rales | 0
white blood cells 5.3 × 10^9/L | 0
neutrophil percentage 78% | 0
lymphocytes 0.9 × 10^9/L | 0
pH 7.45 | 0
PO2 82 mmHg | 0
PCO2 37 mmHg | 0
FIO2 40% | 0
liver and kidney function normal | 0
myocardial enzyme values normal | 0
C reactive protein 52 mg/L | 0
interleukin 6 153 pg/mL | 0
procalcitonin normal | 0
bilateral multi-patchy consolidation | 0
ground-glass opacities | 0
pharyngeal swab nucleic acid test positive | 0
COVID-19 diagnosis | 0
high-flow nasal catheter oxygen therapy | 0
intermittent noninvasive mechanical ventilation | 0
interferon 60 µg twice daily | 0
lopinavir/ritonavir 500 mg twice daily | 0
gamma globulin 10 g once daily | 0
thymalfasin 1.6 mg every 12 h | 0
naltrexone calcium 4100 µg once daily | 0
oxygenation index 200 mmHg | 0
oxygenation index decreased to 150 mmHg | 120
invasive mechanical ventilation | 120
prone position ventilation | 120
oxygenation index 300 mmHg | 120
ribavirin 0.5 intravenous drip twice daily | 120
ceftazidime 2.0 intravenous drip every 8 h | 120
linezolid 600 mg intravenous drip every 12 h | 120
immunoglobulin 300 mL daily | 168
methylprednisolone 60 mg daily | 168
large amount of thin yellow sputum | 168
CT assessment | 168
exudate increased in lungs | 168
C reactive protein 65 mg/L | 168
interleukin 6 56 pg/mL | 168
alveolar lavage fluid galactomannan increased | 168
blood galactomannan increased | 168
1,3 β-glucan level increased | 168
secondary pulmonary aspergillosis suspected | 168
voriconazole 200 mg every 12 h | 168
prone position ventilation stopped | 216
tracheal intubation removed | 216
nucleic acid test negative | 504
discharged from ICU | 504
chest CT showed resolution of infiltrates | 936
discharged | 936