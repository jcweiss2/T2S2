33 years old | 0
male | 0
admitted to the hospital | 0
abdominal pain | -672
distension | -672
bowel obstruction | -672
enterolysis | -672
omentum majus biopsy | -672
exploratory laparotomy | -672
bypass operation | -672
hydrothorax | -672
bilateral thoracentesis | -672
open abdomen | -672
severe intra-abdominal infection | -672
intermittent high fever | 0
cachexia | 0
anti-infection therapy | 0
acid suppression therapy | 0
digestive juices secretion suppression therapy | 0
total parenteral nutrition | 0
double-pipe drainage | 0
enteroatmospheric fistula | 0
high flow of enteric fistula effluent | 0
corrosion on surrounding tissue | 0
corrosion on incision | 0
water electrolyte imbalance | 0
acid-base imbalance | 0
gastrointestinal dysfunction | 0
contamination of exposed wound | 0
exacerbation of infection | 0
sepsis | 0
prolonged hospital stay | 0
increased medical expense | 0
increased mortality | 0
fistula stent implantation | 216
contrast-mediated fistula angiography | 216
decrease in enteric fistula effluent | 216
increase in stool frequency | 216
increase in stool capacity | 216
enteral nutrition restoration | 240
no abnormal discomfort | 240
no obstruction around fistula orifice | 216
drainage fluid reduction | 216
frozen abdomen formation | 432
skin grafting | 432
granulation around EAF | 432
orifice of fistulous tract decrease | 432
orifice enlargement due to position change | 432
butterfly-shaped adhesive application | 432
waiting for definitive intestinal anastomosis | 432
waiting for abdominal closure | 432
hypoalbuminemia | 0
severe intra-abdominal infection diagnosis | 0
enteroatmospheric fistula diagnosis | 0
treatment with fistula stent | 216
skin grafting outcome | 432
patient in good condition | 432
passed crisis | 432
