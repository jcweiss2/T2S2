37 years old | 0
pregnant | 0
G3P2 | 0
admitted to the hospital | 0
breathlessness | -216
feeling generally unwell | -216
non-productive cough | -216
tested positive for COVID-19 | -216
increased work of breathing | -72
denied chest pain | 0
denied calf tenderness | 0
denied orthopnoea | 0
denied paroxysmal nocturnal dyspnoea | 0
asthma | -672
gastric sleeve surgery | -672
hyperemesis gravidarum | -1008
respiratory rate 32 breaths/min | 0
oxygen saturations 95% | 0
heart rate 105 beats/minute | 0
blood pressure 100/60 mmHg | 0
apyrexial | 0
Kussmaul breathing | 0
ketotic breath | 0
unable to complete full sentences | 0
bi-basal crepitations | 0
no wheeze | 0
clinically dehydrated | 0
normal oral glucose tolerance test | -1008
normal glycated haemoglobin A1c | -1008
ECG sinus tachycardia | 0
Chest X-ray COVID-19 pneumonitis | 0
CT pulmonary angiography no pulmonary emboli | 0
WCC 8.4 × 10^9/L | 0
CRP 149 mg/L | 0
urea and electrolytes and liver function tests | 0
arterial blood gas | 0
metabolic acidosis | 0
elevated ketones | 0
high anion gap | 0
diagnosis of starvation ketosis of pregnancy | 0
treatment with intravenous 20% dextrose | 0
treatment with 0.9% sodium chloride | 0
treatment with 1.6% bicarbonate | 0
variable rate insulin infusion | 0
potassium replacement | 0
Pabrinex | 0
resolution of metabolic ketoacidosis | 24
improved work of breathing | 24
RR 26 breaths/min | 24
oxygen saturations 96% | 24
HR 100 beats/min | 24
BP 110/64 mmHg | 24
apyrexial | 24
stopped intravenous 20% dextrose | 24
stopped 0.9% sodium chloride | 24
stopped 1.6% bicarbonate | 24
stopped variable rate insulin infusion | 24
stopped potassium replacement | 24
stopped Pabrinex | 24
commenced low molecular weight heparin | 24
deteriorated oxygen saturations | 144
worsening pneumonitis | 144
pneumomediastinum | 144
right apical pneumothorax | 144
decision to deliver the baby | 144
commenced on ECMO | 144
delivered | 144
baby admitted to special care baby unit | 144
mother decannulated from ECMO | 168
mother discharged from hospital | 192
follow-up 3 months later | 744
mother and baby well | 744