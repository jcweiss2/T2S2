64 years old | 0
male | 0
admitted to the hospital | 0
penetrating abdominal trauma | -22*24
intra-abdominal exsanguinating bleeding | -22*24
duodenal disruption | -22*24
multiple small bowel perforation | -22*24
duodenojejunostomy | -22*24
resection of small bowel | -22*24
anastomosis | -22*24
bleeding control | -22*24
reanastomosis | -22*24
anastomosis failure | -22*24
sepsis | -22*24
multiorgan failure | -22*24
referred to our institution | -22*24
surgical reexploration | 0
duodenojejunal disruption | 0
enteroenteric anastomosis failure | 0
bile-stained fluid in the abdomen | 0
enteroenterostomy | 0
duodenal primary repair | 0
feeding tube placement | 0
massive irrigation | 0
drain tube placement | 0
ventilator weaning | 0
transferred to general ward | 0
enteral feeding | 0
severe retraction of the duodenum | 0
duodenal disruption gap | 0
abdominal wall defect | 0
impossible to close duodenum primarily | 0
impossible to close abdominal wall defect primarily | 0
free flap to repair abdominal wall defect | 0
persistent leakage of gastric, bile, and pancreatic juice | 0
pancreatic duct and bile duct drainage tubes placement | 0
endoscopic retrograde cholangiopancreaticography | 0
covered expandable metallic stent placement | 0
duodenal continuity reestablished | 0
bile and pancreatic juices diverted | 0
stent migration | 5
stent removal | 5
second stent placement | 5
debridement | 12
closure of abdominal wall defect with free flap | 12
duodenostomy | 12
drainage tube placement | 12
endoscopic images | 84
granulation tissue formation | 84
stent removal | 112
pancreatic duct and bile duct drainage tubes removal | 125
oral food intake | 112
abdominal wall defect healed | 112
small enterocutaneous fistula | 112
upper gastrointestinal water-soluble contrast study | 234
good passage of contrast | 234
small enterocutaneous fistula | 234
no significant obstruction | 234