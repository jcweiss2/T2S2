65 years old | 0
male | 0
admitted to the hospital | 0
melena | -24
altered mental status | -24
confusion | -24
incoherent speech | -24
progressive somnolence | -24
profuse diarrhea | -24
dark tarry stools | -24
chronic hepatitis C | 0
polysubstance abuse | 0
chronic alcoholism | 0
binge drinking | -72
blood pressure, 125/100 mmHg | 0
pulse, 135 beats per minute | 0
temperature, 99.2ºF | 0
O2 saturation, 91% on room air | 0
respiratory rate, 18 breaths per minute | 0
mucous membranes were dry | 0
partially healed wound with surrounding erythema on the right knee | 0
no jaundice | 0
no significant findings on the abdominal examination | 0
Murphy’s sign was negative | 0
Glasgow Coma Scale of 8 | 0
intubated in the emergency room | 0
increase in creatinine to 1.5 mg/dL | 0
drop in hemoglobin to 6.7 g/dL | 0
hepatic cirrhosis | 0
heterogeneous and nodular liver | 0
portal hypertension | 0
gastric varices | 0
cellulitis without abscess or gas formation | 0
IV infusion of octreotide | 0
packed red blood cells and platelets | 0
broad-spectrum antibiotics | 0
tachycardia | 0
leukocytosis | 0
systemic inflammatory response syndrome (SIRS) | 0
elevated lactate | 0
hepatic encephalopathy | 0
respiratory failure | 0
concern for bleeding varices | 0
decompensated cirrhosis | 0
admitted to the intensive care unit (ICU) | 0
emergent upper endoscopy | 24
diffuse non-bleeding esophageal and gastric varices | 24
band ligation | 24
octreotide infusion | 0
no further episodes of melena | 48
extubated | 72
return to baseline mentation | 72
bitten by a dog below his right knee | -504
subjective fevers and chills | -504
blood culture collected on admission returned positive for gram-negative rods | 0
Pasteurella multocida | 0
IV ceftriaxone | 120
discharged home | 360