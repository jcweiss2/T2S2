50 years old | 0
male | 0
admitted to the hospital | 0
tick bite on right leg | -168
generalized myalgias | -168
lethargy | -168
dizziness | -168
mitral valve prolapse | 0
chronic anxiety | 0
hyperlipidemia | 0
peak temperature of 101.5 °F | -24
systolic blood pressure of 80 mm Hg | -24
white blood cell count 23.6 10E3/μL | -24
hemoglobin 21.3 g/dL | -24
hematocrit 63.4% | -24
erythrocyte sedimentation rate 1 mm/h | -24
venous doppler without deep vein thrombosis | -24
computed tomography of chest without pulmonary embolism or pneumonia | -24
transthoracic echocardiogram with ejection fraction 56.4% | -24
electrocardiogram showing normal sinus rhythm | -24
Lyme titer negative | -24
admitted to medical intensive care unit | -24
intravenous aztreonam | -24
vancomycin | -24
levofloxacin | -24
pulseless electrical activity arrest | -12
intubated | -12
return of spontaneous circulation | -12
dusky mottling of distal extremities | 0
cool extremities | 0
full and firm extremities | 0
lower extremity pulses with Doppler ultrasound | 0
capillary refill time >3 seconds | 0
right leg lesion concerning necrosis/vasculopathy | 0
vancomycin | 0
tazobactam-piperacillin | 0
doxycycline | 0
norepinephrine drip | 0
vasopressin drip | 0
hemoglobin 22.4 g/dL | 0
hematocrit 65.1% | 0
white blood cell count 34.5 10E3/μL | 0
platelets 167 10E3/μL | 0
lactic acid 7.5 mEq/L | 0
creatinine 2.49 mg/dL | 0
aspartate aminotransferase 433 IU/L | 0
alanine aminotransferase 477 IU/L | 0
alkaline phosphatase 26 IU/L | 0
total bilirubin 0.4 mg/dL | 0
direct bilirubin 0.0 mg/dL | 0
serum albumin <1.5 g/dL | 0
albumin infusions | 0
serum calcium 5.1 mg/dL | 0
intravenous calcium supplementation | 0
fibrinogen 118 mg/dL | 0
D-dimer 16.17 μg/ml | 0
fibrin split products >40 μg/ml | 0
worsening diffuse edema of extremities | 24
inability to perform ankle-brachial index | 24
arterial doppler of bilateral lower extremities | 24
four-compartment right lower extremity fasciotomy | 48
right lateral thigh fasciotomy | 48
right forearm fasciotomy | 48
vacuum-assisted closures applied | 48
compartment syndrome of bilateral lower legs, thighs, forearms | 48
below-knee amputation of right lower extremity | 192
wound VAC changes | 192
closure of wounds | 720
creatine phosphokinase 735 IU/L | -24
creatine phosphokinase 1360 IU/L | 0
creatine phosphokinase peak 33786 IU/L | 24
creatinine 1.2 mg/dL | -24
creatinine 2.5 mg/dL | 0
creatinine 6.61 mg/dL | 24
acute kidney injury | 24
rhabdomyolysis | 24
acute tubular necrosis | 24
continuous renal replacement therapy | 24
transition to intermittent hemodialysis | 336
renal function recovery | 504
furosemide drip | 504
creatinine 1.03 mg/dL | 504
negative infectious workup | 24
low complements C3 31.4 mg/dL | 24
low complements C4 5.5 mg/dL | 24
normalized C3 62.4 mg/dL | 168
normalized C4 14.6 mg/dL | 168
low IgG 148 mg/dL | 24
low IgA 32 mg/dL | 24
low IgM 19 mg/dL | 24
normalized immunoglobulins | 168
serum protein electrophoresis with restriction in gamma region | 24
immunofluorescence showing IgG kappa faint band | 24
monoclonal gammopathy of unknown significance | 24
anti-nuclear antibody titer 1:640 | 24
negative connective tissue disorder workup | 24
hemoglobin 8.5 g/dL | 720
hematocrit 26.7% | 720
fungemia with Candida albicans | 720
treated with micafungin | 720
discharge to acute rehab | 720
idiopathic systemic capillary leak syndrome | 24
no prophylactic therapy | 720
