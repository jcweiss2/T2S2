57 years old | 0
    male | 0
    hepatitis B virus | -3168
    alcoholic liver cirrhosis | -3168
    hepatic failure | -3168
    hospitalized for esophageal varix bleeding | -3168
    hepatic encephalopathy (Child-Pugh grade C) | -3168
    hospitalized again due to variceal bleeding | -2400
    hepatic coma | -2400
    left femoral neck fracture | -2400
    left bipolar hemiarthroplasty | -2400
    decompensated liver cirrhosis aggravated | -2400
    listed as liver transplant candidate (MELD score 28) | -2400
    visited emergency room with painful anal swelling | -2400
    dysuria | -2400
    severe icteric sclera | -2400
    serious abdominal distension | -2400
    hepato&SHORTFORM;renal syndrome | -2400
    admitted to ICU | -2400
    painful anal swelling progressed | -2400
    necrosis progressed | -2400
    diagnosed with Fournier’s gangrene | -2400
    wide debridement of wound | -2400
    T-colostomy performed | -2400
    bleeding control surgery performed | -2400
    norepinephrine administered | -2400
    vasopressin administered | -2400
    bleeding control repeated | -2400
    deceased donor liver transplantation (DDLT) performed | 0
    Enterococcus faecium detected in blood | 0
    Candida albicans detected in blood | 0
    gangrene wound debris studied | 0
    vancomycin-resistant Enterococcus (VRE) present in blood | 0
    C. albicans present in blood | 0
    Achromobacter xylosoxidans present in wound | 0
    Pseudomonas aeruginosa present in wound | 0
    VRE present in wound | 0
    varix bleeding continued | 0
    wound bleeding continued | 0
    coagulopathy | 0
    hemoglobin level dropped to 3 g/dL | 0
    repeated blood transfusions | 0
    bacterial infections improved with antibiotics | 0
    necrotic wound care | 0
    infection status controlled | 0
    tazocin administered | -2400
    meropenem administered | -2400
    vancomycin added after transplantation | 0
    tazocin administered post-surgery | 0
    teicoplanin administered post-surgery | 0
    amphotericin B administered | 0
    micafungin administered | 0
    C-reactive protein levels decreased | 0
    recovered after DDLT | 0
    immunosuppressant regimen (FK-506, mycomofetil, steroids) | 0
    FK-506 trough level adjusted (4-6 ng/mL) | 0
    