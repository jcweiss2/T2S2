40 years old | 0
female | 0
admitted to the hospital | 0
facial and neck swelling | 0
abdominal discomfort | 0
chief complaint of facial and neck swelling and abdominal discomfort | 0
clindamycin treatment | -48
presumed tooth abscess | -48
swelling of face and neck worsened | 0
endotracheally intubated | 0
mechanical ventilation | 0
CT scan of neck | 0
necrotizing fasciitis | 0
soft tissue edema | 0
gas formation | 0
retropharyngeal abscess | 0
tachycardic | 0
tachypneic | 0
blood pressure of 89/41 mmHg | 0
MAP of 69 mmHg | 0
WBC count of 6.7 | 0
H&H of 12.5/37.2 | 0
creatinine of 1.8 | 0
lactic acid level of 2.9 | 0
central venous line placement | 0
3 liters of IV fluids infused | 0
consultation with ENT and Pulmonology | 0
transferred to ICU | 0
fluid resuscitated | 0
sedated on Versed | 0
physical examination | 0
marked swelling of the neck | 0
rhonchorous breath sounds | 0
severe sepsis | 0
multiple organ dysfunction syndrome | 0
Intravenous Fentanyl initiated | 0
additional 1 liter of 0.9% Sodium Chloride | 0
clindamycin started | 0
piperacillin-tazobactam started | 0
vancomycin started | 0
heparin started | 0
pantoprazole started | 0
Levophed infusion started | 0
ENT surgically debrided the neck region | 0
submandibular and anterior neck incisions packed | 0
two teeth removed | 0
right radial arterial line placed | 0
CT chest showed small pericardial effusion | 24
moderate bilateral pleural effusions | 24
loculation on the left side | 24
ground glass opacities | 24
nodular consolidation | 24
acute lung injury/ARDS | 24
bilateral chest tubes placed | 24
tracheostomy performed | 96
percutaneous enterogastrostomy (PEG) tube placed | 96
pericardiocentesis performed | 240
PICC line placed | 240
aerobic and anaerobic culture results | 240
Clostridium subterminale isolated | 240
pleural fluid culture results | 336
sensitivity to ampicillin-sulbactam | 336
sensitivity to cefoxitin | 336
sensitivity to meropenem | 336
sensitivity to metronidazole | 336
sensitivity to penicillin | 336
infectious disease consultation | 336
piperacillin-tazobactam treatment | 336
maintenance enteral antibiotic therapy | 336
chest tubes removed | 624
discharged to subacute rehab | 888