47 years old | 0
    male | 0
    admitted to the hospital | 0
    chest pain | -27
    worked at a lobster catering company | 0
    heart stent implantation | - (assumed prior event, timestamp unknown)
    hypertension | - (assumed prior event, timestamp unknown)
    smoking index of 500 | 0
    dull pain in left chest | -27
    shortness of breath after activity | -27
    chest pain aggravated upon deep inhalation | -27
    chest pain aggravated upon turning over | -27
    symptoms relieved by nitroglycerin | -27
    symptoms reappeared 1-2 hours later | -27
    electrocardiogram normal | 0
    troponin T normal | 0
    referred to department of cardiology | 0
    chest CT revealed inflammation in lower lobes of both lungs | 0
    chest CT revealed inflammation in inferior lingular segment of left lung | 0
    chest CT revealed left pleural effusion | 0
    intravenous ceftazidime administered | 0
    consciousness clear | 0
    left lower lung dullness on percussion | 0
    left lung breath sounds low | 0
    no rales heard in both lungs | 0
    transferred to department of respiratory and critical care medicine | 48
    intravenous levofloxacin administered | 48
    ultrasound-guided thoracentesis drainage | 96
    pleural effusion ADA 50.3 U/L | 96
    pleural effusion LDH 2523 U/L | 96
    pleural effusion protein 49.64 g/L | 96
    no bacteria in pleural fluid | 96
    no tumor cells in pleural fluid | 96
    antibiotics adjusted to ceftazidime and moxifloxacin | 120
    peak body temperature rise | 120
    antibiotics adjusted to meropenem and moxifloxacin | 192
    re-examination chest CT showed pleural effusion increased | 216
    CRP reexamined | 216
    ESR reexamined | 216
    blood routine reexamined | 216
    no significant changes in reexamination | 216
    bronchoscopy performed | 336
    alveolar lavage collected | 336
    mNGS analysis performed | 336
    fever disappeared | 336
    mNGS revealed Gardnerella vaginalis infection | 384
    mNGS revealed Corynebacterium urealyticum infection | 384
    sputum culture negative | 0
    blood culture negative | 0
    urine culture negative | 0
    discharged from hospital | 432
    chest CT before discharge showed pleural effusion wrapped | 432
    chest CT before discharge showed effusion slightly reduced | 432
    ornidazole prescribed post-discharge | 432
    chest CT follow-up showed inflammation absorbed | 960
    chest CT follow-up showed pleural effusion reduced | 960
    ornidazole regimen extended | 960
    chest tightness absent | 2400
    discomfort absent | 2400
    chest CT follow-up showed inflammation absorbed | 2400
    <|eot_id|>
    