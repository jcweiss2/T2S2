70 years old | 0
female | 0
admitted to the Plastic Surgery department | 0
fever | -24
dizziness | -24
unstable angina | -3360
diabetes mellitus | -3360
skin flap operation | -192
third-degree burn | -336
sore at the sacral area | -720
osteomyelitis | -720
fever | 0
temperature of 38.2℃ | 0
intermittent fever | 0
blood pressure 110/80 mmHg | 0
pulse 78/min | 0
respiratory rate 20/min | 0
peripheral white blood cell count 8,730/µL | 0
hemoglobin level 8.6 g/dL | 0
platelet count 261,000/µL | 0
AST/ALT 7/11 U/L | 0
alkaline phosphatase 77 U/L | 0
blood urea nitrogen/creatinine 23.4/1.42 mg/dL | 0
total protein/albumin 5.6/2.9 g/dL | 0
erythrocyte sedimentation rate increased | 0
C-reactive protein increased | 0
urine yellow and turbid | 0
WBC in urine positive | 0
protein in urine positive | 0
WBCs in urine >60 | 0
yeast organisms in urine | 0
right pleural thickening | 0
collapse of the right lower lung | 0
cystitis | 0
fluid collection in abdomen and pleural cavity | 0
blood culture negative | 0
urine culture positive for Candida albicans | 0
fever | 768
blood culture negative | 768
urine culture positive for K. pneumoniae | 768
treated with ertapenem | 0
treated with tigecycline | 768
treated with colistin | 1344
expired | 2160
septic shock | 2160
multiorgan failure | 2160