87 years old|0
female|0
hypertension|0
paroxysmal atrial fibrillation|0
diabetes mellitus type I|0
hypothyroidism|0
sick sinus syndrome|0
pacemaker placement|0
total abdominal hysterectomy|0
multiple caesarean deliveries|0
cholecystectomy|0
hernia repair|0
presented with signs and symptoms of left knee septic arthritis|0
bilateral conjunctivitis|0
swelling in one of her hand joints|0
swelling in the first metatarsophalangeal joint of her left foot|0
fevers|-96
episodic altered mental status|-96
denied sore throat|0
denied dysphagia|0
denied odynophagia|0
denied hoarseness|0
denied other esophageal symptoms|0
bilateral conjunctival erythema|0
mild mucopurulent discharge|0
irregular heart rhythm|0
left knee swollen|0
left knee erythematous|0
left knee tender on passive extension and flexion|0
elevated white blood cell count|0
high erythrocyte sedimentation rate|0
elevated C-reactive protein|0
inconclusive transthoracic echocardiography|0
transesophageal echocardiography performed|0
intravenous sedation with midazolam|0
pharyngeal local anesthesia with benzocaine|0
esophageal transducer introduced blindly|0
diagnostic images obtained|0
moderate distress|0
nausea|0
vomiting|0
severe chest pain|0
severe back pain|0
urgent chest radiography|0
Gastrografin study performed|0
upper third esophageal perforation|0
contrast seen immediately above the gastroesophageal junction|0
esophagogastroduodenoscopy performed|0
mucosal tear confirmed|0
moderate to severe inflammation throughout the esophagus|0
no obvious bleeding|0
WallFlex stent placed|0
transferred to intensive care unit|0
Diflucan started|0
broad-spectrum antibiotics started|0
repeat Gastrografin esophagram after 2 days|48
no leakage|48
liquid diet started|48
respiratory failure|168
multiorgan failure|168
palliative care decided|168
expired|168
