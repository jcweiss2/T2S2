43 years old | 0
female | 0
admitted to the hospital | 0
right upper quadrant pain | 0
fevers | 0
vomiting | 0
raised inflammatory markers | 0
raised bilirubin | 0
cholelithiasis | -672
choledocholithiasis | -672
ERCP | 24
cannulation of common bile duct | 24
sphincterotomy | 24
CBD stent placement | 24
laparoscopic cholecystectomy | 168
repeat ERCP | 2160
stent removal | 2160
balloon sweep | 2160
CBD stones removal | 2160
right shoulder tip pain | 2160
worsening RUQ pain | 2164
tachycardia | 2164
subcapsular hepatic hematoma | 2164
mass effect on inferior vena cava | 2164
CT scan | 2164
close observation | 2164
repeat hemoglobin testing | 2164
non-operative management | 2164
stable subcapsular hematoma | 2172
discharged | 2172
re-presented to emergency department | 2177
shortness of breath | 2177
new fevers | 2177
malaise | 2177
lethargy | 2177
sepsis | 2177
new oxygen requirement | 2177
repeat CT imaging | 2177
pleural effusion | 2177
admitted to intensive care | 2177
treated for infected subcapsular hematoma | 2177
IR guided drainage | 2177
no improvement | 2184
laparoscopic washout | 2191
necrosectomy | 2191
de-roofing | 2191
drainage of purulent liquid | 2191
necrotic debris | 2191
old blood | 2191
partial necrosectomy | 2198
liver capsule | 2198
thorough irrigation | 2198
no bile leak | 2198
sump drain placement | 2198
Blake drains placement | 2198
continued irrigation | 2198
IV antibiotics | 2198
Klebsiella oxytoca | 2198
Escherichia coli | 2198
acute kidney injury | 2208
antibiotic toxicity | 2208
supratherapeutic antibiotic level | 2208
acute tubular necrosis | 2208
AKI resolved | 2216
discharged | 2216
sump drain in situ | 2216
regular follow-up | 2224
sump drain removal | 2232
no long-term complications | 2232