58 years old | 0  
    woman | 0  
    hypertension | 0  
    diabetes mellitus | 0  
    hypothyroidism | 0  
    Hodgkin lymphoma | -87600  
    radiation therapy | -87600  
    metformin | 0  
    aspirin | 0  
    levothyroxine | 0  
    metoprolol | 0  
    dyspnea on exertion | -336  
    blood pressure 96/60 mmHg | 0  
    heart rate 110 beats per minute | 0  
    oxygen saturation 96% | 0  
    clear lung fields | 0  
    elevated jugular venous pressure | 0  
    faint and distant heart sounds | 0  
    weak peripheral pulses | 0  
    low voltage on ECG | 0  
    sinus tachycardia | 0  
    cardiomegaly on chest X-ray | 0  
    large circumferential pericardial effusion | 0  
    end diastolic right ventricular compression | 0  
    swing sign | 0  
    pericardiocentesis | 0  
    drainage of 2200 mL serous fluid | 0  
    minimal hemodynamic improvement | 0  
    worsening dyspnea | 24  
    hypotension 72/40 mmHg | 24  
    labored breathing | 24  
    diffuse bilateral pulmonary edema | 24  
    intubation | 24  
    hypoxic respiratory failure | 24  
    dobutamine | 24  
    norepinephrine | 24  
    resolved pericardial effusion | 24  
    low-normal LVEF 50% | 24  
    mild to moderately dilated right ventricle | 24  
    mild RV hypokinesis | 24  
    septal shift towards left ventricle | 24  
    intravenous saline bolus | 24  
    vasopressors | 24  
    inotropes | 24  
    diuresed with intravenous lasix | 24  
    hemodynamic improvement | 72  
    extubation | 72  
    normalized ventricular function | 120  
    trivial/minimal pericardial effusion | 120  
    discharged | 144  
    pericardial decompression syndrome | 24  
    pulmonary edema | 24  
    respiratory failure | 24  
    transient ventricular dysfunction | 24  
    supportive management | 24  
    spontaneous gradual improvement | 72  
    hemodynamic support weaned | 72  
    CT-chest angiography | 24  
    no pulmonary embolism | 24  
    interval improvement in pulmonary edema | 24