36 years old | 0
    male | 0
    admitted to the emergency room | 0
    abdominal pain | 0
    vomiting | 0
    septic shock | 0
    norepinephrine application | 0
    peripheral ischemia of four extremities | -120
    right knee disarticulation | -1320
    left trans-femoral amputation | -1320
    right elbow disarticulation | -1320
    skin flap operation of right knee | -1464
    left hand skin defect area operation | -1464
    joint range of motion exercise | -1464
    isometric exercise | -1464
    admitted to Severance Rehabilitation Hospital | 0
    prostheses measurement | 0
    rehabilitation program initiation | 0
    depression | -720
    antidepressant medication | -720
    anorexia | -720
    sociophobia | -720
    right elbow disarticulation site club shape | 0
    right knee disarticulation cylindrical shape | 0
    left trans-femoral amputation conical shape | 0
    phantom pain | 0
    phantom sensation | 0
    left hand 2nd, 3rd, 4th, 5th distal interphalangeal joint disarticulation | 0
    skin flap fragility | 0
    blisters due to friction | 0
    passive range of motion left wrist flexion 40° | 0
    passive range of motion left wrist extension 30° | 0
    1st web space length 2 cm | 0
    left hand stretching exercise | 0
    contracture of left hand | 0
    weakness of left hand | 0
    inability to do opposition | 0
    tip pinch using thumb and 2nd finger | 168
    MMT grade 4 bilateral shoulder joints | 0
    MMT grade 3 left elbow and wrist joints | 0
    MMT grade 2 left hand | 0
    MMT grade 3 hip joints | 0
    left hand muscle power improved to grade 3 | 168
    hip joint muscle power improved to grade 4 | 168
    Cybex isokinetic training | 168
    deconditioning | 0
    impaired pulmonary function | 0
    VC 3,480 mL | 0
    PCF 450 mL | 0
    Ambu bag training | 168
    air stacking exercise | 168
    VC improved to 5,300 mL | 168
    PCF improved to 650 mL | 168
    right elbow disarticulation prosthesis fitting | 336
    elbow flexion device control unit | 336
    elbow lock control cable | 336
    outside locking hinge | 336
    constant friction wrist unit | 336
    figure of 8 harness | 336
    artificial hand use | 336
    bimanual activity training | 336
    sound left hand as dominant hand plan | 336
    left hand pinch power 1.8 kg | 336
    Box and Block Test 33 points | 336
    left wrist flexion 50° | 336
    left wrist extension 50° | 336
    skin fragility | 336
    contracture remaining | 336
    right hand as dominant hand plan | 504
    wheelchair measurement | 504
    ADL training with prostheses | 504
    sitting balance good | 0
    FIM self care subunit 6 points | 0
    intensive ADL training | 504
    don upper prosthesis by himself | 504
    dressing minimal assistance | 504
    eating minimal assistance | 504
    grooming minimal assistance | 504
    spoon use training | 504
    drinking with a cup training | 504
    buttoning and unbuttoning training | 504
    FIM score improved to 12 after 1 month | 672
    FIM score improved to 25 on discharge | 1344
    upper dressing by himself | 1344
    dominant leg right leg decision | 672
    height reduced to 162 cm | 672
    right knee disarticulation prosthesis fitting | 1008
    left trans-femoral amputation prosthesis fitting | 1344
    parallel bar weight shift training | 1512
    gait training with anterior walker | 1680
    walked 100 m without pause | 1680
    left leg dragged on swing phase | 1680
    left leg shortened | 1680
    multidisciplinary team meetings | 168
    cane gait difficulty | 1680
    walker indoors | 1680
    electronic wheelchair outdoors | 1680
    stump site management education | 1680
    ADL training for work | 1680
    car rental for disabled | 1680
    driver's seat movement training | 1680
    short distance driving training | 1680
    computer mouse use | 1680
    universal cuff for typing | 1680
    FIM score 90 on discharge | 1680
    Modified Barthel Index 56 on discharge | 1680
    absolute bed rest status | 0
    sit by himself | 1680
    discharge | 1680
    follow-up after discharge | 1680
    back to work | 1680
    ADL independency on wheelchair level | 1680

<|eot_id|>
