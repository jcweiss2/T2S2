43 years old | 0
male | 0
adrenocorticotrophic hormone (ACTH)-secreting pituitary carcinoma | -672
cerebellar and cervical drop metastases | -672
surgery | -672
radiotherapy | -672
ketoconazole | -672
pasireotide | -672
cabergoline | -672
bilateral (subtotal) adrenalectomy | -672
temozolomide chemotherapy | -672
ipilimumab | -24
nivolumab | -24
maintenance therapy with nivolumab | -24
residual endogenous cortisol production | -24
upper respiratory tract symptoms | -168
progressive dyspnoea | -72
consulted emergency department | 0
severe respiratory complaints | 0
tested positive for SARS-CoV-2 | -24
O2 saturation 72% | 0
tachypnoea (40/min) | 0
bilateral pulmonary crepitations | 0
temperature 37.2°C | 0
blood pressure 124/86 mmHg | 0
pulse rate 112 bpm | 0
high-flow oxygen therapy | 0
insufficient improvement | 0
intubated | 0
type 1 respiratory insufficiency | 0
PaO2 of 52.5 mmHg | 0
PaCO2 of 33.0 mmHg | 0
pH of 7.47 | 0
P/F ratio of 65.7 | 0
C-reactive protein level of 275.7 mg/L | 0
white blood cell count of 7.1 × 10⁹ per L | 0
neutrophils 72.3% | 0
plasma ACTH-cortisol level 213 ng/L | -24
plasma cortisol level 195 µg/L | -24
dexamethasone therapy | 0
broad-spectrum antibiotics | 0
thromboprophylaxis with low molecular weight heparin | 0
ketoconazole restarted | 264
hydrocortisone | 0
block-replacement regimen | 0
multiple organ involvement | 24
metabolic acidosis | 24
acute renal failure | 24
continuous venovenous hemofiltration | 24
acute coronary syndrome type 2 | 24
septic thrombophlebitis of the right jugular vein | 24
critical illness polyneuropathy | 24
readmitted to ICU | 168
ventilator-associated pneumonia | 168
central line-associated bloodstream infection | 168
discharged from hospital | 720
rehabilitation | 720
plasma cortisol level 547 µg/L | 504
plasma ACTH level 130 ng/L | 504