17 years old | 0
female | 0
admitted to hospital | 0
abdominal pain | 0
fever | 0
severe sideropenic anemia | 0
diarrhea | 0
ulcerative colitis | 0
mesalamine treatment | 0
discharged home | 168
fever | 216
sore throat | 216
right neck swelling | 216
right neck tenderness | 216
Group A streptococcal rapid antigen test | 216
viral pharyngitis diagnosis | 216
neck swelling enlarged | 222
pain severe | 222
came to emergency department | 240
physical examination | 240
right sided supraclavicular edema | 240
reduced neck movement | 240
red tonsils | 240
spleen palpable | 240
elevated leukocytes | 240
elevated platelets count | 240
inflammatory markers elevated | 240
coagulation test results slightly out of reference range | 240
neck ultrasound | 240
complete thrombosis of right external and internal jugular veins | 240
thrombus within right subclavian vein | 240
neck magnetic resonance imaging | 240
MRI venography | 240
thrombosis of right subclavian vein | 240
thrombosis of right jugular veins | 240
thrombosis of truncus brachiocephalicus | 240
partial thrombosis of right sigmoid and transverse sinus | 240
bilateral pleural effusion | 240
apical pericardial effusion | 240
normal contractility of heart | 240
Lemierre syndrome diagnosis | 240
intravenous antibiotics treatment | 240
subcutaneous low-molecular-weight heparin | 240
paired blood cultures | 240
throat swabs | 240
became afebrile | 312
comprehensive thrombophilia testing | 312
factor V Leiden normal | 312
protein C normal | 312
protein S normal | 312
factor VIII normal | 312
antithrombin III normal | 312
antinuclear antibodies negative | 312
anticardiolipin antibodies negative | 312
homocysteine levels normal | 312
F2 gene mutation not found | 312
FV Leiden mutation not found | 312
discharged from hospital | 720
anticoagulation therapy at home | 720
low-molecular-weight heparin replaced by apixaban | 4320
follow-ups showed amelioration of neck edema | 4320
neck ultrasound and color doppler showed regression of thrombosis | 4320
recanalization of jugular vein | 4320
ulcerative colitis in clinical remission | 4320
Paediatric Ulcerative Colitis Activity Index 0 | 4320
normal calprotectin levels | 4320
no signs of anemia | 4320