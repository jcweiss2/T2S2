48 years old | 0
male | 0
admitted to the hospital | 0
toothache | -96
dyspnea | -96
chest pain | -96
sweating | -96
tachyarrhythmia | -96
sore throat | -96
fever | -96
gross swelling of the lower right cheek | 0
submandibular and mental regions erythematous and warm on palpation | 0
difficulties in opening the jaw | 0
inflammatory changes of the mucous membrane of the oral cavity | 0
treated with ceftriaxone-steroids-based | -96
ineffective treatment | -48
worsened condition | -48
dyspnea | -48
chest pain | -48
increased WBC count | 0
neutrophils | 0
C-reactive protein | 0
orotracheal intubation | 0
left pleural effusion | 0
mediastinitis | 0
right parapharyngeal abscess | 0
drainage of the right neck | 0
left chest drain | 0
intravenous antibiotic therapy with piperacillin sodium plus tazobactam sodium | 0
worsened clinical condition | 48
transferred to Intensive Care Unit | 48
air collection in the right submandibular | 48
air collection in the left carotid | 48
air collection in the retroesophageal and pretracheal spaces | 48
cervical necrotizing fasciitis with DNM | 48
bilateral pleural effusions | 48
additive pleural drain | 72
abscesses in the cervical spaces | 72
extensive mediastinal empyema | 72
left pleural effusion | 72
right hydropneumothorax | 72
aggressive mediastinal debridement | 72
VATS | 72
incision and drainage of the neck abscesses | 72
oral tooth extraction | 72
purulent fluid drainage | 72
Streptococcus anginosus | 72
Gemella morbillorum | 72
Staphylococcus lugdunensis | 72
antibiotic therapy with amoxicillin | 72
antibiotic therapy with metronidazole | 72
dismissed in better health conditions | 168