41 years old | 0
    woman | 0
    admitted to the hospital | 0
    ischemic stroke over the left corona radiata | -2160
    ischemic stroke over the bilateral frontal lobe | -2160
    ischemic stroke over the parietal lobe | -2160
    bilateral internal carotid artery occlusion (BICAO) | -2160
    right hemiplegia | -2160
    Broca’s aphasia | -2160
    T1DM (Type 1 Diabetes Mellitus) | -26208
    hypertension | -43824
    hyperlipidemia | -35064
    hyperthyroidism | -26304
    methimazole | -2160
    aspirin | -2160
    atorvastatin | -2160
    regular subcutaneous insulin injections | -2160
    transferred for further rehabilitation | 0
    right hemiplegia (persisted) | 0
    ambulate with quad cane | 0
    consciousness alert | 0
    Broca’s aphasia (persisted) | 0
    body temperature 36.1 °C | 0
    pulse 84 beats/min | 0
    blood pressure 125/78 mmHg | 0
    breathing 18 breaths per minute | 0
    right central facial palsy | 0
    Brunnstrom stage III/III (upper limb) | 0
    Brunnstrom stage IV (lower limb) | 0
    self-feeding | 0
    dizziness | 24
    vomiting | 24
    Kussmaul breathing | 24
    lowered response to verbal commands | 24
    hyperglycemia (344 mg/dL) | 24
    arterial blood gas metabolic acidosis (pH 7.255) | 24
    ketone 3+ | 24
    DKA (Diabetic Ketoacidosis) | 24
    transferred to ICU | 24
    aggressive hydration | 24
    insulin pump | 24
    bicarbonate infusion | 24
    electrolyte correction | 24
    serum ketone body 5.5 mmol/L | 72
    consciousness alert (post DKA) | 72
    metabolic acidosis with respiratory compensation | 24 to 120
    comatose | 144
    hemodynamic instability | 144
    acute infarction over bilateral MCA and ACA territories | 144
    brain swelling | 144
    midline shift | 144
    occlusion of bilateral ICA | 144
    glycerol administration | 144
    endotracheal intubation | 144
    normal left ventricle contractility | 144
    no thrombus or vegetation | 144
    respiratory failure | 144
    severe hyperglycemia | 144
    coma (day 6 to 29) | 144 to 696
    mechanical ventilation | 144
    compassionate extubation | 696
    expired | 696
    WBC 8600/μL | 24
    neutrophil 61.2% | 24
    hemoglobin 14.3 g/dL | 24
    platelet 250000/μL | 24
    sodium 134 mmol/L | 24
    potassium 4.3 mmol/L | 24
    creatinine 0.75 mg/dL | 24
    CRP 1.345 mg/dL | 24
    WBC 16600/μL | 96
    neutrophil 89% | 96
    hemoglobin 13.5 g/dL | 96
    platelet 356000/μL | 96
    sodium 148 mmol/L | 96
    potassium 3.1 mmol/L | 96
    creatinine 0.74 mg/dL | 96
    WBC 32510/μL | 144
    neutrophil 87% | 144
    sodium 146 mmol/L | 144
    potassium 3.4 mmol/L | 144
    WBC 19890/μL | 192
    neutrophil 70.8% | 192
    hemoglobin 13.8 g/dL | 192
    platelet 181000/μL | 192
    sodium 166 mmol/L | 192
    potassium 3.8 mmol/L | 192
    creatinine 1.59 mg/dL | 192
    WBC 18930/μL | 336
    neutrophil 75% | 336
    hemoglobin 11.7 g/dL | 336
    sodium 152 mmol/L | 336
    potassium 4.3 mmol/L | 336
    creatinine 2.94 mg/dL | 336
    WBC 13520/μL | 408
    neutrophil 81.3% | 408
    hemoglobin 10.3 g/dL | 408
    platelet 472000/μL | 408
    sodium 154 mmol/L | 408
    potassium 3.6 mmol/L | 408
    creatinine 2.49 mg/dL | 408
    WBC 13870/μL | 528
    neutrophil 59.2% | 528
    hemoglobin | 528
    sodium | 528
    potassium | 528
    creatinine 1.55 mg/dL | 528
    Free T4 1.04 ng/dL | 24
    TSH 2.58 μIU/mL | 24
    T3 53.5 ng/dL | 24
    Complement C3 70.9 mg/dL | 168
    Complement C4 21 mg/dL | 168
    ANA 1:80X | 168
    Anti-dsDNA 62.33 IU/mL | 168
    ANCA negative | 168
    no recurrent stroke | -2160 to 0
    no urinary tract infection | -2160 to 0
    no pneumonia | -2160 to 0
    no new limb weakness | 24
    no pyuria | 0
    normal thyroid function | 24
    no bacteremia | 24 to 144
    no urinary tract infection | 24 to 144
    no gastroenteritis | 24 to 144
    no pneumonia | 24 to 144
    no drop in blood pressure | 144
    no moyamoya disease | 144
    no sinus rhythm (ECG) | 144
    no vegetations (echocardiogram) | 144
    no autoimmune-related stroke | 168
    no diet control issues | -26208 to 0
    no glycemic control issues | -26208 to 0
    no regular aerobic exercise | -26208 to 0
    no prior infection | -2160 to 0
    no trauma | -2160 to 0
    no myocardial infarction | -2160 to 0
    no pancreatitis | -2160 to 0
    no psychological stress | -2160 to 0
    no inadequate insulin treatment | -2160 to 0
    no noncompliance | -2160 to 0
    no cerebral edema | 24 to 696
    no noncardiogenic pulmonary edema | 24 to 696
    no hypoglycemia episodes | -26208 to 0
    no alternative stroke etiologies | 144

    41 years old | 0
    woman | 0
    admitted to the hospital | 0
    ischemic stroke over the left corona radiata | -2160
    ischemic stroke over the bilateral frontal lobe | -2160
    ischemic stroke over the parietal lobe | -2160
    bilateral internal carotid artery occlusion (BICAO) | -2160
    right hemiplegia | -2160
    Broca’s aphasia | -2160
    T1DM (Type 1 Diabetes Mellitus) | -26208
    hypertension | -43824
    hyperlipidemia | -35064
    hyperthyroidism | -26304
    methimazole | -2160
    aspirin | -2160
    atorvastatin | -2160
    regular subcutaneous insulin injections | -2160
    transferred for further rehabilitation | 0
    right hemiplegia (persisted) | 0
    ambulate with quad cane | 0
    consciousness alert | 0
    Broca’s aphasia (persisted) | 0
    body temperature 36.1 °C | 0
    pulse 84 beats/min | 0
    blood pressure 125/78 mmHg | 0
    breathing 18 breaths per minute | 0
    right central facial palsy | 0
    Brunnstrom stage III/III (upper limb) | 0
    Brunnstrom stage IV (lower limb) | 0
    self-feeding | 0
    dizziness | 24
    vomiting | 24
    Kussmaul breathing | 24
    lowered response to verbal commands | 24
    hyperglycemia (344 mg/dL) | 24
    arterial blood gas metabolic acidosis (pH 7.255) | 24
    ketone 3+ | 24
    DKA (Diabetic Ketoacidosis) | 24
    transferred to ICU | 24
    aggressive hydration | 24
    insulin pump | 24
    bicarbonate infusion | 24
    electrolyte correction | 24
    serum ketone body 5.5 mmol/L | 72
    consciousness alert (post DKA) | 72
    metabolic acidosis with respiratory compensation | 24 to 120
    comatose | 144
    hemodynamic instability | 144
    acute infarction over bilateral MCA and ACA territories | 144
    brain swelling | 144
    midline shift | 144
    occlusion of bilateral ICA | 144
    glycerol administration | 144
    endotracheal intubation | 144
    normal left ventricle contractility | 144
    no thrombus or vegetation | 144
    respiratory failure | 144
    severe hyperglycemia | 144
    coma (day 6 to 29) | 144 to 696
    mechanical ventilation | 144
    compassionate extubation | 696
    expired | 696
    WBC 8600/μL | 24
    neutrophil 61.2% | 24
    hemoglobin 14.3 g/dL | 24
    platelet 250000/μL | 24
    sodium 134 mmol/L | 24
    potassium 4.3 mmol/L | 24
    creatinine 0.75 mg/dL | 24
    CRP 1.345 mg/dL | 24
    WBC 16600/μL | 96
    neutrophil 89% | 96
    hemoglobin 13.5 g/dL | 96
    platelet 356000/μL | 96
    sodium 148 mmol/L | 96
    potassium 3.1 mmol/L | 96
    creatinine 0.74 mg/dL | 96
    WBC 32510/μL | 144
    neutrophil 87% | 144
    sodium 146 mmol/L | 144
    potassium 3.4 mmol/L | 144
    WBC 19890/μL | 192
    neutrophil 70.8% | 192
    hemoglobin 13.8 g/dL | 192
    platelet 181000/μL | 192
    sodium 166 mmol/L | 192
    potassium 3.8 mmol/L | 192
    creatinine 1.59 mg/dL | 192
    WBC 18930/μL | 336
    neutrophil 75% | 336
    hemoglobin 11.7 g/dL | 336
    sodium 152 mmol/L | 336
    potassium 4.3 mmol/L | 336
    creatinine 2.94 mg/dL | 336
    WBC 13520/μL | 408
    neutrophil 81.3% | 408
    hemoglobin 10.3 g/dL | 408
    platelet 472000/μL | 408
    sodium 154 mmol/L | 408
    potassium 3.6 mmol/L | 408
    creatinine 2.49 mg/dL | 408
    WBC 13870/μL | 528
    neutrophil 59.2% | 528
    hemoglobin | 528
    sodium | 528
    potassium | 528
    creatinine 1.55 mg/dL | 528
    Free T4 1.04 ng/dL | 24
    TSH 2.58 μIU/mL | 24
    T3 53.5 ng/dL | 24
    Complement C3 70.9 mg/dL | 168
    Complement C4 21 mg/dL | 168
    ANA 1:80X | 168
    Anti-dsDNA 62.33 IU/mL | 168
    ANCA negative | 168
    no recurrent stroke | -2160 to 0
    no urinary tract infection | -2160 to 0
    no pneumonia | -2160 to 0
    no new limb weakness | 24
    no pyuria | 0
    normal thyroid function | 24
    no bacteremia | 24 to 144
    no urinary tract infection | 24 to 144
    no gastroenteritis | 24 to 144
    no pneumonia | 24 to 144
    no drop in blood pressure | 144
    no moyamoya disease | 144
    no sinus rhythm (ECG) | 144
    no vegetations (echocardiogram) | 144
    no autoimmune-related stroke | 168
    no diet control issues | -26208 to 0
    no glycemic control issues | -26208 to"