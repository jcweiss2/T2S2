abdominal pain | -120
abdominal distension | -120
constipation | -120
admitted to hospital | -120
managed conservatively | -120
evaluated by surgical team | 0
evaluated by obstetric team | 0
dehydrated | 0
hypotension | 0
tachycardia | 0
tachypnea | 0
abdomen asymmetrically distended | 0
tenderness all over abdomen | 0
rectum empty on digital examination | 0
foetal viability assessed | 0
vaginal examination not suggestive of threatened preterm labour | 0
laboratory investigations within normal ranges | 0
elevated white cell count | 0
urine analysis clear | 0
ultrasound scan of abdomen and pelvis | 0
distended bowel loop | 0
moderate amount of free fluid in peritoneal cavity | 0
single viable foetus | 0
clinical diagnosis of IO proposed | 0
abdominal X-ray | 2
dilated large bowel | 2
abnormal gas pattern | 2
coffee bean appearance | 2
sigmoid volvulus suspected | 2
gastroenterology team consulted | 4
emergency sigmoidoscopy | 4
twisted sigmoid colon confirmed | 4
obstruction not negotiated | 4
foetal distress | 6
deceleration in heart rate | 6
concomitant caesarean section decided | 6
patient taken to emergency theatre | 8
laparotomy | 8
enormously distended sigmoid loop found | 8
ischemic and gangrenous changes | 8
no signs of perforation | 8
necrotic colon posteriorly displaced by pregnant uterus | 8
lower segment caesarean section | 10
preterm infant delivered | 10
male preterm infant | 10
infant weighed 750g | 10
infant admitted to neonatal ICU | 10
infant on mechanical ventilation | 10
gangrenous sigmoid colon resected | 12
Hartmann’s procedure | 12
end colostomy fashioned | 12
rectal stump closed | 12
patient discharged home | 216
child discharged home | 720
reversal of Hartmann’s | 1296
bowel continuity restored | 1296
colo-rectal anastomosis | 1296