81 years old | 0
female | 0
multiple myeloma | -6720
dexamethasone | -6720
zoledronic acid | -6720
breast cancer | -18240
lumpectomy | -18240
radiation therapy | -18240
hypertension | 0
hypothyroidism | 0
admitted to the hospital | 0
7-day history of cough | -168
cough | -168
runny nose | -168
sore throat | -168
denied fever | -168
denied shortness of breath | -168
denied chest pain | -168
denied skin rashes | -168
denied abdominal pain | -168
denied diarrhea | -168
tachypneic | 0
no pharyngeal erythema | 0
no tonsil exudates | 0
no respiratory accessory muscle use | 0
lungs clear to auscultation | 0
no skin rashes | 0
white blood cell count of 15.1 × 10^9/L | 0
95% segmented neutrophils | 0
bicarbonate of 17 mmol/L | 0
lactate of 1.5 mmol/L | 0
procalcitonin of 0.28 ng/mL | 0
chest radiograph showed no consolidations | 0
computed tomography chest showed small airway disease | 0
RSV polymerase chain reaction from a nasopharyngeal swab was positive | 0
required 2 L of oxygen by nasal cannula | 0
ribavirin | 24
oxygen requirements increased | 24
required high-flow oxygen | 24
transferred to the Intensive Care Unit | 120
intubated | 120
extubated | 192
bilateral lower extremity weakness | 192
absent lower extremity deep tendon reflexes | 192
paresthesias of her feet | 192
upper extremities were involved | 216
normal electrolytes | 216
normal complete blood count with differential | 216
normal procalcitonin | 216
alkaline phosphatase was 62 U/L | 216
alanine aminotransferase 22 U/L | 216
aspartate aminotransferase 57 U/L | 216
creatine kinase 198 U/L | 216
bedside lumbar puncture was attempted | 216
plasmapheresis | 216
received five total of treatment | 240
minimal improvement in quadriparesis and sensory nerve deficit | 240
electromyography showed low amplitude motor responses | 240
axonal sensorimotor peripheral neuropathy | 240
extraocular movements diminished | 264
gag reflex became absent | 264
pupil asymmetry appeared | 264
intubated again | 264
care was withdrawn | 264