56 years old | 0
male | 0
breathlessness on exertion | -8760
breathlessness at rest | -8760
prolonged cough | -8760
bloody sputum production | -8760
hoarseness | -8760
decline in performance impact | -8760
reduced tolerance to physical activity | -8760
admitted to the hospital | 0
significant decrease of blood oxygenation | 0
NYHA III-IV condition | 0
stridor | 0
respiratory distress | 0
giant ascending aorta | 0
aortic arch aneurysm | 0
partial-thrombosed ampullary false aneurysm | 0
left main bronchus compression | 0
left pulmonary artery compression | 0
trachea compression | 0
recurrent pneumonia | 0
multivessel coronary artery disease | 0
surgery | 0
cardiopulmonary bypass | 0
tracheal intubation | 0
bronchoscopy | 0
distal anastomoses of the coronary artery bypass grafting | 0
aneurysmal sac separation | 0
ascending aorta transection | 0
blood antegrade cardioplegia | 0
brachiocephalic trunk clamping | 0
visceral arrest | 0
monohemispheral perfusion of the brain | 0
aneurysmal sac opening | 0
intimal rupture | 0
thrombotic masses | 0
aorta-tracheal fistula | 0
aortic arch replacement | 0
supracoronary replacement of ascending aorta | 0
coronary arteries bypass grafts | 0
trachea repair | 0
extubation | 48
discharged | 336
satisfactory echocardiography | 336
no respiratory failure | 336
no heart failure | 336
no coronary failure | 336
follow-up | 8760
NYHA I | 8760
CT scan | 2160
patency of the trachea and main bronchus restored | 2160
histological examination | 0
atherosclerosis | 0
thinning and inflammation of the aortic wall tissue | 0