41 years old | 0
female | 0
smoker | 0
15 pack-year history | 0
admitted for endoscopic resection of submucous uterine myoma | 0
second surgery for same myoma | 0
preoperative examination normal | 0
laboratory test results normal | 0
baseline blood pressure 120/70 mmHg | 0
baseline heart rate 80 beats per minute | 0
intravenous catheter placed | 0
normal saline administered | 0
general anesthesia induced with fentanyl | 0
general anesthesia induced with propofol | 0
I-gel laryngeal mask No. 4 inserted | 0
anesthesia maintained with desflurane in 40% oxygen | 0
lithotomy position | 0
hysteroscopy with bipolar 9-mm resectoscope | 0
0.9% saline as distention/irrigation medium | 0
end-tidal CO2 drop from 35 to 25 mmHg | 50
pulse oximetry (SpO2) drop from 100% to 90% | 50
blood pressure stable | 50
heart rate stable | 50
crackling sounds from base of lungs | 50
pulmonary edema suspected | 50
irrigated saline volume checked | 50
9000 mL saline used | 50
4000 mL saline collected | 50
surgery stopped | 50
generalized edema noticed | 50
marked distended abdomen | 50
cervical edema with tissue tension | 50
inspired fraction of oxygen increased to 100% | 50
arterial blood analysis performed | 50
pH 7.09 | 50
PaCO2 41 mmHg | 50
PO2 70 mmHg | 50
HCO3+ 12.4 mEq/L | 50
Na+ 145 mEq/L | 50
K+ 2.3 mEq/L | 50
Ca2+ 0.76 mEq/L | 50
hemoglobin 5.9 g/dL | 50
O2 sat 89% | 50
blood glucose level 50 mg/dL | 50
100 mL sodium bicarbonate 8.4% administered | 50
20 mg furosemide administered | 50
laryngeal mask replaced by tracheal tube | 50
airway edema observed in arytenoid region | 50
intubation of 6.5-mm tracheal tube | 50
arterial line put | 50
central line put | 50
10 mEq potassium chloride administered | 50
2 g calcium chloride administered | 50
2 g magnesium sulfate administered | 50
20 mL dextrose 30% administered | 50
supine position | 50
laparoscopy performed to exclude uterus perforation | 50
no uterine rupture | 50
prominent edema of intestinal loops | 50
small amount of peritoneal free fluid observed | 50
bladder catheter inserted | 50
auricular temperature 33°C | 50
admitted to ICU | 50
postoperative chest X-ray showing bilateral pulmonary edema | 50
serious electrolyte disturbances corrected | 50
acidosis corrected | 50
hemoglobin increased to 9.3 g/dL | 50
pre-procedure hemoglobin level 11.9 g/dL | -50
no coagulation abnormalities | 50
temperature returned to normal | 50
generalized edema resolved | 50
urine output 3000 mL | 50
extubation possible six hours after ICU admission | 56
oxygen supplementation for 12 hours with nasal cannula | 60
transferred to general ward approximately 24 hours after ICU admission | 74
stayed in general ward another day | 98
discharged | 120
