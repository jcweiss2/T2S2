61 years old | 0
    male | 0
    type II diabetes mellitus | -4320
    hypothyroidism | -4320
    respiratory failure | -4320
    perforated duodenal ulcer | -4320
    septic shock | -4320
    ventilator | -4320
    antibiotics | -4320
    PEG placement | -4320
    discharged to nursing home | -4320
    levothyroxine | -4320
    insulin | -4320
    ipratropium-albuterol nebulizer | -4320
    morphine | -4320
    intralipid | -4320
    clinimix/dextrose amino acid infusion | -4320
    scopolamine patch | -4320
    pulse oximetry 86% | -6
    high fraction supplemental oxygen | -6
    saturation 94% | -6
    three episodes coffee-ground emesis | -6
    denied NSAID use | -6
    denied cough | -6
    denied fever | -6
    denied hemoptysis | -6
    denied hematemesis | -6
    supplemental oxygen | 0
    saturation 96-100% | 0
    frail | 0
    communicating in complete sentences | 0
    blood pressure 113/63 mm Hg | 0
    temperature 97.9 F | 0
    pulse 110 beats/min | 0
    respiratory rate 22 breaths/min | 0
    diminished breath sounds | 0
    inspiratory wheezing | 0
    non-distended abdomen | 0
    normal bowel sounds | 0
    no stigmata of blood | 0
    no secretions from PEG tube | 0
    elevated blood urea nitrogen 54 mg/dl | 0
    creatinine 0.9 mg/dl | 0
    hemoglobin 10.9 g/dl | 0
    leukocytosis 29.4 × 103/mm3 | 0
    bandemia 11% | 0
    hypoalbuminemia 2.4 g/dl | 0
    elevated alanine aspartate 61 u/L | 0
    INR 1.1 | 0
    X-ray air-bronchogram right lower lobe | 0
    possible pneumonia | 0
    intravenous hydration | 0
    broad-spectrum antibiotics | 0
    intravenous pantoprazole | 0
    EGD severe esophagitis | 0
    diffuse dark mucosal discoloration | 0
    erosion | 0
    profound ulceration entire esophagus | 0
    ischemic necrosis | 0
    resolution GI bleeding | 0
    hypoxia episode | 24
    intensive care monitoring | 24
    cardiac arrest | 72
    death | 72
    