55 years old | 0 | 0 
male | 0 | 0 
morbidly obese | 0 | 0 
diabetes mellitus | 0 | 0 
end-stage renal disease | 0 | 0 
hemodialysis | 0 | 0 
peripheral vascular disease | 0 | 0 
left below knee amputation | 0 | 0 
right above knee amputation | 0 | 0 
right extra anatomical axillobifemoral bypass graft | 0 | 0 
admitted to the hospital | 0 | 0 
right-sided abdominal pain | -48 | 0 
vomiting | -48 | 0 
fever | -48 | 0 
conscious | 0 | 0 
alert | 0 | 0 
oriented | 0 | 0 
pale | 0 | 0 
sick | 0 | 0 
temperature 37.8°C | 0 | 0 
blood pressure 150/90 mmHg | 0 | 0 
oxygen saturation 95% | 0 | 0 
abdomen distended | 0 | 0 
tympanic | 0 | 0 
right upper quadrant tenderness | 0 | 0 
right flank tenderness | 0 | 0 
total leukocyte count 20 × 10^3 | 0 | 0 
hemoglobin 10.7 gm% | 0 | 0 
acidotic pH 7.33 | 0 | 0 
end-stage renal disease | 0 | 0 
chest X-ray | 0 | 0 
air under the right hemi-diaphragm | 0 | 0 
evaluated by general surgeon | 0 | 0 
impression of perforated viscous | 0 | 0 
CT scan with contrast | 0 | 0 
right perinephric collection | 0 | 0 
extension into the right sub-phrenic region | 0 | 0 
gas in the right collecting system | 0 | 0 
gas in the urinary bladder | 0 | 0 
no gas in the renal parenchyma | 0 | 0 
right atrial thrombus | 0 | 0 
started on parenteral antibiotics | 0 | 0 
admitted to intensive care unit | 0 | 0 
percutaneous drainage | 0 | 12 
failed percutaneous drainage | 12 | 12 
evaluated by anesthetist | 12 | 12 
not fit for general anesthesia | 12 | 12 
open drainage | 12 | 24 
epidural anesthesia | 12 | 24 
sedation | 12 | 24 
loculated perinephric and sub-phrenic collection | 12 | 24 
cystoscopy | 24 | 24 
abnormal bladder mucosa | 24 | 24 
multiple cystic lesions | 24 | 24 
air “bubbles” all over the bladder | 24 | 24 
ureteric Double J stent | 24 | 24 
urethral catheter | 24 | 24 
reasonably well during the procedure | 24 | 24 
condition started to deteriorate | 24 | 48 
culture of the collection | 24 | 48 
Klebsiella pneumonia extended-spectrum β-lactamase | 24 | 48 
condition continued to deteriorate | 48 | 72 
severe sepsis | 48 | 72 
multiple organ failure | 48 | 72 
died | 72 | 72