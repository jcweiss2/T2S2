42 years old | 0
male | 0
admitted to the hospital | 0
testicular pain | -192
fever | -48
abdominal tenderness | 0
pulmonary ground-glass opacification | 0
pneumonia | 0
colitis | 0
COVID-19-positive status | 48
attended a biotechnology conference | -336
accidental exposure to SARS-CoV-2 | -336
asymptomatic | -672
respiratory symptoms | -672
cardiac manifestations | 0
acute cardiac injury | 0
myocardial infarction | 0
myocarditis | 0
arrhythmia | 0
cardiogenic shock | 0
heart failure | 0
cardiac tamponade | 0
myopericarditis | 0
neuromuscular manifestations | 0
dizziness | 0
headache | 0
impaired consciousness | 0
acute cerebrovascular disease | 0
ataxia | 0
seizure | 0
taste impairment | 0
smell impairment | 0
vision impairment | 0
nerve pain | 0
myalgia | 0
elevated creatine kinase level | 0
absence of dyspnea | 0
viral encephalitis | 0
acute hemorrhagic necrotizing encephalopathy | 0
Guillain-Barre syndrome | 0
gastrointestinal symptoms | 0
anorexia | 0
diarrhea | 0
nausea/vomiting | 0
abdominal pain | 0
digestive symptoms only | 0
abnormal liver tests | 0
virus detected in stool | 0
gastrointestinal bleeding | 0
renal manifestations | 0
AKI | 0
massive albuminuria | 0
proteinuria | 0
hematuria | 0
elevated blood urea nitrogen | 0
kidney inflammation | 0
edema | 0
ocular manifestations | 0
watery eyes | 0
increased secretions | 0
chemosis | 0
ocular irritation | 0
foreign body sensation | 0
follicular conjunctivitis | 0
conjunctivitis | 0
keratoconjunctivitis | 0
hematological abnormalities | 0
hypercoagulable state | 0
venous thromboembolism | 0
pulmonary embolism | 0
deep vein thrombosis | 0
catheter-associated thrombosis | 0
thrombocytopenia | 0
antiphospholipid antibodies | 0
psychiatric manifestations | 0
anxiety | 0
depression | 0
panic attacks | 0
somatic symptoms | 0
posttraumatic stress disorder | 0
delirium | 0
psychosis | 0
suicidality | 0
dermatological manifestations | 0
maculopapular exanthem | 0
papulovesicular rash | 0
urticaria | 0
painful acral red-purple papules | 0
livedo reticularis lesions | 0
petechiae | 0
discharged | 24