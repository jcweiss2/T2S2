44 years old | 0
male | 0
American Caucasian | 0
hypothyroidism | -672
bronchial asthma | -672
low mood | -216
anxiety | -216
social withdrawal | -216
difficulty sleeping | -216
change in employment status | -216
sought medical advice | -216
brain biopsy | -672
craniotomy | -672
dexamethasone | -672
discharged home | -672
weaker on the right side | -96
worse in the leg | -96
readmitted | -72
denied fever | -72
denied weight loss | -72
denied night sweats | -72
denied nausea | -72
denied vomiting | -72
denied raw milk ingestion | -72
denied smoking | -72
denied drug and alcohol use | -72
history of contact with sick cats | -72
normal higher mental functions | -72
normal language | -72
normal speech | -72
normal cranial nerve function | -72
minimally spastic muscle tone | -72
weak elbow and wrist flexion | -72
weak right lower limb | -72
normal power on the left | -72
normal reflexes | -72
could stand and sit with support | -72
brain MRIs | -72
multiple intracranial focal mass lesions | -72
rim enhancement | -72
restricted diffusion | -72
perilesional vasogenic edema | -72
dexamethasone | -72
levetiracetam | -72
escitalopram | -72
quetiapine | -72
infectious diseases team consulted | -72
laboratory investigations | -72
autoimmune and paraneoplastic auto-antibodies | -72
lymphoma | -72
zoonoses | -72
Brucella | -72
Bartonella | -72
Q-fever | -72
Treponema | -72
Histoplasma | -72
HIV | -72
no systemic malignancy | -72
lumbar puncture | -72
normal opening pressure | -72
normal cytology | -72
normal flow cytometry | -72
first brain biopsy | -72
necroinflammatory process | -72
no acid-fast bacilli | -72
no fungi | -72
no toxoplasma | -72
lymphocytic infiltrate | -72
CD3-positive T-lymphocytes | -72
second brain biopsy | -24
external consultation | -24
workup for occult malignancy | -24
tumor markers | -24
CT of the chest | -24
CT of the abdomen | -24
CT of the pelvis | -24
enlarged mesenteric lymph nodes | -24
thyroid ultrasound | -24
scrotum ultrasound | -24
whole-body FDG-PET scan | -24
postoperative changes | -24
right frontal hypometabolic lesion | -24
pulse steroids | 0
intravenous methylprednisolone | 0
improvement in mood | 24
improvement in power on the right side | 24
walking with a cane | 24
foot orthosis | 24
anxiety | 24
hyper-alertness | 24
low mood | 24
right distal leg weakness | 24
foot drop | 24
polyuria | 24
rituximab infusion | 24
chest infection | 48
focal seizures | 48
encephalopathic | 48
follow-up brain MRI | 48
increasing vasogenic edema | 48
histopathology findings | 48
necrotic brain tissue | 48
atypical lymphoproliferative process | 48
small to medium-sized lymphocytes | 48
pleomorphic nuclei | 48
clumped chromatin | 48
CD2 | 48
CD3 | 48
CD7 | 48
granzyme B | 48
TIA 1 | 48
negative for CD4 | 48
negative for CD5 | 48
negative for CD8 | 48
negative for CD56 | 48
negative for TCR beta F1 | 48
negative for TCR delta | 48
EBV-encoded RNA | 48
pulmonary embolism | 144
sepsis | 144
disseminated intravascular coagulation | 144
multiorgan failure | 144
large left frontoparietal intraparenchymal hematoma | 144
vasogenic edema | 144
midline shift | 144
diffuse loss of gray-white differentiation | 144
effacement of sulci | 144
cardiopulmonary arrest | 216
death | 216