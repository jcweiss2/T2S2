48 years old | 0
    male | 0
    seizure disorder | -131400
    antiepileptics | -131400
    valproic acid | 0
    carbamazepine | 0
    clobazam | 0
    type-2 diabetes mellitus | -87600
    oral hypoglycemic agents | -87600
    hypertension | -52560
    impaired level of consciousness | -24
    admitted to critical care unit | 0
    blood pressure 160/100 mmHg | 0
    heart rate 96/min | 0
    respiratory rate 22/min | 0
    Glasgow coma score 11 | 0
    poor coughing | 0
    coarse crepts on right base | 0
    worsening of sensorium | 0
    inability to protect airway | 0
    intubated | 0
    mechanical ventilation | 0
    suspicion of antiepileptic overdose | 0
    antiepileptics stopped | 0
    intravenous infusion of propofol | 0
    elevated creatinine 4.5 mg/dl | 0
    BUN 40 mg/dl | 0
    blood sugar 176 mg/dl |*0
    total leukocyte count 11,400 | 0
    82% polymorphs | 0
    total protein 5 g/dl | 0
    albumin 2.3 g/dl | 0
    total bilirubin 0.25 mg/dl | 0
    AST 27 U/L | 0
    ALT 16 U/L | 0
    Alk. Phosphatase 125 | 0
    increased cortical echotexture | 0
    poorly maintained corticomedullary differentiation | 0
    medical renal disease | 0
    serum creatinine 2.1 mg/dl | -3600
    septic ruled out | 0
    dyselectrolytemias ruled out | 0
    MRI head no abnormality | 0
    cerebrospinal fluid analysis no abnormality | 0
    electroencephalogram continuous generalized slowing | 0
    BUN level 68 mg/dl | 0
    hemodialysis | 0
    no improvement in sensorium | 0
    BUN 21 mg/dl | 0
    serum antiepileptic drugs within therapeutic ranges | 0
    ammonia level 274 μmol/L | 0
    valproate-induced hyperammonemic encephalopathy | 0
    L-carnitine started | 0
    urea cycle enzyme abnormality not evaluated | 0
    no history of drugs leading to hyperammonia | 0
    no hematological disease | 0
    sensorium improved | 168
    weaning trial planned | 168
    refractory septic shock | 168
    ICU-acquired multidrug resistant infection | 168
    succumbed to death | 168
    <|eot_id|>
    