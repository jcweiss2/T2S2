40 years old | 0
male | 0
poorly controlled diabetes mellitus | 0
admitted to ICU | 0
right thigh cellulitis | 0
diabetic ketoacidosis | 0
inferior wall myocardial infarction | 0
right ventricular dysfunction | 0
altered sensorium | 0
hemodynamically unstable | 0
respiratory distress | 0
management of DKA | 0
management of acute coronary syndrome | 0
invasive mechanical ventilation | 0
central line placement | 0
IV fluid resuscitation | 0
vasoactive drugs | 0
anti-platelets | 0
therapeutic heparinization | 0
IV insulin infusion | 0
glycemic control | 0
electrolytes management | 0
neuromuscular weakness | 1008
nosocomial infections | 1008
ischemic cardiomyopathy | 1008
grade III sacral bedsore | 1008
high-grade fever | 1008
S. multivorum cultured from peripheral blood | 1008
bacteremia | 1008
piperacillin/tazobactam sensitive | 1008
levofloxacin sensitive | 1008
ceftazidime resistant | 1008
amikacin resistant | 1008
imipenem resistant | 1008
carbapenem resistant | 1008
aztreonam resistant | 1008
trimethoprim/sulfamethoxazole sensitive | 1008
treated with trimethoprim/sulfamethoxazole | 1008
discharged | unknown