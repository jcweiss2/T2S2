61 years old | 0
male | 0
Indigenous | 0
admitted to the hospital | 0
fever | -96
malaise | -96
cough | -96
breathlessness | -96
seropositive rheumatoid arthritis | -0
cutaneous lupus erythematosus | -0
emphysema | -0
ischaemic heart disease | -0
functional hyposplenism | -0
etanercept | -1296
methotrexate | -0
hydroxychloroquine | -0
allergy to sulfanilamide | -8760
cigarette smoker | -0
no alcohol consumption | -0
no intravenous drugs | -0
no recent gardening | -0
no soil exposure | -0
heart rate 104 beats per minute | 0
respiratory rate 24 breaths per minute | 0
blood pressure 101/56 mmHg | 0
oxygen saturation 97% | 0
temperature 39.7 °C | 0
hypopigmented rash | 0
bronchial breath sounds | 0
crepitations | 0
mild left flank tenderness | 0
normocytic anemia | 0
leucocytosis | 0
neutrophilia | 0
acute kidney injury | 0
right upper lobe opacification | 0
left heart border opacification | 0
community-acquired pneumonia | 0
intravenous ceftriaxone | 0
intravenous gentamicin | 0
oral doxycycline | 0
deterioration | 12
hypoxia | 12
hypotension | 12
hyperlactatemia | 12
oxygen via high-flow nasal-prongs | 12
intravenous noradrenaline | 12
intravenous meropenem | 12
intravenous vancomycin | 12
oral azithromycin | 12
transfer to ICU | 12
pulmonary infiltrates | 24
Gram-negative bacilli | 48
Acinetobacter baumannii complex | 48
sensitive to meropenem | 48
sensitive to ceftazidime | 48
sensitive to co-trimoxazole | 48
sensitive to gentamicin | 48
Burkholderia pseudomallei | 72
sensitive to meropenem | 72
sensitive to co-trimoxazole | 72
sensitive to doxycycline | 72
improved clinically | 96
discharged from ICU | 96
no ongoing oxygen requirement | 96
subsequent blood cultures showed no growth | 120
intravenous ceftazidime | 168
CT scan of abdomen and pelvis | 168
L3/L4 discitis | 168
vertebral osteomyelitis | 168
peripherally inserted central catheter | 168
etanercept withheld | 168
inflammatory arthritis managed | 168
oral trimethoprim/sulfamethoxazole | 168
fixed drug eruption | 240
cessation of TMP/SMX | 240
doxycycline | 240
oral TMP/SMX for six months | 336 
discharged | 720