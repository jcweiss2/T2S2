24 weeks + 3 days | -672
female | -672
breech presentation | -672
cord prolapse | -672
birth weight 645 g | -672
HIV negative | -672
Apgar score 4 | -672
Apgar score 8 | -672
mechanical ventilation | 0
central umbilical catheters | 0
total parenteral nutrition | 0
empiric antibiotics | 0
skin sensors | 0
late-onset sepsis | 216
Escherichia coli bacteremia | 216
cefepime | 216
adhesive patch | 432
skin abrasion | 432
erythema | 432
induration | 432
plaque | 432
necrotic center | 432
ulcer | 480
subcutaneous cell tissue | 480
necrotic area | 480
thermic instability | 480
metabolic acidosis | 480
hyperglycemia | 480
hypotension | 480
cutaneous mucormicosis | 480
skin biopsy | 480
liposomal amphotericin B | 480
refractory shock | 528
renal failure | 528
death | 528
Rhizopus spp. | 528
broad aseptate hyphae | 528
right angle branching | 528
Rhizopus arrhizus | 528