36 years old | 0
    male | 0
    severe lower abdominal pain | -4
    discomfort | -4
    fever | -4
    admitted to the emergency room | 0
    ulcerative colitis | -35040
    mesalazine | -35040
    hepatic dullness upward shift | 0
    abdominal tenderness | 0
    left lower abdominal tenderness | 0
    mild abdominal muscle tension | 0
    no hepatic percussion pain | 0
    no renal percussion pain | 0
    leukocytosis (13.62×10^9/L) | 0
    neutrophils 90.10% | 0
    c-reactive protein 176.50 mg/L | 0
    glucose 10.6 mmol/L | 0
    lactate 3.0 mmol/L |# Import Error: No module named '0'
    coagulation routine: prothrombin time 16.1S | 0
    international normalized ratio 1.43 | 0
    activated partial thromboplastin time 32.0S | 0
    plasma fibrinogen 2.5 g/L | 0
    calcitoninogen 8.967 ng/mL | 0
    abdominal CT: enlarged spleen | 0
    abdominal CT: abnormally thick spleen | 0
    gastrointestinal perforation | 0
    rehydration | 0
    imipenem cilastatin (1.0 g q8h) | 0
    emergency surgery | 0
    pelvic abscess cavity | 0
    dense adhesions (lower abdomen, pelvic ileum, sigmoid colon, peritoneum) | 0
    omental necrosis | 0
    adhesions (ileum, sigmoid colon) | 0
    pelvic abscess | 0
    intestinal wall edema | 0
    thickened intestinal wall | 0
    gray-white attachments (intestinal wall) | 0
    appendix occlusion | 0
    appendix swelling | 0
    pus moss (appendix) | 0
    partial sigmoid resection | 0
    pelvic-abdominal adhesion release | 0
    incidental appendectomy | 0
    pelvic abscess incision | 0
    pelvic abscess drainage | 0
    partial omentum resection | 0
    temporary colostomy | 0
    perforation repair | 0
    postoperative pathology: sigmoid colon rupture | 0
    postoperative pathology: hemorrhage | 0
    postoperative pathology: necrosis | 0
    postoperative pathology: acute and chronic inflammation | 0
    postoperative pathology: inflammatory exudate | 0
    postoperative pathology: granulation tissue | 0
    postoperative pathology: glandular hyperplasia | 0
    postoperative pathology: thrombosis | 0
    postoperative pathology: negative margins | 0
    postoperative CT: enlarged spleen (8 rib units) | 24
    postoperative CT: heterogeneous density | 24
    postoperative CT: large air shadow | 24
    splenic abscess (diagnosis) | 24
    blood culture (negative) | 24
    imipenem cilastatin (1.0 g q8h) continuation | 24
    ultrasound-guided splenic abscess drainage | 24
    infection index not decreased | 24
    platelet count decreased | 24
    prothrombin time decreased | 24
    coagulation routine: prothrombin time 15.4S | 24
    international normalized ratio 1.36 | 24
    activated partial thromboplastin time 48.9S | 24
    prothrombin time 21.6S | 24
    intermittent fever | 24
    abdominal pain | 24
    hypoproteinemia | 48
    coagulopathy | 48
    splenectomy | 48
    abdominal drainage | 48
    splenic gangrene | 48
    red-brown purulent effusion | 48
    peripheral yellow-brown effusion | 48
    yellow-brown pelvic effusion | 48
    postoperative pathology: splenic necrosis | 48
    postoperative pathology: splenic hemorrhage | 48
    symptomatic treatment continuation | 48
    fever improvement | 72
    abdominal discomfort improvement | 72
    imaging normalization | 168
    test indexes normalization | 168
    discharged | 168
    