70 years old | 0
male | 0
admitted to the hospital | 0
hypertension | 0
insulin-dependent diabetes mellitus | 0
hyperlipidemia | 0
statin therapy | 0
sickle cell trait | 0
bilateral upper- and lower-extremity weakness | -2160
difficulty rising from a sitting position | -2160
fatigue | -2160
subjective weight loss | -2160
decreased appetite | -2160
no skin changes | -2160
no previous trauma | -2160
no sick contacts | -2160
no recent immobilization/hospitalization | -2160
no dysphagia | -2160
no discoloration of urine | -2160
3/5 strength in all 4 extremities | 0
no fever | 0
no rash | 0
no tenderness | 0
no swelling | 0
elevated AST | 0
elevated ALT | 0
elevated CPK | 0
Hgb 10 g/dl | 0
MCV of 95 fl | 0
eosinophilia 10% | 0
statin therapy discontinued | -2880
severe myalgia | -2880
right quadriceps muscle biopsy | -2880
elevated HMGCR levels | -2880
autoimmune necrotizing myopathy | -2880
long-standing inflammatory myopathy | -2880
weekly methotrexate | -2880
prednisone twice daily | -2880
intravenous immunoglobulin | -2880
discharged | -2880
prednisone 20 mg twice daily | -2880
oral methotrexate 7.5 mg weekly | -2880
readmitted | 0
lethargy | 0
inability to speak | 0
inability to follow commands | 0
dry cough | -2160
occasional fever | -2160
occasional diarrhea | -2160
deterioration in overall condition | 0
febrile | 0
temperature 39.3°C | 0
tachypnea | 0
tachycardia | 0
blood pressure 109/56 mmHg | 0
crackles | 0
reduced breath sounds | 0
oral thrush | 0
Na+ 122 mmol/l | 0
hemoglobin 8 g/dl | 0
leukopenia | 0
eosinophilia | 0
CPK 163U/L | 0
ABG pH 7.57 | 0
ABG pCO2 27 | 0
ABG pO2 89 | 0
lactic acid 4.5 mmol/L | 0
CT head normal | 0
cerebro-spinal fluid normal | 0
chest X-ray bilateral infiltrates | 0
blood cultures obtained | 0
broad-spectrum antibiotics | 0
hypoxic | 24
cardiopulmonary arrest | 24
intubated | 24
hypoxic respiratory failure | 24
ABG pH 7.18 | 24
ABG PCO2 43 | 24
ABG PO2 67 | 24
ABG HCO3 15 | 24
return of spontaneous circulation | 24
chest X-ray worsening bilateral lower lobe infiltrates | 24
CT chest bilateral consolidation | 24
acute respiratory distress syndrome | 24
PaO2/FiO2 96 | 24
CT negative for pulmonary embolism | 24
bronchoscopy | 24
bronchoalveolar lavage | 24
BAL positive for Strongyloides stercoralis larvae | 24
serology Strongyloides negative | 24
HIV negative | 24
initial stool sample negative | 24
second stool sample positive for rhabditiform larvae | 48
steroids suspended | 24
Ivermectin 200 mg/kg | 24
Albendazole 400 mg | 24
blood cultures positive for Klebsiella pneumoniae | 24
antibiotics continued | 24
died | 456
