44 years old | 0
male | 0
hepatitis B | 0
primary hepatocellular carcinoma | 0
chronic viral hepatitis B without cirrhosis | 0
multiphasic contrast-enhanced MRI showed 9.8 cm × 7.9 cm mass in the right hepatic lobe | 0
arterial hypervascularity | 0
AFP greater than 3,630 ng/mL | 0
BCLC stage B | 0
first TACE (May 8, 2018) | 0
fever | 24
maximum temperature 39.3 °C | 24
severe liver damage | 24
WBC 8.5×10^9/L | 24
GRAN 91.4% | 24
ALT 2.6 ULN | 24
AST 7.9 ULN | 24
TBIL 1.9 ULN | 24
liver preservation treatment | 24
one month after first TACE: ALT, AST, TBIL normal | 744
WBC 9.2×10^9/L | 744
GRAN 82.7% | 744
abdominal MRI showed significant necrosis of lesions | 744
AFP dropped to 1,708 ng/mL | 744
repeated fever | 1272
cough | 1272
maximum temperature 39 °C | 1272
chest CT showed pneumonia in right lung | 1272
pneumorachis with iodine oil deposition | 1272
hepatic abscess | 1272
anti-infection treatment (Tazobactam/Piperacillin) | 1272
pigtail catheter drainage | 1272
bacteria culture negative | 1272
July 31, 2018: enhanced MRI showed reduction in original lesion | 2088
new lesions in liver increased | 2088
AFP rose to more than 3,630 ng/mL | 2088
three more TACE (August to November 2018) | 2544, 2880, 3264
fifth TACE (November 30, 2018) | 3264
fever | 3264
maximum temperature 39.6 °C | 3264
WBC 14.1×10^9/L | 3264
GRAN 98.5% | 3264
ALT 163 U/L | 3264
AST 249 U/L | 3264
TBIL 73 µmol/L | 3264
anti-infection treatment | 3264
liver protection treatment | 3264
three days after fifth TACE: fainted | 3336
difficulty breathing | 3336
enhanced CT showed HPVG | 3336
Streptococcus anginosus culture positive | 3336
died two hours after ICU admission | 3352
