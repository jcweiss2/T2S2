54 years old | 0
female | 0
Latin American | 0
type 2 diabetes mellitus | -8760
end-stage renal disease | -8760
history of headache | -240
history of photophobia | -240
history of chronic cough | -240
history of weight loss | -240
history of low-grade fever | -240
close contact with a person with pulmonary tuberculosis | -8760
admitted to the emergency department | 0
febrile | 0
tachycardic | 0
mild impairment of alertness | 0
diffuse crackles mainly of the left lung | 0
WBC 4800 cells/μL | 0
absolute lymphocyte count 816 cells/μL | 0
hemoglobin 10.3 g/dL | 0
blood sugar 111 mg/dL | 0
liver function tests were normal | 0
creatinine 7.2 mg/dL | 0
blood urea nitrogen 59 mg/dL | 0
bilateral interstitial infiltrates | 0
multiple ring-shaped lesions in posterior areas of both hemispheres | 0
acid-fast bacilli sputum culture was positive | 0
Mycobacterium tuberculosis complex (MTB) | 0
no evidence of antibacterial resistance | 0
HIV1/2 and toxoplasma serologies were negative | 0
lumbar puncture | 0
opening pressure was 30 cm H2O | 0
red blood cell count 1000 cells/μL | 0
WBC 114 cells/μL | 0
lymphocytes 92% | 0
glucose 30 mg/dL | 0
proteins 161 mg/dL | 0
CSF neurocysticercosis serology and cryptococcal antigen were negative | 0
CSF Mycobacterium tuberculosis stain and culture were negative | 0
adenosine deaminase were negative | 0
polymerase chain reaction (PCR) was positive for MTB | 0
anti-TB therapy was started | 0
rifampin | 0
isoniazid | 0
pyrazinamide | 0
ethambutol | 0
pyridoxine | 0
dexamethasone | 0
admission to the intensive care unit | 72
initiation of hemodialysis | 72
uremia | 72
clinical improvement | 120
acute abdominal pain | 504
hematemesis | 504
loculated multiseptated gas and fluid collection along the posterior aspect of the gastric fundus | 504
free intra-abdominal air | 504
gastric perforation | 504
exploratory laparotomy | 504
complete stomach necrosis | 504
total gastrectomy | 504
intestinal discontinuity | 504
cervical esophagostomy | 504
jejunostomy tube (J-tube) placement | 504
oral anti-TB therapy was switched to intravenous treatment | 504
amikacin | 504
linezolid | 504
levofloxacin | 504
rifampin | 504
septic shock | 504
intubation | 504
mechanical ventilation | 504
empiric broad-spectrum antibacterial therapy | 504
piperacillin-tazobactam | 504
intra-abdominal infection | 504
vascular thrombosis | 504
broad, irregularly branched, rarely septate hyphae | 504
angio-invasive gastric mucormycosis | 504
liposomal amphotericin B | 504
TB treatment with levofloxacin, rifampin, isoniazid, and linezolid | 504
posaconazole | 1008
clinical stabilization | 1008
improvement | 1008
returned to her country of origin | 1008
finalized treatment | 1008