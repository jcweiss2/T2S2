64 years old | 0
male | 0
hypertension | -672
arthritis | -672
seizure disorder | -672
Parkinson's disease | -672
hiatal hernia | -672
chronic anemia | -672
non-bloody and non-bilious vomiting | -216
decreased oral intake | -216
progressive generalized weakness | -168
new-onset dyspnea | -168
excessive NSAIDs | -168
gastritis | -3024
severe diverticulosis | -3024
tubular adenoma of the splenic flexure | -3024
hemorrhoids | -3024
unstable blood pressure | 0
low blood pressure | 0
tachypneic | 0
labored breathing | 0
decreased breath sounds on the right side | 0
mild elevations in ALT/AST | 0
normal bilirubin levels | 0
right-sided pneumothorax | 0
moderate right-sided pleural effusion | 0
metabolic acidosis | 0
respiratory compensation | 0
high anion gap | 0
elevated white cell count | 0
elevated neutrophils | 0
low RBC | 0
low hemoglobin | 0
low hematocrit | 0
elevated platelets | 0
elevated PT/INR | 0
elevated APTT | 0
elevated lactate | 0
elevated troponin | 0
hypernatremia | 0
hyperkalemia | 0
hypochloremia | 0
low bicarbonate | 0
elevated anion gap | 0
hyperglycemia | 0
hypocalcemia | 0
elevated creatinine | 0
low eGFR | 0
elevated BUN | 0
low protein | 0
low albumin | 0
elevated lactate dehydrogenase | 0
volume resuscitation | 0
packed red blood cells | 0
transfer to intensive care | 0
blood cultures | 0
sputum cultures | 0
urine cultures | 0
cefepime | 0
coverage of pneumonia | 0
parapneumonic effusion | 0
chest tube placement | 0
drainage of air and purulent fluid | 0
respiratory status decline | 0
intubation | 24
Candida Tropicalis | 24
Candida Glabrata | 24
Stenotrophomonas maltophilia | 24
broadened antibiotic coverage | 24
meropenem | 24
caspofungin | 24
polymicrobial flora | 24
elevated amylase | 24
esophageal tear | 24
upper endoscopy | 48
posterior distal esophagus defect | 48
Boerhaave syndrome | 48
gastric ulcers | 48
tissue fibrosis | 48
friability | 48
esophageal stenting | 48
biopsies | 48
acute inflammation | 48
fungal organisms | 48
candida species | 48
echocardiogram | 48
ejection fraction | 48
moderate to severe tricuspid regurgitation | 48
mitral regurgitation | 48
moderate pulmonary hypertension | 48
clinical improvement | 192
extubation | 192
CT-guided catheter placement | 192
pleural cavity drainage | 192
decompensation | 216
Lactobacillus | 216
Staphylococcus lugdunensis | 216
vancomycin | 216
ceftazidime | 216
metronidazole | 216
caspofungin | 216
worsening infiltrates | 216
mediastinitis | 216
acute respiratory distress syndrome | 216
re-intubation declined | 240
death | 240