19 years old | 0
female | 0
admitted to the department of internal medicine | 0
history of pancreatitis | -336
pancreatitis of unclear nature | -336
computed tomography | -336
portal vein thrombosis | -336
tumor mass located at the pancreatic head | -336
suspicious for pancreatic cancer | -336
explorative laparotomy | -336
tumor mass regarded as unresectable | -336
tumor infiltration of the mesenteric root | -336
biopsies of the tumor mass | -336
portal venous stent placed | -336
dismissed with the diagnosis of chronic pancreatitis | -336
abdominal pain | -1560
imaging confirmed the diffuse and large tumor mass | -1560
intra- and extrahepatic cholestasis | -1560
occlusion of the portal vein stent | -1560
portal-systemic collateralization | -1560
varices | -1560
dislocated portal vein stent | -1560
perforation into the stomach | -1560
Carbohydrate-Antigen 19.9 (CA19.9) slightly elevated | -1560
admitted to our surgical clinic | -1560
pancreatic tumor with unsolved dignity | -1560
compression of the duodenum | -1560
cholestasis | -1560
interdisciplinary meeting | -1560
surgical approach decided | -1560
explorative laparotomy | 0
exposed the portal vein and the mesenteric root | 0
transecting all varices | 0
mesenterico-caval shunt | 0
release portal hypertension | 0
alleviate esophageal varices | 0
ensure biliary drainage | 0
gastro-intestinal passage | 0
recovery of the dislocated stent | 0
dissected the hepatoduodenal ligament | 0
identified the portal vein, hepatic artery and central bile duct | 0
removed the dislocated and stomach-penetrating stent | 0
ligated the portal vein | 0
partial duodenopancreatectomy | 0
resection of the distal stomach | 0
hepatico-jejunostomy | 0
gastro-jejunostomy | 0
pancreatic duct could not be identified | 0
pancreatic stump oversewn with non-absorbable sutures | 0
blindly closed by stitches | 0
monitored on intensive care unit | 24
pathological analysis | 24
pancreatitis with acinar atrophy | 24
ductal ecstasy | 24
inflammatory exudate | 24
no evidence for malignancy | 24
granulocytic epithelial lesion (GELs) | 24
type-2 autoimmune pancreatitis (AIP) | 24
steroid treatment initiated | 24
clinical response | 24
decreasing cholestasis | 24
supported the diagnosis of AIP | 24
postoperative follow-up | 168
all symptoms vanished | 168
good quality of life | 168