37 years old|0
    male|0
    transferred to tertiary care ICU|0
    acute on chronic pancreatitis|0
    severe epigastric pain|0
    progressive lower limbs paresis|0
    alcohol-related acute pancreatitis history|-72
    heart rate 70 beats/minute|0
    blood pressure 126/76 mmHg|0
    saturation 99% at FiO2=0.21|0
    body temperature 38°C|0
    Cullen’s sign|0
    tender abdomen|0
    no signs of peritonitis|0
    absent deep tendon reflexes|0
    weakened middle and lower cutaneous reflexes|0
    attenuation of all sensations below umbilicus|0
    complete loss of sensation below knees|0
    increased amylase (234 U/L)|0
    leukocytosis (12×103/uL)|0
    giant pancreatic pseudocyst (20×14×18 cm)|0
    impaired contrast enhancement left kidney|0
    subcapsular ischemic foci kidneys|0
    central hyper-intense signal on T2 MRI|0
    medullary infarction suspected|0
    LMWH prophylaxis|0
    empiric antimicrobial therapy|0
    mild anemia (hemoglobin 11.7 g/dL)|0
    thrombocytopenia (146×103/uL)|0
    general condition deteriorated|24
    acute renal failure|24
    hemodialysis|24
    acute liver failure|24
    paresis transformed to paraplegia|24
    anemia (6.5 g/dL)|24
    thrombocytopenia (61×103/uL)|24
    decreased fibrinogen (135 mg/dL)|24
    increased D-dimers (29.1 ug/mL)|24
    INR 2.1|24
    prolonged aPTT (40.7 seconds)|24
    intracystic bleeding|24
    FFP administered|24
    packed RBC administered|24
    transferred in critical condition|72
    hypotensive|72
    vasopressors use|72
    septic shock|72
    negative cultures|72
    emergency laparotomy|72
    omentectomy|72
    cholecystectomy|72
    external drainage pancreatic cyst|72
    coagulative necrosis gallbladder mucosa|72
    inflammatory infiltrate|72
    fresh thrombosis intramuscular vessel|72
    ischemic foci liver and spleen|168
    necrotic tissue pancreatic head and body|168
    relaparotomy|168
    pancreatic necrosectomy|168
    lesser sac drainage|168
    rectovesical pouch drainage|168
    pancreatobiliary fistula|168
    amylase-rich fluid output|168
    total parenteral nutrition|168
    somatostatin|168
    hemodiafiltration sessions (8)|168
    hemodialysis sessions (4)|168
    RBC transfusion (4 packs)|168
    packed platelets|168
    FFP transfusion|168
    platelets normalized|216
    hemoglobin normalized|288
    transferred to surgical ward|312
    MRI persistent hyperintense T2 signal|504
    patchy contrast enhancement|504
    persistent pancreatic fistula|504
    scheduled ERCP|504
    atrial fibrillation|624
    cardiac arrest|624
    ERCP complication|624
    ERCP stents introduced|960
    discharged|1368
    lower-limb muscle atrophy|8760
    contractures talocrural regions|8760
    no deep tendon reflexes|8760
    no middle and lower cutaneous reflexes|8760
    no sensation below knees|8760
    regained hip flexion/extension|8760
    urinary retention|8760
    erectile dysfunction|8760
    MRI medullary cone atrophy|8760
    central gliosis|8760
