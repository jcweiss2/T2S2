60 years old | 0
    female | 0
    nursing home patient | 0
    bipolar affective disorder | 0
    hypertension | 0
    hypothyroidism | 0
    paraplegia | 0
    increasing confusion | 0
    admitted to senior behavioral facility | 0
    unable to communicate | -168
    tachycardia | -168
    tachypnea | -168
    flushing | -168
    diaphoresis | -168
    fevers greater than 38°C | -168
    transferred to NCCU | -168
    encephalopathic | 0
    tachypneic | 0
    tachycardic | 0
    hypoxemic | 0
    generalized rigidity | 0
    hyperreflexia | 0
    leukocytosis | 0
    acute kidney injury | 0
    elevated serum creatinine phosphokinase | 0
    procalcitonin elevated | 0
    C-reactive protein within normal limits | 0
    episodes of hypotension | 0
    episodes of hypertension | 0
    possible sepsis | 0
    NMS | 0
    serotonin syndrome | 0
    non-convulsive status epilepticus | 0
    CNS pathology | 0
    blood cultures obtained | 0
    urine cultures obtained | 0
    sputum cultures obtained | 0
    lumbar puncture considered | 0
    medical records obtained | 0
    receiving increasing doses of ziprasidone | -168
    haloperidol | -168
    lithium | -168
    duloxetine | -168
    oxybutynin | -168
    baclofen | -168
    treated with IV bromocriptine | 0
    treated with IV dantrolene | 0
    discontinuation of causative agents | 0
    cooling blanket | 0
    antipyretics | 0
    IV fluids | 0
    SS considered | 0
    escalating doses of ziprasidone | 0
    unaltered use of duloxetine | 0
    unaltered use of lithium | 0
    administer bromocriptine | 0
    dantrolene scheduled | 0
    electroencephalography showed generalized slowing | 0
    no seizure activity | 0
    MRI brain no acute finding | 0
    afebrile | 72
    improved leukocytosis | 72
    no antibiotics | 72
    no lumbar puncture | 72
    autonomic dysregulation resolved | 96
    cessation of labile blood pressures | 96
    supplemental oxygen requirements ceased | 96
    more awake | 96
    less rigid in extremities | 96
    unable to participate in meaningful interview | 96
    dantrolene increased to 100 mg TID | 96
    stable | 120
    transferred out of NCCU | 120

    60 years old | 0
    female | 0
    nursing home patient | 0
    bipolar affective disorder | 0
    hypertension | 0
    hypothyroidism | 0
    paraplegia | 0
    increasing confusion | 0
    admitted to senior behavioral facility | 0
    unable to communicate | -168
    tachycardia | -168
    tachypnea | -168
    flushing | -168
    diaphoresis | -168
    fevers greater than 38°C | -168
    transferred to NCCU | -168
    encephalopathic | 0
    tachypneic | 0
    tachycardic | 0
    hypoxemic | 0
    generalized rigidity | 0
    hyperreflexia | 0
    leukocytosis | 0
    acute kidney injury | 0
    elevated serum creatinine phosphokinase | 0
    procalcitonin elevated | 0
    C-reactive protein within normal limits | 0
    episodes of hypotension | 0
    episodes of hypertension | 0
    possible sepsis | 0
    NMS | 0
    serotonin syndrome | 0
    non-convulsive status epilepticus | 0
    CNS pathology | 0
    blood cultures obtained | 0
    urine cultures obtained | 0
    sputum cultures obtained | 0
    lumbar puncture considered | 0
    medical records obtained | 0
    receiving increasing doses of ziprasidone | -168
    haloperidol | -168
    lithium | -168
    duloxetine | -168
    oxybutynin | -168
    baclofen | -168
    treated with IV bromocriptine | 0
    treated with IV dantrolene | 0
    discontinuation of causative agents | 0
    cooling blanket | 0
    antipyretics | 0
    IV fluids | 0
    SS considered | 0
    escalating doses of ziprasidone | 0
    unaltered use of duloxetine |0
    unaltered use of lithium | 0
    administer bromocriptine | 0
    dantrolene scheduled | 0
    electroencephalography showed generalized slowing | 0
    no seizure activity | 0
    MRI brain no acute finding | 0
    afebrile | 72
    improved leukocytosis | 72
    no antibiotics | 72
    no lumbar puncture | 72
    autonomic dysregulation resolved | 96
    cessation of labile blood pressures | 96
    supplemental oxygen requirements ceased | 96
    more awake | 96
    less rigid in extremities | 96
    unable to participate in meaningful interview | 96
    dantrolene increased to 100 mg TID | 96
    stable | 120
    transferred out of NCCU | 120

    60 years old | 0
    female | 0
    nursing home patient | 0
    bipolar affective disorder | 0
    hypertension | 0
    hypothyroidism | 0
    paraplegia | 0
    increasing confusion | 0
    admitted to senior behavioral facility | 0
    unable to communicate | -168
    tachycardia | -168
    tachypnea | -168
    flushing | -168
    diaphoresis | -168
    fevers greater than 38°C | -168
    transferred to NCCU | -168
    encephalopathic | 0
    tachypneic | 0
    tachycardic | 0
    hypoxemic | 0
    generalized rigidity | 0
    hyperreflexia | 0
    leukocytosis | 0
    acute kidney injury | 0
    elevated serum creatinine phosphokinase | 0
    procalcitonin elevated | 0
    C-reactive protein within normal limits | 0
    episodes of hypotension | 0
    episodes of hypertension | 0
    possible sepsis | 0
    NMS | 0
    serotonin syndrome | 0
    non-convulsive status epilepticus | 0
    CNS pathology | 0
    blood cultures obtained | 0
    urine cultures obtained | 0
    sputum cultures obtained | 0
    lumbar puncture considered | 0
    medical records obtained | 0
    receiving increasing doses of ziprasidone | -168
    haloperidol | -168
    lithium | -168
    duloxetine | -168
    oxybutynin | -168
    baclofen | -168
    treated with IV bromocriptine | 0
    treated with IV dantrolene | 0
    discontinuation of causative agents | 0
    cooling blanket | 0
    antipyretics | 0
    IV fluids | 0
    SS considered | 0
    escalating doses of ziprasidone | 0
    unaltered use of duloxetine | 0
    unaltered use of lithium | 0
    administer bromocriptine | 0
    dantrolene scheduled | 0
    electroencephalography showed generalized slowing | 0
    no seizure activity | 0
    MRI brain no acute finding | 0
    afebrile | 72
    improved leukocytosis | 72
    no antibiotics | 72
    no lumbar puncture | 72
    autonomic dysregulation resolved | 96
    cessation of labile blood pressures | 96
    supplemental oxygen requirements ceased | 96
    more awake | 96
    less rigid in extremities | 96
    unable to participate in meaningful interview | 96
    dantrolene increased to 100 mg TID | 96
    stable | 120
    transferred out of NCCU | 120

    60 years old | 0
    female | 0
    nursing home patient | 0
    bipolar affective disorder | 0
    hypertension | 0
    hypothyroidism | 0
    paraplegia | 0
    increasing confusion | 0
    admitted to senior behavioral facility | 0
    unable to communicate | -168
    tachycardia | -168
    tachypnea | -168
    flushing | -168
    diaphoresis | -168
    fevers greater than 38°C | -168
    transferred to NCCU | -168
    encephalopathic | 0
    tachypneic | 0
    tachycardic | 0
    hypoxemic | 0
    generalized rigidity | 0
    hyperreflexia | 0
    leukocytosis | 0
    acute kidney injury | 0
    elevated serum creatinine phosphokinase | 0
    procalcitonin elevated | 0
    C-reactive protein within normal limits | 0
    episodes of hypotension | 0
    episodes of hypertension | 0
    possible sepsis | 0
    NMS | 0
    serotonin syndrome | 0
    non-convulsive status epilepticus | 0
    CNS pathology | 0
    blood cultures obtained | 0
    urine cultures obtained | 0
    sputum cultures obtained | 0
    lumbar puncture considered | 0
    medical records obtained | 0
    receiving increasing doses of ziprasidone | -168
    haloperidol | -168
    lithium | -168
    duloxetine | -168
    oxybutynin | -168
    baclofen | -168
    treated with IV bromocriptine | 0
    treated with IV dantrolene | 0
    discontinuation of causative agents | 0
    cooling blanket | 0
    antipyretics | 0
    IV fluids | 0
    SS considered | 0
    escalating doses of ziprasidone | 0
    unaltered use of duloxetine | 0
    unaltered use of lithium | 0
    administer bromocriptine | 0
    dantrolene scheduled | 0
    electroencephalography showed generalized slowing | 0
    no seizure activity | 0
    MRI brain no acute finding | 0
    afebrile | 72
    improved leukocytosis | 72
    no antibiotics | 72
    no lumbar puncture | 72
    autonomic dysregulation resolved | 96
    cessation of labile blood pressures | 96
    supplemental oxygen requirements ceased | 96
    more awake | 96
    less rigid in extremities | 96
    unable to participate in meaningful interview | 96
    dantrolene increased to 100 mg TID | 96
    stable | 120
    transferred out of NCCU | 120

    60 years old | 0
    female | 0
    nursing home patient | 0
    bipolar affective disorder | 0
    hypertension | 0
    hypothyroidism | 0
    paraplegia | 0
    increasing confusion | 0
    admitted to senior behavioral facility | 0
    unable to communicate | -168
    tachycardia | -168
    tachypnea | -168
    flushing | -168
    diaphoresis | -168
    fevers greater than 38°C | -168
    transferred to NCCU | -168
    encephalopathic | 0
    tachypneic | 0
    tachycardic | 0
    hypoxemic | 0
    generalized rigidity | 0
    hyperreflexia | 0
    leukocytosis | 0
    acute kidney injury | 0
    elevated serum creatinine phosphokinase | 0
    procalcitonin elevated | 0
    C-reactive protein within normal limits | 0
    episodes of hypotension | 0
    episodes of hypertension | 0
    possible sepsis | 0
    NMS | 0
    serotonin syndrome | 0
    non-convulsive status epilepticus | 0
    CNS pathology | 0
    blood cultures obtained | 0
    urine cultures obtained | 0
    sputum cultures obtained | 0
    lumbar puncture considered | 0
    medical records obtained | 0
    receiving increasing doses of ziprasidone | -168
    haloperidol | -168
    lithium | -168
    duloxetine | -168
    oxybutynin | -168
    baclofen | -168
    treated with IV bromocriptine | 0
    treated with IV dantrolene | 0
    discontinuation of causative agents | 0
    cooling blanket | 0
    antipyretics | 0
    IV fluids | 0
    SS considered | 0
    escalating doses of ziprasidone | 0
    unaltered use of duloxetine | 0
    unaltered use of lithium | 0
    administer bromocriptine | 0
    dantrolene scheduled | 0
    electroencephalography showed generalized slowing | 0
    no seizure activity | 0
    MRI brain no acute finding | 0
    afebrile | 72
    improved leukocytosis | 72
    no antibiotics | 72
    no lumbar puncture | 72
    autonomic dysregulation resolved | 96
    cessation of labile blood pressures | 96
    supplemental oxygen requirements ceased | 96
    more awake | 96
    less rigid in extremities | 96
    unable to participate in meaningful interview | 96
    dantrolene increased to 100 mg TID | 96
    stable | 120
    transferred out of NCCU | 120

    60 years old | 0
    female | 0
    nursing home patient | 0
    bipolar affective disorder | 0
    hypertension | 0
    hypothyroidism | 0
    paraplegia | 0
    increasing confusion | 0
    admitted to senior behavioral facility | 0
    unable to communicate | -168
    tachycardia | -168
    tachypnea | -168
    flushing | -168
    diaphoresis | -168
    fevers greater than 38°C | -168
    transferred to NCCU | -168
    encephalopathic | 0
    tachypneic | 0
    tachycardic | 0
    hypoxemic | 0
    generalized rigidity | 0
    hyperreflexia | 0
    leukocytosis | 0
    acute kidney injury | 0
    elevated serum creatinine phosphokinase | 0
    procalcitonin elevated | 0
    C-reactive protein within normal limits | 0
    episodes of hypotension | 0
    episodes of hypertension | 0
    possible sepsis | 0
    NMS | 0
    serotonin syndrome | 0
    non-convulsive status epilepticus | 0
    CNS pathology | 0
    blood cultures obtained | 0
    urine cultures obtained | 0
    sputum cultures obtained | 0
    lumbar puncture considered | 0
    medical records obtained | 0
    receiving increasing doses of ziprasidone | -168
    haloperidol | -168
    lithium | -168
    duloxetine | -168
    oxybutynin | -168
    baclofen | -168
    treated with IV bromocriptine | 0
    treated with IV dantrolene | 0
    discontinuation of causative agents | 0
    cooling blanket | 0
    antipyretics | 0
    IV fluids | 0
    SS considered | 0
    escalating doses of ziprasidone | 0
    unaltered use of duloxetine | 0
    unaltered use of lithium | 0
    administer bromocriptine | 0
    dantrolene scheduled | 0
    electroencephalography showed generalized slowing | 0
    no seizure activity | 0
    MRI brain no acute finding | 0
    afebrile | 72
    improved leukocytosis | 72
    no antibiotics | 72
    no lumbar puncture | 72
    autonomic dysregulation resolved | 96
    cessation of labile blood pressures | 96
    supplemental oxygen requirements ceased | 96
    more awake | 96
    less rigid in extremities | 96
    unable to participate in meaningful interview | 96
    dantrolene increased to 100 mg TID | 96
    stable | 120
    transferred out of NCCU | 120

    60 years old | 0
    female | 0
    nursing home patient | 0
    bipolar affective disorder | 0
    hypertension | 0
    hypothyroidism | 0
    paraplegia | 0
    increasing confusion | 0
    admitted to senior behavioral facility | 0
    unable to communicate | -168
    tachycardia | -168
    tachypnea | -168
    flushing | -168
    diaphoresis | -168
    fevers greater than 38°C | -168
    transferred to NCCU | -168
    encephalopathic | 0
    tachypneic | 0
    tachycardic | 0
    hypoxemic | 0
    generalized rigidity | 0
    hyperreflexia | 0
    leukocytosis | 0
    acute kidney injury | 0
    elevated serum creatinine phosphokinase | 0
    procalcitonin elevated | 0
    C-reactive protein within normal limits | 0
    episodes of hypotension | 0
    episodes of hypertension | 0
    possible sepsis | 0
    NMS | 0
    serotonin syndrome | 0
    non-convulsive status epilepticus |