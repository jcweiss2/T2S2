30 years old | 0
woman | 0
history of intravenous drug use (IVDU) | 0
admitted to outside hospital | 0
bacterial pneumonia | 0
infective endocarditis suspected | 0
computed tomography chest revealed septic pulmonary emboli | 0
transesophageal echocardiography (TEE) confirmed infective endocarditis | 0
ravaged tricuspid valve with fenestrations | 0
wide-open tricuspid regurgitation with flail segments | 0
multiple mobile tricuspid valve vegetations | 0
preserved left ventricular ejection fraction | 0
consultations with cardiology | 0
consultations with cardiac surgery | 0
consultations with infectious disease | 0
decision to proceed with tricuspid valvulectomy | 0
blood cultures confirmed methicillin-susceptible Staphylococcus aureus | 0
valve cultures confirmed methicillin-susceptible Staphylococcus aureus | 0
postoperative refractory hypoxemia | 0
partial pressure of oxygen 60 mmHg on 100% FiO2 with mechanical ventilation | 0
chest radiography showed no hemopneumothorax | 0
chest radiography showed no pulmonary edema | 0
chest radiography showed no lung consolidation | 0
attempts to aggressively diurese | 0
inhaled epoprostenol initiated | 0
neuromuscular blockade initiated | 0
prone positioning | 0
venovenous extracorporeal membrane oxygenation (ECMO) cannulation | 0
partial pressure of oxygen 145-165 mmHg on ECMO | 0
ECMO specialty transport team retrieval | 0
transthoracic echocardiography performed | 0
TEE performed | 0
ventricularization of the right heart | 0
wide-open systolic regurgitant flow from right ventricle to right atrium | 0
dilated right ventricle | 0
interatrial septum bowing from right to left | 0
ECMO cannulas correctly positioned | 0
return cannula at junction of right atrium and superior vena cava | 0
outflow jet directed into right atrium near interatrial septum | 0
drainage cannula at junction of right atrium and inferior vena cava | 0
reversal of hepatic vein flow | 0
new interatrial communication (patent foramen ovale) | 0
significant right-to-left flow | 0
taken to operating room for PFO closure | 24
tricuspid valve replacement with 31-mm St. Jude Epic porcine bioprosthetic valve | 24
intraoperative TEE showed no residual tricuspid regurgitation | 24
no residual right-to-left shunt by bubble study | 24
deccannulated from ECMO | 24
extubated | 24
remained in hospital for 19 days | 24
IV antibiotic therapy | 24
treatment with addiction specialist | 24
left hospital against medical advice | 456
lost to follow-up | 456
opioid dependence | 0
