68 years old | 0
male | 0
admitted to the hospital | 0
chest pain | 0
acute dyspnea | 0
type 2 diabetes mellitus | -672
hypertension | -672
oral metformin hydrochloride | -672
valsartan | -672
poorly controlled diabetes | -672
hemoglobin A1c 7.7% | -672
white blood cell count high | 0
C-reactive protein high | 0
myocardial enzymes lactate dehydrogenase elevated | 0
aspartate aminotransferase elevated | 0
troponin-T positive | 0
anti-human immunodeficiency virus antibody test negative | 0
percutaneous coronary intervention | 0
intubated | 0
invasive mechanical ventilation | 0
intravenous antibiotics | 0
levofloxacin | 0
ampicillin/sulbactam | 0
vasodilators | 0
diuretics | 0
progressive respiratory failure | 0
fraction of inspired oxygen 80% | 0
positive end expiratory pressure 15 cmH2O | 0
ARDS | 120
extracorporeal membrane oxygenation | 120
intravenous methylprednisolone | 120
prednisolone | 120
respiratory condition improved | 192
blood in stool | 192
dual antiplatelet therapy | 192
monitor closely | 192
condition stabilized | 240
discontinued extracorporeal membrane oxygenation | 240
extubated | 288
prednisolone dose tapered | 408
respiratory condition worsened | 432
re-intubated | 432
intravenous methylprednisolone | 432
respiratory condition improved | 504
prednisolone reduced | 504
bloody diarrhea worsened | 528
colonoscopy | 528
multiple large ulcers in sigmoid colon and rectum | 528
biopsied | 528
histopathological examination | 528
infiltration of neutrophils and lymphocytes | 528
CMV-positive cells | 528
CMV pp65 antigenemia positive | 528
diagnosed with CMV enterocolitis | 528
ganciclovir | 600
improved peripheral blood C7-HRP test results | 600
bloody diarrhea continued | 1080
abdominal pain | 1080
abdominal computed tomography | 1080
free air | 1080
gastrointestinal perforation | 1080
poor general condition | 1080
no surgical treatment | 1080
died | 1080
autopsy | 1080
full-thickness necrotic intestinal wall tissue | 1080
severe infiltration of necrotic tissue with ameba | 1080
Entamoeba histolytica trophozoites | 1080
fulminant amebic colitis | 1080
CMV enterocolitis | 1080