65 years old | 0
female | 0
liver cirrhosis | -6720
chronic hepatitis B | -6720
hepatocellular carcinoma | 0
admitted to the hospital | 0
premedication with glycopyrrolate | 0
general anesthesia induced | 0
intubated and ventilated mechanically | 0
monitored by electrocardiography | 0
monitored by arterial blood pressure | 0
monitored by central venous pressure | 0
monitored by SpO2 | 0
stable vital signs | 0
hepatectomy started | 0
CUSA used | 0
sudden decrease in arterial blood pressure | 1
systolic blood pressure <40 mmHg | 1
end-tidal carbon dioxide <26 mmHg | 1
SpO2 <50% | 1
tachycardia | 1
ST elevation on EKG | 1
resuscitation with colloid and catecholamines | 1
intraoperative ultrasonography | 1
massive air emboli in left and right heart | 1
diagnosed with VAE and PAE | 1
arterial blood gas analysis | 1
catecholamine administration | 1.17
systolic blood pressure maintained | 1.17
heart rate maintained | 1.17
central venous pressure maintained | 1.17
end-tidal carbon dioxide restored | 1.17
ABGA at 30 minutes after episode | 1.5
norepinephrine infusion continued | 1.5
fluid resuscitation continued | 1.5
air emboli in left heart disappeared | 2.17
hepatectomy restarted | 2.17
hepatectomy completed | 5
mechanical ventilation | 5
intensive care unit | 5
intubated | 5
ventilated mechanically | 5
responded to intense pain | 5
systolic pressure maintained | 5
norepinephrine infusion | 5
postoperative laboratory findings | 5
abnormal PT/PTT | 5
abnormal fibrinogen | 5
abnormal d-dimer | 5
abnormal antithrombin III | 5
abnormal CK-MB | 5
abnormal troponin-T | 5
postoperative EKG | 5
ST elevation | 5
POD 1 | 24
EKG findings recovered | 24
trans-thoracic echocardiogram | 24
vital signs stable | 24
norepinephrine infusion tapered out | 24
POD 5 | 120
mental status unchanged | 120
brain CT | 120
brain MRI | 120
multiple acute cerebral infarctions | 120
POD 11 | 264
weaned to spontaneous ventilation | 264
extubated | 264
POD 15 | 360
vital signs unstable | 360
intravenous administration of catecholamines | 360
panperitonitis confirmed | 360
gram (+) cocci on peritoneal culture | 360
POD 31 | 744
cardiac arrest | 744
septic shock | 744
expired | 744