66 years old | 0
female | 0
referred to urology department | -4320
lower abdominal pain | -4320
vital signs within normal range | -4320
unremarkable urine/blood investigations | -4320
CT abdomen/pelvis | -4320
large 35mm right sided PUJ calculus | -4320
xanthogranulomatous pyelonephritic (XGP) kidney | -4320
mild abdominal pain | -4320
lack of flank pain | -4320
lack of urinary symptoms | -4320
unremarkable blood investigations | -4320
outpatient management | -4320
plan for elective surgery | -4320
discussed management options | -4320
consented for endoscopic procedure | -4320
ureteropyeloscopy and lasertripsy surgery | -2160
urine culture with mixed growth | -2160
observed polyps in right ureter | -2160
pus in renal pelvis | -2160
poor visibility | -2160
increased risk of sepsis | -2160
discontinued procedure | -2160
plan for repeat procedure | -2160
intraoperative retrograde pyelogram (RPG) | -2160
no evidence of fistula | -2160
ureteric stent insertion | -2160
recovered well post-operatively | -2160
discharged with oral antibiotics | -2160
ureteric biopsies of polyps | -2160
inflammatory changes | -2160
repeat pyeloscopy procedure | -1728
small volume of renal calculi | -1728
treated with lasertripsy | -1728
no reportable complications | -1728
ureteric stent insertion | -1728
unremarkable intraoperative RPG | -1728
ureteric stent removed | -1680
severe sepsis | -1440
hypothermia | -1440
hypotension | -1440
tachycardia | -1440
tachypnoea | -1440
elevated inflammatory markers | -1440
moderate renal impairment | -1440
positive urinalysis | -1440
leukocytes positive | -1440
nitrites positive | -1440
blood positive | -1440
urine culture with mixed growth | -1440
Proteus mirabilis in blood cultures | -1440
CT KUB | -1440
right sided peri-nephric stranding | -1440
previous findings | -1440
initial resuscitation | -1440
treatment for sepsis | -1440
emergency cystoscopy | -1440
RPG and stent insertion | -1440
RPG revealed uretero-duodenal fistula | -1440
contrast tracking to duodenum | -1440
transfer to tertiary hospital ICU | -1440
right sided nephrectomy | -1440
laparoscopic approach | -1440
bowel mobilisation | -1440
identification of ureter | -1440
conversion to open surgery | -1440
adhesiolysis | -1440
haemostasis | -1440
no duodenum resection | -1440
post-operative management | -1440
tolerating fluids by Day 3 | -1440
full diet by Day 5 | -1440
uneventful recovery | -1440
discharged home | -1440
follow-up appointment | 4320
nil urinary symptoms | 4320
nil pain issues | 4320
CT abdomen/pelvis | 4320
no abnormal collections | 4320
