66 years old | 0
male | 0
admitted to the hospital | 0
intermittent high-grade fever | -216
generalized dull-aching abdominal pain | -216
passing turbid urine | -240
decrease in urine output | -240
swelling of both feet | -240
treated with intravenous medications | -168
type II diabetes mellitus | -2628
conscious | 0
afebrile | 0
tachycardic | 0
heart rate of 136/min | 0
blood pressure was 110/70 mmHg | 0
renal angle tenderness bilaterally | 0
high total leukocyte counts | 0
elevated urea and creatinine levels | 0
pyuria with leukocyte esterase positivity | 0
activated partial thromboplastin time was prolonged | 0
sepsis-induced coagulopathy | 0
enlarged kidneys with bilateral renal abscesses | 0
emergency ultrasound-guided drainage of renal abscesses | 0
transfusion of blood products | 0
coagulopathy | 0
pus smear from renal abscesses showed septate fungal hyphae | 0
intravenous meropenem | 0
intravenous voriconazole | 0
intravenous amphotericin B | 0
cultures from both renal abscesses revealed growth of Aspergillus fumigatus | 0
worsening renal function | 24
acute pulmonary edema | 24
hyperkalemia | 24
metabolic acidosis | 24
hemodialysis | 24
noninvasive ventilation | 24
sudden cardiac arrest | 216
aspiration | 216
succumbed to his illness | 216