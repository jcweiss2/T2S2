47 years old | 0
female | 0
Caucasian | 0
altered mental status | -24
agitation | -24
confusion | -24
fever | -24
respiratory distress | -24
sinusitis | -24
chronic sinusitis | 0
nasal polyp removal | 0
diabetes mellitus type II | 0
no tobacco use | 0
no alcohol use | 0
no illicit drug use | 0
rectal temperature of 106.2 °F | 0
heart rate of 141 beats per minute | 0
blood pressure of 107/59 mmHg | 0
respiratory rate of 32 breaths per minute | 0
alert but not oriented to time, place and person | 0
respiratory distress using accessory muscles of respiration | 0
diaphoretic skin | 0
agitated | 0
pupils equal and reactive to light | 0
no lesions in the nares or nasal drainage | 0
nuchal rigidity | 0
photophobia | 0
right upper quadrant tender to palpation | 0
distended right upper quadrant | 0
rebound tenderness | 0
unremarkable cardiac examination | 0
sodium of 135 mmol/L | 0
potassium of 3.3 mmol/L | 0
chloride of 98 mmol/L | 0
bicarbonate of 23 mmol/L | 0
blood urea nitrogen of 12 mg/dL | 0
creatinine of 0.6 mg/dL | 0
glucose of 542 mg/dL | 0
white blood cell count of 35.1 × 10^9 cells/L | 0
granulocytes of 95.7% | 0
hemoglobin of 12.1 mg/dL | 0
MCV of 75.5 fL | 0
hematocrit of 40.3% | 0
platelets of 258,000/mcL | 0
started on empiric antibiotics with ceftriaxone, vancomycin and acyclovir | 0
lumbar puncture | 0
opening pressure of 46 mm H2O | 0
cloudy and bloody cerebrospinal fluid | 0
WBC count of 820/mm^3 in CSF | 0
red blood cell count of 5500/mm^3 in CSF | 0
glucose concentration of 177 mg/dl in CSF | 0
protein concentration of 672 mg/dl in CSF | 0
Gram stain showed gram-positive cocci in chains | 0
CSF glucose to blood glucose ratio of 0.375 | 0
unremarkable head CT | 0
negative blood cultures | 0
admitted to the intensive care unit | 0
CSF culture grew S. agalactiae | 24
sensitive to gentamicin and ampicillin | 24
antibiotics changed to gentamicin and ampicillin | 24
no change in mental status after 4 days | 96
repeat CT of the head showed a 4 cm acute intracerebral hemorrhage | 96
intracerebral hemorrhage in the right frontal convexity | 96
surrounding edema and mass effect | 96
extubated after a week | 168
opening eyes to verbal stimuli but not following commands | 168
went in respiratory distress and was reintubated | 168
repeat head CT showed intraparenchymal hematoma increased in size | 168
new 1.7 cm hematoma in the left frontal lobe | 168
diffuse cerebral edema and a right to left midline shift | 168
neurosurgery did not recommend draining the hemorrhages | 168
developed Clostridium difficile associated diarrhea | 168
treated with metronidazole | 168
antibiotics course for meningitis was successfully completed | 336
mental status improved significantly | 336
developed a health care associated pneumonia | 336
treated for pneumonia | 336
discharged at her baseline mental status | 720