72 years old | 0
male | 0
admitted to hospital | 0
gastric cancer | -672
distal gastrectomy | -672
right hepatic lobectomy | -672
lymph node metastases | -672
combination chemotherapy | -336
paclitaxel | -336
S-1 | -336
paraaortic lymph node metastases | -168
docetaxel | 0
methyl predonine | 0
high-grade fever | 24
low blood pressure | 24
white blood cell count of 13,550/L | 24
red blood cell count of 2,420,000/L | 24
blood platelet count of 109,000/L | 24
aspartate aminotransferase of 1,112 IU/L | 24
alanine aminotransferase of 774 IU/L | 24
CRP of 4.6 mg/dl | 24
septicemia unknown etiology | 24
dopamine infusion | 24
broad-band antibiotics | 24
liver and renal dysfunction | 48
leucocytosis | 48
high value of C-reactive protein | 48
hemodialysis | 48
respiratory support | 48
death | 120
blood bacterial culture revealed E. coli | 120
autopsy | 120
bone marrow histology | 120
residual lymph node metastases | 120
multiple occult liver abscesses | 120
gram-negative rods | 120
fungi | 120
fatal E. coli septicemia | 120
immuno compromised host | 120
anti-cancer drug treatment | 0