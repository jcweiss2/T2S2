30 years old | 0
female | 0
homozygous sickle cell disease (SCD) | 0
respiratory failure | 0
neurological deterioration | 0
vaso-occlusive crisis | 0
admitted to intensive care unit (ICU) | 0
transfer from outside hospital | 0
acute vaso-occlusive crisis | -72
fever | -72
