81 years old | 0
female | 0
admitted to the hospital | 0
coronary artery disease | -8760
type 2 diabetes mellitus | -8760
endometrial carcinoma | -26280
aseptic meningitis | -17520
syncope | -168
seizure | -168
dysarthria | -168
runny nose | -168
nausea | -168
diarrhea | -168
ciprofloxacin | -168
profound lethargy | -120
bilateral weakness | -120
cranial nerve abnormalities | -120
viral encephalitis | -120
intravenous acyclovir | -120
right frontal brain mass | -120
brain CT | -120
CT imaging of the chest | -120
CT imaging of the abdomen | -120
CT imaging of the pelvis | -120
transferred to the institution | 0
stuporous | 0
left gaze preference | 0
anisocoric pupils | 0
right upper extremity flaccid | 0
right lower extremity flaccid | 0
minimal withdrawal in left lower extremity | 0
hyponatremia | 0
hyperglycemia | 0
mild anemia | 0
brain MRI | 0
high FLAIR signal | 0
tubular/lobulated/ring enhancement | 0
lumbar puncture | 0
CSF studies | 0
elevated protein level | 0
ampicillin | 0
meropenem | 0
vancomycin | 0
voriconazole | 0
pyrimethamine/sulfadiazine | 0
intravenous dexamethasone | 0
open brain biopsy | 72
Gram-positive rods | 72
L. monocytogenes infection | 72
discontinued antibiotics | 72
steroids tapered off | 72
transferred to the regular floor | 240
percutaneous endoscopic gastrostomy | 240
transferred to a rehabilitation facility | 768
completed antibiotic treatment | 1344
eye opening to verbal stimuli | 768
command-following with left upper extremity | 768
incomprehensible sounds | 768
pupils 4 mm bilaterally | 768
reactive to light | 768
partial left third cranial nerve palsy | 768
left nasolabial fold flattening | 768
persistent significant weakness | 768