59 years old | 0
female | 0
mitral valve insufficiency | -12000
MVR surgery | -12000
prosthetic mitral valve dysfunction | -240
redo MVR | 0
hemolysis | 0
decrease in hemoglobin level | 0
acute renal failure | 0
urgent-start hemodialysis | 0
severe mitral valve dysfunction | 0
PRBC transfusion | 0
weak | -720
lethargic | -720
admitted to hospital | 0
exacerbation of symptoms | 0
Hb level 6.3 | 0
HCT 19.7 | 0
RBC 2.27 | 0
WBC 3700 | 0
PLT 235000 | 0
MCHC 32 | 0
MCV 86.8 | 0
MCH 27.8 | 0
PT 15.8 | 0
PTT 54.4 | 0
INR 1.2 | 0
Na 140 | 0
K 4 | 0
BUN 86 | 0
Cr 1.3 | 0
Uric Acid 9.1 | 0
LDH 3418 | 0
AST 64 | 0
ALT 46 | 0
Alph 230 | 0
Bill total 9.6 | 0
Bill direct 2.4 | 0
Bill indirect 7.5 | 0
candidate for blood transfusion | 0
blood transfusion initiated | 0
fever | 0
headache | 0
chills | 0
back pain | 0
urine discoloration | 0
blood transfusion stopped | 0
therapeutic measures | 0
aerobic and anaerobic blood culture | 0
blood smear | 0
antibody screening test | 0
Coombs test | 0
Coombs Wright test | 0
anti-E positive | 0
anti-c positive | 0
anti-Kell positive | 0
PRBC transfusion | 0
Hb level raised to 10.5 | 0
surgery | 0
tricuspid valve repair | 0
aortic valve replacement | 0
MVR | 0
ICU admission | 0
extubated | 48
postoperative lab tests | 48
no evidence of hemolysis | 48
Hb level acceptable | 48
sepsis | 504
expired | 504