43 years old | 0
female | 0
admitted to the hospital | 0
fever | -240
dry cough | -240
mild respiratory distress | -72
peripheral capillary oxygen saturation 88%-89% | -72
diagnosed with COVID-19 | -72
polycystic ovarian disease | 0
blood pressure 140/90 mmHg | 0
pulse rate 88 beats/min | 0
respiratory rate 20 breaths/min | 0
SpO2 92% | 0
bilateral decrease in air entry | 0
total leucocyte count 11650 cells/µL | 0
neutrophils 88% | 0
lymphocytes 8% | 0
C-reactive protein 16.44 mg/L | 0
procalcitonin 9.52 ng/mL | 0
lactate dehydrogenase 282 IU/L | 0
ferritin 158 ng/mL | 0
D-dimer 775.84 ng/mL | 0
interleukin-6 18.55 pg/mL | 0
elevated liver enzymes | 0
arterial oxygen partial pressure 39.0 mmHg | 0
severe hypoxia | 0
non-rebreather mask with 15 L/min of oxygen | 0
100% oxygen saturation | 0
echocardiography | 0
ejection fraction 60% | 0
chest physiotherapy | 0
incentive spirometry | 0
intravenous remdesivir | 0
intravenous dexamethasone | 0
oral doxycycline | 0
low molecular weight heparin | 0
multivitamins | 0
antibiotics | 0
nebulization | 0
oxygen requirement decreased | 168
chest CT | 192
CT severity index score 12/25 | 192
weaned off oxygen | 288
discharged | 456
procalcitonin level persistently elevated | 456
investigating the persistently elevated procalcitonin level | 456
neck examination | 456
ultrasonography of the neck | 456
nodule in the left lobe of the thyroid gland | 456
fine-needle aspiration cytology | 456
malignant epithelial neoplasm | 456
metastatic carcinoma | 456
calcitonin level 406 pg/mL | 456
carcinoembryonic antigen not elevated | 456
positron emission tomography-CT | 456
fluorodeoxyglucose-avid nodule | 456
medullary thyroid carcinoma | 456
total thyroidectomy | 1400
central lymph node dissection | 1400
histological examination | 1400
lymphovascular invasion | 1400
eleven lymph nodes positive | 1400
second radical neck dissection | 1680
six positive nodes | 1680
procalcitonin level dropped | 1680
calcitonin level dropped | 1680
multiple endocrine neoplasia type II syndrome ruled out | 1680
levothyroxine supplementation | 2160
external beam radiotherapy | 2160
no evidence of recurrence | 2160