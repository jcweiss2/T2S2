55 years old | 0
    female | 0
    hepatitis C | 0
    intravenous drug use | 0
    alcohol abuse | 0
    Child-Pugh B liver cirrhosis | 0
    abdominal pain | 0
    diarrhea | 0
    fevers | 0
    confusion | 0
    no history of colonic disease | 0
    computed tomography abdomen | 0
    mildly dilated proximal large bowel | 0
    no fat stranding | 0
    no colonic wall thickening | 0
    stool PCR positive for campylobacter species | 0
    treatment with azithromycin | 0
    treatment with ceftriaxone | 0
    treatment with metronidazole | 0
    intravenous fluids | 0
    electrolyte replacement | 0
    deterioration | 0
    long admission to intensive care unit | 0
    aspiration pneumonitis | 0
    type 2 myocardial infarction | 0
    renal failure | 0
    metabolic acidosis | 0
    intubation | 0
    vasopressors | 0
    dialysis | 0
    transthoracic echocardiography | 0
    lumbar puncture | 0
    blood cultures | 0
    CT scan head | 0
    CT scan chest | 0
    CT scan abdomen | 0
    CT scan pelvis | 0
    no alternative source of sepsis | 0
    antibiotics escalated to piperacillin/tazobactam | 0
    bloody diarrhea | 16*24
    ongoing refractory multi-organ dysfunction | 16*24
    CT abdomen | 16*24
    colonic wall thickening | 16*24
    most prominent in sigmoid and rectum | 16*24
    no gross dilatation | 16*24
    no intramural gas | 16*24
    no free gas | 16*24
    no obvious bleeding points | 16*24
    upper endoscopy | 16*24
    excluded varices | 16*24
    excluded ulcers | 16*24
    transfer to tertiary hospital | 16*24
    ongoing intensive care management | 16*24
    surgical review | 16*24
    emergent laparotomy | 16*24
    viable mildly dilated colon | 16*24
    clear ascites | 16*24
    no evidence of ischemia | 16*24
    no necrosis | 16*24
    no perforation | 16*24
    nodular liver | 16*24
    remainder of bowel normal | 16*24
    flexible sigmoidoscopy | 16*24
    discontinuous areas of non-bleeding ulcerated mucosa | 16*24
    biopsies taken | 16*24
    discussed with intensive care team | 16*24
    discussed with infectious diseases team | 16*24
    findings consistent with infective colitis | 16*24
    septic shock | 16*24
    MODS | 16*24
    returned to ICU | 16*24
    antibiotics changed to daptomycin | 16*24
    antibiotics changed to ciprofloxacin | 16*24
    antibiotics changed to fluconazole | 16*24
    antibiotics changed to metronidazole | 16*24
    deterioration over next 12 hours | 16*24+12
    worsening hemodynamic instability | 16*24+12
    increasing noradrenaline | 16*24+12
    increasing vasopressin | 16*24+12
    re-look laparotomy | 16*24+12
    grossly dilated colon | 16*24+12
    no perforation | 16*24+12
    no full thickness ischemia | 16*24+12
    subtotal colectomy | 16*24+12
    end ileostomy | 16*24+12
    distal sigmoid mucous fistula | 16*24+12
    immediate postoperative improvement | 16*24+12
    vasopressin ceased | 16*24+12
    noradrenaline infusion halved | 16*24+12
    continued improvement until postoperative day 3 | (16*24+12) + 3*24
    escalating vasopressor requirements | (16*24+12) + 3*24
    acidosis | (16*24+12) + 3*24
    liver failure | (16*24+12) + 3*24
    respiratory failure | (16*24+12) + 3*24
    death | (16*24+12) + 4*24
    histology showed infectious colitis | (16*24+12) + 4*24
    histology showed ischemia | (16*24+12) + 4*24
    macroscopic mucosal ulceration | (16*24+12) + 4*24
    no infarcted bowel | (16*24+12) + 4*24
    no pseudomembranes | (16*24+12) + 4*24
    microscopic congestion | (16*24+12) + 4*24
    neutrophilic infiltration | (16*24+12) + 4*24
    fibrin thrombi | (16*24+12) + 4*24
    no architectural distortion | (16*24+12) + 4*24
    no cryptitis | (16*24+12) + 4*24
    no crypt abscesses | (16*24+12) + 4*24
    absence of inflammatory bowel disease features | (16*24+12) + 4*24
    toxic megacolon | 16*24
    Campylobacter colitis | 0
    septic shock | 16*24
    MODS | 16*24
    Child-Pugh B cirrhosis | 0
    alcohol abuse | 0
    intravenous drug use | 0
    hepatitis C | 0
    death due to comorbidities | (16*24+12) + 4*24
    colectomy performed | 16*24+12
    postoperative improvement | 16*24+12
    subsequent deterioration | (16*24+12) + 3*24
    no corticosteroid use | 0
    no inflammatory bowel disease | 0
    no colonic perforation | 16*24+12
    no uncontrolled bleeding | 16*24+12
    no alternative sepsis source | 0
    initial laparotomy findings | 16*24
    second laparotomy findings | 16*24+12
    histopathological confirmation of infectious colitis | (16*24+12) + 4*24
    