60 years old| 0
male | 0
history of dysphagia | 0
barium swallow study | 0
aspirated a large amount of barium | -24
dyspneic | -24
labored breathing | -24
respiratory rate >35 breaths/min | -24
tachycardia (heart rate >120 beat/min) | -24
blood pressure 160/100 mmHg | -24
SPO2 <90% despite oxygen flow 15lit/min by mask | -24
hypoxemia (PO2 86.7 mmHg on oxygen flow 15 lit/min) | -24
crepitation in both lung bases | -24
chest X-ray findings: barium sulfate aspiration involving right and left main stem bronchi, bronchus intermedius, lower lobe basal, and segmental bronchi resembling a tree-in-bud appearance | -24
shifted to intensive care unit (ICU) | -24
intubation | -24
positive pressure mechanical ventilation | -24
bronchioalveolar lavage (BAL) | -24
large amount of barium particles suctioned | -24
postural drainage techniques | -24
developed shock | 4
fluid resuscitation | 4
inotropic support (infusion noradrenaline) | 4
injection hydrocortisone 100 mg thrice daily | 4
broad-spectrum antibiotics with coverage of gut flora | 4
nebulization with N-acetylcystein | 4
hemodynamically stable | 24
extubated | 24
oxygen saturation of 99% on 5 litres of oxygen | 24
shifted to ward | 72
aspirated oral feed and gastric contents | 144
shifted to ICU | 144
succumbed to sepsis | 336
