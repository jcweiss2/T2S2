25 years old | 0
male | 0
athlete | 0
admitted to the hospital | 0
heat stroke | -1
rhabdomyolysis | -1
ischaemic hepatitis | -1
severely hypotensive | 0
unrecordable blood pressure | 0
confused | 0
Glasgow Coma Score of 10 | 0
temperature of 105.4°F | 0
sweaty | 0
tachycardic | 0
heart rate of 160 bpm | 0
systolic blood pressure of 90 mm Hg | 0
intravenous fluids | 0
inotropic support with ephedrine | 0
CT scan of brain | 0
normal CT scan of brain | 0
intravenous co-amoxiclav | 0
elevated creatinine phosphokinase level | 24
rhabdomyolysis | 24
serum alanine aminotransferase rising | 24
ALT level of 143 U/l | 24
transferred from intensive care to general medical ward | 24
ALT peaked | 48
liver screen normal | 48
negative viral screen | 48
negative autoimmune screen | 48
mildly raised ferritin levels | 48
normal ultrasound of liver | 48
intravenous N-acetyl cysteine | 48
discharged home | 72
CPK improving | 72
ALT improving | 72
follow-up | 168
heat stroke associated with rhabdomyolysis and ischaemic hepatitis | -1
running the final stages of a marathon | -1
collapse | 0
seizure | -24
hypoglycaemia | -24
myalgia | -24
deranged liver function | -24
hypoxic hepatitis | 0
vasopressor therapy | 0
liver injury | 0
NAC limits liver injury | 48
NAC started | 48
transplant-free survival | 168
orthotopic liver transplantation | 168
grade 1 or 2 encephalopathy | 168
better 1-year survival | 720
ALT level peaked at 2,912 U/l | 48
CPK level peaked at 178,850 U/l | 24
random glucose | 0
INR | 0
lactate | 0
drugs of abuse screen negative | 0
urine myoglobin test negative | 0
hepatitis B surface antigen negative | 48
hepatitis B core IgM antibody negative | 48
hepatitis A IgM antibody negative | 48
hepatitis C antibody negative | 48
anti-smooth muscle antibody negative | 48
anti-mitochondrial antibody negative | 48
anti-nuclear antibody negative | 48
ferritin | 48
White blood cells | 0
Neutrophils | 0
Haemoglobin | 0
Platelets | 0
Creatinine | 0
Urea | 0
Potassium | 0
Random glucose | 0
INR | 0
CPK | 0
ALP | 0
ALT | 0
GGT | 0
Bilirubin | 0
Lactate | 0