73 years old | 0
    female | 0
    admitted with new-onset atrial flutter | 0
    fatigue | 0
    dizziness | 0
    dyspnoea | 0
    atrial flutter | 0
    rapid regular pulse rate | 0
    normal lung sounds | 0
    normal heart sounds | 0
    no peripheral oedema | 0
    transthoracic echocardiography | 0
    transoesophageal echocardiography | 0
    heterogeneous isoechoic immobile mass | 0
    lobulated margins | 0
    attached to free anterior wall of right atrium | 0
    base of tricuspid valve | 0
    circular hypoechoic pericardial effusion | 0
    compression of right atrium | 0
    pericardiocentesis | 0
    cell-rich pericardial fluid | 0
    protein-rich pericardial fluid | 0
    lactate hydrogenase-rich pericardial fluid | 0
    reactively changed cell population | 0
    histiocytes | 0
    mesothelial cells | 0
    no atypical cell populations | 0
    haemoglobin 11.9 g/dL | 0
    LDH 322 U/L | 0
    C-reactive protein 6.3 mg/dL | 0
    pro-BNP II 2834 pg/mL | 0
    serum protein 5.9 g/dL | 0
    normal carcinoembryonic antigen | 0
    normal CA 125 | 0
    normal CA 15-3 | 0
    normal CA 19-9 | 0
    normal alpha-fetoprotein | 0
    cardiac MRI | 0
    tumourous myocardial isointense mass | 0
    diffuse infiltration of myocardium | 0
    extension into pericardium | 0
    computed tomography of skull | 0
    computed tomography of thorax | 0
    computed tomography of abdomen | 0
    computed tomography of pelvis | 0
    breast sonography | 0
    mammography | 0
    dermatologic screening | 0
    gynaecologic screening | 0
    endoscopy of upper gastrointestinal tract | 0
    endoscopy of lower gastrointestinal tract | 0
    no extracardiac disease | 0
    no enlarged lymph nodes | 0
    referred to cardiac surgery centres | -720
    deemed inoperable | -720
    active surveillance | -720
    best supportive therapy | -720
    fatigue | -504
    dizziness | -504
    AV block II type Mobitz 2 | -504
    transthoracic echocardiography | -504
    massive progression of tumour mass | -504
    transoesophageal echocardiography | -504
    subtotal obstruction of tricuspid valve | -504
    cardiac MRI | -504
    infiltration of cardiac base adjacent to atrial septum | -504
    suspected transpericardial infiltration of diaphragm | -504
    bilateral axillary lymph nodes | -504
    extracardiac metastases | -504
    epicardial right ventricle single lead pacemaker | -504
    axillary lymph node excision | -504
    diffuse large B-cell non-Hodgkin lymphoma | -504
    port catheter insertion | -504
    chemotherapy with pre-phase treatment | -504
    rituximab | -504
    prednisolone | -504
    R-mini-CHOP | -504
    chemotherapy continuation | -504
    R-CHOP | -504
    complete remission | 720
    no remaining cardiac mass | 720
    no extracardiac disease | 720
    no AV conduction disorder | 720
    18F-FDG-PET/CT | 720
    PM-control | 720
    last echocardiography | 720
    axial diaphragma hernia | -36000
    sigma diverticulosis | -36000
    no cardiologic medical history | -36000
    