63 years old | 0
male | 0
farm worker | 0
admitted to the hospital | 0
complaining of weakness | 0
complaining of headache | 0
complaining of fever | 0
working in a farm | -168
developed generalized myalgia | -168
developed malaise | -168
developed vomiting | -168
denied any contact with animals | 0
positive surgical history | 0
no history of consumption of dairy products | 0
no recent travel to endemic areas | 0
alert and oriented | 0
pyrexial | 0
conjunctival suffusion | 0
no scleral jaundice | 0
skin normal | 0
heart normal | 0
lung normal | 0
bladder not felt | 0
liver not felt | 0
rectal examination normal | 0
neurological examination normal | 0
kerning sign negative | 0
brudzinski sign negative | 0
headache increased | 48
hiccup | 120
photophobia | 120
diplopic vision | 120
ptosis | 120
right side preorbital edema | 120
deviation of the right eye to the medial site | 144
brainstem involvement | 144
ataxic | 144
dysarthric | 144
uvula deviated to the left site | 144
lack of gag reflex | 144
right side facial paresis | 144
decreased consciousness | 168
hemoptysis | 168
gastrointestinal bleeding | 168
abdominal sonography normal | 168
serum sample sent for laboratory evaluation | 168
L. Serjoe hardjo equal to 1/1600 | 168
neurological consultation | 168
magnetic resonance imaging/magnetic resonance venography prescribed | 168
cavernous sinus thrombosis syndrome | 168
axial computed tomography scan | 168
increased intensity with conversity in right cavernous sinus | 168
loss of flow in both sides of cavernous sinus | 168
right cavernous sinus expansion | 168
longitudinal filling defect | 168
parietal irregularities with superior sagittal sinus | 168
transverse, sigmoid, and internal jugular vein normal | 168