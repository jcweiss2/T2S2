66 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
intermittent high-grade fever | -216 | 0 | Factual
generalized dull-aching abdominal pain | -216 | 0 | Factual
passing turbid urine | -240 | 0 | Factual
decrease in urine output | -240 | 0 | Factual
swelling of both feet | -240 | 0 | Factual
treated with intravenous medications | -168 | -168 | Factual
type II diabetes mellitus | -2628 | 0 | Factual
regular medication for diabetes | -2628 | 0 | Factual
conscious | 0 | 0 | Factual
afebrile | 0 | 0 | Factual
tachycardic | 0 | 0 | Factual
heart rate of 136/min | 0 | 0 | Factual
blood pressure was 110/70 mmHg | 0 | 0 | Factual
renal angle tenderness bilaterally | 0 | 0 | Factual
high total leukocyte counts | 0 | 0 | Factual
left shift | 0 | 0 | Factual
elevated urea and creatinine levels | 0 | 0 | Factual
pyuria | 0 | 0 | Factual
leukocyte esterase positivity | 0 | 0 | Factual
possibility of pyelonephritis/renal abscess | 0 | 0 | Possible
possibility of acute kidney injury | 0 | 0 | Possible
activated partial thromboplastin time was prolonged | 0 | 0 | Factual
sepsis-induced coagulopathy | 0 | 0 | Possible
enlarged kidneys | 0 | 0 | Factual
bilateral renal abscesses | 0 | 0 | Factual
emergency ultrasound-guided drainage of renal abscesses | 24 | 24 | Factual
transfusion of blood products | 24 | 24 | Factual
coagulopathy | 0 | 24 | Factual
pus smear from renal abscesses showed septate fungal hyphae | 24 | 24 | Factual
intravenous meropenem | 0 | 24 | Factual
intravenous voriconazole | 24 | 24 | Possible
intravenous amphotericin B | 48 | 216 | Factual
cultures from both renal abscesses revealed growth of Aspergillus fumigatus | 48 | 48 | Factual
worsening renal function | 72 | 216 | Factual
acute pulmonary edema | 120 | 120 | Factual
hyperkalemia | 120 | 216 | Factual
metabolic acidosis | 120 | 216 | Factual
hemodialysis | 120 | 216 | Factual
noninvasive ventilation | 120 | 216 | Factual
sudden cardiac arrest | 216 | 216 | Factual
aspiration | 216 | 216 | Possible
death | 216 | 216 | Factual