37 years old | -672
male | -672
rheumatic mitral stenosis | -672
mild aortic insufficiency | -672
pulmonary hypertension | -672
referred to surgical treatment | -672
heart failure | -240
signs of endocarditis | -240
sepsis | -240
excessive organ failure | -240
urgent surgery | -240
mechanical mitral valve implantation | -240
minor commissurotomy of the aortic valve cusps | -240
double valve re-endocarditis | -48
prosthetic mitral valve endocarditis | -48
native aortic valve endocarditis | -48
aortic root abscess | -48
biological mitral valve implantation | 0
full root implantation of Medtronic Freestyle bioprosthesis | 0
reimplantation of the coronary ostia | 0
atrial fibrillation | 0
diabetes mellitus type 2 | 0
warfarin prescription | 0
enalapril prescription | 0
metformin prescription | 0
metoprolol prescription | 0
follow-up transoesophageal echocardiography | 41
well-functioning FB valve | 41
non-ST-elevation myocardial infarction | 1920
chest oppression | 1920
pain in the left arm and hand | 1920
shortness of breath | 1920
discrete heart murmur | 1920
irregular rhythm | 1920
normal vesicular breath sounds | 1920
no oedema | 1920
atrial fibrillation | 1920
ST depressions | 1920
T-wave inversions | 1920
ST elevation | 1920
increasing troponin T concentration | 1920
contrast-enhanced cardiac computed tomography | 1920
significant left- and right coronary ostial stenosis | 1920
no sign of atherosclerosis | 1920
preoperative coronary angiography | 1920
90% stenosis in both ostia | 1920
normal coronary arteries | 1920
emergent reoperation | 1920
coronary artery bypass grafting | 1920
pseudointimal glass-like membranes | 1920
intraoperative findings | 1920
acetylsalicylic acid prescription | 1920
metoprolol reduction | 1920
histological examination | 1920
fibro-intimal thickening | 1920
inflamed granulation tissue | 1920
no sign of acute inflammation | 1920
no calcifications | 1920
no foreign bodies | 1920
no amyloidosis | 1920
follow-up cardiac CT | 1920
follow-up transthoracic echocardiography | 1920
small pseudoaneurysm | 1920
partial rupture of the distal anastomosis | 1920
conservative strategy | 1920
repeat follow-up cardiac CT | 1980
reduction of the pseudoaneurysm | 1980
exercise-induced chest pains | 2160
myocardial perfusion scintigraphy | 2160
exercise-induced myocardial ischaemia | 2160
coronary angiography | 2160
complete revascularization | 2160
mild-moderate stenosis of the FB valve | 2160
well-functioning biological mitral valve | 2160