65 years old | 0
female | 0
diabetes mellitus | 0
systemic arterial hypertension | 0
transesophageal echocardiography | 0
suspected diagnosis of atrial septal defect | 0
topical anesthesia | 0
difficulties in progression of the probe into the esophagus | 0
retching | 0
inability to collaborate with the exam performance | 0
neck pain | 0
oropharyngeal pain | 0
dysphagia | 4
edema | 24
hyperemia | 24
local pain | 24
systemic symptoms | 24
weakness | 24
malaise | 24
admitted to the hospital | 72
blood pressure 150/100 mmHg | 72
pulse rate 100 beats per minute | 72
subcutaneous emphysema | 72
intense hyperemia | 72
computed tomography scan | 72
fistula of the posterior esophageal wall | 72
upper gastrointestinal endoscopy | 72
marked vascular congestion | 72
edema of the hypopharynx | 72
pyriform sinuses | 72
upper esophageal sphincter | 72
esophageal wall perforation | 72
purulent secretion | 72
ceftriaxone | 72
clindamycin | 72
cervicotomy | 72
drainage of pus | 72
septic shock | 72
norepinephrine | 72
mechanical ventilatory support | 72
esophageal fistula | 168
improved clinical status | 168