64 years old | 0
woman | 0
admitted to intensive care unit | 0
confusion | 0
fever | 0
temperature of 38.8°C | 0
blood pressure 105/73 mmHg | 0
heart rate 129 bpm | 0
significant agitated behavior | 0
abdominal sensitivity | 0
WBC 14,000/mm3 | 0
elevated CRP 160.6 mg/l | 0
creatinine 126 μmol/l | 0
all blood cultures negative | 0
HIV negative | 0
HCV negative | 0
HBV negative | 0
syphilis negative | 0
MRI head | 0
cerebellar lesion 28 mm | 0
frontal right lesion 15 mm | 0
parietal lesion 17 mm | 0
occipital lesion 15 mm | 0
lumbar puncture | 0
WBC 275/mm3 | 0
PNN 4% | 0
lymphocytes 89% | 0
no germ retrieved | 0
total body scan imaging | 0
liver abscess 11 cm | 0
right-sided pleural effusion | 0
thoracentesis cultures negative | 0
liver drain cultures negative | 0
intravenous Ceftriaxone | 0
oral Metronidazole | 0
clinical improvement | 0
biological improvement | 0
afebrile | 120
neurological symptoms resolved | 120
transferred to infectious diseases unit | 120
cerebral MRI at 3 weeks | 504
no major difference in brain abscess size | 504
ultrasound | 504
stagnation in liver abscess size | 504
craniotomy recommended | 504
brain biopsy | 504
mixed inflammatory reaction | 504
macrophagic infiltrate | 504
granulomas | 504
no evident pathogenic microorganism | 504
aerobic cultures negative | 504
anaerobic cultures negative | 504
PCR positive for Fusobacterium nucleatum | 504
Ceftriaxone changed to Clindamycine | 504
Metronidazole continued | 504
FDG-PET | 504
no other infection sites | 504
MRI brain at 12 weeks | 2016
cerebellar lesion decreased to 8 mm | 2016
frontal right lesion decreased to 6.5 mm | 2016
parietal lesion decreased to 6.5 mm | 2016
occipital lesion decreased to 6.5 mm | 2016
decrease in ring enhancing intensity | 2016
decrease in surrounding edema | 2016
oral Metronidazole continued | 2016
total treatment duration 20 weeks | 3360
brain imaging at 6 months | 4320
hepatic imaging at 6 months | 4320
pulmonary imaging at 6 months | 4320
brain images stable | 4320
hepatic abscesses complete recovery | 4320
pleural effusion complete recovery | 4320
good clinical recovery | 4320
neuro cognitive function improved | 4320
CRP 3.7 mg/l | 4320
no fever | 4320
intra-uterine device present | -?
intra-uterine device removed | ?
device culture negative | ?
FDG-PET no malignancies | 504
PCR performed | 504
16S ribosomal RNA sequencing | 504
intra2-uterine device removed | ?
blood pressure 105/73 mmHg |/tmp/verse_20240610_235952_9g4d5g/out.txt 0
