21 years old | 0
male | 0
MNGIE | -1320
energy loss | -1320
foot-drop | -1320
difficulty swallowing | -1320
weight loss | -1320
duodenojejunostomy operation | -720
SMA syndrome | -720
TPN | -720
central venous catheterization | -720
catheter changed | -720
catheter changed | -624
catheter changed | -528
catheter changed | -432
catheter inserted | -24
fever | -24
palpitation | -24
body temperature 38.5° | -24
blood pressure 120/77 mmHg | -24
pulse 157 beats/min | -24
elevated sedimentation | -24
elevated CRP | -24
MRSA in blood cultures | -24
catheter-related infection | -24
echocardiography | -24
mobile thrombus | -24
heparin treatment | -18
antibiotic treatment | -18
prothrombin time 12.9 second | -18
INR 1.1 | -18
platelet count 380.000/mm3 | -18
open heart surgery | 0
ECG monitoring | 0
SpO2 monitoring | 0
invasive arterial catheterization | 0
systemic arterial pressure 120/80 mmHg | 0
heart rate 130/min | 0
SpO2 97% | 0
midazolam | 0
thiopental | 0
fentanyl | 0
rocuronium | 0
intubation | 0
central venous catheterization | 0
extracorporeal circulation | 0
thrombus removal | 0
hemoglobin 10.9 g/dl | 0
hemoglobin 7.1 g/dl | 0
blood transfusion | 0
RBC transfusion | 0
FFP transfusion | 0
extubation | 5
transport to Cardiovascular Surgery Department | 72
catheter culture sterile | 72
pathology report infected thrombus | 72
discharged | 120
recommendation for enteral nutrition | 120
recommendation for supportive peripheral nutrition | 120