46 years old | 0
male | 0
sickle cell disease | 0
admitted to the hospital | 0
abdominal pain | -24
acute cholecystitis | -24
laparoscopic cholecystectomy (LC) | -24
discharged home | -24
worsening abdominal pain | 24
abnormal liver function studies | 24
imaging suggesting common bile duct transection | 24
attempted endoscopic retrograde cholangiopancreatogram (ERCP) | 24
aborted ERCP | 24
transferred to neighboring hospital | 24
severe respiratory distress | 48
sickle cell crisis | 48
sinus tachycardia | 48
heart rate 156 | 48
blood pressure 173/87 | 48
pulse oximetry 92% | 48
high flow nasal cannula at 30 l/min | 48
transferred to intensive care unit | 48
total bilirubin 15.1 mg/dl | 48
creatinine 1.1 mg/dl | 48
AST 150 U/l | 48
ALT 434 U/l | 48
alkaline phosphatase 175 U/l | 48
white blood cells 15.3 × 10^3/cm2 | 48
hematocrit 26% | 48
hemoglobin 9.1 g/dl | 48
platelets 216 × 10^3/cm2 | 48
INR 1.5 | 48
CT angiogram of abdomen significant for multifocal pneumonia | 48
free peritoneal fluid | 48
chest CT negative for pulmonary embolism | 48
repeat ERCP confirmed wide-open distal common bile duct | 72
inability to pass a wire distally | 72
percutaneous transhepatic cholangiography (PTC) | 72
PTC study confirmed completely transected duct | 96
wire traversed ductal injury into distal ductal orifice | 96
entry into duodenum | 96
open surgical repair | 96
over 2 l of bilious fluid consistent with bile peritonitis | 96
portal dissection performed | 96
exposed PTC catheter exiting proximal hepatic hilum | 96
entered distal common bile duct | 96
remainder of common bile duct necrosed or resected | 96
multiple surgical clips removed | 96
identified cystic artery | 96
preserved right and left hepatic arteries | 96
PTC catheter pulled from distal common bile duct | 96
orifice closed using 3-0 prolene sutures | 96
retrocolic Roux-en-Y hepaticojejunostomy performed | 96
interrupted 5-0 PDS sutures | 96
PTC catheter placed into roux limb | 96
drain placed under repair | 96
abdomen closed | 96
transferred back to ICU | 96
PTC catheter placed to gravity drainage | 96
extubated | 168
episodes of oxygen desaturations | 168
hemoglobin electrophoresis significant for elevated HgbS and C | 168
red blood cell exchange transfusion performed | 168
goal hemoglobin S and C combined percentage <30% | 168
discharged home | 240
total bilirubin 4.1 mg/dl | 240
normal transaminases | 240
stable hematocrit 30% | 240
normal renal function | 240
seen in clinic 4 weeks post-op | 672
total bilirubin 1.0 mg/dl | 672
cholangiogram showing no evidence of leak or stricture | 672
cholangiogram catheter removed | 672
discharged from clinic | 672
