15 years old | 0
    male | 0
    admitted to the general ward | 0
    vomiting | -24
    lethargy | -24
    left thigh swelling | -336
    fell from bed | -336
    left femur shaft fracture | -336
    underwent orthopedic surgery | -288
    discharged seven days after surgery | -240
    poor oral intake | -48
    refused solid foods | -48
    only took liquids | -48
    body temperature elevated to 38.0°C | -48
    bilious vomiting | -24
    became lethargic | -24
    decreased urine output | -24
    dark urine appearance | -24
    dehydration | 0
    admitted for supportive care and evaluation | 0
    cerebral palsy | 0
    HSAN-IV | 0
    recurrent orthopedic diseases (femur fractures, septic arthritis, osteomyelitis) | 0
    mutilated fingertips | 0
    recurrent cellulitis | 0
    septic arthritis of fingers | 0
    recurrent trauma due to impulse control disorder | 0
    unstable body temperature | 0
    unstable blood pressures | 0
    autonomic dysregulation | 0
    severe dry skin | 0
    hyperkeratosis | 0
    fissuring | 0
    xerotic eczema | 0
    wheelchair-bound | 0
    mentally retarded | 0
    hypokalemia | 0
    hypomagnesemia | 0
    Gitelman syndrome | 0
    taking anti-psychotics | 0
    taking psychostimulants | 0
    taking spironolactone | 0
    alert | 0
    cachectic | 0
    wearing hip spica cast | 0
    height <3rd percentile | 0
    weight <3rd percentile | 0
    blood pressure 130/88 mmHg | 0
    pulse rate 97 beats/minute | 0
    respiratory rate 21 times/minute | 0
    body temperature 37.3°C | 0
    no anemia | 0
    no icteric sclera | 0
    slightly dehydrated lips and mucous membranes | 0
    intact tympanic membranes | 0
    no palpable cervical lymph nodes | 0
    symmetrical chest expansion | 0
    clear breath sounds | 0
    regular heartbeat without murmur | 0
    soft and flat abdomen | 0
    no abdominal tenderness | 0
    no rebound tenderness | 0
    hyperactive bowel sounds | 0
    no shifting dullness | 0
    non-palpable liver or spleen | 0
    no peripheral edema | 0
    no digital clubbing | 0
    no cyanosis | 0
    dry skin | 0
    no rash | 0
    no petechia | 0
    sodium 138 mmol/L | 0
    potassium 3.2 mmol/L | 0
    AST 23 IU/L | 0
    ALT 12 IU/L | 0
    total bilirubin 1.0 mg/dL | 0
    BUN 29 mg/dL | 0
    creatinine 0.41 mg/dL | 0
    CRP <0.03 mg/dL | 0
    serum magnesium 1.6 mg/dL | 0
    supportive treatment initiated | 0
    high fever 41.8°C | 72
    blood pressure dropped to 50/17 mmHg | 72
    seizure-like movements (upward eyeball deviation, loss of consciousness, clonic movement) | 72
    fixed pupils 2 mm diameter | 72
    WBC 19.4×10³/µL | 72
    hemoglobin 9.6 g/dL | 72
    platelets 90×10³/µL | 72
    sodium 137 mmol/L | 72
    potassium 2.6 mmol/L | 72
    AST 454 IU/L | 72
    ALT 258 IU/L | 72
    total bilirubin 4.3 mg/dL | 72
    direct bilirubin 2.6 mg/dL | 72
    amylase 228 IU/L | 72
    lipase 888 IU/L | 72
    creatinine phosphate kinase 1258 IU/L | 72
    lactate dehydrogenase 985 IU/L | 72
    BUN 49 mg/dL | 72
    creatinine 1.62 mg/dL | 72
    CRP 0.6 mg/dL | 72
    plasma hemoglobin 27.5 mg/dL | 72
    serum ferritin 250 ng/mL | 72
    weakly positive antinuclear antibody (1:40) | 72
    AST 492 IU/L | 72
    ALT 545 IU/L | 72
    total bilirubin 10.8 mg/dL | 72
    direct bilirubin 5.1 mg/dL | 72
    amylase 520 IU/L | 72
    lipase 5071 IU/L | 72
    PT INR 3.1 | 72
    aPTT 52.7 seconds | 72
    fibrinogen 160 mg/dL | 72
    D-dimer 17.62 µg/mL | 72
    alkaline phosphatase 126 IU/L | 72
    γ-glutamyltranspeptidase 98 IU/L | 72
    fluid resuscitation | 72
    intravenous inotropes (dopamine, norepinephrine) | 72
    antibiotics | 72
    gabexatemesilate | 72
    transferred to PICU | 72
    ventilator care | 72
    seizure-like movements | 72
    lorazepam injection | 72
    mannitol initiated | 72
    abdominal CT negative for acute pancreatitis | 72
    multiple kidney filling defects | 72
    hypoxic ischemic encephalopathy | 72
    low serum ceruloplasmin 5.5 mg/dL | 72
    increased 24-hour urine copper 1028 µg/dL | 72
    liver biopsy with copper deposition | 72
    centrilobular confluent necrosis | 72
    liver copper deposit 74 µg/g | 72
    no Kayser-Fleischer rings | 72
    NTRK1 gene mutations (c.2002G>T, c.360-1G>A) | 72
    SLC12A3 gene mutation (c.1216A>C) | 72
    ATP7B gene negative | 72
    trientine started 25 mg/kg/day | 72
    low copper diet | 72
    WBC 8.66×10³/µL | 360
    hemoglobin 12.9 g/dL | 360
    platelets 364×10³/µL | 360
    sodium 137 mmol/L | 360
    potassium 4.0 mmol/L | 360
    AST 128 IU/L | 360
    ALT 127 IU/L | 360
    total bilirubin 1.3 mg/dL | 360
    BUN 25 mg/dL | 360
    creatinine 0.1 mg/dL | 360
    PT INR 1.15 | 360
    aPTT 52.3 seconds | 360
    tracheostomy | 360
    percutaneous endoscopic gastrostomy | 360
    trientine continued | 360
    copper restriction diet | 360
    discharged | 360
    <|eot_id|>
    