66 years old | 0
    female | 0
    admitted to the hospital | 0
    cough | 0
    tachypnoea | 0
    chills | 0
    weakness | 0
    reduced oxygen saturation | 0
    diabetes mellitus | -infinity
    hypertension | -infinity
    dyslipidemia | -infinity
    hypothyroidism | -infinity
    hypoxic respiratory failure | 0
    intubated | 0
    ventilated | 0
    septic shock | 0
    acute kidney injury | 0
    haemodialysis | 0
    high white blood cell count (14.5 K/dl) | 0
    low platelets (145 K) | 0
    high activated partial thromboplastin time (64.4 seconds) | 0
    normal international normalized ratio (1) | 0
    normal prothrombin time (11.2 seconds) | 0
    high fibrinogen (5 g/l) | 0
    high D-dimer (2.6 mg/l) | 0
    high C-reactive protein (67.8 mg/l) | 0
    high creatinine (217 μmol/L) | 0
    high alanine aminotransferase (60 U/l) | 0
    high aspartate aminotransferase (40 U/l) | 0
    high alkaline phosphatase (175 U/l) | 0
    recent travel history | -infinity
    tested positive for COVID-19 | 0
    CT scan of the head | 504
    feverish | 504
    drop in level of consciousness | 504
    left parietal centrum semiovale vasogenic oedema | 504
    MRI head | 504
    intracranial magnetic resonance angiography | 504
    microbleeds predominantly involving juxtacortical white matter | 504
    larger bleeding foci in left parietal region | 504
    perilesional oedema | 504
    tiny foci of microbleeds in internal capsules | 504
    critical illness-associated cerebral microbleeds | 504
    vasogenic oedema in left parietal region | 504
    discharged | 504