31 years old | 0
male | 0
admitted to the hospital | 0
bilateral joint pains | -24
bilateral joint swelling | -24
ankle joint pain | -24
wrist joint pain | -24
coryzal symptoms | -24
sore throat | -24
fever | -24
polyarthralgia | -24
no symptoms suggestive of meningism | -24
no headache | -24
no photophobia | -24
no neck stiffness | -24
born in the U.K. | 0
received the U.K. childhood vaccination scheme | 0
full-time bus driver | 0
heterosexual relationship for the last 16 years | 0
no significant medical or family history | 0
no foreign travel | 0
alert and orientated in time, place and person | 0
temperature 36.9 °C | 0
heart rate 101 bpm | 0
blood pressure 125/85 mmHg | 0
respiratory rate 16 breaths per minute | 0
oxygen saturations 99 % in room air | 0
qSOFA score of zero | 0
bilateral swelling and pain in the small joints of the hands and wrist joints | 0
reduced range of movement | 0
mild purpuric rash | 0
no cardiac murmurs | 0
metabolic acidosis | 0
raised lactate of 9.29 mmol/L | 0
cryptic shock | 0
hyperlactataemia | 0
cellular and metabolic stress | 0
normal radiographs of the chest, abdomen, wrist, knee, and ankle joints | 0
significant inflammatory response | 0
C reactive protein 223 mg/L | 0
erythrocyte sedimentation rate 45 mm/h | 0
white cell count 4.9 × 109/L | 0
coagulopathy | 0
international normalised ratio 2 | 0
prothrombin time 24.9 s | 0
D-dimer 42,011 ng/mL | 0
mild liver dysfunction | 0
alanine aminotransferase 58 U/L | 0
alkaline phosphatase 81 U/L | 0
haematuria | 0
proteinuria | 0
negative leucocytes and nitrites | 0
provisional diagnosis of ‘sepsis of unknown source with associated DIC’ | 0
blood cultures taken | 0
commencement of broad-spectrum intravenous antibiotics | 0
piperacillin/tazobactam | 0
intravenous fluids | 0
intravenous vitamin K | 0
ankle joints aspirated | 0
joint fluid negative for organisms and crystals | 0
further blood tests sent | 0
anti-neutrophil cytoplasmic antibodies | 0
anti-nuclear antibodies | 0
anti-Streptolysin O titre | 0
rheumatoid factor | 0
lupus anticoagulant | 0
Human Immunodeficiency Virus test | 0
hepatitis B test | 0
hepatitis C test | 0
mildly raised rheumatoid factor | 0
lupus anticoagulant | 0
urine total protein: creatinine ratio markedly raised | 0
blood cultures grew gram-negative diplococcus | 48
N. meningitidis group W135 | 48
sensitive to penicillin | 48
antibiotic regime tailored to the identified pathogen | 48
benzylpenicillin | 48
Public Health England informed | 48
household contacts given prophylactic ciprofloxacin | 48
fever persisted | 216
inflammatory markers continued to rise | 216
CRP 354 mg/L | 216
extensive ecchymosis | 216
purpuric macules | 216
large bullous lesions | 216
soft tissue induration | 216
cutaneous lesions | 216
purpura fulminans | 216
vasculitic element | 216
CT scan of the chest, abdomen and pelvis | 216
transthoracic echocardiogram | 216
no secondary foci of infection | 216
magnetic resonance imaging scan of all four limbs | 240
necrotising fasciitis excluded | 240
failure to defervesce | 240
new skin lesions | 240
post-infectious, immune-driven complications | 240
immune-complex hypersensitivity reactions | 240
type three immune reactions | 240
antibody and antigen complex | 240
inflammation and activation of the complement pathway | 240
leukocytes recruitment | 240
tissue damage | 240
skin necrosis | 240
ibuprofen 400 mg three times per day | 240
pulsed intravenous methylprednisolone | 240
fever lysis | 264
clinical and biochemical improvement | 264
antibiotics stopped | 336
convalescence complicated by recrudescence of fever | 360
re-introduction of intravenous antibiotics | 360
Meropenem 1 g three times per day | 360
oral steroids | 360
prednisolone 40 mg once daily | 360
cutaneous lesions regressed | 360
tissue loss persisted | 360
CT angiogram | 360
macrovascular ischaemia excluded | 360
MRI scan of the right foot | 360
extensive, deep-seated soft tissue collection | 360
inflammatory aetiology | 360
soft tissue fat necrosis | 360
skin grafting attempted | 360
surgical debridement | 360
flap cover unsuccessful | 360
right above-knee amputation | 360