23 years old|0
    man|0
    presented to the emergency department with abdominal pain, nausea, vomiting, and diarrhea|0
    abdominal pain|0
    nausea|0
    vomiting|0
    diarrhea|0
    developed pulseless electrical activity cardiac arrest|0
    started on peripheral venoarterial (VA) extracorporeal membranous oxygenation (ECMO)|0
    healthy individual without a past medical history|0
    septic shock|-1
    hypovolemic shock|-1
    pulseless electrical activity arrest|0
    cardiovascular failure|0
    transthoracic echocardiogram (TTE) performed|0
    near cardiac standstill|0
    moderate posterior pericardial effusion|0
    systolic blood pressure was 30 mm Hg|0
    ECMO flow was low|0
    checked bridge circuit for thrombus|0
    no change in ECMO flow|0
    decision to augment venous drainage|0
    right internal jugular venous cannula inserted|0
    venovenous (VV)-arterial ECMO started|0
    blood pressure improved|0
    increased venous drainage|0
    better ECMO flow|0
    remained hemodynamically unstable|0
    pericardial effusion enlarged|0
    emergent pericardiotomy performed|0
    400 ml of clear fluid removed|0
    severe myocardial edema|0
    near cardiac standstill noted|0
    left ventricle (LV) nonpulsatile|0
    competing with retrograde ECMO flow|0
    severe LV dilation|0
    pulmonary edema|0
    taken to cardiac catheterization lab for Impella CP heart pump placement|0
    aortic pressure was 72/64 mm Hg|0
    LV end-diastolic pressure was 25 mm Hg|0
    LV cavity size decreased|0
    improved unloading from Impella CP|0
    lower extremities became tense|0
    creatinine kinase level rose to >100,000 U/l|0
    severe fulminant skeletal myositis|0
    H3N2 viremia|0
    rhabdomyolysis|0
    required bilateral leg fasciotomies|0
    removal of Impella device|0
    treated empirically with oseltamivir|0
    treated with broad-spectrum antibiotics|0
    respiratory swab resulted positive for influenza A (H3N2)|0
    blood cultures grew Streptococcus viridans|0
    shock precipitated by fulminant myocarditis from influenza A infection|0
    intravenous immunoglobulin added|0
    ECMO flow requirement decreased|24
    cardiac contractility increased|24
    TTE on hospital day 12|288
    estimated LV ejection fraction of 30% to 35%|288
    improvement in cardiac contractility|288
    lungs remained severely damaged|288
    developed differential upper extremity hypoxemia|288
    concerns for North-South syndrome|288
    ECMO circuit rearranged to VA-venous configuration|288
    oxygenated blood returned to upper and lower body|288
    oxygenation improved|288
    significant facial swelling due to right internal jugular cannula|288
    superior vena cava syndrome|288
    cannula removed|288
    facial swelling resolved|288
    ECMO configuration switched to VA through left femoral artery and vein|288
    hemodynamic improvement|288
    vasopressor requirements decreased|288
    ECMO circuit decannulated on hospital day 18|432
    fought multiple infections over next 6 months|432
    extensive wound debridement of lower extremities|432
    tracheostomy placed|432
    tracheostomy decannulated before discharge|432
    weaned off hemodialysis|432
    TTE before discharge showed LV ejection fraction of 55%|432
    fulminant myocarditis from influenza A (H3N2) infection|0
    complexity of mechanical circulatory support management with ECMO|0