35 years old | 0
male | 0
no significant chronic degenerative history | 0
surgical history of autograft | 0
left upper limb | 0
left lateral region of the neck | 0
left lateral aspect of the thorax | 0
secondary to a third-degree burn | 0
radius and ulna fracture | 0
treated with a splint | 0
without sequelae | 0
family history of hypertension | 0
type 2 diabetes mellitus | 0
unspecified gastric carcinoma | 0
maternal branch | 0
intermittent crampy abdominal pain | -168
predominantly in the hypogastrium | -168
progressed to diffuse abdominal pain | -168
weight loss | -168
approximately 10.5 kg | -168
in 3 months | -168
stools decreased in consistency | -168
abdominal ultrasound | -30
multiple heterogeneous liver lesions | -30
splenomegaly | -30
carcinoembryonic antigen | -30
197.31 ng/mL | -30
CA 19-9 antigen | -30
10,386 ng/mL | -30
computerized axial tomography | -30
metastatic lesions in the liver | -30
thickening of the hepatic angle of the colon | -30
tumor of the descending colon | -30
outpatient colonoscopy | -30
abdominal pain | 0
unquantified fever | 0
unstable vital signs | 0
tendency to hypotension | 0
tachycardia | 0
respiratory distress | 0
cardiopulmonary without apparent compromise | 0
abdominal distension | 0
generalized pain | 0
involuntary muscular resistance | 0
positive rebound | 0
bowel sounds of metallic hue | 0
leukocytes | 0
15.10 × 10e3/μL | 0
neutrophils | 0
14.6 × 10e3/μL | 0
hemoglobin | 0
6.7 g/dL | 0
platelets | 0
623.00 × 10e3/μL | 0
glucose | 0
108 mg/dL | 0
urea | 0
95.3 mg/dL | 0
creatinine | 0
2.26 mg/dL | 0
uric acid | 0
11.3 mg/dL | 0
total cholesterol | 0
67 mg/dL | 0
triglycerides | 0
135 mg/dL | 0
direct bilirubin | 0
1.27 mg/dL | 0
indirect bilirubin | 0
0.58 mg/dL | 0
aspartate aminotransferase | 0
1442 U/L | 0
alanine aminotransferase | 0
714 U/L | 0
albumin | 0
2.49 g/dL | 0
total proteins | 0
5 g/dL | 0
lactic dehydrogenase | 0
1592 U/L | 0
sodium | 0
123 mEq/L | 0
chlorine | 0
84 mEq/L | 0
potassium | 0
5.7 mEq/L | 0
calcium | 0
7.83 mg/dL | 0
magnesium | 0
2.8 mg/dL | 0
phosphorus | 0
7.2 mg/dL | 0
prothrombin | 0
20.6 s | 0
INR | 0
1.9 | 0
activated partial thromboplastin | 0
40.9 s | 0
fibrinogen | 0
628 mg/dL | 0
procalcitonin | 0
43.5 ng/dL | 0
pH | 0
7.3 | 0
pCO2 | 0
22.8 mm Hg | 0
pO2 | 0
17.9 mm Hg | 0
HCO3 | 0
11.1 mmol/L | 0
BE | 0
15.2 mmol/L | 0
lactate | 0
15.92 mmol/L | 0
abdominal X-ray | 0
dilation of intestinal loops | 0
up to 12 cm | 0
inter-loop edema | 0
chest radiograph | 0
subdiaphragmatic free air | 0
emergency exploratory laparotomy | 0
perforation in a tumor of the left colon | 0
splenic angle | 0
tumor measuring approximately 12 × 10 × 8cm | 0
proximal third of the ascending colon | 0
locally advanced to the para-aortic ganglionic chain | 0
evidence of necrosis | 0
free intestinal fluid | 0
approximately 600 mL | 0
multiple firms and lax loop-loop adhesions | 0
multiple liver metastases | 0
abscesses | 0
radical total colectomy | 0
resection at the level of the R2 ileocolic artery | 0
formation of a Brooke-type terminal ileostomy | 0
duration of the surgical procedure | 0
1 h 16 min | 0
anesthetic time | 0
2 h | 0
total bleeding | 0
estimated at 500 mL | 0
transferred to the intensive care unit | 0
hemodynamic instability | 0
septic shock | 0
multiple organ failure | 0
adequate ileostomy functioning | 12
after 12 h after surgery | 12
refractory septic shock | 48
cardiorespiratory arrest | 48
without response to advanced maneuvers | 48
death | 48
malignant neoplastic lesion | 0
epithelial lineage | 0
glandular and in loose nests pattern | 0
replaces the mucosa | 0
infiltrates the lamina propria | 0
muscularis mucosas | 0
submucosa | 0
muscularis propria | 0
subserosa | 0
loss of continuity | 0
perforation | 0
neoplastic cells | 0
hyperplasia | 0
mesothelial inflammation | 0
intestinal phenotype glands | 0
pseudostratified simple columnar epithelium | 0
nucleus: cytoplasm ratio | 0
2-3:1 | 0
clear cytoplasm | 0
round nuclei | 0
moderate atypia | 0
membrane reinforcement nuclear | 0
salt and pepper chromatin | 0
evident nucleolus | 0
few mitosis | 0
fibrovascular tissue | 0
segmented mononuclear inflammatory infiltrate | 0
stage IVc | 0
T4c | 0
N2b | 0
M1c | 0
TNM classification | 0
American Joint Committee on Cancer | 0
eighth edition | 0
2017 | 0