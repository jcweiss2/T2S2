9 years old | 0
male | 0
spina bifida | 0
hydrocephalus | 0
imperforate anus | 0
scoliosis | 0
solitary kidney | 0
multiple urinary tract infections | 0
abdominal pain | -12
nonbilious vomiting | -12
no fever | -12
normal stool output via colostomy | -12
ventriculoperitoneal shunt | -672
colostomy | -672
titanium rib placement | -672
Monti procedure | -210
catheterization schedule every 3 hours | -210
little blood with catheterization | -210
intermittent difficulty catheterizing | -168
mild difficulty inserting catheter | -168
good output | -168
heart rate of 166 beats/min | 0
blood pressure of 132/90 | 0
respiratory rate of 25 breaths/min | 0
temperature of 99.6 | 0
oxygen saturation of 98% | 0
alert and talkative | 0
comfortable in sitting position | 0
pain when placed supine | 0
abdominal distension | 0
white blood cell count of 32.1 × 10^3/mm^3 | 0
77% neutrophils | 0
14% bands | 0
serum bicarbonate of 12 mEq/L | 0
blood urea nitrogen of 24 mg/dL | 0
cloudy, blood-tinged fluid | 0
malodorous urine | 0
50-100 red blood cells per high power field | 0
50-100 white blood cells per high power field | 0
nitrite negative | 0
leukocyte esterase 3+ | 0
CT scan of abdomen and pelvis | 0
ascitic fluid | 0
worsening hydronephrosis | 0
CT cystogram | 0
urine extravasation | 0
perforation of continent ileovesicostomy | 0
neurosurgery and urology consulted | 0
CT scan of brain | 0
cerebrospinal fluid clear | 0
mild increase in ventricular size | 0
fracture in shunt tubing | 0
externalization of proximal shunt | 0
removal of indwelling shunt | 0
urology consulted | 0
bladder neck reconstruction | -840
right ureteral implant | -840
construction of Monti channel vesicostomy | -840
fluid bolus | 0
cefepime | 0
admitted to PICU | 0
worsening tachycardia | 12
diminished pulses | 12
compensated septic shock | 12
vancomycin | 12
additional fluid bolus | 12
surgery | 24
proximal shunt externalized | 24
distal catheter removed | 24
purulent material aspirated | 24
endoscopy of catheterizable stoma | 24
large posterior false passage | 24
catheter placed across stoma | 24
cystoscopy | 24
cystogram | 24
no bladder perforation | 24
Foley catheter placed | 24
mechanical ventilation | 24
low-dose norepinephrine | 24
urine culture grew Escherichia coli | 48
shunt and peritoneal fluid cultures negative | 48
removal of retained fractured piece of shunt catheter | 144
peritoneal catheter removed | 144
original shunt converted to ventriculocardiac shunt | 264
discharged | 336
intravenous antibiotics | 336
urethral and vesicostomy catheters to gravity drainage | 336
Monti catheter left in place | 336
cystoscopy for perceived difficulty in catheterization | 672
no stenosis or false passage | 672
catheterization difficulty and urinary retention | 840
cystoscopy revealed false passage | 840
Monti revision for stenosis | 1008