56 years old | 0
male | 0
obese | 0
smoker | 0
occasional alcohol drinker | 0
admitted to the Intensive Care Unit | 0
community-acquired bacterial meningitis | 0
neurological emergency |3
early diagnosis |3
targeted treatment |3
Streptococcus suis infection |0
zoonotic origin bacterial meningitis |0
auditory complications |0
labyrinthitis |0
septic shock |0
pig cattle exposure |-120
outbreak |0
epidemic |0
meningitis |0
secondary bacteremia |0
oppressive holocranial headache |-120
strong intensity |-120
fever |-120
duration five days |-120
hearing loss |-120
vomiting |-120
dysthermic sensation |-120
onset of disease after preparation of roast pork |-120
handling of roast pork |-120
intake of roast pork |-120
treatment with diazepam |-120
treatment with metamizole |-120
treatment with tramadol |-120
treatment with metoclopramide |-120
referred to Hospital Emergency Department |-120
persistent headache |-120
oxygen saturation 85% |0
diaphoresis |0
signs of meningeal irritation |0
progressive state of agitation |0
cranial computed tomography scan |0
no pathological findings |0
lumbar puncture |0
cloudy-whitish cerebrospinal fluid |0
CSF bacteriological culture |0
CSF cytochemical study |0
blood culture |0
white blood cell count 18.7 x 10³/µL |0
hemoglobin 15.2 g/dL |0
platelet count 115 x 10³/µL |0
glucose 141 mg/dL |0
creatinine 0.8 mg/dL |0
lactate 15.7 mg/dL |0
C-reactive protein 7 mg/dL |0
procalcitonin 0.45 ng/mL |0
CSF glucose <10 mg/dL |0
CSF total protein 950 mg/dL |0
CSF leukocytes 13,720/µL |0
polymorphonuclear neutrophils 98% |0
Gram-positive diplococci |0
differential diagnosis |0
purulent meningitis |0
septic encephalopathy |0
administration of dexamethasone |0
broad-spectrum antimicrobial therapy |0
ampicillin |0
ceftriaxone |0
vancomycin |0
acyclovir |0
alpha-hemolytic streptococci isolation in CSF |24
alpha-hemolytic streptococci isolation in blood cultures |24
identified as S. suis |24
antibiotic susceptibility to penicillin |24
antibiotic susceptibility to cefotaxime |24
antibiotic susceptibility to levofloxacin |24
antibiotic susceptibility to vancomycin |24
targeted treatment with cefotaxime |24
referred to Internal Medicine Service |144
stayed for three weeks |144
hearing loss at admission |0
inter-consultation with otorhinolaryngology |0
audiometry |0
complementary tests |0
normal test results |0
exacerbation of hearing loss |0
appearance of tinnitus |0
discharged after four weeks |672
treatment with amoxicillin/clavulanic acid |672
scheduled follow-up |672
S. suis infection due to contact with pigs |0
consumption of contaminated meat |0
occupational disease |0
use of metaphylactic agents |0
vaccination |0
improvement in hygienic conditions |0
instruction of pig workers |0
training of pig workers |0
barrier methods during handling |0
hand washing |0
proper cooking of meat |0
early use of dexamethasone |0
reduced incidence of hearing loss |0
reduced neurological sequelae |0
