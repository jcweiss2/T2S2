70 years old | 0
    female | 0
    Diabetes Mellitus | -672
    chronic renal disease | -672
    hypertension | -672
    pacemaker | -672
    anticoagulants | -672
    admitted to the hospital | 0
    left deep ear pain | 0
    gradual decrease in hearing | 0
    facial asymmetry | -168
    no tinnitus | 0
    no discharge | 0
    no itching | 0
    febrile | 0
    left ear edema | 0
    left ear pain on touch | 0
    tympanic membrane not visible | 0
    ear pack inserted | 0
    polypoidal mass in left external canal | 0
    inflammatory mass | 0
    right ear unremarkable | 0
    facial nerve weakness | 0
    oral asymmetry | 0
    forehead asymmetry | 0
    unable to raise right eyebrow | 0
    incomplete eye closure | 0
    mouth drop on smiling | 0
    grade 2 left facial palsy | 0
    hypoglossal nerve palsy | 0
    mild bulging in fossa of Rusenmuller | 0
    COVID-19 nasopharyngeal swab negative | 0
    IV Tazocin | 0
    IV Fortum | 0
    slurred speech | 24
    CT scan of ear and skull base | 24
    left nasopharyngeal mass | 24
    bone erosion | 24
    skull base destruction | 24
    suspected jugular thrombosis | 24
    left middle ear opacity | 24
    left mastoid opacity | 24
    left sphenoidal sinus mucosal thickening | 24
    surgical debridement | 48
    biopsy of nasopharynx | 48
    biopsy of left ear mass | 48
    fungal hyphae with right angle branching | 48
    mucormycosis | 48
    discontinued IV Tazocin | 48
    discontinued IV Fortum | 48
    started liposomal amphotericin B | 48
    insulin therapy | 48
    Eliquis administered | 48
    hypothermia | 96
    AKI on CKD | 96
    hyponatremia | 96
    discontinued liposomal amphotericin B | 96
    started Posaconazole | 96
    septic shock | 120
    WBC 39 109/L | 120
    hypotension | 120
    tachycardia | 120
    shifted to ICU | 120
    levophid infusion | 120
    death | 144