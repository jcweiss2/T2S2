54 years old | 0
female | 0
admitted to the hospital | 0
type 2 diabetes mellitus | -7776
basal insulin 20 IU per day | -7776
home-based capillary blood glucose monitoring 300 mg/dL | -7776
urinary symptoms | -72
nausea | -72
diffuse abdominal pain | -72
fatigue | -72
increased urinary frequency | -72
urgency | -72
acute urinary retention | -72
Foley catheter | -72
fevers 39 °C | -48
vomiting | -48
blood pressure 58/36 mmHg | 0
pulse 77 beats per minute | 0
respiration rate 26 breaths per minute | 0
body temperature 36 °C | 0
room-air oxygen saturation 92 % | 0
capillary blood glucose 337 mg/dL | 0
altered mental status | 0
Glasgow Coma Scale 12 points | 0
capillary refill 3 s | 0
normal lung examination | 0
abdomen without signs of peritoneal irritation | 0
vesical globus | 0
bilateral costovertebral angle tenderness | 0
hematuria | 0
resuscitation with IV fluids | 0
vasopressor agents | 0
third-generation cephalosporins | 0
leukocytes 35.7 × 10^3/uL | 0
total neutrophils 33.4 × 10^3/uL | 0
hemoglobin 11.7 g/dl | 0
platelets 138 × 10^3/uL | 0
fibrinogen 981 mg/dL | 0
creatinine 4.3 mg/dL | 0
glucose 334 mg/dL | 0
urea 132 mg/dL | 0
corrected sodium 136 mEq/L | 0
potassium 5 mEq/L | 0
chloride 94 mEq/L | 0
calculated serum osmolality 282 mOsm/L | 0
pH 7.31 | 0
PCO2 25 mmHg | 0
PO2 37 mmHg | 0
HCO3 12.37 mmol/L | 0
base excess -13.7 mmol/L | 0
leukocyte esterase test positive | 0
nitrite test negative | 0
500 leukocytes per high-power field | 0
ketones | 0
ESBL-producing E. coli | 0
meropenem-sensitive | 0
levofloxacin-resistant | 0
non-contrast abdominal CT scan | 0
loss of anatomy | 0
gas in the perirenal space | 0
pneumoperitoneum | 0
septic shock | 0
grade IV emphysematous pyelonephritis | 0
mild diabetic ketoacidosis | 0
stage 3 acute kidney injury | 0
carbapenem antibiotics | 0
fluid resuscitation | 0
IV insulin | 0
total bilateral nephrectomy | 24
appendectomy | 24
necrosis greater than 90 % | 24
parenchymal abscesses | 24
septic thrombi | 24
acute appendicitis | 24
Intensive Care Unit | 24
continuous veno-venous hemofiltration | 24
death | 192