29 years old | 0
    women | 0
    presented to hospital | -4032
    self-inflicted gunshot injury to abdomen | -4032
    three wounds (epigastrium, left hypochondrium, left lumbar area) | -4032
    underwent laparotomy | -4032
    perforation in antrum of stomach | -4032
    multiple small bowel perforations | -4032
    primary surgical repair | -4032
    bilateral lateral (zone 2) retroperitoneal hematomas | -4032
    non-expanding hematomas | -4032
    non-pulsatile hematomas | -4032
    transferred to ICU | -4032
    developed pulmonary embolism | -4032
    developed DIC | -4032
    managed with blood products | -4032
    recovered over one month | -4032
    discharged home | -4032
    presented two weeks later to local health center | -2688
    left iliac fossa pain | -2688
    watery stool | -2688
    reduced hemoglobin level | -2688
    raised serum CRP | -2688
    underwent abdominal CT scan | -2688
    left-sided retroperitoneal collection | -2688
    contrast extravasation into retroperitoneal space | -2688
    left ureteral injury | -2688
    urinoma formation | -2688
    colonic fistula | -2688
    referred to trauma center | -2688
    underwent cystoscopy | 0
    retrograde pyelogram | 0
    complete transection of left upper ureter | 0
    contrast extravasation into retroperitoneal space | 0
    underwent left percutaneous nephrostomy | 0
    left-sided pigtail drain inserted | 0
    treated with antibiotics | 0
    sepsis workup showed multi-drug-resistant coliform | 0
    clear urine draining from urinoma | 0
    repeat CT scan one week later | 168
    reduction in size of left-sided urinoma | 168
    peripherally enhancing collection in right pelvis | 168
    compression of urinary bladder | 168
    underwent pigtail drain insertion | 168
    minimal dark reddish fluid drained | 168
    drain removed after 48 hours | 216
    discharged | 216
    brought back three weeks later | 720
    elective surgery | 720
    cystoscopy prior to surgery | 720
    extra-luminal compression of bladder | 720
    intraoperative dense fibrosis in upper ureter | 720
    complete ureteral transection | 720
    mobilized ureter | 720
    left end-to-end ureteric anastomosis | 720
    excision of injured ureter | 720
    ureteroureterostomy | 720
    spatulation of ends | 720
    tension-free waterproof anastomosis over DJS | 720
    colonoscopy intraoperatively | 720
    methylene blue instillation through pigtail drain | 720
    negative methylene blue testing | 720
    spontaneous fistula healing | 720
    discharged on third post-operative day | 792
    seen in OPD two months later | 3600
    flexible cystoscopy | 3600
    removal of left DJS | 3600
    failed follow-up | 3600