41 years old | 0
male | 0
presented with lower extremity edema | -504
presented with fatigue | -504
presented with shortness of breath | -504
pale appearance | 0
melenic stool on rectal examination | 0
admitted to ICU | 0
resuscitation | 0
urgent endoscopy | 0
multiple gastric ulcers | 0
diffuse lymphadenopathy | 0
suspected metastatic lymphoma | 0
excisional biopsy | 0
Hodgkin lymphoma | 0
acute renal failure | 0
temporary hemodialysis | 0
acute respiratory failure | 0
intubation | 0
septic shock | 0
vasopressor support with norepinephrine | 0
sedation with propofol | 0
sedation with fentanyl | 0
ventilator use | 0
sudden onset of ST-segment elevations | 0
significant abdominal distention | 0
no murmurs on cardiac auscultation | 0
blood pressure 101/57 mmHg | 0
heart rate 112 beats/min | 0
respiratory rate 23 breaths/min | 0
oxygen saturation 99% | 0
sinus tachycardia | 0
ST-segment elevations in precordial leads | 0
deep T-wave inversions | 0
J-point depression in inferior leads | 0
marked QT prolongation | 0
ECG interpreted as STEMI | 0
emergency cardiology consultation | 0
troponin-T <0.01 ng/ml | 0
potassium 4.3 mEq/l | 0
calcium 7.6 mg/dl | 0
anion gap 12 mEq/l | 0
hemoglobin 10.1 g/dl | 0
hematocrit 29.4% | 0
pH 7.40 | 0
bicarbonate 21 mmol/l | 0
lactate 3.1 mmol/l | 0
LVEF 60-65% | 0
no regional wall motion abnormalities | 0
no pericardial effusion | 0
abrupt resolution of ST-segment elevations with ultrasound probe | 0
no significant abdominal compression during ultrasound | 0
resolution of ST-segment elevations with abdominal palpation | 0
significant gastric distention | 0
ileus | 0
gastric decompression with nasogastric tube | 0
resolution of ST-segment elevations post-decompression | 0
deferred coronary angiography | 0
no further ST-segment changes | 0
new-onset seizures | 0
focal neurological deficits | 0
leptomeningeal enhancement | 0
metastatic spread | 0
comfort care | 0
death | 0
