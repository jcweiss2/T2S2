64 years old | 0
male | 0
admitted to the hospital | 0
fever | -336
back pain | -336
no gastro-intestinal symptoms | -336
blood culture showed Salmonella enterica infection | -336
sensitive to Ampicillin/Sulbactam | -336
sensitive to Doripenem | -336
sensitive to Doxycycline | -336
sensitive to Imipenem | -336
sensitive to Amoxicillin/Clavulanic acid | -336
sensitive to Ampicillin | -336
sensitive to Cefepime | -336
sensitive to Cefotaxime | -336
sensitive to Ceftazidime | -336
sensitive to Ceftriaxone | -336
sensitive to Meropenem | -336
sensitive to Ertapenem | -336
sensitive to Piperacillin/Tazobactam | -336
received meropenem 1g daily for 7 days | -336
history of coronary artery bypass grafting surgery | -2628
history of steroid-induced diabetes mellitus | -2628
history of chronic kidney disease | -2628
readmitted to the emergency ward | 0
hypotension | 0
persistently high fever | 0
severe back pain | -168
paraplegia | -168
pain centered in the upper back | -168
pain radiating to the chest wall | -168
Visual Analogue Scale (VAS) 7 | -168
weakness of both lower extremities | -168
sensory loss below the chest | -168
no history of recent trauma | -168
lost 1 kg of weight in the past one month | -168
blood sample for hematology and coagulation profile | 0
blood culture | 0
urinary sample | 0
no leukocytosis | 0
increase in neutrophils | 0
decrease in lymphocytes | 0
C-Reactive Protein high | 0
procalcitonin 0.27 ng/mL | 0
Mantoux test negative | 0
IGRA negative | 0
HIV testing negative | 0
CD4 cell count 504 cells/mm3 | 0
referred to the intensive care unit | 0
septic shock | 0
given high dose meropenem injection | 0
renal function normal | 0
maximum level of 37 mg/dL for ureum | 0
maximum level of 1.23 mg/dL for creatinine | 0
critical condition subsided | 120
re-assessed for neurological deficit | 120
consulted an orthopedic spine surgeon | 120
midline tenderness over the upper thoracic spine region | 120
spinal cord compression | 120
signs of upper motor neuron involvement | 120
decreased sensation from Th5 dermatome | 120
Medical Research Council Scale for muscle power of 0/5 from L2-S1 | 120
Magnetic resonance imaging (MRI) of the spine | 120
wedging on the 5th and 6th thoracal | 120
intrathecal infiltration of hyperintensity mass in T2 weighted images | 120
posterior stabilization with pedicle screws and rods system | 168
transpedicular biopsy on 6th vertebra | 168
purulent discharge from the 6th thoracal body | 168
tissue samples for culture and pathological exam | 168
debridement | 168
decompression by laminectomy and flavectomy | 168
granulation tissue found underneath the laminae and yellow ligament | 168
postoperatively sent back to ICU | 168
pathological exam revealed chronic inflammation | 168
no tuberculoma and caseous necrotic formation | 168
no malignant cells | 168
tissue culture revealed Salmonella enterica infection | 168
same sensitivity profile as the previous blood culture | 168
changed antibiotic regimen to ciprofloxacin | 168
ciprofloxacin 400 mg IV twice daily for two weeks | 168
ciprofloxacin 500 mg twice daily for 6 weeks | 168
total of 8 weeks therapeutic antibiotic | 168
discharged | 504
significant improvement of neurological condition | 504
excellent motoric strength (ASIA E) | 504
free of fever | 504
slight discomfort over the surgical scar | 504
pain significantly subsided | 504
independently ambulated with a spinal brace | 504
symptom-free at 3 month follow-up | 936
began exercises to strengthen the back | 936