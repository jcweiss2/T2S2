26 years old | 0
male | 0
previously diagnosed with restrictive subaortic ventricular septal defect | -6480
previously diagnosed with mild pulmonary hypertension | -6480
no history of drug abuse | 0
presented to the hospital in critical condition | 0
hypochromic anemia | -6480
fatigue | -6480
effort limitation | -6480
exertional dyspnea | -6480
ascites | -6480
persistent inflammatory syndrome | -6480
weight loss of 20 kg | -6480
increased blood cell count | 0
C-reactive protein 76 mg/L | 0
procalcitonin 0.77 ng/mL | 0
anemia | 0
thrombocytopenia | 0
echocardiography revealing infective endocarditis | 0
mobile vegetations | 0
severe regurgitation of aortic valve | 0
severe regurgitation of tricuspid valve | 0
severe regurgitation of pulmonary valve | 0
aortic annulus abscess | 0
restrictive ventricular septal defect | 0
severely dilated left ventricle | 0
dilated right ventricle | 0
severe biventricular dysfunction | 0
left ventricle ejection fraction 25% | 0
tricuspid annular plane systolic excursion 11 mm | 0
severe pulmonary hypertension | 0
broad-spectrum antibiotics initiated | 0
antifungals initiated | 0
septic shock | 0
multiple organ dysfunction syndrome | 0
hypotension | 0
hypoxemia | 0
severe metabolic acidosis | 0
oliguria | 0
neurologic dysfunction | 0
mechanical ventilation | 0
hemodynamic support with dobutamine | 0
hemodynamic support with norepinephrine | 0
continuous venovenous hemodiafiltration | 0
cytokine removal filter | 0
gram-negative bacilli found on blood cultures | 0
meropenem prescribed | 0
gradual clinical improvement | 168
weaning of norepinephrine | 168
weaning of mechanical ventilation | 168
organ functions recovered | 168
ventricular function improved | 168
LV ejection fraction 30% | 168
TAPSE 16 | 168
elevated pulmonary artery pressure | 168
dobutamine-dependent | 168
paroxysmal supraventricular tachycardia | 384
septic discharge | 384
fever >39°C | 384
WBC increase | 384
recurrence of septic shock | 384
hemodynamic deterioration | 384
lactate increase | 384
transient hepatic cytolysis | 384
oliguria | 384
clinical improvement after electrical conversion | 384
administration of dobutamine | 384
administration of levosimendan | 384
surgery performed | 432
bicaval-aortic cardiopulmonary bypass | 432
Custodiol cardioplegia | 432
aortic valve replaced | 432
tricuspid valve replaced | 432
pulmonary valve replaced | 432
aortic annular abscess debrided | 432
VSD closed with bovine pericardial patch | 432
sinus rhythm recovered | 432
dobutamine used post-CPB | 432
norepinephrine used post-CPB | 432
inhaled nitric oxide | 432
ultrafiltration with cytokine removal | 432
postoperative outcome good | 432
stable hemodynamics | 432
no arrhythmias | 432
extubation | 456
Milrinone infusion | 456
levosimendan administration | 576
inotrope withdrawal | 576
LVEF below 35% | 576
sacubitril/valsartan started | 576
valve cultures positive for Rhizobium radiobacter | 432
intravenous meropenem continued | 576
levofloxacin started | 576
co-trimoxazole started | 576
resumed work | 4320
normally functioning valves | 4320
improved ventricular function | 4320
no sign of infection | 4320
asymptomatic at 18 months | 12960
LVEF 50% | 12960
