13 years old | 0
female | 0
admitted to the hospital | 0
fever | -72
loss of appetite | -72
appendectomy | -72
dehydrated | 0
tachycardia | 0
tachypnea | 0
fever (axillary temperature was 38.8 °C) | 0
blood pressure was 120/70 mmHg | 0
cardiac examination was normal | 0
pulmonary examination was normal | 0
abdomen was diffusely tender | 0
rebound test was painful | 0
intestinal sounds were present and normal | 0
surgical scar was hyperemic | 0
abdominal ultrasound examination showed a pericolic image consistent with abscess | 0
abdominal secretion culture was positive for multisensitive E. coli and group G, β-hemolytic Streptococcus sp | 0
ceftriaxone and metronidazole were prescribed | 0
abdominal pain | 72
fever relapsed | 72
antibiotics were changed to vancomycin, ceftazidime and amikacin | 72
fever remained intermittently present | 72
abdominal computed tomography (CT) ruled out any surgical complication | 120
broad-spectrum antibiotic regimen, to which fluconazole was added | 120
hypotensive | 288
tachycardic | 288
temperature rose to 39.4 °C | 288
vasoactive drugs were required for hemodynamic stabilization | 288
blood and urine cultures were negative | 288
transthoracic echo Doppler Cardiogram was normal | 288
progressive respiratory failure | 288
referred to the ICU | 288
hemodialysis | 432
frequent blood transfusions | 432
died | 576
autopsy was performed | 576
Bogota bag closing the peritoneotomy | 576
mild serohemorrhagic effusion was drained | 576
non-dehiscent surgical sutures were revealed joining the distal ileum with the ascending colon | 576
liver was enlarged | 576
liver weighed 1280 g | 576
extensive poorly defined yellowish parenchyma areas were evident intermingled with winy-colored areas consistent with infarction | 576
extensive ischemic lobular necrosis was present | 576
macro and microvesicular steatosis | 576
spleen was enlarged | 576
spleen weighed 271 g | 576
cut surface was winy, friable, and consistent with a reactive pattern | 576
white pulp was depleted | 576
red pulp was congested | 576
numerous histiocytes, phagocytizing red blood cells, and lymphocytes were present | 576
pancreas weighed 70 g | 576
purplish areas at the cut surface | 576
steatonecrosis and ischemic necrosis | 576
adrenal glands exhibited extensive cortical ischemic necrosis | 576
petechiae were evident on both lung surfaces and pericardium | 576
heart weighed 191 g | 576
myocardial hemorrhagic suffusions mainly on the left ventricle | 576
recent pericardial and myocardial hemorrhage | 576
lungs presented increased volume | 576
cut surface was winy-colored | 576
parenchyma was not friable | 576
alveolar spaces were filled by numerous macrophages, fibrin, and red blood cells | 576
no hemophagocytosis was found at this site | 576
numerous mediastinal and intra-abdominal lymph nodes were detected | 576
sinusal histiocytosis lymphadenitis pattern with associated lymphocytic depletion and histiocytes with erythrocytes phagocytosis | 576
histiocytes were phenotypically CD68-positive, S100-negative | 576
bone marrow showed evident hypercellularity | 576
granulocytic series elements associated with the presence of numerous histiocytes with hemophagocytosis | 576
hypoxic-ischemic encephalopathy | 576
acute tubular necrosis | 576
hemophagocytic syndrome | 576
hemophagocytic lymphohistiocytosis (HLH) | 576
febrile illness | 0
multiple organ involvement | 0
hepatomegaly | 0
lymphadenopathy | 0
edema | 0
jaundice | 0
rash | 0
neurological symptoms | 0
cytopenias | 0
hypofibrinogenemia | 0
hyperferritinemia | 0
hemophagocytosis | 0
sustained fever | 0
elevated ferritin | 288
low fibrinogen | 288
thrombocytopenia | 480
hyperbilirubinemia | 480
enlarged prothrombin time | 480
altered liver enzymes | 480
exploratory laparotomy | 528
loose peritoneal adhesions | 528
no purulent secretion, nor intestinal perforation or bowel necrosis | 528
multiple organ failure | 576
hemophagocytic syndrome triggered by acute appendicitis | 576