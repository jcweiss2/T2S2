47 years old | 0
    male | 0
    presented to the emergency department | 0
    fever | -72
    sore throat | -72
    left-sided neck swelling | -72
    generalized fatigue | -72
    myalgia | -72
    no other symptoms | 0
    blood pressure 100/65 mmHg | 0
    heart rate 115 beats/min | 0
    temperature 38.9°C | 0
    respiratory rate 20 breaths/min | 0
    oxygen saturation 100% | 0
    throat congestion | 0
    left-sided mild posterior lymphadenopathy | 0
    remainder systemic examination insignificant | 0
    high C-reactive protein | 0
    slight rise in serum creatinine | 0
    high international normalized ratio | 0
    initial chest x-ray unremarkable | 0
    SARS-CoV-2 infection confirmed by RT-PCR | 0
    received hydroxychloroquine | 0
    received azithromycin | 0
    received cefuroxime | 0
    transferred to quarantine facility | 0
    developed diarrhea | 48
    developed vomiting | 48
    mild diffuse abdominal pain | 48
    abdominal pain became severe | 48
    abdominal pain localized to right lower quadrant | 48
    transferred back to hospital | 48
    looked sick | 48
    alert | 48
    not oriented | 48
    blood pressure 84/52 mmHg | 48
    heart rate 102 beats/min | 48
    temperature 38.1°C | 48
    oxygen saturation 96% | 48
    diffuse abdominal tenderness | 48
    right iliac fossa guarding | 48
    acute kidney injury | 48
    transaminitis | 48
    worsening CRP | 48
    worsening procalcitonin | 48
    repeat chest x-ray bilateral reticular infiltrates | 48
    shifted to intensive care unit | 48
    started on meropenem | 48
    resuscitated with crystalloid fluids | 48
    CT scan abdomen no bowel perforation | 48
    CT scan abdomen no appendiceal inflammation | 48
    diffuse paracolic gutters fat stranding | 48
    mild free fluid | 48
    bilateral mild pleural effusion | 48
    consolidations | 48
    filling defect at superior mesentery vein | 48
    CT angiogram abdomen suboptimal venous system opacification | 48
    no acute thrombosis detected | 48
    patent major abdominal arterial system | 48
    high serum lipase >600 U/L | 48
    high serum amylase 451 U/L | 48
    sepsis workup unremarkable | 48
    surgical causes ruled out | 48
    treated conservatively | 48
    pain settled within few days | 48
    kidney injury improved | 48
    liver injury improved | 48
    inflammatory markers trending down | 48
    discharged | 48
    asymptomatic follow-up | 48
<|eot_id|>
    
47 years old | 0
male | 0
presented to the emergency department | 0
fever | -72
sore throat | -72
left-sided neck swelling | -72
generalized fatigue | -72
myalgia | -72
no other symptoms | 0
blood pressure 100/65 mmHg | 0
heart rate 115 beats/min | 0
temperature 38.9°C | 0
respiratory rate 20 breaths/min | 0
oxygen saturation 100% |$0
throat congestion | 0
left-sided mild posterior lymphadenopathy | 0
remainder systemic examination insignificant | 0
high C-reactive protein | 0
slight rise in serum creatinine | 0
high international normalized ratio | 0
initial chest x-ray unremarkable | 0
SARS-CoV-2 infection confirmed by RT-PCR | 0
received hydroxychloroquine | 0
received azithromycin | 0
received cefuroxime | 0
transferred to quarantine facility | 0
developed diarrhea | 48
developed vomiting | 48
mild diffuse abdominal pain | 48
abdominal pain became severe | 48
abdominal pain localized to right lower quadrant | 48
transferred back to hospital | 48
looked sick | 48
alert | 48
not oriented | 48
blood pressure 84/52 mmHg | 48
heart rate 102 beats/min | 48
temperature 38.1°C | 48
oxygen saturation 96% | 48
diffuse abdominal tenderness | 48
right iliac fossa guarding | 48
acute kidney injury | 48
transaminitis | 48
worsening CRP | 48
worsening procalcitonin | 48
repeat chest x-ray bilateral reticular infiltrates | 48
shifted to intensive care unit | 48
started on meropenem | 48
resuscitated with crystalloid fluids | 48
CT scan abdomen no bowel perforation | 48
CT scan abdomen no appendiceal inflammation | 48
diffuse paracolic gutters fat stranding | 48
mild free fluid | 48
bilateral mild pleural effusion | 48
consolidations | 48
filling defect at superior mesentery vein | 48
CT angiogram abdomen suboptimal venous system opacification | 48
no acute thrombosis detected | 48
patent major abdominal arterial system | 48
high serum lipase >600 U/L | 48
high serum amylase 451 U/L | 48
sepsis workup unremarkable | 48
surgical causes ruled out | 48
treated conservatively | 48
pain settled within few days | 48
kidney injury improved | 48
liver injury improved | 48
inflammatory markers trending down | 48
discharged | 48
asymptomatic follow-up | 48