60 years old | 0
female | 0
hepatitis B virus-induced liver cirrhosis | 0
hepatocellular carcinoma (HCC) | 0
diagnosed with hepatitis B virus-induced liver cirrhosis and hepatocellular carcinoma (HCC) | -52512
trans&shy;arterial chemoembolization | -52512
palliative radiotherapy | -52512
albuterol inhaler use once a month for asthma | 0
umbilical hernia repair | -17520
total thyroidectomy for papillary thyroid carcinoma | -35040
antiviral agent for hepatitis B virus | 0
warfarin for portal vein thrombosis | 0
diuretics for ascites | 0
refractory ascites | 0
preoperative hematocrit 0.283% | 0
preoperative hemoglobin 9.2 g/dl | 0
preoperative platelet count 63000 /μl | 0
preoperative prothrombin time INR 1.17 | 0
preoperative sodium 133 mmol/L | 0
preoperative MELD score 15 points | 0
vital signs within normal range | 0
preoperative chest radiography confirmed no active lung lesion | 0
preoperative elevated diaphragm | 0
preoperative pulmonary function test showed severe obstructive and moderate restrictive pattern | 0
transthoracic echocardiography showed diastolic dysfunction grade 1 | 0
esophagogastroduodenoscopy revealed esophageal varices | 0
portal hypertensive gastropathy | 0
gastric varices at cardia | 0
ABO-incompatible living donor liver transplantation (ABO-i LDLT) planned | 0
son's AB blood type | 0
rituximab (525 mg) administered two weeks prior to LT | -336
isoagglutinin IgM and IgG titers against B antigen measured before rituximab injection | -336
isoagglutinin titers measured daily for 7 days before surgery | -168
plasmapheresis with AB FFP | -168
target isoagglutinin titer < 1 : 16 | 0
two consecutive plasmaphereses | -168
RBC antibody screen negative 1 day prior to operation | -24
preoperative preparation of 5 units of packed RBCs of blood group A | 0
albuterol administered | 0
anesthesia induced with thiopental sodium, rocuronium, and sevoflurane | 0
radial artery cannulation | 0
bispectral index (BIS) monitoring | 0
RBC antibody screen positive 2 days prior to surgery | -48
packed RBCs cross&shy;matched | 0
femoral artery and vein catheter insertion | 0
central catheter placement via left internal jugular vein | 0
IVC reconstruction | 0
methylprednisolone infusion during portal vein anastomosis | 0
basiliximab infusion after reperfusion | 0
hepatic artery bleeding controlled | 0
diaphragm repair | 0
chest tube insertion | 0
open abdomen transfer to ICU | 0
total anesthesia time 16 h 30 min | 0
crystalloid administration 17,500 ml | 0
5% albumin administration 1,200 ml | 0
6% hydroxyethyl starch administration 1,500 ml | 0
pre-storage leukocyte&shy;reduced RBCs 5 units | 0
leukocyte&shy;depleted RBCs 5 units | 0
Cell Saver blood 4,872 ml | 0
AB FFP 9 units | 0
AB SDP 2 units | 0
AB cryoprecipitate 12 units | 0
intraoperative blood loss 4,123 ml | 0
urine output 1,320 ml | 0
wound closure on POD 2 | 48
wedge biopsy of transplanted liver | 48
biopsy showing centrilobular hemorrhagic necrosis | 48
graft dysfunction with hepatic vein stricture | 48
tracheostomy on POD 7 | 168
IgM and IgG antibodies increased | 168
IgM titer 1 : 4 | 168
IgG titer 1 : 8 | 168
no further plasmapheresis | 168
re&shy;transplantation planned | 168
sepsis | 744
expired on POD 31 | 744
RBC antibody screen conversion | 0
first SDP transfusion 3 years prior | -26280
first RBC antibody screen negative | -26280
second SDP transfusion 2 years prior | -17520
second RBC antibody screen positive | -17520
anti-C (Rh system) identified | -17520
anti-M (MNS system) identified | -17520
electronic medical record system marking 'Ab' | 0
RBC antibody screen result window revision needed | 0
