59 years old | 0
female | 0
Vietnamese | 0
admitted to the hospital | 0
syncopal episode | 0
motor vehicle accident | 0
gastrointestinal illness | -48
vomiting | -48
abdominal pain | -48
received COVID-19 vaccine | -336
thalassaemia | 0
sinus rhythm | 0
fixed ST elevation | 0
low QRS voltages | 0
cardiac troponin I elevated | 0
c-reactive protein elevated | 0
erythrocyte sedimentation rate elevated | 0
calcified granuloma | 0
left ventricular ejection fraction 30% | 0
moderate-severe global systolic dysfunction | 0
mild concentric increase in wall thickness | 0
severely reduced tissue Doppler velocities | 0
mild-moderate aortic regurgitation | 0
moderate pericardial effusion | 0
symptomatic hypotension | 24
bradycardia | 24
new bundle branch blocks | 24
high grade atrioventricular block | 24
left bundle branch block | 24
isoprenaline infusion | 24
transferred to coronary care unit | 24
permanent pacemaker insertion | 48
persistently hypotensive | 48
oliguric | 48
dopamine infusion | 48
conscious, symptomatic episodes of brief accelerated idioventricular rhythm | 48
transferred to intensive care unit | 48
severe LV dysfunction | 72
ejection fraction 10% | 72
global hypokinesis | 72
severely impaired RV systolic function | 72
dilated inferior vena cava | 72
endomyocardial biopsy | 96
florid infiltrate of lymphocytes | 96
histiocytes | 96
plasma cells | 96
scattered eosinophils | 96
marked oedema | 96
cardiomyocyte necrosis | 96
poorly formed granulomas | 96
giant cell myocarditis | 96
intravenous methylprednisone | 96
cyclosporin | 96
progressively worsening lactic acidosis | 120
intubated | 120
transferred to cardiac transplant centre | 120
biventricular assist device inserted | 144
haemorrhage | 144
coagulopathy | 144
massive transfusion | 144
thoracic washout | 144
multiorgan failure | 168
hepatic encephalopathy | 168
anuric renal failure | 168
dialysis | 168
distal ischaemia of limbs | 168
digital gangrene | 168
bowel ischaemia | 168
immune thrombocytopaenia | 168
intravenous immunoglobulin | 168
plasma exchange | 168
polymicrobial sepsis | 168
Pseudomonas aeruginosa bacteraemia | 168
Candidaemia | 168
meropenem | 168
vancomycin | 168
caspofungin | 168
LV assist device explanted | 432
redo-sternotomy | 432
tissue aortic valve replacement | 432
RV assist device explanted | 600
cerebral infarction | 600
unresponsive off sedation | 600
palliated | 648
passed away | 648