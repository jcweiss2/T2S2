21 years old | 0 | 0 
male | 0 | 0 
obese | 0 | 0 
admitted to the hospital | 0 | 0 
cough | -72 | 0 
fever | -72 | 0 
shortness of breath | -72 | 0 
pleuritic chest pain | -72 | 0 
light-headedness | -24 | 0 
near syncope | -24 | 0 
dyspnoea | -24 | 0 
COVID-19 | 0 | 0 
sub-massive pulmonary embolism | 0 | 0 
unfractionated heparin | 0 | 12 
hypotensive | 12 | 12 
massive pulmonary embolism | 12 | 12 
catheter-directed thrombolysis | 12 | 18 
improved clinically | 18 | 24 
planned discharge | 24 | 24 
acute respiratory failure | 72 | 72 
hypotension | 72 | 72 
intubated | 72 | 72 
cardiac arrest | 72 | 72 
return of spontaneous circulation | 72 | 72 
vasopressors | 72 | 120 
extracorporeal membrane oxygenation | 72 | 240 
recurrent massive pulmonary embolism | 72 | 120 
repeat catheter-directed thrombolysis | 120 | 126 
ventilation parameters improved | 120 | 240 
vasopressors discontinued | 120 | 240 
weaning of extracorporeal membrane oxygenation | 120 | 240 
deep venous thrombus | 168 | 168 
inferior vena cava filter | 168 | 168 
low-molecular-weight heparin | 168 | 504 
septic shock | 240 | 240 
treated with broad spectrum antibiotics | 240 | 240 
right thigh haematoma | 360 | 360 
compartment syndrome | 360 | 360 
surgical debridement | 360 | 360 
transitioned to rivaroxaban | 360 | 504 
discharged | 504 | 504 
anticoagulated on rivaroxaban | 504 | 1008 
no major adverse events | 1008 | 1008 
returned home | 1008 | 1008 
performing activities of daily living independently | 1008 | 1008