74 years old | 0 | 0 
male | 0 | 0 
admitted to the hospital | 0 | 0 
hypertension | 0 | 0 
diabetes mellitus | 0 | 0 
intermittent subjective fever | -96 | 0 
rigors | -96 | 0 
generalized headache | -96 | 0 
altered mentation | -96 | 0 
body malaise | -96 | 0 
nausea | -96 | 0 
vomiting | -96 | 0 
no history of loss of consciousness | -96 | 0 
no abdominal pain | -96 | 0 
no change in stool habits/urine color | -96 | 0 
no recent trauma or falls | -96 | 0 
febrile | 0 | 0 
tachypneic | 0 | 0 
disoriented | 0 | 0 
good nutritional status | 0 | 0 
not jaundiced | 0 | 0 
not cyanosed | 0 | 0 
pulse rate of 103 beats/min | 0 | 0 
respiratory rate of 23 breaths/min | 0 | 0 
blood pressure of 96/60 mmHg | 0 | 0 
saturating at 98% on room air | 0 | 0 
normal vesicular breath sounds | 0 | 0 
normal abdominal examination | 0 | 0 
IV resuscitation | 0 | 0 
analgesia | 0 | 0 
WBC of 8.2 × 103/μL | 0 | 0 
hemoglobin of 11.5 g/dL | 0 | 0 
thrombocytopenia of 46,000/mm3 | 0 | 0 
elevated creatinine 117 μmol/L | 0 | 0 
BUN 10.5 mmol/L | 0 | 0 
slightly low sodium of 131 mmol/L | 0 | 0 
normal serum electrolytes | 0 | 0 
normal liver | 0 | 0 
normal coagulation profile | 0 | 0 
normal Chest X-ray | 0 | 0 
P. falciparum with high parasitemia | 0 | 0 
admitted to the ICU | 0 | 72 
intravenous artesunate-based regimen | 0 | 72 
supportive measures | 0 | 72 
improvement in clinical status | 72 | 72 
improvement in lab parameters | 72 | 72 
shifted to the general ward | 72 | 72 
acute abdomen | 120 | 120 
progressive, dull, constant generalized abdominal pain | 120 | 120 
nausea | 120 | 120 
non-bilious vomiting | 120 | 120 
anxious | 120 | 120 
afebrile | 120 | 120 
diaphoretic | 120 | 120 
tachycardic | 120 | 120 
tachypneic | 120 | 120 
hypotensive | 120 | 120 
saturating well on room air | 120 | 120 
slightly distended abdomen | 120 | 120 
tender on superficial palpation | 120 | 120 
inaudible bowel sounds | 120 | 120 
low Hb of 7.1 g/dL | 120 | 120 
hypoechoic nodular cystic area | 120 | 120 
hyperdense intrasplenic hematoma | 120 | 120 
hypodense subcapsular hematoma | 120 | 120 
splenic laceration | 120 | 120 
intraperitoneal free fluid | 120 | 120 
grade 3 splenic injury | 120 | 120 
blood products mobilized | 120 | 120 
adequate resuscitation | 120 | 120 
explorative laparotomy | 120 | 120 
splenectomy | 120 | 120 
2.5 L of frank blood evacuated | 120 | 120 
enlarged spleen | 120 | 120 
long laceration on the upper pole | 120 | 120 
uneventful postoperative period | 120 | 168 
discharged home | 168 | 168 
fully recovered | 168 | 168 
post-splenectomy care | 168 | 168