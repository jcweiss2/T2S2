49 years old | 0
male | 0
alcohol abuse | 0
esophageal rupture | 0
severe retrosternal chest pain | -40
vomiting | -40
dyspnea | -40
intubated | -40
admitted to the medical intensive care unit | -40
small left pneumothorax | -40
subcutaneous emphysema | -40
chest tube placed | -40
hypotensive | -40
vasopressor support | -40
septic shock | -40
CT of the chest | -24
oral contrast material through the nasogastric tube | -24
esophageal perforation | -24
EGD | -24
3-cm linear perforation in the distal esophagus | -24
EndoVAC therapy | 0
nothing by mouth | 0
Dobhoff tube | 0
PEG-J | 0
EndoVAC procedure repeated | 72
EndoVAC sessions | 72
granulation tissue | 168
fourth EndoVAC | 168
follow-up EGDs | 216
chest CT | 216
barium swallow | 216
complete healing of the esophageal perforation | 216
discharged | 504 
life-flighted to our tertiary care medical center | -40
nasogastric feeding tube | -24
gastrojejunal feeding tube | 168
healthy granulation tissue | 216
healed esophageal perforation | 216
no leakage of contrast material | 216