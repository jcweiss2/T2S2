48 years old | 0
female | 0
G6P2042 | 0
admitted to the hospital | 0
fever | -360
chills | -360
diffuse abdominal pain | -360
abnormal uterine bleeding | -720
dysmenorrhea | -720
large uterine fibroids | -720
underwent UAE | -360
hypertension | 0
obesity class III | 0
cholecystectomy | -10000
thyroidectomy | -10000
left knee meniscal repair | -10000
two term uncomplicated vaginal deliveries | -10000
four spontaneous abortions | -10000
temperature of 101.5F | 0
heart rate of 110 beats per minute | 0
respiratory rate of 24–37 breaths per minute | 0
normal blood pressure | 0
abdomen was distended | 0
diffusely tender | 0
scant blond‑tinged vaginal discharge | 0
white blood cell count was 26,300 | 0
91% neutrophils | 0
CT scans of the abdomen and pelvis | 0
distended uterus | 0
multiple intra-cavitary uterine masses | 0
large amount of gas | 0
air–fluid level | 0
broad-spectrum intravenous antibiotics | 0
fluid resuscitation with lactated ringers | 0
exploratory laparotomy | 12
possible hysterectomy | 12
abscess drainage | 12
purulent material in the pelvis | 12
enlarged uterus | 12
inflamed, necrotic uterine fundus | 12
adherent to severely inflamed small bowel | 12
total hysterectomy | 12
bilateral salpingectomy | 12
small bowel resection | 12
primary end-to-end anastomosis | 12
frozen section of the uterus | 12
negative for malignancy | 12
ovaries were spared | 12
transferred to the surgical intensive care unit | 12
prolonged course of antibiotics | 12
discharged from the hospital | 504
poorly differentiated serous carcinoma of the fallopian tube | 720
staging procedure | 720
stage 1a fallopian tube carcinoma | 720
following up with the oncology service | 720