14 years old | 0
male | 0
admitted to the hospital | 0
near-drowning incident | -1
cardiopulmonary resuscitation (CPR) | -1
abdominal pain | 0
diffuse abrasions on torso | 0
hemodynamically stable | 0
fully conscious | 0
pneumoperitoneum | 0
pneumomediastinum | 0
intraabdominal free fluid | 0
hollow viscus perforation | 0
taken to the operating room | 1
gross contamination with food debris | 1
total gastroesophageal junction (GEJ) disruption | 1
patient became hemodynamically labile | 1
damage control procedure | 1
distal esophagus and proximal stomach stapled closed | 1
discontinuity | 1
four drains placed | 1
mediastinal drain | 1
gastrostomy (G) tube | 1
large bore nasogastric (NG) tube | 1
septic shock | 24
respiratory failure | 24
prolonged intubation | 24
deep venous thrombosis | 24
pulmonary embolism | 24
bilateral pleural effusions | 24
general deconditioning | 24
parenteral nutrition | 24
extubated | 432
fluoroscopic evaluation | 432
leak in the esophagus | 432
stomach negative for leak | 432
enteral nutrition via G tube | 432
discharged | 1200
Ivor-Lewis distal esophagectomy | 2160
gastric pull-up for esophagogastric anastomosis | 2160
partial left lateral decubitus position | 2160
midline abdominal incision | 2160
gastric conduit | 2160
right thoracotomy | 2160
distal esophagus identified | 2160
tubularized portion of stomach advanced | 2160
esophagogastric anastomosis | 2160
leak test | 2160
jejunostomy tube | 2160
extubated | 2163
nutritionally supported with jejunostomy enteral feeds | 2167
esophagram | 2167
no leak at the anastomosis | 2167
initiated on liquid diet | 2167
discharged | 2170
tolerate regular diet | 2700
gaining weight | 2700
recovering well | 2700