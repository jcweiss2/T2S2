67 years old | 0
male | 0
Asian | 0
attended the emergency room | 0
nausea | -24
vomiting | -24
diarrhoea | -24
fever | -24
lower abdominal pain | -24
no haematemesis | -24
no melena | -24
no urinary complaints | -24
passed eight watery bowel motions | -24
no previous febrile illness | 0
no sweating | 0
no weight loss | 0
no STD | 0
no allergies | 0
non-smoker | 0
does not drink alcohol | 0
came to Saudi Arabia to perform Umrah | 0
looked sick | 0
dry mucous membranes | 0
temperature 38.7°C | 0
pulse rate 112/min | 0
blood pressure 140/90 | 0
oxygen saturation 98% | 0
severe tenderness at the right iliac fossa | 0
no rebound | 0
normal bowels sounds | 0
unremarkable heart and chest examinations | 0
WBC count 24,000×10^9/l | 0
90% neutrophils | 0
haemoglobin 10 g/dl | 0
normal MCV | 0
normal platelets | 0
serum creatinine 190 μmol/l | 0
urea nitrogen 12.5 mmol/l | 0
normal electrolytes | 0
normal liver function tests | 0
normal coagulation profile | 0
normal lactic acid | 0
stool analysis showed WBCs >20/hpf | 0
RBCs 3–5/hpf | 0
no ova or parasites | 0
blood culture negative | 72
stool culture negative | 72
Clostridium difficile PCR negative | 0
C-reactive protein high at 70 mg/l | 0
received saline | 0
received paracetamol | 0
received ciprofloxacin 500 mg intravenously | 0
CT scan of the abdomen and pelvis | 0
AAA arising just above the origins of both renal arteries | 0
hyper-dense retroperitoneal haematoma | 0
intramural thrombus | 0
AAA measured 74 mm at the maximum sagittal diameter | 0
aortic leak | 0
transferred to the vascular surgery team | 0
empirical antibiotics continued | 0
fever resolved | 24
inflammatory markers improved | 24
RPR serology normal | 24
chest x-ray normal | 24
underwent exploratory laparotomy | 48
large leaking juxtarenal AAA 10×7 cm in diameter | 48
aneurysm extended from the level of the renal artery down to the level of the iliac bifurcation | 48
intramural thrombus removed | 48
bifurcated silver-coated 20×10 mm Dacron graft applied | 48
postoperatively moved to the ICU | 48
received ventilation | 48
received inotropes | 48
correction of anaemia | 48
taken off the ventilator | 72
taken off inotropes | 72
renal functions normalized | 120
transferred to a normal ward | 120
started rehabilitation | 120
discharged | 504
flew back home | 504