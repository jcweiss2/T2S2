52 years old | 0
male | 0
presented to the Emergency Department | 0
septic shock | 0
right sided abdominal pain | 0
cardiac arrest | 0
cardiopulmonary resuscitation (CPR) | 0
return of spontaneous circulation (ROSC) | 10
broad spectrum intravenous antibiotics with cefuroxime and metronidazole | 0
intubation | 0
ventilation | 0
computer tomography (CT) scan of the abdomen | 0
moderate volume of free fluid | 0
locules of gas within the pelvis | 0
hollow viscus perforation | 0
calcified structure within the appendix | 0
foreign body causing perforated appendicitis | 0
laparotomy | 0
perforated appendicitis | 0
four-quadrant purulent peritonitis | 0
appendicectomy | 0
firm foreign body causing luminal obstruction | 0
decaying tooth containing a metallic filling | 0
washout with copious irrigation | 0
abdomen closed | 0
transferred to the intensive care unit (ICU) | 0
multi-organ failure | 36
sepsis | 36
death | 36
ingested teeth and dental prostheses causing appendicitis | -672
obstruction of the appendix lumen due to an exogenous foreign body | -672 
faecolith | -672 
appendicitis | -72 
impacted molar tooth | -72 
luminal obstruction | -72 
mucus production | -72 
gas production | -72 
distension of the distal appendix | -72 
pain | -72 
inflammation | -72 
impaired venous return | -72 
ischaemia | -72 
perforation | -72