67 years old | 0
female | 0
Caucasian | 0
admitted to the intensive care unit | 0
elective posterior spinal instrumentation and fusion with laminectomy | 0
chronic back pain | -720
obesity | -720
hypertension | -720
gastritis | -720
HSV1 | -720
tobacco use | -720
completed six courses of prednisone | -2160
desaturated to SpO2 of 85% | 24
oxygenation improved with continuous positive airway pressure | 24
bilateral lower lobe infiltrates | 24
glucocorticoid taper with dexamethasone and hydrocortisone | 0
hydrocortisone 100 mg | 0
dexamethasone 10 mg twice daily | 0
dexamethasone 8 mg twice daily | 24
dexamethasone 6 mg once | 48
hydrocortisone 50 mg every 6 h | 72
hydrocortisone 25 mg every 6 h | 120
acute kidney injury | 48
febrile episodes | 48
vancomycin | 48
piperacillin–tazobactam | 48
hemodynamically unstable | 120
hypercapnic respiratory failure | 120
intubated | 120
norepinephrine | 120
hemodialysis | 120
white blood cell count doubled | 144
procalcitonin elevated | 144
antimicrobials broadened to vancomycin and meropenem | 144
acute respiratory distress syndrome (ARDS) | 144
Candida albicans | 144
fluconazole | 144
concerns for immunosuppression | 144
β-D-Glucan not performed | 144
sputum negative for Pneumocystis jirovecii | 144
immunostaining showed many nuclear and cytoplasmic cells positive for HSV | 144
disseminated HSV1 infection confirmed with DNA PCR | 144
acyclovir | 144
history of oral HSV1 | -720
recurrent oral infections | -720
bloody output from the orogastric tube | 360
esophagogastroduodenoscopy | 360
diffuse esophageal and gastric ulcerations | 360
HSV esophagitis | 360
vasopressors discontinued | 384
extubated | 384
transferred out of the ICU | 672
improvement of renal function | 672
discontinuation of dialysis | 672
discharged | 936