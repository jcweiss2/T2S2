66 years old | 0
female | 0
admitted to the hospital | 0
haematuria | 0
nausea | 0
elevated calcium | 0
elevated alkaline phosphatase | 0
elevated amylase | 0
elevated lipase | 0
elevated creatinine | 0
elevated troponin T | 0
elevated C-reactive protein | 0
elevated white blood cell count | 0
septic shock | 0
admitted to the intensive care unit | 0
noradrenaline administration | 0
adrenaline administration | 0
calcitonin administration | 0
isotonic fluids administration | 0
severe pancreatitis | 0
parathyroid tumour | 0
thyroid or parathyroid tumour | 0
intact parathyroid hormone level | 24
ultrasound imaging | 24
hypoechoic heterogeneous tumour | 24
ill-defined borders | 24
parathyroid carcinoma | 24
hypercalcaemia | 24
hyperparathyroidism | 24
circulatory function decline | 24
respiratory function decline | 24
altered mentation | 24
ventilator support | 24
ECMO-assisted surgery | 48
elcatonin administration | 48
zoledronic acid administration | 48
evocalcet administration | 48
CHDF | 48
parathyroidectomy | 72
left thyroidectomy | 72
left recurrent laryngeal nerve resection | 72
tumour resection | 72
ECMO termination | 96
circulatory function improvement | 96
calcium levels decrease | 96
pancreatitis treatment | 96
i.v. fluids administration | 96
antibiotics administration | 96
dialysis | 96
noradrenaline administration | 96
discharged from ICU | 720
rehabilitation | 720
ventilatory support weaning | 720
respiratory muscles weakening | 720
transferred to another hospital | 720