Here is the table of events and timestamps:

14 years old | 0
male | 0
near-drowning incident | -24
trapped against a large suction intake drain | -24
loss of consciousness | -24
rescued | -24
bystander CPR | -24
hemodynamically stable | -24
fully conscious | -24
abdominal pain | -24
diffuse abrasions on torso | -24
square configuration | -24
pneumoperitoneum | -24
chest x-ray | -24
CT scan | -24
pneumomediastinum | -24
intraabdominal free fluid | -24
GE junction disruption | -24
gross contamination with food debris | -24
hemodynamically labile | -24
damage control procedure | -24
distal esophagus and proximal stomach stapled closed | -24
mediastinal drain and gastrostomy tube placed | -24
nasogastric tube placed | -24
intraabdominal and mediastinal drains placed | -24
fascia closed | -24
transferred to ICU | -24
septic shock | -24
respiratory failure | -24
prolonged intubation | -24
deep venous thrombosis | -24
pulmonary embolism | -24
bilateral pleural effusions | -24
general deconditioning | -24
parenteral nutrition started | -24
extubated | -18
fluoroscopic evaluation | -18
leak in the esophagus | -18
mediastinal drain controlled the leak | -18
enteral nutrition initiated | -18
nasogastric tube and mediastinal drain | -18
discharged | -18
Ivor-Lewis distal esophagectomy | -18
partial left lateral decubitus position | -18
midline abdominal incision | -18
gastric conduit made | -18
right thoracotomy | -18
distal esophagus identified | -18
tubularized portion of the stomach advanced into the chest | -18
esophagogastric anastomosis | -18
leak test via upper endoscopy | -18
jejunostomy tube placed | -18
extubated | -15
jejunostomy enteral feeds | -15
esophagram | -15
no leak at the anastomosis | -15
immediate stomach emptying | -15
liquid diet initiated | -15
discharged | -15
tolerates regular diet | -5
gaining weight and recovering well | -5