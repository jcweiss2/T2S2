22 years old | 0
male | 0
Afghan | 0
migrant worker | 0
admitted to the hospital | 0
dysphagia | -168
chest pain | -168
fever | -168
chills | -168
BMI 16 | 0
symptoms started | -168
worsening of symptoms | -24
emergency room visit | 0
past medical history unremarkable | 0
past surgical history unremarkable | 0
no recent upper endoscopy | 0
history of prolonged fever | -432
history of weight loss | -432
history of dealing with suspected TB patient | -432
drug history negative | 0
allergy history negative | 0
febrile | 0
tachycardic | 0
tachypneic | 0
oxygen saturation 89% | 0
chest X-ray showed left side effusion | 0
CT scan reconfirmed effusion | 0
CT scan showed left side pneumothorax | 0
CT scan showed pneumomediastinum | 0
extraluminal contrast observed | 0
distal esophageal perforation | 0
chest tube inserted | 0
purulent fluid | 0
aggressive resuscitation | 0
transferred to operating room | 0
thoracotomy | 0
large perforation in distal esophagus | 0
esophagectomy | 0
cervical esophagostomy | 0
gastrostomy | 0
transferred to surgical intensive care unit | 0
septic shock | 0
multi-organ failure | 96
passed away | 96
detection of mycobacterial DNA by PCR | 0
surgical pathology of esophagus | 0
diagnosis of mycobacterium tuberculosis | 0
granuloma | 0
exudative inflammation | 0 
TB treatment not started | 0 
TB treatment should have been started | -168 
antibiosis | 0 
isoniazid | 0
rifampin | 0
pyrazinamide | 0
ethambutol | 0
streptomycin | 0 
surgery for complications | 0 
thoracic lavage | 0
drainage | 0
esophagostomy | 0
gastrostomy | 0 
damage control surgery | 0