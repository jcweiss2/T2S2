79 years old | 0
male | 0
admitted to the hospital | 0
lower abdominal pain | -24
pyrexia | -24
pain at the peri-umbilical region | -24
pain migrated to right lower quadrant | -24
history of hypertension | 0
history of type 2 diabetes mellitus | 0
history of hyperlipidaemia | 0
recently admitted for bronchoscopy | -168
recently admitted for biopsy of a left bronchial mass | -168
diagnosed with bronchial carcinoid tumour | -168
generalized lower abdominal tenderness | 0
maximal tenderness around the periumbilical and right lower quadrant | 0
mild guarding | 0
active bowel sounds | 0
tachycardia | 0
tachypnea | 0
mild hypertension | 0
pyrexia | 0
normal oxygen saturations | 0
no acute confusion | 0
no neurological deficit | 0
raised white cell count | 0
raised neutrophils | 0
C-reactive protein within normal range | 0
CT of the abdomen and pelvis with contrast | 0
dilated tubular structure with mild fat stranding | 0
increased enhancement | 0
preliminary diagnosis of acute appendicitis | 0
laparoscopic appendectomy | 24
intact and mildly erythematous appendix resected | 24
clear ascitic fluid drained | 24
acute deterioration | 24
increasing oxygen requirements | 24
concomitant acute changes of consolidation on chest radiograph | 24
further review of CT scans | 24
fine fishbone of 1.4 cm in length | 24
microperforation at the inferior border of the 3rd segment of the duodenum | 24
formation of an abscess | 24
associated fat stranding along the right pararenal fascia | 24
exploratory laparotomy | 36
broad-spectrum intravenous antibiotics | 24
Meropenam | 24
localized retroperitoneal abscess drained | 36
10 mL of pus aspirated | 36
manual pressure applied at the presumed site of microperforation | 36
area washed out | 36
retroperitoneal drain inserted | 36
transferred to the intensive care unit | 36
feeding jejunostomy inserted | 36
enteral feeding | 36
prevent recurrence of retro-peritonitis | 36
decreasing amounts of ventilatory support | 36
oxygen saturations improved | 36
changes on chest radiograph resolved | 36
pain well controlled with analgesia | 36
stepped down to the wards | 48
antibiotics converted to oral form | 48
levofloxacin | 48
retroperitoneal drain removed | 48
regular oral feeding re-introduced | 48
discharged | 264
follow-up | 264
jejunostomy tube removed | 264
no further follow-up | 264
pathological examination of the resected appendix | 24
minimal infiltration of neutrophils | 24
excluded acute appendicitis | 24
cultures from the abscess isolated intestinal coliforms | 24
infection from a GI source | 24
oxygen desaturation secondary to pulmonary haemorrhage | 24
pulmonary haemorrhage from traumatic suctioning during anaesthesia | 24
incidental and not related to intrabdominal sepsis | 24
fishbone ingestion a week ago | -168
consumption of fish soup as a traditional remedy | -168
following recent biopsy for bronchial carcinoid tumour | -168
no awareness of fishbone ingestion | -168