76 years old | 0
female | 0
admitted to the hospital | 0
atrial fibrillation | -672
rheumatic heart disease | -672
congestive heart failure | -672
digoxin | -672
coumadin | -672
generalized malaise | -168
shortness of breath | -168
lower extremity swelling | -168
subjective fever | -168
denies chest pain | -168
denies orthopnea | -168
denies paroxysmal nocturnal dyspnea | -168
blood pressure 79/54 mmHg | 0
oral temperature 38.3°C | 0
heart rate 55 beats/min | 0
crackles up to the mid-lung fields bilaterally | 0
irregularly irregular heart rhythm | 0
2+ pitting edema up to the knees | 0
congestion in the bilateral lower lung fields | 0
cardiomegaly | 0
sodium level 126 | 0
potassium 5.2 | 0
blood urea nitrogen 33 | 0
creatinine 2.77 | 0
white blood count 4.9 | 0
INR 2.8 | 0
signs of digoxin toxicity | 0
peak troponin level 0.20 ng/mL | 0
digoxin level 3.6 ng/mL | 0
given digoxin immune fab | 0
ejection fraction 45% to 49% | 0
possible vegetation on the mitral valve | 0
severe eccentric mitral and tricuspid regurgitation | 0
mitral valve vegetation measuring 1.2×0.7 cm | 0
severe biatrial enlargement | 0
left atrium volume 101.40 mL/m2 | 0
right atrium volume 233.80 mL/m2 | 0
blood cultures positive for Pasteurella multocida | 0
ceftriaxone started | 0
head computed tomography revealed numerous chronic infarctions | 0
septic emboli | 0
owns 4 cats | -672
evaluated for multi-valve replacement surgery | 0
biopsy of the vegetation | 0
classified as high risk for surgery | 0
chose conservative treatment | 0
condition stabilized | 24
discharged to a skilled nursing facility | 24
6-week course of ceftriaxone | 24
readmitted for congestive heart failure exacerbation | 720
elected for hospice care | 720