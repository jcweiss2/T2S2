40 years old | 0
female | 0
visited the emergency department | 0
fever | -72
minor headache | -72
abdominal pain | -72
living in a postpartum care center | -504
cesarean section | -504
front of neck swollen | -264
needle aspiration | -264
thyroid gland no specific findings | -264
no relevant medical history | 0
denied family history of malignant tumors | 0
body temperature 40.6 ℃ | 0
blood pressure 100/48 mmHg | 0
heart rate 100 bpm | 0
respiratory rate 18 breaths/min | 0
no specific findings in thyroid gland | 0
no neck stiffness | 0
no tonsil hypertrophy | 0
no abdominal tenderness | 0
no abnormal breath sounds | 0
no costal spine angle tenderness | 0
no signs of infection at cesarean section site | 0
no signs of infection at thyroid fine-needle aspiration site | 0
colposcopy | 0
bicytopenia | 0
hemoglobin 14.0 g/dL | 0
platelets 133000/μL | 0
absolute neutrophil count 2512/μL | 0
total bilirubin 0.3 mg/dL | 0
aspartate transaminase 65 U/L | 0
alanine transaminase 35 U/L | 0
thyroid function test T3 65.1 ng/dL | 0
thyroid function test free T4 0.88 ng/dL | 0
urinalysis one white blood cell/high-powered field | 0
C-reactive protein 4.46 mg/dL | 0
chest radiograph normal | 0
abdominal computed tomography | 0
elevated CRP levels | 0
intermittent post-delivery abdominal pain | 0
no prominent infectious focus | 0
antipyretic drug administration | 0
fever subsided | 0
vital signs stable | 0
discharged | 96
broad-spectrum antibiotics prescription | 96
referral to infectious disease outpatient department | 96
returned to ED | 144
fever 38 ℃ | 144
blood pressure 60/30 mmHg | 144
thrombocytopenia | 144
platelets 94000/μL | 144
total bilirubin 3.1 mg/dL | 144
aspartate transaminase 202 U/L | 144
alanine transaminase 444 U/L | 144
blood urea nitrogen 42.1 mg/dL | 144
creatinine 3.35 mg/dL | 144
ferritin 3429.0 μg/L | 144
triglyceride 957 mg/dL | 144
admitted to ICU | 144
treated with broad-spectrum antibiotics | 144
treated with steroids | 144
no high-dose steroid regimen | 144
bone marrow biopsy not confirmed | 144
thrombocytopenia worsened | 168
serum ferritin increased | 168
condition rapidly deteriorated | 168
died | 168
hematochezia due to disseminated intravascular coagulation | 168
HLH diagnosis confirmed | 168
HLH etiology unclear | 168
