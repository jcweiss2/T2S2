70 years old | 0
male | 0
emergency esophageal diversion | 0
injury to the cervical esophagus | 0
spinal surgery | 0
retrosternal gastric pull-up procedure | -4320
postoperative anastomotic leakage | -4320
endoscopy | -4320
discharged with fully covered esophageal stent | -4320
local cervical infection | -3864
sepsis | -3864
transfer to tertiary university hospital | -3864
arterial hypertonus | 0
non-active smoking status | 0
ischemic stroke | 0
incomplete senso-motoric hemiparesis | 0
thyroidectomy | 0
open prostatectomy | 0
prostate cancer | 0
malnutrition | 0
systemic inflammation | 0
jugular phlegmon | 0
cervical phlegmon | 0
hemoglobin level 6.7 g/dL | 0
white blood cell count 6400 cells/μL | 0
platelet count 210 × 10³/μL |B0
creatinine level 0.76 mg/dL | 0
unremarkable liver parameters | 0
unremarkable cholestasis parameters | 0
albumin level 2.8 g/dL | 0
chest computed tomography scan | 0
endoscopy | 0
dislodged esophageal stent | 0
extraesophageal air-filled cavity | 0
extraesophageal fluid-filled cavity | 0
partially epithelialized esophageal perforation | 0
infected cavity | 0
5 cm-long stenosis of the remaining esophagus | 0
secondary injury due to dislocated cervical stent tulip | 0
calculated antibiotic treatment | 0
intensive care unit transfer | 0
stent removal | 0
pus evacuation | 0
debridement of the fistula | 0
insertion of fully covered self-expanding metal stent | 0
percutaneous jejunal feeding catheter insertion | 0
stent slippage | 0
stent position correction | 0
stent dislocation | 0
endoscopic management switch to endoscopic vacuum therapy | 0
EsoSponge system placement | 0
jugular phlegmon resolution | 336
cervical phlegmon resolution | 336
repeated endoscopic balloon dilatation | 336
persistence of broad and rigid fistula | 336
partially obliterated esophagus | 336
interdisciplinary discussion | 336
therapeutic aim redefinition | 336
profound consolidation of cervical infection | 336
salvage surgery | 336
subtotal esophageal resection | 336
reconstruction using free-jejunal graft interposition | 336
CT angiography | 336
partial sternotomy | 336
cervical esophagus resection | 336
fistula resection | 336
laparotomy | 336
jejunal segment harvesting | 336
left carotid artery as recipient vessel | 336
left jugular vein as recipient vessel | 336
graft implantation in isoperistaltic position | 336
cervical anastomosis end-to-end fashion | 336
upper mediastinal gastro-jejunostomy side-to-side fashion | 336
partial upper sternum resection | 336
sternocleidomastoid muscle flap coverage | 336
end-to-end jejunojejunostomy | 336
oral alimentation reestablishment | 336
daily speech therapy | 336
anastomotic healing confirmation | 336
transfer to rehabilitation clinic | 336
good clinical condition | 336
