42 years old | 0
female | 0
Systemic Lupus Erythematosus | 0
disease modifying drugs | 0
acute calculous cholecystitis | 0
open cholecystectomy | 0
transient leukocytosis | 0
abnormal gall bladder imaging | 0
sepsis | 72
multiorgan dysfunction | 72
catheter-related blood stream infection | 72
preoperative right subclavian CVC placement | -72
CVC removal | 72
left IJV CVC placement | 72
free flow of blood from all ports | 72
normal chest x-ray | 72
correct CVC positioning | 72
absence of pneumothorax | 72
left neck swelling | 96
fluctuant swelling | 96
non-tender swelling | 96
local hematoma | 96
left CVC removal | 96
right IJV CVC placement | 96
rapidly worsening dyspnea | 120
desaturation | 120
diminished breath sounds | 120
bilateral pleural effusion | 120
bilateral pleurocentesis | 120
milky effusion | 120
increased triglycerides | 120
bilateral chylothorax | 120
thoracic duct injury | 120
intra pleural drainage tubes | 120
underwater seals | 120
chyle drainage | 120
nil per mouth | 120
subjective improvement | 120
reduced chest tube drainage | 168
chest drain removal | 216
