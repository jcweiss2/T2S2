57 years old | 0
male | 0
right postauricular tingling | -72
discharge-like pain in the right postauricular region | -72
pain intense | -72
pain severely affected life | -72
no nausea | -72
no vomiting | -72
no cough | -72
no diarrhea | -72
no limb weakness | -72
no fever | -72
right postauricular occipital nerve distribution area acupuncture-induced hypersensitivity | 0
normal nervous system examination | 0
neutrophils 84.6% | 0
ESR 25 mm/h | 0
sodium 131.0 mmol/L | 0
normal coagulation tests | 0
normal thyroid function tests | 0
normal liver function tests | 0
normal kidney function tests | 0
normal ASO | 0
normal rapid detection of infectious diseases | 0
normal urine analysis | 0
normal stool analysis | 0
normal glycosylated hemoglobin | 0
normal serum homocysteine levels | 0
right lesser occipital nerve hypersensitive | 0
H7N9 virus PCR positive | 0
H7N9 virus positive at Beijing CDC and CNIC | 0
fever occurred afternoon of admission | 0
temperature 39.2 °C | 0
cough | 0
headache relieved after oxcarbazepine | 0
persistent moderate to high fever | 0
cough and sputum | 0
pharyngeal pain | 0
yellow phlegm with blood filaments | 0
pneumonia | 0
transferred to Respiratory Department | 18
wheezing | 18
dyspnea | 18
oxygenation decreased to 50% | 18
widely flooded bubbles in both lungs | 18
temperature 39.5 °C | 18
cyanosis of the lip | 18
spots on the trunk and lower extremities | 18
administered lysine aspirin | 18
noninvasive ventilator-assisted ventilation | 18
oxygenation increased to 80% | 18
dyspnea not improved | 18
respiratory frequency 40 breaths/min | 18
ventilator parameters adjusted | 18
administered imipenem and moxifloxacin | 18
administered oseltamivir | 18
heart rate 190 beats/min | 18.75
blood oxygen level 80% | 18.75
bilateral lung infection worsened | 18.75
propofol sedation | 18.75
tracheal intubation | 18.75
hemorrhagic secretions from oral cavity and tracheal cannula | 18.75
treated with invasive ventilator | 18.75
reduced left ventricular systolic and diastolic functions | 18.75
administered tolasemide | 18.75
administered morphine | 18.75
pH 7.08 | 19.25
PO2 60 mmHg | 19.25
PCO2 55 mmHg | 19.25
sodium bicarbonate administered | 19.25
concentrated salt supplementation | 19.25
heart rate decreased to normal | 19.25
whole body damp and cold | 19.25
administered noradrenaline | 19.25
administered vasoactive dopamine | 19.25
agitated | 19.25
sedated with propofol and midazolam | 19.25
transferred to ICU |# Table with events and timestamps extracted from the case report.
