47 years old | 0
male | 0
diabetes mellitus | -720
admitted to the hospital | 0
severe headache | -24
right-sided blindness | -24
history of COVID-19 infection | -480
COVID-19 infection confirmed by RT-PCR | -480
pulmonary symptoms | -480
intensive care unit admission | -480
drowsy | 0
oriented to person, place, and time | 0
blood pressure of 170/100 mmHg | 0
dysarthric speech | 0
right homonymous hemianopia | 0
alexia without agraphia | 0
normal systemic examinations | 0
no evidence of petechiae or purpura | 0
intraparenchymal hemorrhage | 0
edema surrounding it in the left occipital lobe | 0
string sign suggesting thrombus or stagnation in the left transverse sinus | 0
D-dimer level of 1030 | 0
platelet count of 20,000 | 0
giant platelets without any evidence of schistocytes | 0
COVID-19 RT-PCR negative | 0
hepatitis C virus (HCV) antibody negative | 0
hepatitis B virus (HBV) antibody negative | 0
human immunodeficiency virus (HIV) antibody negative | 0
received 10 units of platelets | 0
dexamethasone 8 mg three times a day | 0
platelet count increased temporarily to 49,000 | 24
bone marrow aspiration and biopsy demonstrated hypolobulated megakaryocytes | 24
intravenous immunoglobulin (IVIG) 20 g for 5 days | 24
thrombocytopenia responded dramatically after 2 days | 48
platelet count increased to 115,000 | 48
discharged | 192
follow-up | 720
platelet count was 140,000 | 720
neurological symptoms including homonymous hemianopia were improved substantially | 720
difficulties in reading | 720
cerebral venous sinus thrombosis (CVST) | 0
immune thrombocytopenic purpura (ITP) | 0
transverse sinus thrombosis | 0
hemorrhagic venous infarction | 0