53 years old | 0
male | 0
diagnosed with grade II follicular lymphoma | -672
autologous bone marrow transplant | 0
R-CVP treatment | -672
R-ICE treatment | -336
R-DA-EPOCH treatment | -168
conditioning regimen with BEAM | -24
prophylactic antimicrobial treatment with fluconazole | -24
neutropenia | 24
fever | 72
intense myalgia | 72
papular skin lesion | 72
empiric antimicrobial treatment with meropenem, vancomycin, and liposomal amphotericin | 72
skin biopsy | 96
abundant hyphae structures | 96
blood cultures identified Fusarium solani | 96
transferred to intensive care unit | 96
voriconazole treatment | 96
ophthalmologic evaluation | 96
no signs of endophthalmitis | 96
radiographic images unremarkable | 96
heavy myoglobinuria | 96
normal creatine phosphokinase | 96
worsened renal function | 96
increased blood lactate | 96
elevation of C-reactive protein and pro-calcitonin | 96
granulocyte transfusion | 120
refractory septic shock | 168
unresponsive cardiac arrest | 168
no previous history of fungal diseases | 0
no skin or nail lesion before terminal event | 0
fungal susceptibility testing | 168
resistance to fluconazole | 168
susceptibility to voriconazole and amphotericin | 168
investigation of potential source of infection | 168
cultures of tap and shower bath water negative for fungal growth | 168