18 years old | 0
male | 0
admitted to the hospital | 0
pregnancy | -37
spontaneous vaginal delivery | -37
episiotomy | -37
severe pain | -1
shortness of breath | -1
severe pain in the region of her buttocks | -1
severe pain in the region of her buttocks | -1
tachypneic | -1
oxygen saturation of 56% on room air | -1
tachycardia | -1
fever | -1
hypotensive | -1
drowsy | -1
high-flow oxygen supply | -1
noradrenaline infusion | -1
IV heparin 5000 units | -1
IV amoxicillin-clavulanate | -1
septicemic shock | -1
transferred to a tertiary hospital | -1
electively intubated | -1
severe metabolic and lactic acidosis | -1
worsening respiratory distress | -1
crystalloid | -1
persistently hypotensive | -1
adrenaline | -1
vasopressin | -1
dobutamine | -1
grossly swollen right thigh | -1
extensive blistering ecchymotic patches | -1
necrotizing fasciitis of the right thigh | -1
septicemic shock | -1
acute kidney injury | -1
rhabdomyolysis | -1
coagulopathy with thrombocytopenia | -1
ischemic hepatitis | -1
IV meropenem | -1
IV clindamycin | -1
IV vancomycin | -1
high vaginal swab for culture and sensitivity | -1
CT pulmonary angiography | -1
incidental finding of a small pulmonary embolism | -1
bedside echocardiography | -1
good contractility | -1
intravenous immunoglobulin | -1
toxin neutralization | -1
Continuous veno-venous hemofiltration (CVVH) | -1
severe lactic acidosis | -1
lactate ranging from 9.8 to 18 mmol/L | -1
grossly elevated creatinine kinase | -1
condition of the patient remained critical | -3
required 4 inotropes | -3
CVVH was continued | -3
skin lesion spread over her bilateral upper and lower limbs | -3
bluish discoloration | -3
blistering of the bilateral lower limbs | -3
bilateral lower limbs that extended to her right lower abdomen | -3
similar lesion was also noted on her right upper limb | -3
right upper limb that extended to her right elbow | -3
Gram positive cocci in chains on staining | -3
S. pyogenes | -3
blood culture taken at the district hospital | -3
positive for group A beta hemolytic streptococcus | -3
multidisciplinary discussion | -6
diagnosis of group A streptococcal toxic shock syndrome with necrotizing fasciitis | -6
IV clindamycin | -6
high dose of IV crystalline penicillin G | -6
CVVH was continued | -6
surgical intervention was not feasible | -6
skin biopsy was not performed | -6
succumbed to death | -7
cause of death | -7
septic shock with tissue necrosis and toxic shock syndrome secondary to S. pyogenes | -7