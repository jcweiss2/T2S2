44 years old | 0
male | 0
admitted to the hospital | 0
onset of mild-flu like syndrome | -72
fever | -72
chills | -72
headache | -72
myalgia | -72
cough | -72
fatigue | -72
nasopharyngeal specimen was tested for RT-PCR | -72
RT-PCR result was positive | -72
referred to emergency ward | -72
serious respiratory failure | -72
oxygen supply with cPAP | -72
chest computed tomography scan | -72
multiple bilateral ground glass opacities and consolidations | -72
denied other symptoms | -72
tobacco use or abuse | 0
drugs use or abuse | 0
diabetes mellitus type 2 | -672
obesity | -672
mild cognitive impairment | -672
psychotic disorder | -672
transferred to intensive-care unit | 0
severe deterioration of respiratory condition | 0
acute renal failure | 24
bacteric pulmonary sovrainfection | 24
antibiotic treatment | 24
complete atelectasia of left lung | 24
tracheostomy | 24
systemic sepsis | 24
urinary tract infection | 24
antibiotic therapy | 24
high blood pressure levels | 24
antihypertensive therapy | 24
stabilization of clinical conditions | 168
transferred to Rehabilitation ward | 168
normal consciousness | 168
Glasgow Coma Scale | 168
no cranial nerves abnormality | 168
upper and lower limbs strength was evaluated | 168
manual muscle testing | 168
Medical Research Council scale | 168
absent deep tendon reflexes | 168
normal plantar response | 168
no sensitivity alteration | 168
respiratory gas exchanges | 168
good balance | 168
no need for oxygen supply | 168
neurophysiological investigation | 168
axonal polineuropathy | 168
impairment of sensory and motor component | 168
absence of sural nerve sensory action potential | 168
absence of common peroneal nerve compound muscle action potential | 168
decreased tibial nerve velocity | 168
severely decreased CMAP amplitude | 168
decreased SAP amplitude for ulnar nerve | 168
Motricity Index | 168
Timed Up and Go Test | 168
Barthel Index | 168
comprehensive rehabilitation treatment | 168
respiratory and motor rehabilitation | 168
training program | 168
5 sessions per week | 168
60 minutes per session | 168
9 months duration | 168
progressive evolution and intensity | 168
physiotherapy | 168
daily standardized passive or active motion session | 168
active postural changes | 168
breathing exercises | 168
chest expansion | 168
controlled breathing | 168
diaphragmatic re-education | 168
coordination exercises | 336
trunk control | 336
recovery of standing position | 336
reconditioning of walking | 336
functional activities | 336
overground ambulatory training | 504
orthosis | 504
improvement of mobility | 720
TUG test | 720
partial improvement of motor abilities | 720
Motricity Index | 720
complete recovery for upper extremities | 720
lower extremities function remained impaired | 720
Barthel Index score | 720
overall functional abilities improved | 720
self-care activities | 720
feeding | 720
bathing | 720
mobility | 720
postural transfers | 720
ambulatory function | 720
discharged | 2160