30 years old | 0
woman | 0
presented | 0
abdominal pain | -48
nausea | -48
vomiting | -48
fever | -48
medical history of severe pulmonary hypertension | 0
bilateral pulmonary emboli | 0
right heart failure | 0
hypothyroidism | 0
systemic hypertension | 0
classified as WHO functional class III for pulmonary hypertension | 0
tenderness to palpation over the right lower quadrant | 0
no rebound | 0
leukocytosis (18.3 k/µL) | 0
left shift (82.5% neutrophils) | 0
CT scan of the abdomen and pelvis | 0
distended fluid-filled appendix | 0
small appendicoliths | 0
surrounding edema | 0
transferred to our facility | 0
higher level of care requiring cardiopulmonary evaluation | 0
optimization before possible appendectomy | 0
developed respiratory distress | 0
admitted directly to the intensive care unit | 0
right heart catheterization | 0
severe pulmonary hypertension | 0
right ventricular systolic pressure of 120 mm Hg | 0
moderate to severe tricuspid regurgitation | 0
high risk for right ventricular failure | 0
high risk for pulmonary hypertensive crisis | 0
initial aim to optimize medical condition | 0
hope to avoid operative intervention | 0
started on sildenafil | 0
intravenous epoprostenol | 0
titration goal of 20 ng/kg/min | 0
heparin infusion | 0
intravenous piperacillin/tazobactam | 0
medical management of acute appendicitis | 0
worsening leukocytosis (20.7 k/µL) | 24
fever of 39.1°C | 24
tachypnea | 24
worsening focal peritonitis | 24
initiated surgical planning | 24
severe sepsis | 24
impending shock | 24
multidisciplinary preoperative planning | 24
preparation for intraoperative venoarterial extracorporeal membrane oxygenation | 24
femoral vessel cannulation | 24
cardiovascular surgery under local anesthesia | 24
femoral artery cannulated with small sheaths | 24
femoral vein cannulated with small sheaths | 24
planned conversion to large ECMO cannulas | 24
avoid risks of ECMO cannulation | 24
planned open procedure | 24
avoid impairment of venous return | 24
careful induction of general anesthesia | 24
open appendectomy | 24
lower midline laparotomy incision below the umbilicus | 24
purulent peritoneal fluid | 24
necrotic and gangrenous appendix | 24
multiple perforations | 24
appendectomy completed | 24
abdominal cavity irrigated | 24
abdomen closed with Jackson-Pratt drain | 24
extubated | 24
transferred to the intensive care unit | 24
stable condition | 24
no need for ECMO | 24
arterial sheaths removed | 24
venous sheaths removed | 24
septic shock resolved | 24
discharged on postoperative day 18 | 432
sildenafil | 432
bumetanide | 432
macitentan | 432
intravenous epoprostenol | 432
titration goal of 30 ng/kg/min for 30 days | 432
outpatient follow-up | 432
progressing medically | 432
tolerating medication regimen | 432
no significant side effects | 432
