58 years old | 0
male | 0
Japanese | 0
admitted to the hospital | 0
lower abdominal pain | -336
loss of appetite | -336
aortic dissection | -6720
DeBakey IIIb | -6720
conservatively treated | -6720
body temperature 37.3°C | 0
left abdominal tenderness | 0
no swollen superficial lymph nodes | 0
no leg edema | 0
mild thrombocytopenia | 0
hypoalbuminemia | 0
elevated C-reactive protein | 0
elevated alkaline phosphatase | 0
elevated γ-glutamyl transferase | 0
elevated creatinine | 0
elevated fibrinogen | 0
elevated D-dimer | 0
elevated serum soluble interleukin-2 receptor | 0
elevated rheumatoid factor | 0
elevated antinuclear antibody index | 0
elevated anti-Sjögren’s-syndrome-related antigen A antibody index | 0
negative anti-Sjögren’s-syndrome-related antigen B antibody | 0
negative anti-platelet antibody | 0
normal serum β-D-glucan | 0
negative blood cultures | 0
mild proteinuria | 0
no hematuria | 0
small pleural effusion | 0
no other abnormal findings | 0
platelet count decreased | 24
ascites increased | 24
pleural effusion increased | 24
renal insufficiency progressed | 24
blood urea nitrogen 46.7 mg/dL | 24
creatinine 2.16 mg/dL | 24
bone marrow biopsy | 120
severely hypocellular marrow | 120
whole body 18-F-fluorodeoxyglucose-positron emission tomography/computed tomography scan | 264
18-F-fluorodeoxyglucose uptake by the left cervical and submandibular lymph nodes | 264
cervical lymph node biopsy | 384
pulse therapy with methylprednisolone | 384
prophylactic platelet transfusion | 384
lymph node size normal | 384
germinal centers atrophic | 384
high endothelial venules | 384
plasma cell infiltration | 384
diagnosed with TAFRO syndrome | 384
tocilizumab initiated | 504
prednisolone administered | 504
anasarca worsened | 504
renal function worsened | 504
transferred to intensive care unit | 504
ventilator | 504
continuous hemofiltration | 504
gastrointestinal bleeding | 648
methicillin-resistant Staphylococcus aureus sepsis | 648
bacterial peritonitis | 648
Stenotrophomonas maltophilia | 648
antibiotics administered | 648
gastrointestinal perforation | 1104
candidemia | 1224
elevated β-D-glucan | 1224
micafungin administered | 1224
trimethoprim-sulfamethoxazole administered | 1224
died | 1368
disseminated candidiasis | 1368
hemophagocytic lymphohistiocytosis | 1368
large amounts of pleural effusion | 1368
large amounts of ascites | 1368
Candida in blood vessels | 1368
Candida in lungs | 1368
Candida in pleura | 1368
Candida in gastrointestinal tract | 1368
Candida in peritoneum | 1368
Candida in liver | 1368
Candida in kidneys | 1368
Candida in heart | 1368
Candida in diaphragm | 1368
Candida in thyroid gland | 1368
macrophage infiltration | 1368
hemophagocytosis | 1368
ischemic small intestine | 1368
ischemic large intestine | 1368
necrotic small intestine | 1368
necrotic large intestine | 1368
no macroscopic perforation | 1368
lymph node samples normal size | 1368
no TAFRO syndrome features | 1368