55 years old | 0
male | 0
non-alcoholic steatohepatitis (NASH) cirrhosis | 0
admitted to the hospital | 0
shortness of breath | -96
fever | -96
chills | -96
denies urinary symptoms | -96
denies diarrhea | -96
denies nausea | -96
denies vomiting | -96
history of bleeding esophageal varices | -672
history of hepatic encephalopathy | -672
history of ascites | -672
hospitalized at an outside hospital | -240
fever up to 103.4 | -240
sepsis work-up | -240
negative blood cultures | -240
negative urine cultures | -240
chest x-ray | -240
sizeable right sided pleural effusion | -240
treated empirically with intravenous antibiotics | -240
discharged on ten days of oral Levofloxacin | -240
physical exam significant for fever of 102.2 | 0
mild tachypnea | 0
icteric sclera | 0
decreased breath sounds on the right lung base | 0
no crackles or rhonchi | 0
mildly distended abdomen | 0
mild right upper quadrant tenderness | 0
trace bilateral lower extremity edema | 0
leukocytosis 11.55 k/ul | 0
74% neutrophils | 0
hemoglobin 10.5 g/dl | 0
thrombocytopenia 57 k/ul | 0
INR 1.6 | 0
negative blood cultures | 0
negative urinalysis | 0
MELD-Na 23 | 0
Child-Pugh score 10 | 0
class C | 0
chest X-ray showed a large right pleural effusion | 0
no consolidation | 0
chest computed tomography (CT) | 0
large right side pleural effusion | 0
no evolving airspace disease or consolidation | 0
abdominal ultrasound | 0
small amount of ascites | 0
not amenable to paracentesis | 0
thoracentesis | 24
1100 ml of blood-tinged exudative fluid removed | 24
RBC 16000 | 24
WBC 2643 | 24
70% neutrophils | 24
serum/pleural fluid albumin gradient >1.1 g/dL | 24
fluid gram stain showed moderate polymorphonuclear white blood cells | 24
fluid culture was negative | 24
post-thoracentesis chest X-ray | 48
improvement in the right sided pleural effusion | 48
no evidence of airspace disease | 48
diagnosis of spontaneous bacterial empyema | 48
treated with intravenous ceftriaxone | 48
2 gram every 24 hours | 48
for seven days | 120
discharged in a stable condition | 168
on ciprofloxacin prophylaxis | 168
scheduled hepatology outpatient follow-up | 168