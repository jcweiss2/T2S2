55 years old | 0
male | 0
Hodgkin lymphoma | -18240
autologous peripheral blood stem cell transplantation | -1440
chemotherapy | -1440
fever | -168
dyspnea | -168
hospitalization | 0
increased serum lactate dehydrogenase | 0
increased C-reactive protein | 0
hypoxemia | 0
ground-glass opacities in bilateral lower lung fields | 0
extensive consolidation with ground-glass opacities in bilateral lung fields | 0
negative urinary pneumococcal and Legionella antigen tests | 0
no significant bacteria detected in sputum and blood cultures | 0
drug-induced lung injury | 0
methylprednisolone pulse therapy | 0
decreased CRP level | 72
improved lung involvement | 72
second steroid pulse therapy | 240
elevated CRP levels | 240
progressive bilateral diffuse extensive infiltrates | 240
tazobactam/piperacillin treatment | 240
micafungin treatment | 240
respiratory failure | 240
death | 336
Corynebacterium spp. detected in tracheal sputum culture | 240
diffuse alveolar damage | 336
extensive fibrosis | 336
no evidence of bacterial pneumonia | 336
neutrophilic infiltration in the tracheal epithelium | 336
mucosal hemorrhage | 336
acute respiratory distress syndrome | 336
ventilator-associated tracheobronchitis | 336 
vancomycin treatment considered | 240 
severe renal dysfunction | 240 
multiple organ failure | 240