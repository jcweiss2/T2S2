65 years old | 0
female | 0
diabetes mellitus | -131400
glycosylated hemoglobin 6.6% | -672
glimepiride | 0
