74 years old | 0
male | 0
non-traumatic acute subdural hematoma on the right hemisphere | -24
emergency cranial trepanation | -24
mechanical ventilation | -24
ventilator-associated pneumonia | -24
computed tomography scan | -24
soft-tissue infection of the craniotomy wound | 0
purulent secretion | 0
erythema | 0
swelling | 0
2-cm parietal area with cerebral herniation | 0
elevated intracranial pressure | 0
midline shift of 10 mm | 0
external ventricular drain implemented | 0
surgical revision | 0
old hematoma | 0
intracranial abscess formation | 0
empirical antibiotic therapy | 0
meropenem | 0
rifampicin | 0
vancomycin | 0
microbiological samples | 0
intraoperative swabs | 0
blood culture series | 0
bronchoalveolar lavage | 0
diagnosis of intracranial abscess confirmed | 0
leucocyte count 17.48/nL | 0
C-reactive protein 445.2 mg/dL | 0
fever 38.3°C | 0
septic shock | 24
