22 years old | 0
man | 0
hospitalized | 0
fatigue | -432
chest tightness | -432
shortness of breath | -432
inability to walk | -432
gradual aggravation of shortness of breath | -432
muscle weakness | -4032
chest tightness | -4032
shortness of breath | -4032
progressive shortness of breath | 0
respiratory rate 32/min | 0
SpO2 96% | 0
sinus tachycardia (pulse rate 115/min) | 0
pCO2 65 mmHg | 0
blood pressure 16.7/9.04 Kpa | 0
body temperature 36.8 °C | 0
muscle strength in extremities symmetrically reduced | 0
grade 4 muscle strength | 0
no aphasia | 0
abnormal breath sounds | 0
lactate 25 mmol/L | 0
creatinine phosphokinase-MB 385 U/L | 0
N-terminal pro-brain natriuretic peptide 1622 pg/mL | 0
white blood cell count 1.88 × 1010/L | 0
neutrophils 84.4% | 0
procalcitonin 5.6 ng/mL | 0
interleukin-6 32 pg/mL | 0
global heart enlargement | 0
mild mitral valve regurgitation | 0
mild tricuspid valve regurgitation | 0
pulmonary artery pressure 3.86 Kpa | 0
small amounts of pericardial effusion | 0
left ventricular systolic function normal | 0
enlargement of the right heart | 0
no infiltrations | 0
mitochondrial myopathy | 0
mitochondrial crisis | 0
intravenous methylprednisone | 0
intravenous immunoglobulin | 0
high-dose B vitamins | 0
coenzyme Q10 | 0
L-carnitine | 0
adenosine triphosphate | 0
fat emulsion | 0
amino acids | 0
hormones | 0
traditional Chinese medicine | 0
norepinephrine 18.2 µg/kg/min | 0
epinephrine 1 µg/kg/min | 0
lactic acid 31 mmol/L | 0
blood pressure 70/30 mmHg | 0
extracorporeal membrane oxygenation | 0
norepinephrine 10.8 µg/kg/min | 24
epinephrine 0.5 µg/kg/min | 24
lactic acid 27 mmol/L | 24
blood pressure 110/70 mmHg | 24
extracorporeal membrane oxygenation | 24
norepinephrine 3.2 µg/kg/min | 48
epinephrine 0.1 µg/kg/min | 48
lactic acid 15 mmol/L | 48
blood pressure 120/65 mmHg | 48
extracorporeal membrane oxygenation | 48
norepinephrine 1.8 µg/kg/min | 72
epinephrine 0.05 µg/kg/min | 72
lactic acid 11.5 mmol/L | 72
blood pressure 125/73 mmHg | 72
extracorporeal membrane oxygenation | 72
norepinephrine 0.16 µg/kg/min | 96
lactic acid 9.2 mmol/L | 96
blood pressure 130/75 mmHg | 96
extracorporeal membrane oxygenation | 96
norepinephrine 0.04 µg/kg/min | 120
lactic acid 6.8 mmol/L | 120
blood pressure 140/75 mmHg | 120
extracorporeal membrane oxygenation | 120
lactic acid 3.4 mmol/L | 168
blood pressure 120/73 mmHg | 168
cervical muscle paralysis | 168
respiratory muscle paralysis | 168
proximal muscle strength 0 | 168
distal muscle strength 0 | 168
myalgia | 168
cervical muscle paralysis | 240
respiratory muscle paralysis | 240
proximal muscle strength 0 | 240
distal muscle strength 1 | 240
myalgia | 240
cervical muscle paralysis | 480
respiratory muscle paralysis | 480
proximal muscle strength 0 | 480
distal muscle strength 1-2 | 480
myalgia | 480
proximal muscle strength.1-2 | 960
distal muscle strength 3 | 960
myalgia | 960
proximal muscle strength 2-3 | 1440
distal muscle strength 3-4 | 1440
proximal muscle strength 4 | 2160
distal muscle strength 5 | 2160
walk with assistance | 2160
walk independently | 4320
discharged | 4320
