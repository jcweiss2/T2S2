45 years old | 0
female | 0
admitted to the hospital | 0
end-stage heart failure | -720
cardiac cirrhosis | -720
valvular heart disease | -720
mitral valve replacement | -744
tricuspid annuloplasty | -744
ischemic kidney injury | -744
continuous renal replacement therapy | -744
cardiac arrest | -744
ventricular fibrillation | -744
venoarterial extracorporeal membrane oxygenation | -744
admitted to our institution | 0
severe biventricular dysfunction | 0
left ventricular ejection fraction less than 5% | 0
peripheral ECMO converted to central ECMO | 0
heparinization | 0
norepinephrine infusion | 0
progressive hyperbilirubinemia | 0
abdominal computed tomographic images | 0
hepatic fissure widening | 0
irregularity of hepatic contours | 0
heterogeneous enhancement of parenchyma | 0
splenomegaly | 0
moderate amount of ascites | 0
dilated inferior vena cava | 0
congestive hepatopathy | 0
tracheostomy | 0
sedated with remifentanil | 0
new atrial fibrillation | 0
ventricular response of 76 bpm | 0
plain chest X-ray | 0
cardiomegaly | 0
total atelectasis of the left lung | 0
bronchoscopic examination | 0
compression of the left main bronchus | 0
preoperative blood test results | 0
total bilirubin 47.3 mg/dl | 0
direct bilirubin 36.2 mg/dl | 0
aspartate transaminase 92 units/L | 0
alanine transaminase 51 units/L | 0
creatinine 0.91 mg/dl | 0
platelet count 34,000 /µl | 0
prothrombin time international normalized ratio 1.49 | 0
Child-Pugh class C | 0
model for end-stage liver disease score of 26 | 0
emergent CHLT | 0
general anesthesia induced | 0
midazolam | 0
etomidate | 0
atracurium | 0
mechanical ventilation | 0
hemodynamic monitoring | 0
intra-arterial | 0
central venous | 0
inferior vena cava | 0
pulmonary arterial pressures | 0
cardiac output measurements | 0
transesophageal echocardiogram | 0
sequential heart and liver transplant | 0
heart graft immersed in histidine-tryptophan-ketoglutarate solution | 0
liver graft immersed in histidine-tryptophan-ketoglutarate solution | 0
re-sternotomy | 0
left femoral vessels cannulated | 0
superior vena cava cannulated | 0
cardiopulmonary bypass established | 0
heart transplantation performed | 0
temporary pacemaker inserted | 0
liver transplantation initiated | 0
separate incision below the subcostal area | 0
full mobilization of the recipient's liver | 0
substantial hemorrhage | 0
massive volume resuscitation | 0
cardiac surgeon called for bleeding control | 0
piggyback technique applied | 0
transfusion conducted | 0
LDRBC transfused | 0
FFP transfused | 0
single-donor platelets transfused | 0
cryoprecipitate transfused | 0
protamine sulfate administered | 0
heparinization reversed | 0
anesthesia time 13 h and 15 min | 0
postoperative care | 0
dobutamine administered | 0
norepinephrine administered | 0
vasopressin administered | 0
epinephrine administered | 0
ECMO support | 0
ischemic signs in the right hand | 24
thromboembolectomy of the right radial and brachial artery | 24
ECMO removed | 96
norepinephrine infusion tapered | 720
transaminase levels normalized | 720
prothrombin time normalized | 720
bilirubin levels normalized | 720
type II respiratory failure | 720
oliguric acute kidney injury | 720
CRRT | 720
hemodialysis | 720
defective wound healing | 720
transudative ascites | 1440
right pleural effusion | 1440
abdominal computed tomography | 1440
septic shock | 1440
catheter-related infection | 1440
recent echocardiogram | 2160
normal left ventricular function | 2160
slightly reduced right ventricular systolic function | 2160
small amount of pericardial effusion | 2160
discharged | 2160