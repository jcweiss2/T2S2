23 years old | 0
male | 0
modified Fontan operation | -113208
Tausing-Bing syndrome | -113208
atrial septal defect | -113208
ventricular septal defect | -113208
pulmonary artery stenosis | -113208
right ventricular double outlet | -113208
pulmonary orifice sutured | -113208
tricuspid valve sewn closed | -113208
left auricle connected with pulmonary artery | -113208
double outlet in right ventricle | -26160
right atrial enlargement | -26160
aortic valve regurgitation | -26160
ejection fraction 50% | -26160
fever | -120
highest temperature 39.1 °C | -120
cephalosporin antibiotics | -144
chest CT scan | -96
consolidation of lower lobe right lung | -96
consolidation of superior lobe left lung | -96
arterial blood gas analysis (pH 7.476, PCO2 22 mmHg, PO2 54.1 mmHg, HCO3- 20.4 mmol/L) | -96
fraction of inspiration O2 21% | -96
influenza A antigen positive | -96
admitted to ICU | 0
temperature 38.4 °C | 0
blood pressure 86/54 mmHg | 0
respiration rate 40/min | 0
pulse rate 110/min | 0
SPO2 80% | 0
breath sounds thick | 0
moist rales | 0
arrhythmia | 0
dropped-beat pulse | 0
respiratory failure | 0
septic shock | 0
skin wet | 0
skin cold | 0
skin bluish | 0
white blood cell count 11.89 × 109/L | 0
neutrophil percentage 84.94% | 0
hemoglobin 173.10 g/L | 0
hematocrit 48.70% | 0
sodium 128.5 mmol/L | 0
creatinine 279.6 µmol/L | 0
procalcitonin 4.51 ng/mL | 0
C-reactive protein 212.9 mg/L | 0
alanine aminotransferase 48.6 U/L | 0
aspartate aminotransferase 100.4 U/L | 0
total bilirubin 26.2 µmol/L | 0
direct bilirubin 21.4 µmol/L | 0
chest X-ray | 0
Venturi mask | 0
oxygen flow 15 L/min | 0
saturation of pulse oxygen 80% | 0
difficulty breathing | 0
arterial blood gas analysis (pH 7.45, PCO2 30 mmHg, PO2 48.2 mmHg) | 0
intubated | 0
ventilator intermittent positive pressure ventilation | 0
FiO2 100% | 0
tidal volume 560 mL | 0
respiratory frequency 20/min | 0
positive end-expiratory pressure 10 cmH2O | 0
peak airway pressure 23 cmH2O | 0
moxifloxacin hydrochloride | 0
paramivir | 0
cefoperazone-sulbactam sodium | 96
vancomycin hydrochloride | 96
voriconazole | 96
central venous pressure 40 mmHg | 0
noradrenaline | 0
continuous renal replacement therapy | 0
protective lung ventilation strategy | 0
ventilation in prone position | 0
arterial blood gas analysis (pH 7.193, PCO2 48 mmHg, PO2 52 mmHg, base excess -10 mmol/L, lactate 1.34 mmol/L) | 24
venoEvenous extracorporeal membrane oxygenation (VV ECMO) | 24
left femoral vein catheter | 24
right internal jugular vein catheter | 24
rotation speed 3100 turns/min | 24
blood flow 4.3 L/min | 24
oxygen flow 4.5 L/min | 24
FiO2 100% | 24
venoEvenous-arterial extracorporeal membrane oxygenation (VVA ECMO) | 120
right femoral artery catheter | 120
left femoral vein catheter | 120
right internal jugular vein catheter | 120
rotation speed 3800 turns/min | 120
blood flow 4 L/min | 120
oxygen flow 4 L/min | 120
negative liquid equilibrium | 120
negative fluid balance 272 mL | 120
negative fluid balance 345 mL | 120
central venous pressure 28 mmHg | 120
noradrenaline dose 0.7-1.4 ug/kg/min | 120
cumulative positive balance 10000 mL | 144
central venous pressure 35 mmHg | 144
noradrenaline discontinued | 240
oxygenator and circulation line replaced | 408
tracheotomy | 528
venoEvenous-arterial ECMO removed | 648
withdrawn from artificial ventilation | 1344
discharged | 1464
follow-up on October 25, 2021 | 0
light manual labor | 0
