55 years old | 0
male | 0
presented to the ED with weakness | 0
light-headedness | 0
muscle aches | 0
non-productive cough | 0
wheeze | 0
symptoms for 5 days | -120
did not measure temperature at home | -120
frequent shivering | -120
no complaint of shortness of breath | 0
no chest pain | 0
previous ED evaluation 2 days before | -48
symptoms at previous ED visit | -48
discharged after intravenous hydration | -48
Penicillin V prescription | -48
asthma | 0
hypertension | 0
diet-controlled type 2 diabetes | 0
taking lisinopril | 0
taking hydrochlorothiazide | 0
25 pack-year smoking history | 0
quit smoking 16 years ago | -140784
family history non-contributory | 0
syncope in ED | 0
lying supine | 0
blood pressure 109/87 mmHg | 0
no pulsus paradoxus | 0
heart rate 109 bpm | 0
respiratory rate 24 bpm | 0
temperature 36.5°C | 0
oxygen saturation 100% | 0
skin mottling | 0
cyanosis of cheeks | 0
cyanosis of chest | 0
cyanosis of neck | 0
no jugular venous distension | 0
no lymphadenopathy | 0
clear lungs | 0
no distant cardiac sounds | 0
regular heart rate and rhythm | 0
normal S1/S2 | 0
no heart murmur | 0
unremarkable abdomen | 0
unremarkable extremities | 0
portable chest radiograph showed right upper lobe infiltrate | 0
borderline enlarged cardiac silhouette | 0
radiologist noted possible artifactual enlargement | 0
electrocardiogram showed sinus tachycardia | 0
no tall QRS complex | 0
electrical alternans absent | 0
white blood cell count 16.6 103/µL | 0
hemoglobin 13.4 g/dL | 0
sodium 129 mmol/L | 0
potassium 4.2 mmol/L | 0
carbon dioxide 21 mEq/L | 0
creatinine 1.0 mg/dL | 0
glucose 152 mg/dL | 0
cardiac enzymes normal | 0
B-natriuretic peptide 915 pg/mL | 0
lactic acid 3.8 mmol/L | 0
antibiotics started | 0
fluid resuscitation initiated | 0
concern for severe sepsis | 0
3 liters normal saline administered | 0
no improvement in symptoms | 0
no change in blood pressure | 0
no change in heart rate | 0
dusky mottling persisted | 0
no jugular venous distention after fluid resuscitation | 0
intensivist consulted | 0
bedside ultrasound performed | 0
pericardial effusion | 0
diastolic collapse of right atrium | 0
diastolic collapse of right ventricle | 0
normal ejection fraction | 0
suboptimal subcostal view | 0
no precise evaluation of inferior vena cava | 0
another syncopal episode | 0
decision for bedside pericardiocentesis | 0
200 mL bloody pericardial fluid drained | 0
symptoms improved | 0
cyanosis improved | 0
continued symptom free | 24
hemodynamically stable | 24
open pericardiotomy performed | 24
pericardial window placement performed | 24
repeat chest radiograph showed smaller cardiac silhouette | 24
repeat electrocardiogram showed increased QRS voltage | 24
CT scan showed pericardial drainage tube | 24
trace pericardial effusion | 24
right upper pneumonic infiltrate | 24
small bilateral pleural effusion | 24
pericardial biopsy analysis | 24
pericardial effusion fluid analysis | 24
adenocarcinoma diagnosed | 24
immune stain suggested pulmonary primary source | 24
bronchial brushing and washing suggested adenocarcinoma | 24
blood culture negative | 24
urine culture negative | 24
bronchial-alveolar washing cultures negative | 24
discharged to oncology clinic | 24
