31 years old | 0
female | 0
chronic hypertension | 0
systemic lupus erythematosus | 0
hydroxychloroquine | 0
deep venous thrombosis | 0
enoxaparin therapy | 0
presented to the emergency department | 0
heavy vaginal bleeding | 0
4-day postpartum | 0
term pregnancies | -168
postpartum transient ischemic attack | -168
preterm pregnancy | -168
severe preeclampsia | -168
spontaneous abortions | -168
ectopic pregnancy | -168
preeclampsia | -168
diagnosed by week 27 | -168
labetalol | -168
vaginal delivery at 35 weeks | -168
tachycardia | 0
hypotension | 0
fever | 0
anemia | 0
hemoglobin 6.9 g/dl | 0
thrombocytopenia | 0
34,000/μL | 0
liver function tests within normal limits | 0
fibrinogen within normal limits | 0
renal function within normal limits | 0
intravenous fluid resuscitation | 0
red blood cells transfusion | 0
platelet transfusions | 0
broad-spectrum antibiotics | 0
sepsis | 0
enoxaparin discontinued | 0
hydroxychloroquine discontinued | 0
admitted to the surgical Intensive Care Unit | 0
obstetric consultation | 0
intrauterine balloon tamponade | 0
general anesthesia | 0
vaginal bleeding ceased | 0
hemodynamics improved | 0
platelet count decreased to 17,000/μL | 72
anemia persisted | 72
red blood cells transfusions | 72
platelet transfusions | 72
schistocytes present | 72
normal haptoglobin | 72
normal bilirubin | 72
normal reticulocyte count | 72
autoimmune panel evaluation | 168
complement levels | 168
cardiolipin antibodies | 168
antinuclear antibody | 168
anti-Smith | 168
dsDNA | 168
SSA/SSB | 168
ADAMTS-13 activity | 168
ADAMTS-13 antibodies | 168
antibodies against hydroxychloroquine | 168
heparin-induced thrombocytopenia panel | 168
persistent elevated blood pressure | 168
160/100 mmHg | 168
epigastric pain | 168
acute kidney injury | 168
creatinine 2.75 mg/dL | 168
magnesium sulfate initiated | 168
worsening preeclampsia | 168
granular casts | 168
acute tubular necrosis | 168
proteinuria | 168
absent dysmorphic red blood cells | 168
adequate urine output | 168
acute aphasia | 360
altered mental status | 360
negative for stroke | 360
neurologic symptoms resolved | 360
multidisciplinary team conference | 360
initiate daily PLEX | 360
autoimmune panel unremarkable | 360
severe deficiency of ADAMTS13 activity | 360
<5% | 360
diagnosis of TTP | 360
PLEX initiated | 432
clinical improvement within 72 h | 432
thrombocytopenia refractory | 432
methylprednisolone initiated | 672
rituximab initiated | 864
vincristine initiated | 1008
platelet count improved | 1008
discharged to rehabilitation | 1008
