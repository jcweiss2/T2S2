82 years old | 0
female | 0
admitted to ICU | 0
treated arterial hypertension | -8760
septic shock | 0
heart rate at 124/min | 0
blood pressure at 80/45 mmHg | 0
polypnea at 28 cycles/min | 0
abdomen tense and painful | 0
hyperlactatemia-related metabolic acidosis | 0
pH at 7.21 | 0
PCO2 at 24 mmHg | 0
bicarbonate level at 14 mmoL/L | 0
lactate level at 9 mmoL/L | 0
liver abscess | 0
mechanical ventilation | 0
norepinephrine infusion | 0
piperacillin/tazobactam | 0
gentamicin | 0
emergency laparotomy surgery | 0
crepitation of thoracic and cervical region | 12
subcutaneous emphysema | 12
pneumoperitoneum | 12
second CT scan | 12
perforated lesion of transverse colon | 24
second emergency laparotomy | 24
colon removal | 24
colostomy | 24
multiorgan failure | 72
death | 72 
no upper airway injuries | 0
no pneumothorax | 0 
no suggestive medical history | -8760 
alveolar rupture | -8760 
barotrauma | -8760 
colonoscopy | -8760 
colonic ischemia | 12 
septic shock | 0 
liver abscess-associated septic shock | 0 
respiratory failure | 0 
hemodynamic failure | 0 
voluminous liver abscess | 0 
air–fluid level | 0 
massive subcutaneous emphysema | 12 
diffuse subcutaneous emphysema | 12 
pneumomediastinum | -8760 
tense pneumothorax | -8760 
alveolar rupture-related barotrauma | -8760 
recent laparoscopy | -8760 
colonic procedure | -8760 
abdominal CT scan | 0 
EQUATOR Network guidelines | -8760 
CARE guideline | -8760 
Institutional Review Board / Ethics Committee | -8760 
patient consent | -8760 
EQUATOR Network | -8760 
CARE | -8760 
patient's images | -8760 
patient's clinical information | -8760 
patient's name | -8760 
patient's initial | -8760 
conflicts of interest | -8760 
Financial support | -8760 
sponsorship | -8760 
Nil | -8760