47 years old | 0
female | 0
Korean | 0
schizophrenia | -8760
treated with clozapine | -8760
poor adherence to medication | -720
divorced | -720
mother passed away | -120
moved in with son | -72
drowsy and incoherent | -24
admitted to emergency department | 0
azotemia | 0
muscle enzyme elevation | 0
gross hematuria | 0
metabolic acidosis | 0
anuria | 0
rhabdomyolysis | 0
respiratory distress | 0
pulmonary edema | 0
leukocytosis | 0
high acute phase reactant | 0
sustained fever | 0
sepsis | 0
systemic antibiotics | 0
hemodialysis | 0
mechanical ventilation | 0
continuous renal replacement therapy | 24
low blood pressure | 24
inotropic agents | 24
pulmonary edema improved | 48
extubation | 96
drowsiness | 96
generalized tonic-clonic seizure | 96
brain magnetic resonance image | 96
electroencephalogram | 96
cerebrospinal fluid analysis | 96
elevated protein levels | 96
antiepileptic drug | 96
seizure-like movement subsided | 120
urine culture | 120
extended-spectrum beta-lactamase-resistant Escherichia coli | 120
urosepsis | 120
clozapine resumed | 168
leukocytosis worsened | 168
fever reappeared | 168
antipyretic drug | 168
short-term systemic steroids | 192
BCR/ABL1 rearrangement test | 192
suicidal intent | -24
clozapine overdose | -24
NMS suspected | 0
clozapine discontinued | 216
leukocytosis resolved | 216
clozapine resumed at low dose | 240
transferred to general ward | 240
delusional symptoms | 240