60 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
impaired consciousness | -1 | 0 | Factual
atrial fibrillation | -672 | 0 | Factual
dilated cardiomyopathy | -672 | 0 | Factual
oral warfarin | -672 | 0 | Factual
biventricular pacing implantable cardioverter defibrillator | -672 | 0 | Factual
found lying at home | -1 | 0 | Factual
transported to hospital | -1 | 0 | Factual
Japan Coma Scale score II-10 | 0 | 0 | Factual
Glasgow Coma Scale score 14 | 0 | 0 | Factual
no clear neurological deficits | 0 | 0 | Factual
non-contrast head CT | 0 | 0 | Factual
hemorrhage in third and fourth ventricles | 0 | 0 | Factual
hemorrhage in bilateral lateral ventricles | 0 | 0 | Factual
brain 3D-CTA | 0 | 0 | Factual
spot enhancement on lateral wall of anterior horn of left lateral ventricle | 0 | 0 | Factual
blood pressure control | 0 | 72 | Factual
ventricular drainage not performed | 0 | 0 | Negated
cerebral angiograph | 72 | 72 | Factual
aneurysm at distal site of mLSA | 72 | 72 | Factual
embolization | 72 | 72 | Factual
endovascular treatment | 72 | 72 | Factual
N-butyl-2-cyanoacrylate injection | 72 | 72 | Factual
no signs of hemorrhagic complications | 72 | 72 | Factual
no cerebral infarction | 72 | 72 | Factual
sepsis triggered by pneumonia | 120 | 240 | Factual
decrease in muscle strength | 120 | 240 | Factual
disuse | 120 | 240 | Factual
rehabilitation | 240 | 720 | Factual
discharged to home | 720 | 720 | Factual
modified Rankin Scale 1 | 720 | 720 | Factual