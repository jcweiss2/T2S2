36 years old | 0
male | 0
diabetic | 0
admitted to the hospital | 0
high-grade fever | -72
multiple swellings around joints | -72
weight loss of 10 kg | -72
septic shock | -72
recovered from septic shock | -72
fever persisted | -72
swellings did not respond to antibiotics | -72
cefaperazone/sulbactum | -72
amikacin | -72
levofloxacin | -72
sterile blood cultures | -72
proteinuria | -72
chest CT showed patchy infiltrates in lungs | -72
no cough | -72
no dyspnoea | -72
no abdominal pain | -72
granulomatosis with polyangiitis considered | -72
anti-neutrophil cytoplasmic antibody negative | -72
anti-proteinase 3 negative | -72
anti-myeloperoxidase negative | -72
rheumatoid factor negative | -72
anti-nuclear antibody negative | -72
HIV negative | -72
empirical steroids | -72
worsening of symptoms | -72
enlargement of swellings | -72
no past history of tuberculosis | -72
no recurrent infections | -72
no alcoholism | -72
no intravenous drug abuse | -72
no exposure to dust | -72
no bird droppings exposure | -72
no animal handling | -72
no agriculture work | -72
referred to Rheumatology Center | -72
cachectic | 0
bilateral knee joint contractures | 0
diffuse, multiple, tender and firm nodules | 0
deep in muscle plane above left elbow | 0
right wrist | 0
right forearm | 0
right knee | 0
ankles | 0
CT revealed mild hepatosplenomegaly | 0
multiple bilateral lung nodules | 0
musculoskeletal ultrasound showed multiple intramuscular densities | 0
fine needle aspiration from lesions | 0
inconclusive | 0
no organism detected on gram and acid fast stains | 0
high dose of insulin | 0
febrile | 0
nodules developed into abscesses | 0
vancomycin | 0
large volume of pus drained | 24
drank untreated water from a waterfall | -720
review of patient's history | 24
infective aetiology considered | 24
repeat blood culture | 24
sterile | 24
gram/acid fast/potassium hydroxide stains and culture of pus | 24
no organism | 24
melioidosis suspected | 24
discussed with microbiologist | 24
blood culture incubated in special media | 24
isolated Burkholderia pseudomallei | 24
diagnosis of melioidosis confirmed | 24
intravenous ceftazidime | 24
dramatic improvement | 168
fever subsided | 168
pyomyositis resolved | 168
nodules in lungs subsided | 168
eradication phase with oral cotrimoxazole | 168
repeat contrast CT scan of the thorax | 720
clearance of lung nodules | 720
managed diabetes with metformin | 720
physical therapy | 720
relieve contractures | 720
complete resolution of symptoms | 720
return to baseline function | 720