19 years old | 0
    male | 0
    admitted to the hospital | 0
    paraquat ingestion | -2
    suicide attempt | -2
    nausea | -2
    vomiting | -2
    hypothyroidism | 0
    levothyroxine tablets | 0
    nasogastric tube placement | 0
    gastrointestinal washing | 0
    activated charcoal administration | 0
    dithionite test positive | 0
    hemodialysis catheter implantation | 0
    hemodialysis | 0
    N-acetylcysteine administration | 0
    Vitamin C infusion | 0
    Vitamin E injection | 0
    methylprednisolone administration | 0
    pantoprazole administration | 0
    silymarin administration | 0
    chest X-ray | 0
    respiratory recovery condition | 0
    sudden worsening of respiratory condition | 504
    cervical pain | 504
    difficulty breathing | 504
    right cervical emphysema | 504
    chest X-ray | 504
    lateral neck graphy | 504
    surgical consultation | 504
    lung service consultation | 504
    air in soft tissue of neck | 504
    air in frontal area of trachea | 504
    air in mediastinum | 504
    bilateral pneumothorax | 504
    severe emphysema of neck | 504
    severe pneumomediastinum | 504
    bilateral chest tube placement | 504
    transfer to pulmonary ICU | 504
    broad-spectrum antibiotic administration | 504
    fever | 504
    pulmonary infection symptoms | 504
    sepsis | 504
    continued paraquat poisoning treatment | 504
    supportive ICU care | 504
    ALT elevation | 288
    ALT normalization | 552
    ALT increase to 691 U/L | 648
    AST elevation to 1372 U/L | 648
    BUN elevation | 96
    BUN maximum level 54.6 mg/dL | 504
    creatinine elevation | 72
    anemia | 0
    platelet decrease | 504
    INR elevation to 2.29 | 648
    death due to severe pneumomediastinum | 648
    