60 years old | 0
female | 0
newly diagnosed T2b, N1, M0 (Stage IIb) squamous cell carcinoma of the right lung | -216
surgical resection requiring pneumonectomy and mediastinal lymphadenectomy | -216
post-operative discharge on post-operative day 4 | -120
progressive dyspnea | -12
denied cough | -12
denied wheezing | -12
denied chest pain | -12
denied fevers | -12
emergency intubation by paramedics | 0
admitted to intensive care unit | 0
intubated and sedated | 0
hypotensive | 0
tachycardic | 0
healing right pneumonectomy wound site without infection | 0
right thorax dull to percussion | 0
absent right-sided breath sounds |1
cardiac point of maximal impulse shifted toward the left |0
tracheal deviation towards the left |0
normal cardiac auscultation |0
right lower extremity leg swelling |0
central venous pressure 18 cm H2O |0
elevated leukocytes (26.3 ×109/L) |0
mild normocytic anemia (hemoglobin 11.1 g/dL) |0
creatinine 1.8 mg/dL |0
mild hyperkalemia (5.8 mmol/L) |0
lactate elevated (3.7 mmol/L) |0
undetectable troponin |0
chest radiograph showing complete right hemithorax opacification |0
computed tomography pulmonary angiogram showing complete opacification of the right hemithorax |0
moderate left pleural effusion |0
no pulmonary embolus |0
transthoracic echocardiogram showing severe biatrial compression |0
no tamponade |0
no restrictive physiology |0
no pericardial effusion |0
normal right and left ventricular function |0
right distal leg deep venous thromboses |0
urgent bedside decompressive chest tube placement |0
left chest drained |0
milky white pleural fluid with elevated triglycerides (1729 mg/dL) |0
hemodynamics improved |0
off pressors |0
successfully extubated |0
diagnosis of tension chylothorax |0
lymphangiography did not identify thoracic duct leak |0
left chest tube drainage less than 500 cc/day over two days |48
clinical status improved |48
surgical exploration not indicated |48
large right chylothorax |48
pigtail catheter placed in right chest |48
right hemithorax irrigated daily with antibiotic solution |48
chylothorax secondary to mediastinal lymphadenectomy |48
left-sided chylothorax secondary to mediastinal transit of chyle |48
started on complete parenteral nutrition (CPN) |48
chest tube drainage decreased over several days |72
transitioned to medium chain triglyceride diet on hospital day 10 |240
minimal and serous chest tube fluid output on hospital day 10 |240
no increase in chest drain output |240
right pigtail catheter removed on hospital day 13 |312
left chest tube removed on hospital day 14 |336
discharged home on hospital day 17 |408
right leg deep venous thrombosis noted on admission |0
initially treated with intravenous heparin |0
developed pulmonary embolism |24
diagnosed with heparin-induced thrombocytopenia with thrombosis |24
alternative parenteral anticoagulation |24
retrievable inferior vena cava filter placed |24
discharged home on rivaroxaban |408
tolerating regular diet at four-month follow-up |2904
no evidence of recurrent chylothorax |2904
completed adjuvant chemotherapy |2904
