54 years old | 0
male | 0
nausea | -24
vomiting | -24
diarrhea | -24
abdominal pain | -24
generalized skin flushing | 0
blood pressure 60/39 mmHg | 0
heart rate 131/min | 0
temperature 37.8°C | 0
aggressive fluid resuscitation | 0
intravenous ciprofloxacin | 0
intravenous metronidazole | 0
white blood count 18.9 × 10^9/L | 0
neutrophils 17.63 × 10^9/L | 0
hemoglobin 162 g/L | 0
platelets 120 × 10^9/L | 0
creatinine 445 μmol/L | 0
estimated glomerular filtration rate (GFR) 12 mL/min | 0
metabolic acidosis | 0
pH 7.29 | 0
thickened terminal ileum | 0
distended appendix | 0
mild stranding of the surrounding fat | 0
turbid fluid retrieved from the right lower quadrant (RLQ) | 0
Gram stain | 0
culture | 0
necrotic zone at the base of the appendix | 0
appendectomy | 0
peritoneal lavage | 0
intraoperative short colonoscopy | 0
transesophageal echocardiography | 0
support with vasopressors | 0
disseminated intravascular coagulation (DIC) | 24
empirical intravenous treatment with ciprofloxacin and metronidazole | 0
oral amoxicillin/clavulanic acid | 168
flushing syndrome persisted | 0
left the ICU | 144
recovered uneventfully | 240
discharged | 240
R. ornithinolytica | 0
acute inflammation of the appendicular muscularis | 0
periappendicular inflammation of the fatty tissue | 0
no perforation | 0
no inflammation of the mucosa | 0