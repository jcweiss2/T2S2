37 years old | 0
man | 0
presented with complaint of loss of vision in the left eye | 0
COVID-19 infection | -2160
shortness of breath | -2160
difficulty in breathing | -2160
generalized weakness | -2160
fever | -2160
loss of smell | -2160
loss of taste | -2160
real-time reverse transcription-polymerase chain reaction (RT-PCR) for COVID-19 positive | -2160
admitted to the hospital | -2160
inflammatory markers ESR | -2160
CRP | -2160
D-dimers | -2160
ferritin | -2160
interleukin-6 | -2160
electrocardiogram normal | -2160
CT scan of the chest showed ground-glass opacities with reticulations in bilateral lungs | -2160
condition deteriorated | -120
shifted to ICU | -120
intubated | -120
treated with remdesivir | -120
azithromycin | -120
tocilizumab | -120
plasma transfusion | -120
recovered from pneumonia | 0
shifted to the ward | 0
sudden onset of swelling | 0
foreign body sensation | 0
drooping of upper eyelid | 0
diminution of vision of the left eye | 0
ophthalmological opinion sought | 0
no perception of light | 0
ptosis | 0
proptosis | 0
complete ophthalmoplegia | 0
fundus photography showed severe optic disc edema with cherry red spot and retinal whitening | 0
MRI brain and orbit showed CST with left diffuse pre-septal and retro>orbital edema | 0
CT venography demonstrated asymmetric bulging and filling defect of the left cavernous sinus | 0
axial images showed thickened and prominent left optic nerve sheath | 0
ESR | 0
CRP | 0
admitted | 0
managed with intravenous steroids | 0
antibiotics | 0
anticoagulant | 0
symptomatic care | 0
biopsy taken from nasal mucosa | 0
reports unremarkable | 0
no visual recovery | 168
discharged | 168
proptosis recovered | 432
ptosis recovered | 432
ophthalmoplegia recovered | 432
presented with complaints of loss of vision in the left eye | 432
unaided visual acuity of 20/20 in right eye | 432
normal color vision | 432
exodeviation of 15° on Hirschberg’s test | 432
grade four relative afferent pupillary defect | 432
anterior segment of both eyes unremarkable | 432
fundus examination revealed optic disc atrophy with gliosis | 432
macular pucker | 432
intraocular pressure 18 mm Hg in right eye | 432
intraocular pressure 16 mm Hg in left eye | 432
spectral domain optical coherence tomography showed loss of foveal contour with thinning | 432
hyper-reflective internal limiting membrane with vitreomacular traction | 432
few fluid pockets in parafoveal area | 432
visual fields examination of right eye unremarkable | 432
VEP normal in right eye | 432
VEP nearly extinguished in left eye | 432
diagnosis of CST | 432
subsequent CRAO | 432
optic neuropathy | 432
secondary to COVID-19 infection | 432
no cilioretinal sparing | 432
no fungal infection (Aspergillosis) | 432
no visual recovery noticed | 168
