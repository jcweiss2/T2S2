83 years old | 0
male | 0
osteoarthritis | -6048
extreme pain | -72
magnetic resonance imaging | -72
lesions in the medial femoral condyle cartilage | -72
left primary TKA | -1900
incapacitating knee pain | -1900
conservative therapy | -1900
warfarin | -672
paroxysmal AF | -672
smoking history | -768
cholecystectomy | -480
normal femoral, popliteal, and ankle pulses | 0
ankle brachial index | 0
echocardiography | 0
warfarin hold | -72
perioperative bridging anticoagulation therapy | -72
INR | -72
enoxaparine sodium | -72
TKA | 0
spinal anesthesia | 0
tourniquet | 0
anterior parapatellar approach | 0
total blood loss | 0
compressive dressing | 0
motor and sensory functions not checked | 0
lower limb warm | 0
pulsation of the dorsalis pedis artery intact | 0
mental state declined | 1
drowsy | 1
respiration decreased | 1
blood pressure decreased | 1
transferred to the intensive care unit | 1
CT images | 1
supportive therapy | 1
vital signs recovered | 24
unstable mental status | 24
delirium | 24
sedative | 24
restraint bands | 24
drain tube removed | 48
Hemovac drain amount decreased | 48
compressive dressing removed | 48
pulse and temperature of the lower limb not checked | 48
Cnoxane administered | 48
warfarin administered | 48
INR increased | 48
air pressure device used | 48
mechanical prophylaxis | 48
warfarin dosage same as before surgery | 72
necrosis of the foot | 48
no pulsation of the dorsalis pedis artery | 48
capillary filling of the toenail | 48
emergency lower-extremity CT angiography | 48
total occlusion of the right femoral artery | 48
angiography | 48
total embolic occlusion of the right femoral artery | 48
Fogarty thrombectomy attempted | 48
reperfusion of the popliteal and anterior and posterior tibial arteries not satisfactory | 48
no back bleeding | 48
open thrombectomy performed | 48
flow maintenance observed | 48
sepsis suspected | 96
rhabdomyolysis suspected | 96
drowsy | 96
decreased blood pressure | 96
necrosis below the knee deteriorated | 96
above-knee amputation | 408
vital signs stabilized | 408
discharged | 720
wheelchair for ambulation | 720