74 years old | 0
male | 0
referred to outpatient department | 0
intermitted fever | 0
progressive back pain |
