17 years old | 0
female | 0
admitted to the hospital | 0
fever | -504
productive cough | -504
right pleuritic chest pain | -504
respiratory rate was 28 breaths/minute | 0
blood pressure was 87/52 mm Hg | 0
heart rate was 140 beats/minute | 0
temperature was 39.5°C | 0
oxygen saturation was 96% | 0
crepitations bilaterally | 0
reduced breath sounds at the right lower hemithorax | 0
stony dullness on percussion | 0
hemoglobin was 9.0 g/dL | 0
platelet count was 386,000/μL | 0
white blood cell count was 12,140/μL | 0
coagulation profile was normal | 0
large right loculated pleural effusion | 0
chest tube inserted | 0
1.2 L of pus was drained | 0
diagnosed with right loculated empyema thoracis | 0
started on intravenous co-amoxiclav | 0
vital signs returned to normal | 48
chest tube was replaced | 48
chest tube drainage remained poor | 48
intrapleural streptokinase 250,000 units | 72
complained of palpitations | 96
sweating | 96
giddiness | 96
respiratory rate of 25 breaths/minute | 96
blood pressure of 70/50 mm Hg | 96
pulse rate of 140 beats/minute | 96
temperature of 38.3°C | 96
hemoglobin had dropped to 6.5 g/dL | 96
platelet count of 209,000/μL | 96
white cell count of 18,600/μL | 96
International Normalized Ratio was 1.5 | 96
activated partial thromboplastin time was normal | 96
right massive hemothorax | 96
thoracic surgical consult | 96
chest tube was blocked | 96
chest tube was replaced | 96
new chest tube drained 1.1 L of altered blood | 120
transfused with 7 units of packed red blood cells | 120
hemoglobin level was 9.6 g/dL post-transfusion | 168
coagulation profile normalized | 168
transferred to the cardiothoracic center | 336
underwent right lung decortications | 336