68 years old | 0
female | 0
emphysematous cystitis | 0
admitted to the hospital | 0
altered mental status | -96
unresponsive | -96
blood sugar of 498 | -96
type 2 diabetes mellitus | 0
peripheral artery disease | 0
atherosclerosis | 0
coronary artery disease | 0
mesenteric ischemia | 0
gastroparesis | 0
fibromyalgia | 0
stenting procedure | 0
vascular graft | 0
tachycardic with heart rate of 169 | 0
hypotensive to 86/45 | 0
tachypneic to 46 | 0
oxygen saturation of 92% | 0
WBC of 19.4 thous/mm³ | 0
Na 129 Meq/dL | 0
Cl 92 Meq/dL | 0
creatinine 3.63 mg/dL |+0
Co2 10 Meq/L | 0
CRP 40.2 mg/dL | 0
ESR 70 mm/hr | 0
glucose 719 mg/dL | 0
lactic acid 3.6 mmol/L | 0
turbid urine | 0
glucose >1000 | 0
WBCs 10–20 | 0
RBCs 5–10 | 0
4+ bacteria | 0
TNTC of yeast | 0
Candida glabrata infection | 0
IV micafungin initiated | 0
IV cefepime initiated | 0
DKA protocol implemented | 0
absence of ketones | 0
hyperosmolar hyperglycemic state | 0
CT abdomen and pelvis | 0
free air in extraperitoneal space | 0
extraperitoneal bladder perforation | 0
clinical instability | 0
surgical intervention deferred | 0
foley catheter placement | 0
admitted to ICU | 0
intubated | 24
extubated | 168
transferred to hospitalist service | 168
hypoxia | 192
tachypnea | 192
hypertension | 192
ABG PaO₂ in the 40s | 192
reintubated | 192
heparin initiated | 192
suspected pulmonary embolus | 192
fever | 192
intermittent tachycardia | 192
tracheostomy | 192
pressure support | 192
goals of care discussed | 528
transition to comfort care | 528
passed away | 528
multiorgan failure | 528
respiratory failure | 528
cardiac arrest | 528
