62 years old | 0
male | 0
visited hospital | 0
penetrating trauma in right chest | 0
dyspnea | 0
hemoptysis | 0
respiratory rate 23 breaths per minute | 0
oxygen saturation 90% | 0
conscious | 0
fully responsive to questions | 0
blood pressure 150/90 mm Hg | 0
heart rate 100 beats per minute | 0
no inotropic drugs | 0
hemoglobin level 12.2 g/dL | 0
partial oxygen pressure 60 mm Hg | 0
left pneumonectomy | -19008
pulmonary tuberculosis infection | -19008
foreign body in right lower lobe | 0
fracture of right seventh rib | 0
no pneumothorax | 0
no hemothorax | 0
emergent surgery | 0
general anesthesia | 0
intermittent apnea technique | 0
mini-thoracotomy | 0
adhesiolysis | 0
lung retraction | 0
identification of penetration tract | 0
no damage to major vessels | 0
no damage to hilar structure airways | 0
Duval clamps placement | 0
linear stapler placement | 0
stapler firing | 0
hemostasis | 0
airway control | 0
suture ligation | 0
metal fragment extraction | 0
chest tube indwelling | 0
wound closure | 0
surgery time 90 minutes | 0
no transfusion | 0
endotracheal tube removal | 0
recovery from general anesthesia | 0
transfer to general ward | 0
no significant complications | 0
chest tube removal | 72
discharge | 168
penetrating trauma | -1 
symptoms | -1