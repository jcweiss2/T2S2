17 days old | 0
premature | 0
female | 0
transferred to NICU | 0
failure to thrive | 0
severe metabolic derangements | 0
severe intractable diarrhea | 0
34 5/7 wk gestation | 0
African American descent | 0
vaginal delivery | 0
abnormal Penta screen | 0
meconium-stained amniotic fluid | 0
duration of rupture of membranes 5 h | 0
no polyhydramnios | 0
Apgar scores 8 | 0
Apgar scores 9 | 0
birthweight 2.445 kg | 0
length 47 cm | 0
head circumference 34 cm | 0
admitted to NICU | 0
prematurity | 0
respiratory distress | 0
maternal uncle history of gastroschisis | 0
no consanguinity | 0
intubated for surfactant administration | 0
extubated to nasal CPAP | 0
treated with ampicillin | 0
treated with gentamicin | 0
clinical sepsis | 0
started on feeds of breastmilk | -384
feeds fortified | -408
watery diarrhea | -408
down 25% from birthweight | -408
metabolic acidosis | -408
serum CO2 level 6 mmol/L | -408
acute kidney injury | -408
creatinine 3.02 mg/dL | -408
hypernatremia 157 mmol/L | -408
hyperkalemia 9.2 mmol/L | -408
hyperchloremia 128 mmol/L | -408
hyperglycemia 227 mg/dL | -408
unconjugated hyperbilirubinemia | -408
total bilirubin 15.2 mg/dL | -408
direct bilirubin 1.2 mg/dL | -408
started on phototherapy | -408
leukocytosis 25000/µL | -408
I:T ratio 0.10 | -408
made NPO | -408
electrolyte abnormalities corrected | -408
normal saline replacement | -408
sodium bicarbonate replacement | -408
stool culture positive for campylobacter antigen | -408
treated with azithromycin | -408
mother’s breastmilk positive for coagulase negative staph | -408
mother’s breastmilk positive for rare E. coli | -408
blood cultures negative | -408
started on donor expressed breast milk | -504
started on Similac Sensitive | -504
started on Alimentum | -504
relapse of profuse watery stools | -504
relapse of electrolyte derangements | -504
cessation of enteral feeds | -504
transferred to our institution | 0
work-up and management of refractory diarrhea | 0
dehydration | 0
receiving TPN with SMOFlipid | 0
sunken eyes | 0
dry skin | 0
capillary refill 4 s | 0
loose stools approximately 8/d | 0
infectious disease consult | 0
gastrointestinal consult | 0
thought to be consistent with infectious diarrhea | 0
stool studies negative | 0
full sepsis work-up negative | 0
maternal HIV testing negative | 0
GI pathogen PCR panel negative | 0
stool positive for abundant leukocytes | 0
stool positive for occult blood | 0
stool cultures negative | 0
blood cultures negative | 0
stool osmotic gap 30 mOsm/kg | 0
newborn screen positive for G6PD deficiency | 0
confirmed G6PD deficiency | 0
worsening unconjugated hyperbilirubinemia | 0
TPN-induced cholestasis | 0
continued diarrhea despite NPO | 48
suspicion of secretory diarrhea | 48
EGD performed | 48
flexible sigmoidoscopy performed | 48
duodenal biopsy normal | 48
hyponatremia | 48
hypochloremia | 48
stool sodium increased | 48
stool chloride increased | 48
urine sodium decreased | 48
urine chloride decreased | 48
started on Enfalyte | 72
advanced to Elecare | 72
relapse of severe diarrhea | 120
congenital secretory diarrhea genetic panel returned | 456
MYO5B c.1462del mutation | 456
diagnosed with MIVD | 456
supportive IV nutritional support | 456
correction of electrolyte imbalance | 456
transferred to bowel transplant center | 480
transferred back to our institution | 480
maintained on intravenous TPN | 480
nephrocalcinosis | 480
dehydration managed with fluids | 480
bowel transplant evaluation | 480
waiting list for bowel transplant | 480
