86 years old | 0
male | 0
admitted to the ICU | 0
chronic heart failure | -672
atrial fibrillation | -672
septic shock | 0
urinary tract infection | 0
Charlson morbidity score was 7 | 0
respiratory distress | 0
intubation for mechanical ventilation | 0
advanced care | 0
impaired level of consciousness | 0
consent from the patient's family | 0
antibiotic therapy | 0
management of mechanical ventilation | 0
recovery of physical status | 24
reduction in level of consciousness | 36
brain infarction | 36
magnetic resonance imaging | 36
poor prognosis | 36
acute panperitonitis | 48
gastrointestinal perforation | 48
conservative management | 48
oliguria | 49
renal insufficiency | 49
consultation for renal replacement therapy | 49
hemodialysis | 49
systolic blood pressure was barely maintained | 49
sepsis | 49
multiple organ failure | 49
thrombocytopenia | 49
discussion about HD | 49
decision not to practice HD | 49
explanation to the patient's family | 49
consent for NDT | 50
death | 52
family satisfaction with care | 52
NDT as end-of-life care | 0
palliative care | 0
life-sustaining support | 0
end-of-life care in ICU | 0
decision-making in ICU | 0
patient-centered medicine | 0
disease-based medicine | 0
balance between disease-based and patient-centered care | 0
palliative care plan | 0 
informed consent | 0