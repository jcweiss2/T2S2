18 years old | 0
    male | 0
    admitted to the emergency room | 0
    posterior uveitis | -720
    testicular pain | -720
    hypo-echoic lesions in testicles | -720
    massive bleeding from mouth | 0
    cardiac arrest | 0
    cardiopulmonary resuscitation | 0
    intubated | 0
    ventilated | 0
    shifted to intensive care unit | 0
    endotracheal tube drainage of bloody aspirate | 0
    nasogastric tube drainage of bloody aspirate | 0
    asphyxia from aspiration of blood | 0
    esophagogastrodudenoscopy showing coffee ground material | 0
    no active bleeding | 0
    toxicology screening negative | 0
    autoimmune profile negative | 0
    viral serology negative | 0
    Brucella serology negative | 0
    mechanically ventilated | 0
    Glasgow coma scale 7 | 0
    CT chest with contrast negative for pulmonary embolism | 0
    echocardiogram showing probable mass over tricuspid valve | 48
    IV antibiotics (vancomycin and amikacin) | 48
    antifungal (amphotericin B) | 48
    culture negative | 48
    second echocardiography | 48
    no surgical intervention | 48
    afebrile from 3rd post admission day | 72
    antibiotics discontinued after 14 days | 336
    antifungal discontinued after 14 days | 336
    CT brain revealing hypoxic brain injury | 0
    minimal cerebral edema | 0
    resolved cerebral edema | 0
    myoclonic seizures | 0
    phenytoin treatment | 0
    sodium valproate maintenance | 0
    biopsy of testicular lesions considered | 0
    no further workup for testicular lesions | 0
    recurrent oral ulcers | -336
    recurrent genital ulcers | -336
    recurrent joint pains | -336
    Pathergy test inconclusive | 336
    posterior uveitis | 336
    CT chest showing pulmonary arteriovenous malformations | 336
    left small pulmonary infarct | 336
    no thromboembolism | 336
    methylprednisolone pulse therapy | 336
    azathioprine initiated | 336
    cyclophosphamide therapy declined | 336
    steroids tapered over 6 months | 4320
    prednisolone 10 mg | 4320
    azathioprine 75 mg daily | 4320
    osteoporosis prevention medications | 4320
    extubated | 4320
    tracheostomy closed | 4320
    irreversible brain hypoxic injury | 4320
    minimal responsiveness | 4320
    no motor response in limbs | 4320
    testicular lesions resolved | 8760
    tricuspid lesion resolved | 8760
    CT chest showing resolved pulmonary aneurysms | 8760
    discharged | 8760
    home health care | 8760
    bedridden | 8760
    persistent hypoxic brain injury | 8760
    no new lesions | 8760
    no active problems | 8760
    