24 years old | 0
female | 0
Tanzanian | 0
primigravida | 0
gestational age of 26 weeks | 0
persistent abdominal pain | -744
recurrent vaginal bleeding | -744
admitted to local community hospital | -744
abdominal pain | -744
denies previous pelvic inflammatory disease | 0
denies intrauterine contraceptive device use | 0
denies pelvic surgery | 0
suspected abruptio placenta | -48
induced with oxytocin | -48
transferred to hospital | 0
severe pain | 0
pale | 0
afebrile | 0
distended abdomen | 0
uterine fundus of 30 cm | 0
generalized tenderness | 0
fetal heartbeats not detected | 0
closed cervix | 0
uneffaced cervix | 0
firm cervix | 0
posterior cervix | 0
presenting part not found | 0
live intrauterine diamniotic–dichorionic twins | 0
estimated gestational age 26 weeks | 0
enlarged cystic placentas | 0
retro-placental clots | 0
hemoglobin level 7.0g/dl | 0
blood group A | 0
Rhesus positive | 0
diagnosis of concealed abruptio placenta | 0
live twin pregnancy | 0
emergency abdominal delivery | 0
thickened peritoneum | 0
area of hematoma | 0
cystic mass | 0
normal-sized intact uterus | 0
pregnant sac | 0
thickened omentum | 0
live female twins | 0
placenta attached to ceacum and ascending colon | 0
placenta attached to posterior aspect of omentum | 0
profuse bleeding | 0
ligation of placental blood vessels | 0
placentas left in situ | 0
umbilical cords cut | 0
estimated blood loss 2000ml | 0
transfused 4 units of whole blood | 0
first twin weighed 700g | 0
second twin weighed 800g | 0
Apgar score 5 at first minute | 0
Apgar score 6 at fifth minute | 0
no congenital abnormalities | 0
admitted to neonatal intensive care unit | 0
both babies died | 168
postoperative broad spectrum antibiotics | 0
admitted to intensive care unit | 0
septicemia | 72
treated with meropenem | 72
discharged on postoperative day 14 | 336
readmitted with peritonitis | 448
repeat laparotomy | 448
attempt to remove placentas | 448
massive hemorrhage | 448
intra-abdominal packing | 448
transfused 3 units of blood | 448
abdominal packs removed | 496
no active bleeding | 496
fascial dehiscence | 528
exploration | 528
placentas easily detached | 528
no provoking bleeding | 528
discharged from clinic | 1008