55 years old | 0
male | 0
admitted to the hospital | 0
gastrointestinal bleeding | 0
weakness | 0
urinary tract infection | 0
Pseudomonas aeruginosa | 0
tacrolimus | -8760
prednisolone | -8760
azathioprine | -8760
simultaneous pancreas-kidney transplantation | -8760
diabetes type 1 | -8760
end-stage renal disease | -8760
stroke | -8760
coronary artery disease | -8760
dialysis | -10950
pancreas graft | -8760
kidney graft | -8760
arterial anastomosis | -8760
portal vein anastomosis | -8760
enteric exocrine drainage | -8760
duodeno-jejunostomy | -8760
immunosuppression | -8760
tacrolimus | -8760
mycophenolate mofetil | -8760
prednisolone | -8760
anti-thymocyte globulin | -8760
recurring hemorrhages | 0
euglycemia | 0
C-peptide 7.9 ng/ml | 0
renal allograft function impaired | 0
serum creatinine 2.1 mg/dl | 0
anti-infective therapy | 0
imipenem | 0
renal function normalized | 24
esophagogastroduodenoscopy (EGD) | 24
ulcer at the jejuno-duodenal anastomosis | 24
varicose vessels | 24
CT angiography | 48
pantoprazole therapy | 48
recurring low hemoglobin values | 72
multiple transfusions of RBCs | 72
double-balloon endoscopy | 120
colonoscopy | 120
capsule endoscopy | 120
bone marrow biopsy | 168
low peripheral leucocyte counts | 168
septic episodes | 168
immunosuppressive medication reduced | 168
hydrocortisone treatment | 168
liver function impaired | 216
elevated liver enzymes | 216
abdominal ultrasound | 216
no signs of cirrhosis | 216
hepatitis E infection | 240
high viral loads | 240
ascites | 240
CMV reactivation | 240
hemorrhagic shock | 720
EGD | 720
jejunal varices clipped | 720
adrenalin injection | 720
CT scan | 720
stenosis of the porto-caval anastomosis | 720
venous angiography | 720
balloon catheter | 720
dilatation of the stenosis | 720
partial improvement of the stenosis | 744
CT scan | 744
perfusion of the abdominal organs | 744
unremarkable | 744
erythrocyte transfusions | 744
low hemoglobin levels | 744
surgical intervention | 936
end-to-side anastomosis | 936
splenic vein | 936
right iliac vein | 936
pancreatectomy | 936
segmental jejunal re-section | 936
no complications | 936
chronic inflammation | 936
tortuous collateral vessels | 936
bleeding stopped | 936
transfusing more than 70 units of RBCs | 936
follow-up | 10920
no more blood products needed | 10920
patient’s health improved | 10920
hepatitis E infection no longer detected | 10920
CMV reactivation treated | 10920
CD4 T cell count recovered | 10920
immunosuppressive therapy restarted | 10920
tacrolimus | 10920
prednisolone | 10920
donor-specific human leukocyte antigen-antibodies | 10920
single-antigen bead assay | 10920
discharged | 12960
good health | 12960
kidney function good | 12960
follow-up | 15552
good health | 15552
kidney function good | 15552