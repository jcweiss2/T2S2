76 years old | 0
male | 0
married | 0
farmer | 0
rural background | 0
admitted to ER | 0
non-healing wound | -168
fell from a tree | -168
wound on posterior part of left thigh | -168
ulcerated suppurative wound | 0
wound explored | 0
wound debrided | 0
wound dressed | 0
tetanus toxoid given | 0
wound swab sent for culture and sensitivity | 0
discharged on oral Flucloxacillin | 0
discharged on Metronidazole | 0
discharged on analgesics | 0
follow up in outpatient department | 0
sought help at local medical center | -24
wound cleaned | -24
analgesics given | -24
temporary relief of pain | -24
pain returned | -12
swelling | -12
purulent discharge | -12
presented to ER again | -12
increasing white blood cell count | -12
pus cells in urine | -12
discharged home on Ofloxacin | -12
presented to ER with slurring of speech | 0
disoriented | 0
board-like abdominal rigidity | 0
muscle spasms | 0
risus sardonicus | 0
symptoms induced by minor stimuli | 0
bilateral plantar reflexes down going | 0
jaw reflex increased | 0
admitted to ICU | 0
started on IVIG | 0
antibiotics upgraded to Tazobactam-Piperacillin | 0
antibiotics upgraded to Vancomycin | 0
antibiotics upgraded to Metronidazole | 0
lumbar puncture impossible | 0
non-contrast CT head normal | 0
electively intubated | 0
sedated with fentanyl | 0
sedated with midazolam | 0
started on Vecuronium | 0
blood culture sent | 0
blood culture returned with Clostridium tetani | 12
renal function deteriorated | 24
underwent hemodialysis | 24
hemoglobin dropped | 24
received packed red cells | 24
family counseled about course of illness | 24
left ICU against medical advice | 192
succumbed to disease | 216