Here is the table of events and timestamps:

age | 0
sex | 0
breast cancer | -672
chemotherapy | -672
radiation to the chest | -672
severe aortic stenosis | -672
coronary artery disease | -672
90% occlusion of the left anterior descending artery | -672
tissue aortic valve replacement | 0
saphenous vein graft bypass to the left anterior descending artery | 0
induction of anesthesia | 0
intubation | 0
dissection of the left internal mammary artery | 0
use of the greater saphenous vein | 0
decline in cerebral head saturations | 0
use of vasopressors | 0
extubation | 2
persistent lactic acidosis | 0
high-dose vasopressor support | 0
mixed cardiogenic and vasoplegic shock | 0
lethargic | 15
leftward gaze | 15
right upper extremity weakness | 15
symptoms resolved | 30
bilateral tongue ecchymoses | 15
tongue numbness | 15
dysgeusia | 15
CT scan of the head | 15
CT angiogram of the brain and neck | 15
mild calcification at the bifurcation of the right common carotid artery | 15
50% focal stenosis of the distal left common carotid artery | 15
completely occluded right lingual artery | 15
mild distal collateral flow | 15
multifocal irregularities of the left lingual artery | 15
normal postoperative platelet count | 15
normal prothrombin time | 15
normal international normalized ratio | 15
normal fibrinogen | 15
no prior history of known vasculitic disease | 15
ADAMTS13 inhibitor screen returned normal | 15
volume resuscitation | 15
low-dose epinephrine | 15
norepinephrine and vasopressin | 15
persistent high-dose requirement of vasopressors | 15
systemic vascular resistance improved | 48
serial examinations of the patient’s tongue | 15
evaluation with multiple flexible bronchoscopes | 15
persistent tongue numbness and dysgeusia | 15
supportive therapy | 15
examination and symptoms gradually improved | 15
tongue sensation and taste returned to baseline | 672