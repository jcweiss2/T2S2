93 years old | 0
    male | 0
    admitted to the hospital | 0
    syncopal episode | 0
    coronary heart disease | -1296
    percutaneous coronary intervention | -1296
    stent implantation | -1296
    left anterior descending artery | -1296
    dual antiplatelet therapy | -1296
    aspirin | -1296
    clopidogrel | -1296
    atrioventricular pacemaker implantation | -120960
    2:1 atrioventricular block | -120960
    ventricular pacemaker lead replacement | -120960
    LBB pacing lead implantation | -120960
    blood pressure 112/68 mm Hg | 0
    heart rate 60 beats/min | 0
    normal pacemaker function | 0
    atrial stimulation | 0
    ventricular stimulation | 0
    DDD mode | 0
    chest radiography no abnormalities | 0
    normal cardiac marker levels | 0
    ejection fraction 63% | 0
    255 episodes of ventricular noise reversion | 0
    ventricular oversensing | 0
    asystole periods | 0
    ventricular lead change | 0
    RV lead extraction | 0
    LBB pacing lead placement | 0
    arterial hypertension | 0
    severe fall in blood pressure | 0
    pallor | 0
    hypoperfusion | 0
    shock | 0
    atrial sensing | 0
    ventricular-paced rhythm | 0
    selective LBB capture | 0
    inverted T waves | 0
    reduced left ventricular function | 0
    ejection fraction 15% | 0
    apical dyskinesis | 0
    hyperkinesia of basal segments | 0
    LVOT obstruction | 0
    intraventricular pressure gradient 83 mm Hg | 0
    moderate-to-severe mitral regurgitation | 0
    normal coronary arteries | 0
    apical ballooning | 0
    basal hyperkinesia | 0
    intra-aortic balloon pump | 0
    cardiogenic shock | 0
    inotropes avoided | 0
    gradual reduction in LVOT obstruction | 48
    inotropes started | 48
    improved hemodynamics | 120
    IABP removed | 120
    complete resolution of LVOT obstruction | 120
    LV function recovered | 504
    ejection fraction 50% | 504
    regression of inverted T waves | 504
    prolonged mechanical ventilation | 504
    septic shock | 840
    ventilation-associated pneumonia | 840
    death | 840
    