80 years old | 0
male | 0
severe dementia | 0
status post poliomyelitis | 0
prior alcohol overconsumption | 0
epilepsy | 0
chronic urinary catheter | 0
admitted to the Emergency Room | 0
left groin and scrotal infection | 0
12 h history of fever | -12
increasing drowsiness | -12
6 h without passing of urine | -6
missing urinary catheter | 0
multiple prior ER visits | -672
cutting or removing the catheter | -672
urethral stricture | -216
unable to replace catheter | -216
passed urine spontaneously | -216
evaluated urine production | -216
drowsy | 0
blood pressure 90/57 mmHg | 0
pulse 102/min | 0
respiratory rate 21/min | 0
oxygen saturation 95% | 0
afebrile | 0
paracetamol given | -12
swollen, red and tender left groin, scrotum and perineum | 0
no signs of gangrene | 0
lower abdominal pain | 0
no peritonitis | 0
normal rectal examination | 0
residual urinary volume 580 mL | 0
serum creatinine 2.0 mg/dL | 0
CRP 360 mg/L | 0
serum lactate 5.3 mM | 0
white blood cell count 14,000 cells per μl | 0
obstruction in the urethra | 0
12 French suprapubic catheter | 0
blood and urine cultures secured | 0
piperacillin-tazobactam 4 g every 8 h initiated | 0
CT-scan | 0
no hernia | 0
no signs of gas in the tissues | 0
limit care | 0
exclude from intensive care | 0
no operation room | 0
intravenous antimicrobials and fluid treatment | 0
inflamed area examined | 0
borders marked with a pen | 0
systolic blood pressure fluctuated | 24
pulse normalized | 24
no fever | 24
general condition improved | 24
inflamed area did not expand or darken | 24
blood cultures negative | 48
ultrasound showed abscess | 48
abscess 2.5 × 5 × 4 cm | 48
general condition deteriorated | 72
CRP increased to 523 mg/L | 72
admitted for surgical drainage | 72
metronidazole 1.5 g given | 72
surgery with scrotal incision | 96
pus removed | 96
necrotic area removed | 96
left testicle removed | 96
incision extended | 96
necrotic material removed | 96
cultures obtained | 96
perineal urethra exposed | 96
necrotic material cleared | 96
perioperative iatrogenic hole in the urethra sutured | 96
rectoscopy normal | 96
cranial part of wound closed | 96
lower part of wound left open | 96
tissue cultures grew A. urinae | 96
antimicrobial sensitivity results | 96
piperacillin-tazobactam treatment continued | 96
per oral treatment initiated | 216
ciprofloxacin 500 mg twice daily | 216
clindamycin 300 mg three times daily | 216
wound care in the ward | 216
wound closed | 288
cavity with no remnant signs of infection | 288
discharged | 360