45 years old | 0
    male | 0
    admitted to the hospital | 0
    lizard (GOH) bite | -48
    severe pain | -48
    marked swelling of the right leg | -48
    decreased urine output | -48
    conscious | 0
    Glasgow coma scale (E4V5M6) | 0
    stable vitals | 0
    respiratory distress | 24
    respiratory rate (RR) of 34–36/min | 24
    oxygen saturation 85%–90% | 24
    PaO2 64.1 mmHg | 24
    FiO2 0.4 | 24
    PCO2 22.7 mm Hg | 24
    pH 7.29 | 24
    bicarbonate17.2 mmol/L | 24
    BE (−) 15.4 | 24
    invasive mechanical ventilation | 24
    total urine output ≈350 ml over last 24 h | 24
    tea coloured urine | 24
    extensive cellulitis of right leg | 0
    marked oedema extending up to the lower abdomen | 0
    two big hemorrhagic bullae on dorsal aspect of right lower leg | 0
    many smaller bullae on dorsal aspect of foot | 0
    Doppler study ruled out compartment syndrome | 24
    neutrophil leucocytosis | 24
    intravascular haemolysis | 24
    acute kidney injury (AKI) | 24
    intravenous (IV) antibiotics (tigecycline, metronidazole) | 24
    normal saline infusion | 24
    frusemide 40 mg IV | 24
    oliguria | 24
    reddish brown urine | 24
    3+ protein in urine | 24
    urine pH 6 | 24
    positive for blood in urine | 24
    20–25 red blood cells/high-power field | 24
    2–5 white blood cells/high-power field | 24
    AKI due to rhabdomyolysis | 24
    serum creatinine kinase 5340 U/L | 24
    serum myoglobin >500 ng/ml | 24
    haemodialysis initiated | 168
    urine output <30 ml | 168
    deteriorating renal profile | 168
    general condition improved | 168
    weaned off ventilator | 168
    creatine kinase (CK) levels decreasing trend | 168
    serum myoglobin decreasing trend | 168
    creatine kinase (CK) levels returned to normal | 312
    serum myoglobin returned to normal | 312
    15 haemodialysis sessions | 360
    urine output improved to 2 ml/kg/h | 360
    enteral renal formula nutrition | 360
    oral renal diet | 360
    shifted to ward | 432
    discharged from hospital | 504
    
    
    <|eot_id|>
    
  