6 years old | 0
    girl | 0
    admitted to pediatric intensive care unit | 0
    acute hypoxic respiratory failure | -216
    septic shock | -216
    suspected pneumonia | -216
    chest radiograph on admission | 0
    diffuse bilateral interstitial opacities | 0
    acute respiratory distress syndrome | 0
    non-invasive positive pressure ventilation | 0
    tracheal intubation | 6
    empiric broad spectrum antibiotics | 0
    sedation | 0
    initial ventilator settings | 0
    tidal volume 200ml | 0
    respiratory rate 30 | 0
    PEEP 6 cmH2O | 0
    FiO2 1.0 | 0
    mean airway pressure 21 cmH2O | 0
    peak inspiratory pressure 32 cmH2O | 0
    oxygenation index 19.3 | 0
    PaO2:FiO2 ratio 102.3 | 0
    severe PARDS | 0
    arterial blood gas analysis | 0
    pH 7.27 | 0
    PaCO2 49 | 0
    PaO2 87 | 0
    base deficit 4.8 | 0
    prone positioning | 0
    paralysis | 0
    worsening chest x-ray | 0
    transthoracic echocardiogram | 0
    normal LV shortening fraction 54.9% | 0
    no pulmonary hypertension | 0
    esophageal balloon catheter placement | 0
    transpulmonary pressure measurement | 0
    PEEP titration | 0
    tidal volume titration | 0
    PL ≤ 10 cmH2O | 0
    PLexp 0 ± 2 cmH2O | 0
    neuromuscular blockade discontinued | 72
    PEEP weaning | 72
    esophageal balloon removed | 103
    extubated | 155
    weaned off respiratory support | 155
    <|eot_id|>
    