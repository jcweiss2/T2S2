33 years old | 0
woman | 0
admitted to our center for left hemithyroidectomy | 0
papillary thyroid carcinoma | 0
epilepsy | 0
taking medication | 0
laparoscopic distal gastrectomy | -17520
stomach cancer | -17520
preoperative laboratory findings unremarkable | -24
preoperative ultrasonogram | -24
7-mm sized hypoechoic nodule with microcalcifications | -24
left hemithyroidectomy | 0
left central compartment neck node dissection | 0
no antibiotic prophylaxis | 0
no drain placement | 0
no intraoperative events | 0
postoperative fever | 8
pain at surgical site | 8
intravenous antipyretics | 8
postoperative day 1 nausea | 24
postoperative day 1 tachycardia | 24
high fever over 38°C | 42.5
hypotension | 42.5
tachycardia | 42.5
suspected septic shock | 42.5
admitted to surgical ICU | 42.5
empirical antibiotics | 42.5
carbapenem | 42.5
vancomycin | 42.5
massive hydration | 42.5
vasopressors | 42.5
neck CT | 42.5
chest CT | 42.5
abdomen CT | 42.5
deep neck emphysema | 42.5
focal pneumomediastinum | 42.5
infiltration in anterior neck | 42.5
mediastinum with abscess formation | 42.5
explored infected site through thyroidectomy incision | 42.5
edematous changes in entire surgical field | 42.5
no signs of esophageal perforation | 42.5
no signs of tracheal perforation | 42.5
massive irrigation | 42.5
two closed-suction drains inserted | 42.5
bedside thoracostomy | 42.5
ultrasonogram | 42.5
blood culture no bacterial growth | 42.5
wound culture no bacterial growth | 42.5
postoperative day 7 general condition stabilized | 168
postoperative day 7 vital signs stabilized | 168
transferred to general ward | 168
CT scan interval reduction in fluid collection deep neck | 168
minimal changes in mediastinum fluid collection | 168
multidisciplinary approach | 168
planned VATS for mediastinum drainage | 168
esophagogram performed | 168
gastrografin contrast media | 168
no contrast leakage | 168
deep neck infection caused by open thyroidectomy | 168
VATS day bronchospasm | 168
general anesthesia induced | 168
retransferred to surgical ICU | 168
monitoring | 168
extubated | 192
transferred to general ward | 192
empirical antibiotics continued | 192
discharged | 504
no complications | 504
infection status acceptable at 1-year follow-up | 8760
follow-up CT scans no fluid collection | 8760
