35 years old | 0
    male | 0
    fever | -360
    pain in the right thigh | -360
    pain in the right shoulder | -360
    pain progressed to the right foot | -336
    pain progressed to the left foot | -336
    pain progressed to the right index and left ring fingers | -336
    oral amoxicillin-clavulanate | -336
    paracetamol | -336
    fever persisted | -336
    limb pains persisted | -336
    admitted to a private hospital | -336
    neutrophilic leukocytosis | -336
    hyperglycemia | -336
    ultrasonography of the right mid arm | -336
    ultrasonography of the right forearm | -336
    ultrasonography of the right thigh | -336
    echogenic intramuscular collections | -336
    pyomyositis | -336
    early stage of abscess formation | -336
    aspiration of pus | -336
    Gram-negative microorganisms | -336
    intravenous antibiotics (piperacillin-tazobactam and vancomycin) | -336
    subcutaneous insulin therapy | -336
    referred to our hospital | -336
    respiratory distress | 0
    intensive care unit (ICU) admission | 0
    encephalopathy | 0
    septic shock | 0
    impending respiratory failure | 0
    diffuse swellings | 0
    warm swellings | 0
    tender swellings | 0
    APACHE II score 19 | 0
    SOFA score 6 | 0
    intubated | 0
    moderate acute respiratory distress syndrome | 0
    ventilated with lung protective ventilation strategy | 0
    vasopressor support (norepinephrine @ 0.1 mcg/kg/min) | 0
    repeat ultrasound | 0
    inflamed muscle membranes | 0
    lost fibrillary pattern of muscle | 0
    Doppler screen of limbs | 0
    no venous thrombosis | 0
    two-dimensional-echocardiogram | 0
    no infective endocarditis | 0
    empirical antimicrobials (meropenem and vancomycin) | 0
    admission blood cultures positive for B. cepacia | 0
    subsequent blood cultures positive for B. cepacia | 0
    pancytopenia | 0
    hyperferritinemia (serum ferritin 5500 ng/ml) | 0
    hypertriglyceridemia (serum triglycerides 300 mg/dl) | 0
    hepatosplenomegaly | 0
    suspicion of secondary lymphohistiocytosis | 0
    bone marrow examination | 0
    hemophagocytosis | 0
    growth of B. cepacia in bone marrow | 0
    resistance to amikacin | 0
    resistance to gentamicin | 0
    resistance to piperacillin tazobactam | 0
    sensitivity to meropenem | 0
    sensitivity to cotrimoxazole | 0
    sensitivity to levofloxacin | 0
    no granuloma | 0
    no necrosis | 0
    no fungal elements | 0
    cotrimoxazole added | 0
    shock improved | 120
    hypoxemia improved | 120
    febrile (core temperature of 40°C) | 0
    became afebrile | 240
    meropenem stopped | 168
    vancomycin stopped | 168
    cotrimoxazole continued | 168
    transferred to ward | 360
    discharged home | 360
   