50 years old | 0
    man | 0
    presented to the emergency department | 0
    progressively worsening unsteady gait | -48
    weakness | -48
    somnolence | -48
    systolic heart failure | 0
    ejection fraction of 21% | 0
    remote orthotopic liver transplantation | -2928
    alcohol-induced cirrhosis | -2928
    hepatitis C-induced cirrhosis | -2928
    acute renal failure | 0
    hemodialysis | 0
    nonadherence to tacrolimus | -2928
    nonadherence to everolimus | -2928
    creatinine of 6.1 mg/dL | 0
    blood urea nitrogen of 23 mg/dL | 0
    prothrombin time of 15.9 seconds | 0
    partial thromboplastin time of 35 seconds | 0
    international normalized ratio of 1.5 | 0
    leukocytosis of 13.4 × 10^9/L | 0
    diagnostic and therapeutic paracentesis | 0
    bloody ascitic fluid | 0
    drained 2 liters of ascitic fluid | 0
    no spontaneous bacterial peritonitis | 0
    concern for sepsis | 0
    started on vancomycin | 0
    started on piperacillin/tazobactam | 0
    hypotensive to 73/35 mm Hg | 24
    hemoglobin drop from 7.4 to 5.6 gm/dL | 24
    received 3 units of packed red blood cells | 24
    received 1 L of Ringer's lactate | 24
    received 75 g of albumin | 24
    received 1 unit of fresh frozen plasma | 24
    hemoglobin improved to 7.1 mg/dL | 24
    hemodynamics normalized | 24
    no vasopressor initiation | 24
    computed tomography of abdomen and pelvis | 24
    intraperitoneal active extravasation | 24
    right lateral abdomen extravasation | 24
    suspected injury to right inferior epigastric artery | 24
    suspected intercostal artery injury | 24
    taken to interventional radiology suite | 24
    right common femoral artery accessed | 24
    5Fr sheath placed | 24
    right 10th intercostal artery selected | 24
    right 11th intercostal artery selected | 24
    right 12th intercostal artery selected | 24
    arteriograms performed | 24
    11th intercostal artery irregularity | 24
    12th intercostal artery irregularity | 24
    embolization of right 11th intercostal artery | 24
    embolization of right 12th intercostal artery | 24
    gelatin foam slurry used | 24
    successful occlusion on completion angiogram | 24
    hemoglobin decreased to 5.6 mg/dL | 48
    repeat computed tomography | 48
    persistent arterial extravasation | 48
    required 3 units of packed red blood cells | 48
    required 1 unit of platelets | 48
    required 2 units of fresh frozen plasma | 48
    required prothrombin complex concentrate | 48
    no vasopressor initiation again | 48
    discussion of treatment options | 48
    conservative management implemented | 48
    deemed too high risk for surgery | 48
    endovascular success unlikely | 48
    Doppler ultrasound evaluation | 72
    color jet into peritoneum | 72
    vessel not traceable proximally/distally | 72
    attempted clotting-agent injection | 72
    25-gauge needle used | 72
    5000 U bovine thrombin | 72
    saline mixed with thrombin | 72
    ultrasound-guided injection | 72
    3.5 mL thrombin-saline injected | 72
    vascular jet cessation | 72
    hemoglobin stabilization | 72
    hemodynamic improvement over 72 hours | 72
    persistent leukocytosis | 72
    no systemic inflammatory response syndrome | 72
    no identified infection source | 72
    continued on vancomycin | 72
    continued on piperacillin/tazobactam | 72
    restarted on immunosuppressants | 72
    transferred to outside hospital | 72