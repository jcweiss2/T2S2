60 years old|0
    male|0
    benign prostatic hyperplasia|0
    diabetes mellitus type 2|0
    hemoglobin A1c of 7.8|0
    history of urinary tract infections|0
    presented to the emergency department|-168
    abdominal pain|-168
    gross hematuria|-168
    difficulty voiding|-168
    worsening pain|-24
    pneumaturia|-24
    acute urinary retention|-24
    tachycardic|0
    normotensive|0
    febrile to 102°F|0
    rigors|0
    abdominal guarding|0
    rebound tenderness|0
    suprapubic tenderness|0
    bedside bladder scan showed a volume of 50 cc|0
    lactic acid of 3.4 mMol/L|0
    white blood cell count of 7.9 K/μL|0
    hemoglobin of 8.9 g/dL|0
    serum sodium of 132 mEq/L|0
    creatinine of 2.27 mg/dL|0
    urinalysis demonstrated 11–50 WBC/hpf|0
    >100 RBC/hpf|0
    positive nitrates|0
    moderate leukocyte esterase|0
    upright chest x-ray|0
    concern for perforated viscus|0
    free air under the diaphragm|0
    computed tomography (CT) scan of the abdomen and pelvis|0
    extensive pneumoperitoneum|0
    emphysematous cystitis|0
    bilateral hydronephrosis|0
    emphysematous pyelitis|0
    possible abscess near the dome of the bladder|0
    high suspicion for a bowel perforation|0
    differential included enterovesical fistula|0
    possible bladder perforation|0
    general surgery consultation|0
    urology consultation|0
    intravenous fluids administered|0
    broad-spectrum antibiotics administered|0
    taken urgently to the operating room|0
    exploratory laparotomy|0
    cystoscopy|0
    significant amount of cloudy free fluid encountered|0
    sent for culture|0
    full examination of the bowel failed to identify perforation|0
    intraperitoneal portion of the bladder grossly abnormal|0
    fibrotic appearance|0
    devitalized appearance|0
    small 3–4 mm defect identified at the bladder dome|0
    large area of necrosis|0
    concurrent cystoscopy confirmed bladder perforation|0
    diffuse inflammation|0
    trabeculations|0
    diverticula|0
    partial cystectomy performed|0
    removal of a 7×5 cm segment of necrotic bladder tissue|0
    several discrete abscess pockets|0
    bladder edges debrided to healthy tissue|0
    suprapubic catheter placed|0
    urethral catheter placed|0
    bladder closed in two layers|0
    abdomen copiously irrigated|0
    transferred to the Intensive Care Unit (ICU)|0
    sepsis management|0
    lactic acidosis resolved|0
    remained hemodynamically stable|0
    discharged on postoperative day four|96
    two-week course of trimethoprim-sulfamethoxazole|96
    failed voiding trials|96
    scheduled for transurethral resection of the prostate|96
    urine cultures grew Escherichia coli|96
    intra-abdominal cultures grew Escherichia coli|96
    final pathology revealed focal transmural necrosis|96
    acute and chronic inflammation|96
    intramural abscess|96
    serositis with fibrosis|96
    
    
    60 years old|0
    male|0
    benign prostatic hyperplasia|0
    diabetes mellitus type 2|0
    hemoglobin A1c of 7.8|0
    history of urinary tract infections|0
    presented to the emergency department|-168
    abdominal pain|-168
    gross hematuria|-168
    difficulty voiding|-168
    worsening pain|-24
    pneumaturia|-24
    acute urinary retention|-24
    tachycardic|0
    normotensive|0
    febrile to 102°F|0
    rigors|0
    abdominal guarding|0
    rebound tenderness|0
    suprapubic tenderness|0
    bedside bladder scan showed a volume of 50 cc|0
    lactic acid of 3.4 mMol/L|0
    white blood cell count of 7.9 K/μL|0
    hemoglobin of 8.9 g/dL|0
    serum sodium of 132 mEq/L|0
    creatinine of 2.27 mg/dL|0
    urinalysis demonstrated 11–50 WBC/hpf|0
    >100 RBC/hpf|0
    positive nitrates|0
    moderate leukocyte esterase|0
    upright chest x-ray|0
    concern for perforated viscus|0
    free air under the diaphragm|0
    computed tomography (CT) scan of the abdomen and pelvis|0
    extensive pneumoperitoneum|0
    emphysematous cystitis|0
    bilateral hydronephrosis|0
    emphysematous pyelitis|0
    possible abscess near the dome of the bladder|0
    high suspicion for a bowel perforation|0
    differential included enterovesical fistula|0
    possible bladder perforation|0
    general surgery consultation|0
    urology consultation|0
    intravenous fluids administered|0
    broad-spectrum antibiotics administered|0
    taken urgently to the operating room|0
    exploratory laparotomy|0
    cystoscopy|0
    significant amount of cloudy free fluid encountered|0
    sent for culture|0
    full examination of the bowel failed to identify perforation|0
    intraperitoneal portion of the bladder grossly abnormal|0
    fibrotic appearance|0
    devitalized appearance|0
    small 3–4 mm defect identified at the bladder dome|0
    large area of necrosis|0
    concurrent cystoscopy confirmed bladder perforation|0
    diffuse inflammation|0
    trabeculations|0
    diverticula|0
    partial cystectomy performed|0
    removal of a 7×5 cm segment of necrotic bladder tissue|0
    several discrete abscess pockets|0
    bladder edges debrided to healthy tissue|0
    suprapubic catheter placed|0
    urethral catheter placed|0
    bladder closed in two layers|0
    abdomen copiously irrigated|0
    transferred to the Intensive Care Unit (ICU)|0
    sepsis management|0
    lactic acidosis resolved|0
    remained hemodynamically stable|0
    discharged on postoperative day four|96
    two-week course of trimethoprim-sulfamethoxazole|96
    failed voiding trials|96
    scheduled for transurethral resection of the prostate|96
    urine cultures grew Escherichia coli|96
    intra-abdominal cultures grew Escherichia coli|96
    final pathology revealed focal transmural necrosis|96
    acute and chronic inflammation|96
    intramural abscess|96
    serositis with fibrosis|96

    <|eot_id|>
