47 years old | 0  
    man | 0  
    presented to the emergency room | 0  
    pain | -336  
    massive cervical swelling | -336  
    pain started two weeks back | -336  
    oral antibiotic therapy | -336  
    swelling extended through cervical region | 0  
    evident necrotic soft tissue areas | 0  
    pus presence | 0  
    difficulty in breathing | 0  
    difficulty in swallowing | 0  
    routine examination | 0  
    laboratory tests | 0  
    no medical history | 0  
    computed tomography of neck and chest | 0  
    extensive soft tissue emphysema | 0  
    left third molar | 0  
    extraction of third molar | 0  
    drainage | 0  
    extended surgical debridement | 0  
    gauze dressing | 0  
    necrotizing fasciitis | 0  
    postoperative day 1 | 12  
    exudate decreasing | 12  
    fever | 12  
    necrotic tissue on wound margins | 12  
    second-look surgery | 12  
    more aggressive surgical debridement | 12  
    handcrafted vacuum device | 12  
    NPWT | 12  
    drainage tube connected to central negative pressure system | 12  
    negative pressure magnitude 70–100 mmHg | 12  
    changing dressing twice a day | 24  
    additional irrigation with saline solution | 24  
    calcium alginate placement | 24  
    NPWT device installed | 48  
    bacteriological examination | 0  
    antibiogram | 0  
    released from hospital | 0  
    methicillin-sensitive Staphylococcus aureus (MSSA) | 0  
    Clindamycin | 0  
    NPWT unit changed every four days | 168  
    NPWT unit changed every seven or ten days | 336  
    postoperative day 35 | 840  
    wound completely healed | 840  
    wound reduced size enterally | 840  
    healing tissue covered the injure | 840  
    no skin graft | 840  
    no reconstruction surgery | 840  
    silicone scar sheet recommended | 840  
    scar reduced | 840  
    follow-up outpatient after 18 months | 1314  
