60 years old | 0
male | 0
presented to the Emergency Department (ED) | 0
right-sided leg pain | 0
allergic to bee venom | 0
stung on the face and neck by several bees | -24
injected himself with epinephrine auto-injector | -24
anterolateral thigh | -24
no problems for the rest of the day | -24
presented to the ED reporting “the worst pain in my life” | -14
prostate cancer | 0
hypertension | 0
hypothyroidism | 0
eye surgery | 0
ankle surgery | 0
acute distress | 0
morbidly obese | 0
diaphoretic | 0
right anterolateral thigh extreme tenderness | 0
distal pulses intact | 0
skin warm | 0
blood pressure 155/83 mmHg | 0
heart rate 112 beats/min | 0
respiratory rate 16 breaths/min | 0
oxygen saturation 97% | 0
initial temperature 36.6°C | 0
temperature increased to 38.5°C | 1
weight 142.9 kg | 0
ALT 60 U/L | 0
AST 42 U/L | 0
bilirubin 1.5 mg/dL | 0
WBC 9.8 E9/L | 0
neutrophils 93.4% | 0
platelets 120 E9/L | 0
thigh not extremely erythematous | 0
thigh not warm | 0
small induration at injection site | 0
lack of findings on physical exam | 0
stable vital signs | 0
stable laboratory values | 0
ordered computed tomography (CT) scan | 0
prominent gas within anterior compartment of the right thigh | 0
vastus lateralis involvement | 0
rectus femoris involvement | 0
suggesting necrotizing fasciitis | 0
clindamycin 900 mg IV | 0
piperacillin-tazobactam (PTZ) 4.5 g IV | 0
vancomycin 2.5 g IV | 0
clindamycin initiated pre-operatively | 0
PTZ initiated pre-operatively | 0
vancomycin initiated intra-operatively | 0
surgery for right leg debridement | 1.17
anterolateral thigh incision | 1.17
muscle bulged out | 1.17
palpable crepitus | 1.17
visible crepitus | 1.17
dark malodorous liquefied muscle | 1.17
incision extended toward the greater trochanter | 1.17
incision extended toward the knee | 1.17
anterior compartment fasciotomy | 1.17
muscle bulged out confirming compartment syndrome | 1.17
vastus lateralis debrided | 1.17
rectus femoris lateral aspect debrided | 1.17
iliotibial band tendon debrided | 1.17
BUN 39 mg/dL | 24
serum creatinine 2.4 mg/dL | 24
anion gap 17 mmol/L | 24
lactic acid 3.1 mmol/L | 24
C-reactive protein 16.3 mg/dL | 24
total CK 11603 U/L | 24
ALT 61 U/L | 24
AST 180 U/L | 24
bilirubin 5.1 mg/dL | 24
WBC 23.6 E9/L | 24
neutrophils 88.7% | 24
platelets 200 E9/L | 24
acute kidney injury (AKI) | 24
metabolic acidosis secondary to AKI | 24
bicarbonate infusion initiated | 24
wound debrided again | 24
clindamycin discontinued | 24
PTZ 3.375 g IV every 8 h | 24
vancomycin continued | 24
required intermittent hemodialysis | 48
renal function continued to deteriorate | 48
urine output 20 mL | 48
subjectively feeling better | 48
afebrile | 48
hemodynamically stable | 48
no uncontrolled pain | 48
WBC 13.0 E9/L | 48
liver function tests down-trending | 48
bilirubin normalized to 1.0 mg/dL | 48
total CK 12765 U/L | 48
dressings changed wet to dry twice daily | 48
wound in good condition | 48
hyperbaric oxygen therapy initiated | 48
Clostridium perfringens identified from wound cultures | 96
vancomycin discontinued | 96
total CK 2278 U/L | 96
WBC 10.4 E9/L | 96
regaining strength in right leg | 96
moved to medical floor | 96
antibiotics changed to ertapenem 500 mg IV | 120
excisional debridement of fascia and muscle | 120
vacuum-assisted wound closure device placed | 120
tolerating oral diet | 120
debridement | 192
wound vac change | 192
tunneled dialysis catheter placement | 192
discharged | 264
acute kidney injury resolved | 864
dialysis catheter removed | 864
hyperbaric oxygen therapy completed | 864
wound healing very well | 864
able to walk “fairly decently” | 864
no significant pain | 864
