28 years old | 0
male | 0
schizophrenia | 0
admitted to the hospital | 0
impaired vigilance | -1
found in apartment | -1
8 depleted blisters of clozapine | -1
somnolent | 0
reduced Glasgow coma scale | 0
sinus tachycardia | 0
hypertension | 0
cranial computed tomography | 0
pulmonary infiltrates | 0
atelectasis | 0
pneumomediastinum | 0
soft-tissue emphysema | 0
rhabdomyolysis | 0
crush syndrome | 0
acute renal failure | 0
progressive impairment of vigilance | 1
respiratory insufficiency | 1
invasive ventilation | 1
sepsis | 10
Piperacillin/Tazobactam | 10
septic shock | 10
vasopressors | 10
hypertensive | 10
moderate tachycardia | 10
sodium nitroprusside | 10
extubated | 31
anticholinergic syndrome | 31
intravenous physostigmine | 31
drowsiness | 31
tachycardia | 31
hypertension | 31
hyposalivation | 31
physostigmine stopped | 50
follow-up CT | 144
pneumomediastinum regressed | 144
soft-tissue emphysema regressed | 144
pneumonia healed | 144
serum clozapine analysis | 96
clozapine level decreased | 96
transferred to Psychiatry Department | 144
completely awake | 144
oriented | 144
good general condition | 144
good respiratory condition | 144
regression of renal failure | 144
regression of rhabdomyolysis | 144
regression of inflammation | 144