63 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
general body malaise | -48 | 0 | Factual
diarrhea | -48 | 0 | Factual
vomiting | -48 | 0 | Factual
influenza-like symptoms | -48 | 0 | Factual
confused | 0 | 0 | Factual
splenectomy | -7744 | -7744 | Factual
idiopathic thrombocytopenic purpura | -7744 | -7744 | Factual
menometrorhagia | -7744 | -7744 | Factual
vaccinated with PPV23 | -128 | -128 | Factual
antibody response to the vaccine | -128 | -128 | Factual
fever | 0 | 0 | Factual
hypotension | 0 | 0 | Factual
bradycardia | 0 | 0 | Factual
tachypnea | 0 | 0 | Factual
decreased oxygen saturation | 0 | 0 | Factual
cyanosis of the lips and distal extremities | 0 | 0 | Factual
no sign of neck stiffness | 0 | 0 | Negated
no meningeal reactions | 0 | 0 | Negated
normal cardiac and pulmonic auscultations | 0 | 0 | Factual
soft and not tender abdomen | 0 | 0 | Factual
diagnosed with severe sepsis | 0 | 0 | Factual
volume therapy | 0 | 0 | Factual
broad-spectrum antimicrobial therapy | 0 | 0 | Factual
hydrocortisone | 0 | 0 | Factual
white blood cell count | 0 | 0 | Factual
neutrophils | 0 | 0 | Factual
hemoglobin | 0 | 0 | Factual
thrombocytes | 0 | 0 | Factual
C-reactive protein | 0 | 0 | Factual
P-lactate | 0 | 0 | Factual
aB-P-O2 | 0 | 0 | Factual
aB-P-CO2 | 0 | 0 | Factual
aB-pH | 0 | 0 | Factual
Streptococcus pneumococcal urinary antigen test | 0 | 0 | Factual
discrete pulmonic stasis | 0 | 0 | Factual
transferred to the intensive care unit | 0 | 0 | Factual
disseminated intravascular coagulation | 24 | 24 | Factual
microthrombi in the hands and feet | 24 | 24 | Factual
blood cultures showed growth of S. pneumoniae | 48 | 48 | Factual
antimicrobial treatment changed to penicillin G | 48 | 48 | Factual
suspicion of endocarditis | 72 | 72 | Factual
trans-thoracic echocardiography | 72 | 72 | Factual
modest hypokinesia of the apical part of the left ventricle | 72 | 72 | Factual
ejection fraction of 45% | 72 | 72 | Factual
endocarditis dismissed | 72 | 72 | Negated
necrosis of the fingertips and toes | 96 | 96 | Factual
renal insufficiency | 96 | 96 | Factual
hemodialysis | 96 | 96 | Factual
antibiotic therapy altered to ceftriaxone | 96 | 96 | Factual
leucocytes and CRP decreased | 96 | 96 | Factual
fever dissolved | 96 | 96 | Factual
tracheal secret for culture | 96 | 96 | Factual
culture was negative | 96 | 96 | Factual
transferred from the ICU to the medical department | 216 | 216 | Factual
antibiotics stopped | 216 | 216 | Factual
serological analysis of the pneumococcal isolate | 216 | 216 | Factual
serotype 12F | 216 | 216 | Factual
remained afebrile | 216 | 432 | Factual
fluctuating CRP | 216 | 432 | Factual
condition improved clinically | 216 | 432 | Factual
discharged | 528 | 528 | Factual
oral dicloxacillin | 528 | 538 | Factual
raised leucocytes and CRP | 528 | 528 | Factual
necrotic tissue on fingers and toes | 528 | 528 | Factual
wound cultures showed Staphylococcus aureus and haemolytic streptococci group C/G | 528 | 528 | Factual
new TTE | 528 | 528 | Factual
amputated fingers and toes | 744 | 744 | Factual
readmitted with severe sepsis | 1296 | 1296 | Factual
sepsis regimen and ceftriaxone therapy | 1296 | 1296 | Factual
transesophageal echocardiography | 1296 | 1296 | Factual
endocarditis with several moving elements on the aortic valve | 1296 | 1296 | Factual
blood cultures showed growth of S. pneumoniae | 1296 | 1296 | Factual
antimicrobial treatment altered to penicillin G | 1296 | 1296 | Factual
treated conservatively with penicillin G | 1296 | 1476 | Factual
recovered | 1476 | 1476 | Factual
antipneumococcal-12F-antibodies measured | -432 | -432 | Factual
antipneumococcal-12F-antibodies measured | 360 | 360 | Factual
antipneumococcal-12F-antibodies measured | 876 | 876 | Factual