37 years old | 0
male | 0
admitted to the hospital | 0
fever | -72
headache | -72
unilateral, painful neck swelling | -72
no significant medical history | 0
no recent international travel | 0
no known contact with anyone with COVID-19 | 0
area of redness in the posterior palate | 0
tender, non-fluctuant swelling | 0
denied cough | 0
denied neck stiffness | 0
denied pain on swallowing | 0
denied respiratory distress | 0
denied chest pain | 0
febrile at 41°C | 0
tachycardic at 115 beats per minute | 0
normotensive at 119/76 mm Hg | 0
mentally alert | 0
intermittently raised respiratory rate | 0
peripheral oxygen saturation of 100% on room air | 0
sinus tachycardia with moderately flattened T-waves on ECG | 0
unremarkable chest X-ray | 0
respiratory alkalosis | 0
elevated C reactive protein | 0
elevated procalcitonin | 0
normal leucocytes | 0
elevated troponin T | 0
elevated N-terminal pro-B-type natriuretic peptide | 0
good ventricular function on echocardiography | 0
no hypokinesia | 0
no significant valve pathology | 0
subcutaneous oedema on the left side with multiple enlarged lymph nodes on CT of the neck | 0
deterioration of the left ventricular function on echocardiography on day 2 | 48
reduced systolic function of 40% | 48
respiratory distress on day 3 | 72
transferred to intensive care | 72
broad-spectrum antibiotics cefotaxime and clindamycin | 0
acetylsalicylic acid 300 mg | 0
telemetry | 0
CT angiogram planned | 0
cardiac MRI planned | 0
nasopharyngeal swab positive for SARS-CoV-2 | 0
respiratory distress on day 3 | 72
saturating 94% on room air | 72
oxygen therapy | 72
oliguria | 72
hypotension | 72
invasive haemodynamic monitoring | 72
transpulmonary thermodilution measurements | 72
intravenous furosemide | 72
low-dose norepinephrine infusion | 72
continuous positive airway pressure | 72
bibasal consolidations on chest X-ray | 48
elevated TnT and NT-proBNP | 48
cardiac MRI showing diffuse myocardial oedema on day 5 | 120
CT angiogram showing no coronary artery stenosis | 120
discharged on day 11 | 264
readmitted with unilateral, right-sided peripheral facial nerve palsy | 168
cerebral CT scan normal | 168
spinal fluid examination showing elevated protein and IgG | 168
mild mononuclear pleocytosis | 168
empirically treated with doxycycline | 168
discharged | 168
high levels of anti-SARS-CoV-2 IgG antibodies in serum | 168
low levels of anti-SARS-CoV-2 IgG antibodies in spinal fluid | 168
antibody index indicating no definite intrathecal specific antibody production | 168
antiganglioside antibodies detected in serum | 168
cerebral MRI normal | 168
recovered from facial palsy | 168
decreased exercise tolerance | 720 
Note: The time stamps are approximate and based on the information provided in the case report. The events that occurred before admission have negative time stamps, and the events that occurred after admission have positive time stamps. The time stamps are in hours.