66 years old | 0
male | 0
admitted to the hospital | 0
COVID-19 infection | 0
hypertension | -8760
diabetes | -25560
metformin | -25560
angiotensin-converting-enzyme inhibitor | -8760
dyspnea | 0
respiratory rate 25/min | 0
oxygen saturation 83% | 0
temperature 39.7°C | 0
weight 99 kg | 0
height 1.76 cm | 0
body mass index 31.96 kg/m2 | 0
lymphopenia | 0
increased ferritin | 0
CRP | 0
LDH | 0
hypoxemia | 0
Partial Pressure of Oxygen 55 mm Hg | 0
oxygen therapy | 0
nasal cannula | 0
flow rate 7l/min | 0
SpO2% 93% | 0
intensive care unit | 0
Vitamin C | 0
Zinc | 0
corticosteroid therapy | 0
dexamethasone | 0
low-molecular-weight heparin | 0
gastric protection | 0
proton pump inhibitors | 0
difficulty in breathing | 72
SpO2 84% | 72
severe hypoxemia | 72
Partial Pressure of Oxygen 47 mm Hg | 72
contrast-enhanced chest CT | 72
pulmonary involvement more than 75% | 72
high-concentration mask | 72
flow rate 14l/min | 72
prone decubitus sessions | 72
SpO2 90% | 72
palpitations | 120
dyspnea | 120
heart rate 186 bpm | 120
blood pressure 134/80 mm Hg | 120
atrial fibrillation | 120
electrocardiogram | 120
irregular narrow-QRS complex tachycardia | 120
Amiodarone | 120
rhythm control strategy | 120
continuous infusion | 120
initial bolus | 120
heart rate slowed | 122
ventricular response 205 bpm | 122
hemodynamic instability | 122
BP 70/50 mm Hg | 122
alteration of state of consciousness | 122
Glasgow Coma Scale 8/15 | 122
external electric shock | 122
sinus rhythm restored | 122
HR 98 bpm | 122
BP 125/80 mm Hg | 122
stroke suspected | 122
cerebral MRI | 123
brainstem acute ischemic stroke | 123
National Institutes of Health Stroke Scale score 35 | 123
thrombolysis contraindicated | 123
neuro-vegetative disorders | 123
prolonged apnea | 123
extreme bradycardia | 123
tachycardia | 123
cardiac arrest | 128
refractory ventricular fibrillation | 128
resuscitation measures | 128
death | 128