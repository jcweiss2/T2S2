57 years old | 0
male | 0
admitted to the hospital | 0
diarrhea | -504
weight loss | -504
intermittent fever | -504
right loin pain | -504
intermittent abdominal pain | -504
small volume diarrhea | -504
denies fever | 0
denies vomiting | 0
denies cough | 0
denies urinary symptoms | 0
no prior comorbidities | 0
history of tuberculosis | -504
tuberculosis contact | -504
exposure to cattle or pets | -504
consumption of cooked food | -504
no food intolerance | -504
lives in rural South India | -504
walk bare footed in farm | -504
consume alcohol daily | -504
denied intravenous drug abuse | 0
denied high-risk sexual behavior | 0
not on steroids | 0
not on immunosuppressive drugs | 0
married | 0
blessed with two children | 0
family members healthy | 0
bank manager | 0
cachexia | 0
hypotension | 0
blood pressure 80/60 | 0
dry tongue | 0
sunken eyes | 0
oral candida | 0
perioral vitiligo | 0
generalized macular erythematous | 0
purpuric lesion | 0
right loin tenderness | 0
bilateral wheezes | 0
no neck stiffness | 0
cardiac examination normal | 0
provisional diagnosis of chronic diarrhea syndrome | 0
possible sepsis | 0
admitted to medical Intensive Care Unit | 0
started on ertapenem | 0
started on flucanozole | 0
neutrophilic leucocytosis | 0
low protein | 0
low albumin | 0
macrocytic anemia | 0
low mg | 0
low K | 0
low B12 | 0
low folate | 0
normal cortisol | 0
stool sent for GI pathogen multiplex PCR | 0
contrast CT of chest and abdomen | 24
ground glass opacities in lung | 24
ileocaecal thickening | 24
upper GI endoscopy | 24
biopsy | 24
antral gastritis | 24
colonoscopy | 48
biopsy | 48
small ulcers throughout colon | 48
blood grew Klebsiella pneumoniae | 0
stool routine initial sample revealed pinworms | 0
biopsy of duodenal mucosa revealed Strongyloides larval forms | 48
colonic biopsy revealed chronic colitis | 48
repeat stool for Strongyloides was positive | 72
diagnosis of Strongyloides hyperinfection | 72
started on ivermectin | 72
diarrhea settled | 96
developed encephalopathy | 96
switched to meropenem | 96
Bran imaging normal | 96
CSF done | 96
pyogenic meningitis | 96
CSF multiplex PCR revealed Klebsiella | 96
CSF culture grew Enterococcus faecium | 120
improved with meropenem and vancomycin | 120
repeat stool routine revealed persistent Strongyloides worms | 144
albendazole 400 mg twice daily added | 144
skin lesions suggestive of larva migrans | 144
autoimmune workup negative | 144
HIV 1 and 2 antibody negative | 144
CD4 1270 | 144
low IgG | 144
low IgM | 144
low IgE | 144
normal IgA | 144
no evidence of thymoma | 144
no lymph node enlargements | 144
peripheral smear did not reveal abnormal cells | 144
common variable immunodeficiency considered | 144
HTLV serology negative | 144
CD19 and CD20 negative | 144
antiendomysial antibody negative | 144
tissue transglutaminase antibody negative | 144
single dose of 400 mg/kg of IVIg given | 168
cleared stool of Strongyloides | 192
improved remarkably | 192
discharged | 240