36 years old | 0
female | 0
33-week pregnancy | 0
dry cough | -96
shortness of breath | -96
dyspnea when exerting moderate effort | -96
heart palpitations | -96
respiratory distress | -96
dyspnea progressed to orthopnea | -96
generalized malaise | -96
myalgia | -96
arthralgia | -96
tobacco consumption | -40320
suspended tobacco consumption | 0
denied use of controlled substances | 0
denied allergies | 0
denied past blood transfusions | 0
denied travel to endemic regions | 0
denied tattoos and body piercings | 0
no history of lung disease | 0
no history of asthma | 0
no chronic or degenerative diseases | 0
four pregnancies | 0
one delivery | 0
two cesarean surgeries | 0
recumbent position | 0
Glasgow coma score 15 | 0
no focal neurologic deficits | 0
no meningeal signs | 0
aware of environment | 0
diaphoretic | 0
dehydrated skin and mucosae | 0
no head and neck alterations | 0
oral ventilation | 0
tachypnea | 0
thoracic and abdominal dissociation | 0
decreased chest expansion | 0
no vibrations or fremitus | 0
no asymmetries or abnormalities on percussion | 0
bilateral crepitant crackles | 0
bilateral decreased inspiratory breath sounds | 0
tachycardia | 0
heart sounds of good intensity | 0
globous abdomen | 0
live single fetus | 0
fetal heart rate 158 bpm | 0
no visceromegaly | 0
no abdominal abnormalities | 0
filiform pulse | 0
BP 130/90 mm Hg | 0
HR 100 bpm | 0
RR 21 rpm | 0
SO2 74% | 0
temperature 36°C | 0
weight 70 kg | 0
height 165 cm | 0
BMI 25.7 | 0
type 1 respiratory insufficiency | 0
BP 130/85 mm Hg | 0
HR 120 bpm | 0
RR 36 rpm | 0
Temp 36.7°C | 0
arterial blood gas pH 7.4 | 0
PaO2 43 mm Hg | 0
PaCO2 24 mm Hg | 0
HCO3– 16.9 mEq/L | 0
O2 content 78% | 0
base excess -7.0 mmol/L | 0
lactate 0.9 mmol/L | 0
endotracheal tube | 0
emergency cesarean | 0
live newborn male 1940gr | 0
400 cc hemorrhage | 0
admitted to ICU | 0
blood cultures negative | 24
bronchial secretion culture negative | 24
Mycoplasma pneumoniae IgG negative | 24
galactomannan assay negative | 24
procalcitonin 0.02 ng/mL | 24
urinalysis abundant bacteria | 24
erythrocytes 118 per field | 24
leukocytes 163 per high power field | 24
immunoassays negative | 24
extubated | 48
adequate respiratory mechanics | 48
arterial blood gas pH 7.46 | 48
PaO2 74.9 mm Hg | 48
PaCO2 39 mm Hg | 48
HCO3– 28 mEq/L | 48
O2 content 95.6% | 48
base excess 6.0 mmol/L | 48
lactate 0.5 mmol/L | 48
dependent on supplemental oxygen | 48
admitted to Internal Medicine | 48
echocardiogram LVEF 66% | 168
mild diastolic dysfunction | 168
global pericardial effusion 300 cc | 168
no intracavitary thrombi | 168
no valvular pathology | 168
CT-guided lung biopsy | 168
invasive pulmonary adenocarcinoma | 168
lepidic growth pattern | 168
immunohistochemistry confirms diagnosis | 168
pneumothorax >25% | 168
tube thoracostomy | 168
pleural effusion exudate | 168
ECOG 4 | 336
chemotherapy contraindicated | 336
sepsis of unknown origin | 336
negative follow-up cultures | 336
declined further interventions | 336
palliative care initiated | 336
morphine administered | 336
continued orthopnea | 504
temperature 39°C | 504
leukocytosis | 504
extreme bradycardia | 720
asystole | 720
death | 720
