32 years old | 0
female | 0
admitted to neurosurgery outpatient department | 0
weakness in bilateral upper and lower limbs | -336
altered sensorium | -336
pineocytoma | -672
obstructive hydrocephalus | -672
right frontal burr hole with endoscopic third ventriculostomy and ventriculoperitoneal shunting | -4320
admitted for radiotherapy | -720
limb weakness | -720
headache | -720
vomiting | -720
generalized seizures | -48
altered sensorium | -48
difficulty in moving limbs | -48
febrile | 0
conscious | 0
Glasgow Coma Score (GCS) of 4/15 | 0
diminished deep tendon reflexes | 0
heterogeneous lesion with predominantly solid component in pineal recess–residual tumor | 0
obstructive hydrocephalus with trans ependymal CSF seepage | 0
fasting blood sugar 126 mg/dl | 0
random blood sugar 289 mg/dl | 0
shunt tapped | 0
ventricular fluid with 20 RBC/mm3 and 40 WBC/mm3 | 0
glucose of 79 mg/dl | 0
protein of 71.4 mg/dl | 0
gram-positive cocci on gram stain | 0
shunt externalized | 0
extraventricuar device placed | 0
Vitek 2 AST card used for identification and sensitivity | 0
Staphylococcus lugdunensis resistant to penicillin | 0
Staphylococcus lugdunensis susceptible to all other antibiotics tested | 0
IV vancomycin | 0
afebrile after 3 days of IV vancomycin | 72
discharged home | 240
IV oxacillin | 0
reinternalization of VPS | 240
follow-up to neurosurgery OPD | 720