68 years old | 0
female | 0
admitted to the hospital | 0
CLL/SLL | -13104
lymphocytosis | -13104
absolute lymphocyte count greater than 5000/µL | -13104
peripheral smear showing abnormal mature B cells | -13104
FCR therapy | -13104
total thyroidectomy | -4680
chronic lymphocytic thyroiditis | -4680
Hurthle cell adenoma | -4680
basal cell carcinoma | -3120
cervical lymphadenopathy | -936
Rituxan and Bendamustine therapy | -936
FISH performed on the peripheral blood | -936
mono-allelic deletion of 13q14.3 locus | -936
regression of the cervical lymphadenopathy | -936
complete remission | -936
left axillary lymphadenopathy | -120
CT imaging | -120
enlarged retroperitoneal and mesenteric lymph nodes | -120
Gazyva therapy | -120
Venetoclax | -120
clinical improvement | -24
regression of her mesenteric lymphadenopathy | -24
recurrent fever | 0
weakness | 0
abdominal pain | 0
vomiting | 0
elevated alkaline phosphatase | 0
AST 10 | 0
ALT 26 | 0
total bilirubin 1.4 | 0
serological studies negative for hepatitis A, B, and C | 0
serological studies negative for antinuclear antibody (ANA) | 0
serological studies negative for anti-smooth muscle antibody (ASMA) | 0
no duct dilatation | 0
no gallbladder thickening | 0
no peripancreatic ascites | 0
extensive splenomegaly | 0
splenic varicosities | 0
ascites | 0
porta hepatis lymphadenopathy | 0
hepatosplenomegaly | 0
enlarged intra-abdominal lymph nodes | 0
pleural effusion | 0
liver biopsy | 0
periportal fibrosis | 0
histiocytic-predominant inflammation | 0
acute granulomatous hepatitis | 0
hemophagocytosis | 0
no evidence of steatosis | 0
no evidence of cholestasis | 0
no evidence of malignancy | 0
no evidence of infectious agents | 0
peritoneal fluid showed sparse normal-appearing small lymphocytes | 0
peritoneal fluid negative for carcinoma | 0
blood transfusion | 0
consultations by gastroenterology, infectious disease, and hematology/oncology specialists | 0
treatment for neutropenic fever | 0
hypotension | 360
septic shock | 360
death | 432
autopsy | 432
diffuse lymphadenopathy | 432
multi-organ involvement | 432
Reed-Sternberg cells | 432
CD30 positive | 432
CD15 positive | 432
Pax 5 positive | 432
Bcl-2 positive | 432
EBV positive | 432
CD20 negative | 432
ALK negative | 432
CD138 negative | 432
kappa/lambda in situ hybridization negative | 432
granulomatous areas in the liver | 432
CD 68 predominant | 432
CD30/CD15 atypical Reed-Sternberg-rich area | 432
CD30/CD15 abnormal large neoplastic cells | 432
abdominal lymph nodes involvement | 432
para-aortic lymph nodes involvement | 432
mesenteric lymph nodes involvement | 432
perihilar lymph nodes involvement | 432
bilateral lungs involvement | 432
liver involvement | 432
spleen involvement | 432
pancreatic surface involvement | 432
fallopian tubes involvement | 432
bone marrow involvement | 432
Richter transformation | 432
Hodgkin lymphoma | 432
EBV-associated HL | 432
p53 expression | 432
clonal relationship between CLL cells and HL cells | 432
elevated alkaline phosphatase | 432
poor prognostic factor | 432
extranodal involvement | 432
anemia | 432
low albumin | 432
high LDH levels | 432
granulomatous liver disease | 432
elevated LDH levels | 432
noncaseating granulomatous liver disease | 432
infection | 432
autoimmune cholangitis | 432
sarcoidosis | 432
drug toxicity | 432
carcinoma | 432
lymphoma | 432
HLRT | 432
hemophagocytic lymphohistiocytosis | 432
fever | 432
splenomegaly | 432
histiocytic hemophagocytosis | 432
hypertriglyceridemia/hyperfibrinogenemia | 432
bicytopenia | 432
hyperferritinemia | 432
low NK activity | 432
high IL-2 receptor levels | 432
primary HLH | 432
secondary HLH | 432
genetic mutation | 432
abnormal cytokine production | 432
abnormal immune response | 432
treatment of underlying disease process | 432
chemotherapy | 432
EBV-associated HL | 432
fludarabine therapy | 432
Ibrutinib | 432
Venetoclax | 432
targeted therapy | 432
combination chemotherapy | 432
ABVD | 432
MOPP | 432
CVPP | 432
therapeutic transfusion | 432
bone marrow transplant | 432