74 years old | 0
    female | 0
    VATS-LA maze procedure | 0
    general anesthesia | 0
    sequential one lung ventilation | 0
    EZ-Blocker endobronchial blocker | 0
    transesophageal echocardiography (TEE) | 0
    exclusion of the LA appendage | 0
    assessment of flow in the pulmonary veins | 0
    ablation lesions created with bipolar radiofrequency catheter | 0
    no esophageal temperature probe inserted | 0
    presented to the emergency department | -1008
    persistent fever | -1008
    altered mental status | -1008
    left upper extremity weakness | -1008
    CT of the thorax | -1008
    air collected in the posterior LA | -1008
    suspicion for LA wall abscess | -1008
    suspicion for AEF | -1008
    surgical exploration through median sternotomy | -24
    cardiopulmonary bypass (CPB) on standby | -24
    intubated the night prior | -24
    worsening mental status | -24
    9F double-lumen central venous catheter inserted | -24
    poor distal circulation in both upper and lower extremities | -24
    18-G catheter inserted in the right axillary artery | -24
    blood pressure monitoring | -24
    blood sampling | -24
    EGD performed | -24
    no esophageal pathology detected | -24
    severe hypotension | -24
    treated with phenylephrine boluses | -24
    treated with norepinephrine | -24
    treated with epinephrine | -24
    TEE probe replacement | -24
    air visualized within the LA | -24
    air visualized within the left ventricle | -24
    air visualized within the aortic root | -24
    emergent median sternotomy | -24
    institution of CPB | -24
    no obvious lesion identified | -24
    NG tube placed | -24
    air injected through NG tube | -24
    fistula opening identified | -24
    defect patched with bovine pericardium | -24
    integrity of repair assessed | -24
    transferred to surgical intensive care unit | -24
    intubated | -24
    mechanically ventilated | -24
    continued neurological deterioration | 0
    MRI on POD 1 | 24
    punctate and confluent hyperintensities | 24
    hyperintensities in pons | 24
    hyperintensities in caudal midbrain | 24
    hyperintensities in posterior cerebral artery territory | 24
    hyperintensities in middle cerebral artery territories | 24
    hyperintensities in anterior cerebral artery territories | 24
    EEG on POD 3 | 72
    global slowing on EEG | 72
    global disturbance of cortical function | 72
    withdrawal of care on POD 10 | 240
    profound neurologic injury | 240
    poor prognosis | 240
    