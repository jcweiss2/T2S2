39 years old | 0
male | 0
admitted to the emergency department | 0
paraesthesia in all limbs | -48
diplopia | -48
nausea | -48
weakness in both lower and upper limbs | -24
bilateral abducens nerve paralysis | -24
facial diplegia | -24
flaccid areflexic paralysis of the limbs | -24
bowel and bladder not involved | -24
electromyography examination | -24
electromyogram confirmed acute acquired disseminated polyneuropathy syndrome | -24
cerebrospinal fluid examination | -24
elevated protein concentration | -24
normal cell count | -24
anti-ganglioside antibodies negative | -24
intravenous immune globulin administration | -24
weakness progressed rapidly | -12
respiratory muscle weakness | -12
respiratory failure | -12
mechanical ventilation | -12
intensive care unit admission | -12
plasmapheresis | -12
booster intravenous immune globulin | -12
rehabilitation | -12
oral prednisolone administration | -12
pain in both hips | 144
decreased range of motion in both hips | 144
neurogenic heterotopic ossification diagnosis | 144
plain X rays of the pelvis | 144
elevated serum calcium | 144
elevated serum alkaline phosphatase | 144
intravenous ibandronic acid administration | 144
etidronate disodium administration | 144
rehabilitative management | 144
passive and active-assistive ROM exercises | 144
breathing exercises | 144
electrotherapy | 144
discharged from ICU | 720
muscle strengths improved | 720
standing with support | 720
unable to walk or sit in low position | 720
restricted passive ROM of both hips | 720
three-phase bone scan study | 720
corticosteroid injection | 720
pain decreased | 720
increased flexion | 720
rehabilitation program continued | 1296
walking with a walker | 1296
sitting without support | 1296