27 years old | 0
pregnant | 0
G4P2 | 0
28th gestational week | 0
born in Western Africa | -3600
living in Italy | -240
headache | -48
vomiting | -48
diarrhea | -48
pelvic and low back pain | -48
admitted to the hospital | 0
ED laboratory tests | 0
lactic dehydrogenase increased | 0
mild anemia | 0
hemoglobin 9.9 g/dl | 0
renal echography | 0
no morphological abnormalities | 0
discharged | 48
returned to the hospital | 72
persistent symptoms | 72
hyperpyrexia | 72
prophylactic ceftriaxone | 72
peak hyperthermia | 96
loss of consciousness | 96
recovered | 96.25
residual aphasia | 96
cognitive impairment | 96
no rigor nucalis | 96
no focal deficit | 96
head computed tomography scan | 96
no pathological abnormalities | 96
respiratory parameters stable | 96
hemodynamic parameters stable | 96
SpO2 99% | 96
blood pressure 135/70 mmHg | 96
heart rate 95 bpm | 96
C-reactive protein increased | 96
bilirubin increased | 96
lactic dehydrogenase increased | 96
hemoglobin 7.8 g/dl | 96
malaria parasites found | 96
quinine prescribed | 96
clindamycin prescribed | 96
fetal parasitemia suspected | 96
hemolysis suspected | 96
cesarean delivery planned | 96
lactated Ringer's solution administered | 96
ranitidine administered | 96
spinal anesthesia performed | 96
hyperbaric bupivacaine injected | 96
sufentanil injected | 96
surgery initiated | 96
blood pressure decreased | 96
blood pressure stable | 96
baby born | 96
Apgar score 8 | 96
oxytocin administered | 96
postoperative analgesia | 96
patient-controlled analgesia pump | 96
morphine administered | 96
acetaminophen prescribed | 96
surgery uncomplicated | 96
blood loss estimated | 96
Plasmodium falciparum identified | 100
blood parasites decreased | 120
antibiotic therapy continued | 120
symptoms resolved | 120
oxygen therapy discontinued | 120
blood samples drawn from baby | 120
no parasites found | 120
no fetal hemolysis | 120
discharged | 168