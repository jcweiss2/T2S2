78 years old | 0
female | 0
admitted to the hospital | 0
hypertension | -672
hyperlipidemia | -672
renal calculi | -672
trichlormethiazide | -672
warfarin potassium | -672
fluvastatin sodium | -672
re-fabrication of the upper and lower partial dentures | -672
initial examination | -672
lower partial dentures re-fabricated | -336
upper partial dentures re-fabrication planned | -336
intense instability in the upper left molar region | -168
tooth mobility level 3 | -168
marked alveolar bone resorption | -168
spontaneous pain in the upper left molar region | -120
swelling in the upper left molar region | -120
pus discharge from the periodontal pocket | -120
area cleaned and sterilized | -120
loprofen sodium prescribed | -120
swelling spread to the left buccal region | -96
spontaneous pain became more intense | -96
difficulty eating | -96
primary care physician instructed the patient to visit the hospital | -48
Glasgow Coma Scale score 11 | 0
facial pallor | 0
cold hands and fingers | 0
shivering | 0
weak radial artery pulse | 0
axillary temperature 41°C | 0
systolic blood pressure 80-90 mmHg | 0
diastolic blood pressure 40-50 mmHg | 0
pulse rate 130-160 bpm | 0
SpO2 75-85% | 0
oxygen administration at 10 L/min | 0
venous line secured | 0
drip infusion of acetate linger solution | 0
drip infusion of normal saline solution | 0
ampicillin sodium administered | 0
blood examination | 0
malnutrition suspected | 0
severe infection suspected | 0
consciousness level 14 on the Glasgow Coma Scale | 12
axillary temperature 38.5°C | 12
systolic blood pressure 120-130 mmHg | 12
diastolic blood pressure 80-90 mmHg | 12
pulse rate 120-140 bpm | 12
SpO2 100% | 12
transferred to a general hospital | 12
blood examinations performed at the general hospital | 24
high levels of D-dimer | 24
high levels of fibrin degradation products | 24
disseminated intravascular coagulation suspected | 24
systemic management in intensive care unit | 24
condition worsened | 36
death confirmed | 48
pleural effusion | 48
pulmonary infiltration | 48
pulmonary shadow | 48
malignant neoplasm suspected | 48
autopsy not performed | 48
histopathological testing not performed | 48