64 years old | 0
male | 0
hypertension | 0
mild chronic renal insufficiency | 0
diabetes mellitus type 2 | 0
admitted to the intensive care unit | 0
Fournier's gangrene | 0
septic shock | 0
respiratory deterioration | 0
hemodynamic instability | 0
scrotum involvement | 0
perineum involvement | 0
right ischial area involvement | 0
lower abdomen involvement | 0
hemodynamic stabilization | 0
broad-spectrum antibiotic therapy | 0
first surgical debridement | 0
temporary diverting colostomy | 0
second radical debridement | 48
suprapubic cystostomy | 48
negative pressure wound therapy | 48
hyperbaric oxygen therapy | 48
methicillin-resistant Staphylococcus epidermidis | 0
Proteus mirabilis | 0
Enterococcus faecalis | 0
NPWT dressing changed twice a week | 48
healthy granulation tissue | 504
primary delayed closure of lower abdomen | 504
scrotal advancement flaps | 504
Integra dermal regeneration template | 504
split-thickness skin graft | 504
NPWT applied over dermal template | 504
NPWT removed after 5 days | 504
healed | 1392
discharged | 1392
