62 years old | 0
    male | 0
    diabetes mellitus | 0
    hypertension | 0
    fever | -48
    dyspnea | -48
    productive cough | 0
    yellow purulent sputum | 0
    smoked 20 cigarettes a day for 40 years | 0
    worked as a house painter | 0
    visited a hot spring 10 days prior | -240
    no history of immunosuppression | 0
    no recurrent infection | 0
    no chemotherapy | 0
    no steroid use | 0
    blood pressure 118/60 mmHg | 0
    heart rate 130 beats/min | 0
    respiratory rate 28/min | 0
    percutaneous oxygen saturation 95% (10 L/min via reservoir mask) | 0
    body temperature 37.5℃ | 0
    holoinspiratory coarse crackles in right lung | 0
    high anion gap metabolic acidosis | 0
    increased lactate | 0
    leukopenia | 0
    thrombocytopenia | 0
    renal dysfunction | 0
    elevated transaminase | 0
    chest radiograph infiltration right upper and middle lobes | 0
    chest computed tomography consolidation with air bronchogram in right upper and middle lobes | 0
    diagnosed with community-acquired pneumonia | 0
    admitted to hospital | 0
    Gram-negative cocci and coccobacilli on sputum Gram staining | 0
    excellent sputum quality | 0
    suspicion of S. pneumoniae pneumonia | 0
    Gram-positive cocci not present | 0
    consideration of A. baumannii as causative organism | 0
    initiation of meropenem | 0
    initiation of azithromycin | 0
    intubation | 0
    noradrenaline administration | 0
    recuperation from septic shock | 24
    respiratory improvement | 24
    A. baumannii identified in sputum culture | 72
    antibiotic change to ampicillin/sulbactam | 72
    negative blood cultures | 0
    extubation | 96
    nasal high-flow therapy | 96
    transfer out of intensive care unit | 168
    Serratia marcescens identified in sputum culture | 288
    diagnosis of hospital-acquired pneumonia | 288
    antibiotic change to cefepime | 288
    necrotizing pneumonia | 312
    intravenous antibiotics for 42 days | 0
    oral ciprofloxacin for 14 days | 0
    discharge | 1008
    