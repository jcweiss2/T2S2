3 years old | 0
female | 0
admitted to the hospital | 0
fever | -168
cough | -168
respiratory distress | -168
decreased mental status | -168
oseltamivir | -144
difficult breathing | -144
sleepiness | -144
impending respiratory failure | -48
decreased mental status | -48
intubated | 0
chest wall retraction | 0
left lung sounds decreased | 0
drowsy | 0
pancytopenia | 0
elevated C-reactive protein | 0
decreased immunoglobulin G | 0
high dose oseltamivir | 0
intravenous immunoglobulin G | 0
H1N1 influenza virus detected | 0
diffuse haziness in the entire left lung field | 0
right upper lung field infiltration | 0
thoracentesis | 0
turbid chocolate-colored fluid drained | 0
pleural fluid analysis | 0
chest tube inserted | 72
necrotizing pneumonia | 144
persistent high fever | 144
leukocytosis | 144
broad spectrum antibiotics | 144
pneumothorax | 168
chest tube replaced | 168
ventilator support | 168
cefotaxime changed to meropenem | 168
progressive respiratory failure | 216
purulent pleural effusion | 216
recurrent massive pneumothorax | 216
venovenous ECMO support initiated | 216
multidrug resistant Acinetobacter baumannii | 240
bacteremia | 240
tracheal aspirate cultures positive | 240
pleural fluid cultures positive | 264
ECMO support discontinued | 360
ventilator weaning | 888
antimicrobials discontinued | 1,368
left chest tube removed | 1,512
discharged | 1,512
no respiratory symptoms | 1,512
chest radiograph improved | 1,512