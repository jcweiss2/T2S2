27 years old | 0
    male | 0
    admitted to the emergency department | 0
    gingival bleeding | -144
    haematuria | -144
    haematochezia | -144
    pain in the right lower abdomen | -144
    swelling of the left lower limb | -144
    numbness of the left lower limb | -144
    weakness of the left lower limb | -144
    no dizziness | 0
    no fever | 0
    no cough | 0
    no expectoration | 0
    no chest tightness | 0
    no palpitation | 0
    white blood cell count 23.36 × 10^9/l | 0
    neutrophil percentage 68.1% | 0
    haemoglobin 110 g/l | 0
    platelet count 276 × 10^9/l | 0
    urinary protein 3+ | 0
    urinary occult blood 3+ | 0
    occult blood in the stool | 0
    activated partial thromboplastin clotting time 85.4 s | 0
    prothrombin time 16.6 s | 0
    alanine transaminase 86 U/l | 0
    albumin 35 g/l | 0
    creatinine 65 µmol/l | 0
    blood glucose 7.1 mmol/l | 0
    anti-infection treatment | 0
    haemostasis treatment | 0
    symptomatic treatments | 0
    admitted to the intensive care unit | -24
    abdominal CT showed bilateral renal pelvis density increase | -24
    bilateral perirenal fascia thickening | -24
    fat density around bilateral ureteral area increased | -24
    pelvic fascia thickening | -24
    liver morphology irregular | -24
    liver cirrhosis not excluded | -24
    gastrointestinal decompression | -24
    enema | -24
    crystal and colloidal liquid replenishment | -24
    volume expansion | -24
    blood transfusion | -24
    haemostasis | -24
    anti-infection | -24
    nutrition support | -24
    symptomatic support | -24
    white blood cell count 34.24 × 10^9/l | 0
    haemoglobin 66 g/l | 0
    activated partial thromboplastin time 130 s | 0
    transferred to Qilu Hospital emergency department | 0
    hepatitis B virus positive | -4320
    no drug or food allergy | 0
    no trauma history | 0
    no surgery history | 0
    no blood transfusion history | 0
    smoking history 10 years | -87600
    stopped smoking 3 weeks | -504
    father with diabetes mellitus | 0
    father with hypertension | 0
    no family genetic diseases | 0
    no family infections | 0
    body temperature 36.8°C | 0
    heart rate 146 beats/min | 0
    respiration rate 22 breaths/min | 0
    blood pressure 94/66 mmHg | 0
    oxygen saturation 98% | 0
    poor spirit | 0
    drowsiness | 0
    anaemic appearance | 0
    sclera yellow stained | 0
    bilateral pupils equal in size | 0
    pupils sensitive to light reflection | 0
    bleeding at right subclavian vein catheterization | 0
    respiratory sounds thick | 0
    no dry rales | 0
    no wet rales | 0
    heart rhythm uniform | 0
    no pathological murmurs | 0
    abdomen bulging | 0
    no muscle tension | 0
    large areas of ecchymosis on waist | 0
    skin around umbilicus blue-purple | 0
    left lower abdomen tender | 0
    right lower abdomen tender | 0
    no rebound pain | 0
    hard mass in left lower abdomen | 0
    liver not palpable | 0
    spleen not palpable | 0
    left lower limb circumference 72 cm | 0
    right lower limb circumference 62 cm | 0
    bilateral Babinski signs negative | 0
    coagulation factor V 54% | 0
    coagulation factor VII 28% | 0
    coagulation factor VIII 1% | 0
    coagulation factor IX 85% | 0
    double lung inflammation | 0
    pleural effusion | 0
    abdominal effusion | 0
    pelvic effusion | 0
    peritoneal thickening | 0
    omental thickening | 0
    abdominal wall edema | 0
    pelvic wall edema | 0
    bilateral femoral muscle space edema | 0
    subcutaneous fat edema | 0
    soft tissue edema | 0
    preliminary diagnosis of septic shock | 0
    hypovolaemic shock | 0
    anemia to be investigated | 0
    coagulation dysfunction | 0
    gastrointestinal bleeding | 0
    urinary tract bleeding | 0
    chronic HBV | 0
    diet prohibition | 0
    meropenem treatment | 0
    vitamin K1 | 0
    phenolsulfonamethylamine | 0
    aminometrinic acid | 0
    batroxobin haemostatic | 0
    omeprazole | 0
    octreotide | 0
    magnesium isoglycyrrhizin | 0
    reduced glutathione | 0
    entecavir | 0
    plasma supplements | 0
    cold precipitation | 0
    red blood cell infusion | 0
    nutrition support | 0
    symptomatic support | 0
    possible anticoagulant rodenticide poisoning | 0
    transferred to Department of Poisoning and Occupational Diseases | 24
    black stools on day 3 | 72
    red blood cell infusion | 72
    plasma infusion | 72
    glucose water test negative | 120
    acidified serum haemolysis test negative | 120
    plasma free Hb 41.9 mg/l | 120
    direct antiglobulin test negative | 120
    anticoagulant rodenticide not detected | 120
    black stools decreased on day 7 | 168
    no special discomfort | 168
    skin ecchymosis deepened | 168
    blood cultures no anaerobic growth | 168
    blood cultures no bacterial growth | 168
    coagulation factor V 89% | 168
    coagulation factor VII 85% | 168
    coagulation factor VIII 1% | 168
    coagulation factor IX 92% | 168
    ferritin 709 ng/ml | 288
    CA 19-9 294.3 U/ml | 288
    CA 125 306.1 U/ml | 288
    neuron specific enolase 27.27 ng/ml | 288
    immune system no abnormality | 288
    systemic lupus erythematosus excluded | 288
    bone marrow puncture no abnormality | 288
    abdominal CT cholecystitis on day 14 | 336
    retroperitoneal lymph nodes swollen | 336
    multiple low-density shadows in abdomen | 336
    pancreatic area blurred | 336
    peritoneal thickening | 336
    left chest soft tissue swelling | 336
    abdominal wall swelling | 336
    laboratory indices improved on day 21 | 504
    coagulation factor VIII 5.2% | 504
    factor VIII inhibitor 1.5 BU | 504
    PLAT gene p.Y471H mutation | 504
    SERPINE1 gene p.Y244Y mutation | 504
    diagnosed with acquired FVIII deficiency | 504
    prednisone 30 mg daily | 504
    transferred to Department of Haematology | 504
    cryoprecipitate 10 U | 504
    symptoms improved after 2 days | 576
    discharged | 576
    no bleeding at follow-up | 720
    coagulation factor VIII increased | 720
    factor VIII antibody negative | 720
    left iliopsoas muscle swelling | 720
    bleeding cannot be excluded | 720
    <|eot_id|>