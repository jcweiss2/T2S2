56 years old | 0
male | 0
admitted to ICU | 0
chronic kidney disease | -720
maintenance hemodialysis | -720
septic shock | 0
coagulopathy | 0
altered sensorium | 0
hypotension | 0
Glasgow coma scale 7/15 | 0
heart rate 112 beats/min | 0
non-invasive blood pressure 87/48 mmHg | 0
axillary temperature 38.5℃ | 0
dialysis-related septic shock | 0
fluid resuscitation | 0
routine cultures | 0
empirical antibiotic therapy | 0
intubated | 0
mechanical ventilation | 0
leukocyte count 17 × 10^6/cm^3 | 0
sodium levels 122 mEq/L | 0
potassium 3.2 mEq/L | 0
international normalized ratio 3.2 | 0
normal platelet count | 0
vasopressor therapy | 0
dialysis catheter in right internal jugular vein | -720
central venous catheter insertion | 0
ultrasound-guided insertion | 0
catheter formed a loop inside left brachiocephalic vein | 0
catheter tip in left subclavian vein | 0
dialysis catheter removed | 2
new dialysis catheter inserted in femoral vein | 2
central line repositioned | 2
catheter entered right subclavian vein | 2
catheter withdrawn 1-2 cm | 4
catheter tip at junction of great veins | 4
discharged | 24