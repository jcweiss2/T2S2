48 years old | 0
male | 0
paraplegia | 0
spina bifida | 0
admitted to the hospital | 0
long-term indwelling urethral catheter | -6720
temperature of 39°C | -240
urine microbiology revealed Pseudomonas aeruginosa | -240
ciprofloxacin 500 mg twice a day for 7 days | -240
ultrasound examination of urinary tract | -240
bilateral renal calculi | -240
isotope renogram | -240
divided renal function | -240
persistent obstructive pattern | -240
CT revealed large staghorn calculus | -240
flexible uretero-renoscopy | -192
left ureteroscopy with laser lithotripsy | -192
insertion of left ureteric stent | -192
repeat left ureterorenoscopy and laser lithotripsy | -96
ureteroscopy and laser lithotripsy | -96
CT of kidney, ureters, bladder | -72
generalized shrinkage of left kidney | -72
multifocal scarring | -72
ureteric stent in situ | -72
lower pole stones | -72
dilatation of the upper pole pelvicalyceal system | -72
left JJ stent removed | -28
gentamicin 160 mg | -28
stone analysis revealed struvite | -28
blood pressure was recorded as 143/97 mmHg | -14
urine sample sent for microbiology | -14
mixed growth | -14
left rigid ureterorenoscopy | 0
gentamicin 240 mg intravenously | 0
ureter was normal | 0
access sheath of size 13/15, 46 cm | 0
flexible ureteroscopy and laser lithotripsy | 0
fragments removed with a basket | 0
right rigid ureteroscopy | 0
ureter was normal | 0
access sheath of size 13/15, 46 cm | 0
laser lithotripsy | 0
fragments removed with a basket | 0
possible intrarenal mucosal perforation | 0
JJ stent inserted in both ureters | 0
surgery lasted for 2 hours and 40 minutes | 0
blood pressure was 80/40 mmHg | 0
frank hematuria | 0
sinus tachycardia | 0
admitted to the critical care unit | 0
hemodynamically stable | 0
temperature of 39°C | 0
hemoglobin: 116 g/L | 0
white blood cell count: 24.5×10^9/L | 0
neutrophils: 22.6×10^9/L | 0
INR: 1.2 | 0
APTT: 32 seconds | 0
APTT ratio: 1.3 | 0
C-reactive protein: 137 mg/L | 0
creatinine: 64 μmol/L | 0
cefuroxime intravenously nocte and mane | 0
transferred to the spinal unit | 24
temperature of 38°C | 24
urine was dark red | 24
blood tests | 24
INR: 1.1 | 24
hemoglobin: 120 g/L | 24
white blood cell count: 20×10^9 | 24
neutrophils: 17.9×10^9 | 24
C-reactive protein: 168.1 mg/L | 24
gentamicin for 5 days | 24
hematuria subsided | 168
discharged home | 168
ureteric stents removed | 168
gentamicin 160 mg | 168
developed temperature | 192
CT of kidneys | 192
hemoglobin: 128 g/L | 192
white blood cell count: 9.6×10^9 | 192
C-reactive protein: 133.4 mg/L | 192
urine culture: P. aeruginosa | 192
ciprofloxacin 500 mg twice a day for 5 days | 192
CT of urinary tract | 336
subcapsular collection on the left kidney | 336
minor perinephric fat stranding | 336
residual stones/fragments | 336
elevated left hemidiaphragm | 336
minimal atelectasis in the left lower zone | 336
percutaneous drainage not carried out | 336
ciprofloxacin 500 mg twice a day for 5 days | 336
urine sample sent for culture | 336
Pseudomonas aeruginosa resistant to gentamicin and ciprofloxacin | 336
ciprofloxacin discontinued | 336
ferrous sulfate 200 mg daily | 336
isotope renogram | 560
deterioration in the left renal function | 560
left kidney contributed only 17% | 560
right kidney contributed 83% | 560
ultrasound scan of left kidney | 616
residual hematoma 3.3 cm in depth | 616
CT of kidney, ureters, bladder | 784
left renal subcapsular collection much reduced in size | 784
inflammatory stranding in the left perinephric fat | 784
no hydronephrosis | 784
residual calculi | 784
blood pressure was 146/93 mmHg | 784
24-hour mean blood pressure: 130/91 mmHg | 784
ramipril 1.25 mg daily | 784
hemoglobin had increased to 157 g/L | 1344