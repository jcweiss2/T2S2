70 years old | 0
female | 0
admitted to the hospital | 0
constipation | -240
abdominal pain | -240
vomiting | -240
not passed stool or flatus | -240
dehydrated | 0
febrile | 0
temperature of 37.8 centigrade | 0
pulse of 130/minute | 0
blood pressure of 100/70 mm Hg | 0
respiratory rate of 26/min | 0
BMI of 16 kg/m2 | 0
history of asthma | 0
on steroid inhalers | 0
bilateral rhonchi | 0
tense and tender abdomen | 0
generalized guarding | 0
hyperdynamic bowel sounds | 0
inconclusive digital rectal examination | 0
total white cell count of 16×109/L | 0
multiple scattered air fluid levels on x-ray | 0
dilated small bowel loops on ultrasonography | 0
normal peristaltic activity on ultrasonography | 0
provisional diagnosis of acute small bowel obstruction | 0
exploratory laparotomy | 3
strangulated obturator hernia | 3
loop of the ileum in the hernia sac | 3
Meckel diverticulum in the hernia sac | 3
perforation at the base of the Meckel diverticulum | 3
resection of 2.5 feet of the dusky ileum | 3
hernia defect repair with non-absorbable purse string sutures | 3
loop ilestomy creation | 3
abdomen cleansed with 6 liters of normal saline | 3
retention sutures applied | 3
abdomen closed with skin defect left open | 3
transferred to the intensive care unit | 3
ventilator support | 3
expired due to multiple organ dysfunction and overwhelming sepsis | 72
history of multiparity | 0
low BMI | 0
emaciation | 0
protective preperitoneal fat in the pelvis reduced | 0
frequent bouts of forceful coughing | 0
chronic bronchitis | 0
preperitoneal connective tissue and fat entering the pelvic orifice of the obturator canal | -6720
formation of a peritoneal sac | -6720
entrance of an organ into the hernia sac | -6720
CT scan not performed | 0
facility located a considerable distance from the CT scan centre | 0
urgent surgical intervention due to acute peritonitis | 0
transperitoneal approach | 3
importance of early surgical intervention | 0
duration of onset of symptoms to surgery | -240
development of numerous complications | -240
Multi Organ Dysfunction (MODS) | -240
patient belonged to a family with low literacy and socio-economic status | 0
delay in seeking medical attention | -240
Meckel’s diverticulum in the hernia sac | 3
mixed Littré’s hernia | 3
true Littré’s hernia | 0
Meckel’s diverticulum perforation | 3
compromised circulation | 0
narrow neck | 0
peptic ulceration | 0
ectopic gastric tissue | 0
Littré’s hernia in femoral, sciatic, paraumbilical, lumbar, and laparoscopic port site hernias | 0
Meckel’s diverticulum in an obturator hernia | 3
Howship Romberg sign | 0
CT scan or laparotomy for accurate diagnosis | 0
early diagnosis and surgical intervention | 0
high morbidity and mortality | 0