58 years old | 0
male | 0
admitted to the hospital | 0
fecal occult blood | -48
underwent partial endoscopic mucosal resection | -72
electrocoagulation electro resection | -72
cold resection | -72
polyps in the cecum and colon | -72
broad-based or pedicled polyps | -72
diameters of 0.5-2.0 cm | -72
removed polyps by EMR | -72
cold resection | -72
electrocoagulation and electro resection | -72
shock | -72
dyspnea | -72
sweating | -72
BP decreased to 79/44 mmHg | -72
oxygen saturation decreased to 77% | -72
HR increased to 133 beats/min | -72
transferred to the ICU | -71
stable vital signs | -48
normal coagulation function | -48
underwent colonoscopy-guided polypectomy | 144
ulcerative foci scattered in the transverse colon and descending colon | 144
wound of the first surgery | 144
three 0.8-1.2 cm polyps scattered in the descending colon and sigmoid colon | 144
removed by EMR | 144
wound surface closed with titanium clips | 144
BP suddenly decreased to 76/42 mmHg | 144
HR increased to 133 beats/min | 144
SpO2 dropped to 90% | 144
mental irritability | 144
gastrectomy | -7300
surgical treatment for oral cancer | -365
hospitalized for oral cancer | -1096
painless colonoscopy | -1096
polyps found in the colon | -1096
denies family genetic history | 0
vital signs and physical examination changed rapidly | 0
blood gas analysis | -72
pH 7.33 | -72
partial pressure of carbon dioxide 37 mmHg | -72
partial pressure of oxygen 211 mmHg | -72
lactate levels 4.8 mmol/L | -72
bicarbonate radical concentration 19.5 mmol/L | -72
base excess 5.8 mmol/L | -72
potassium ion concentration 2.9 mmol/L | -72
PaO2/FiO2 221 mmHg | -72
WBC count 3.29 × 10^9/L | -72
neutrophil percentage 87.8% | -72
platelet count 142 × 10^12/L | -72
PCT concentration 1.66 ng/mL | -72
IL-6 concentration > 5000 pg/mL | -72
PT 36.2 s | -72
INR 3.6 | -72
PTA 21% | -72
APTT 69.1 s | -72
fibrinogen concentration < 0.6 g/L | -72
FDP concentration > 360 μg/mL | -72
D-dimer concentration > 40 μg/mL | -72
AT III level 69% | -72
blood culture negative | -72
blood gas analysis | 144
pH 7.23 | 144
PaCO2 33 mmHg | 144
PaO2 149 mmHg | 144
lactate level 7.1 mmol/L | 144
bicarbonate radical concentration 13.8 mmol/L | 144
BE -12.7 mmol/L | 144
potassium ion concentration 6.5 mmol/L | 144
PaO2/FiO2 186 mmHg | 144
leukocytosis | 144
elevated concentrations of infection markers | 144
coagulopathy | 144
WBC count 12.38 × 10^9/L | 144
neutrophil percentage 86.4% | 144
hemoglobin concentration 84 g/L | 144
platelet count 192 × 10^12/L | 144
PCT concentration 1.26 ng/mL | 144
IL-6 concentration > 5000 pg/mL | 144
PT 36.5 s | 144
INR 3.64 | 144
PTA 20% | 144
APTT 62 s | 144
fibrinogen concentration < 0.6 g/L | 144
FDP concentrations > 360 μg/mL | 144
D-dimer concentration > 40 μg/mL | 144
AT III 65% | 144
thromboelastography | 144
comprehensive coagulation index -9.9 | 144
fibrinogen function α-angle 17.8 | 144
K-time exceeding the upper limit | 144
maximum amplitude 19.2 mm | 144
blood gas analysis | 216
pH 7.23 | 216
PaCO2 33 mmHg | 216
PaO2 149 mmHg | 216
lactate level 7.1 mmol/L | 216
bicarbonate radical concentration 13.8 mmol/L | 216
BE -12.7 mmol/L | 216
potassium ion concentration 6.5 mmol/L | 216
PaO2/FiO2 186 mmHg | 216
WBC count 20.46 × 10^9/L | 216
hemoglobin concentration 62 g/L | 216
PCT concentration 5.72 ng/mL | 216
platelet count and coagulation function normal | 216
abdominal CT | 216
superior mesenteric artery CT angiography | 216
no intestinal perforation or lumbar lesion | 216
no vascular damage | 216
sepsis | -72
septic shock | -72
SOFA score 4 | -72
Respiration 2 | -72
Coagulation 1 | -72
Cardiovascular 1 | -72
elevated PCT | -72
infection | -72
PPS with sepsis and septic shock | -72
SOFA score 5 | 144
Respiration 3 | 144
Cardiovascular 2 | 144
elevated PCT and IL-6 | 144
infection | 144
septic shock with Sepsis-3 | 144
blood culture results | 216
Moraxella osloensis | 216
discharged | 288
sepsis and septic shock caused by PPS | 288
gastrointestinal bleeding | 288
coagulopathy | 288
abdominal pain | -72
fever | -72
inflammatory markers | -72
abnormal coagulation | -72
life-threatening sepsis | -72
septic shock | -72
gastrointestinal bleeding | -72
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 0
gastrointestinal bleeding | 0
PPS without abdominal pain | 0
severe coagulopathy | 0
gastrointestinal bleeding | 0
sepsis | 0
septic shock | 0
PPS | 0
abdominal pain | 0
fever | 0
inflammatory markers | 0
abnormal coagulation | 0
life-threatening sepsis | 0
septic shock | 