term male neonate | 0
born by normal spontaneous vaginal delivery | 0
membranes spontaneously ruptured for 13 h | -13
pregnancy with gestational diabetes | -672
hydronephrosis | -672
stent placement | -672
multiple urinary tract infections secondary to Klebsiella sp | -672
transferred to neonatal ICU | 0
temperature instability | 0
respiratory distress | 0
increasing supplemental oxygen requirement | 0
appeared dusky | 0
oxygen saturations of 80% | 0
placed on 2 L nasal cannula at 21% FiO2 | 0
continued respiratory distress | 0
grunting | 0
tachypnea | 0
FiO2 increased to 40% | 0
serum glucose unremarkable | 0
blood gas unremarkable | 0
complete blood count unremarkable | 0
renal function panel unremarkable | 0
C-reactive protein unremarkable | 0
chest radiograph mild diffuse ground glass opacities | 0
blood culture drawn | 0
empirically started on ampicillin | 0
gentamicin | 0
ceftazidime | 0
respiratory failure on day 2 | 48
intubation | 48
copious purulent drainage from left eye | 48
ophthalmologic examination | 48
diffuse fleshy red pseudomembrane coating bulbar conjunctiva | 48
pseudomembrane coating tarsal conjunctiva | 48
pseudomembrane debrided | 48
purulent drainage | 48
serosanginous drainage | 48
bacterial culture from left eye grew E. coli | 48
viral culture sent | 48
blood culture negative | 48
urine culture negative | 48
cerebral spinal fluid studies negative | 48
placental pathology normal | 48
mother hospitalized for urosepsis secondary to E. coli | 48
sensitivities mirrored | 48
extubated to nasal cannula | 72
repeat ophthalmologic examinations | 72
significant clinical improvement | 72
intravenous antimicrobials | 72
topical antimicrobials | 72
completed 14-day course of ampicillin | 336
pneumonia | 0
sepsis | 0
completed 11 days of moxifloxacin eye drops | 264
weaned to room air | 120
discharged home | 336
follow-up eye examination normal | 432
complete resolution of conjunctivitis | 432
