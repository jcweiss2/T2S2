18 years old | 0
male | 0
admitted to the hospital | 0
shortness of breath | 0
severe right-sided chest pain | 0
fever | -336
sore throat | -336
dysphagia | -336
fatigue | -336
cervical lymphadenopathy | -336
pharyngitis | -336
splenomegaly | -336
infectious mononucleosis | -336
EBV infection | -336
admitted to hospital for tonsillitis | -144
discharged from hospital | -120
Penicillin V | -144
dyspnoeic | 0
respiratory rate 30 breaths per minute | 0
peripheral oxygen saturations 94% | 0
temperature 37.4°C | 0
pulse rate 120 beats per minute | 0
blood pressure 100/70 mmHg | 0
bilateral symmetrical tonsillar swelling | 0
white exudate | 0
bilateral cervical lymphadenopathy | 0
leucocytosis | 0
atypical lymphocytes | 0
elevated C-reactive protein | 0
elevated liver enzymes | 0
alkaline phosphatase 147 IU/l | 0
alanine aminotransferase 76 IU/l | 0
pneumomediastinum | 0
mediastinal fat stranding | 0
pockets of fluid in the anterior mediastinum | 0
right pleural effusion | 0
inflammatory consolidation in the right lung | 0
reactive lymph nodes | 0
splenomegaly | 0
enlarged lymphoid tissue in the posterior nasopharynx | 0
no oesophageal perforation | 0
no peritonsillar or retropharyngeal abscesses | 0
IV opioid analgesia | 0
fluid resuscitation | 0
amoxicillin and clavulanic acid | 0
cardiothoracic surgery consultation | 0
increased chest pain | 4
worsening physiology | 4
antibiotics changed to IV Piperacillin and tazobactam with clindamycin | 4
video-assisted thoracoscopic surgery | 4
drainage and decortication of a right pleural empyema | 4
drainage of multiple mediastinal abscesses | 4
debridement of mediastinal necrotic tissue | 4
insertion of a right-sided intercostal drain | 4
Fusobacterium necrophorum detected | 4
Dialister pneumosintes detected | 4
Peptostreptococcus anaerobius detected | 4
admitted to intensive care unit | 4
supportive care | 4
discharged home | 528