29 years old | 0
    male | 0
    metformin overdose | -5.5
    suicide attempt | -5.5
    ethanol ingestion | -5.5
    no diabetes | 0
    psychosis | 0
    depression | 0
    prior suicide attempts | 0
    discontinued olanzapine | -720
    discontinued sertraline | -720
    daily ethanol use | 0
    daily tobacco use | 0
    vomiting | -5.5
    diarrhea | -5.5
    thirst | -5.5
    abdominal pain | -5.5
    bilateral leg pain | -5.5
    agitation | -5.5
    fingerstick glucose 180 mg/dL | -5.5
    temperature 35.2°C | 0
    pulse 113 beats/min | 0
    blood pressure 129/59 mmHg | 0
    respirations 28 breaths/min | 0
    oxygen saturation 100% | 0
    awake and oriented x4 | 0
    confusion | 0
    GCS=14 | 0
    pupils equal and reactive | 0
    dry oral mucous membranes | 0
    tachycardia | 0
    unremarkable heart exam | 0
    unremarkable lung exam | 0
    mild diffuse abdominal tenderness | 0
    soft abdomen | 0
    no guarding | 0
    no rebound | 0
    fecal incontinence | 0
    guaiac-negative stool | 0
    normal rectal tone | 0
    sinus tachycardia | 0
    fingerstick glucose 364 mg/dL | 0
    combative behavior | 0
    attempted biting | 0
    attempted spitting | 0
    soft restraints | 0
    respiratory protection mask | 0
    lorazepam 2 mg | 0
    dolasetron 12.5 mg | 0
    morphine sulfate 4 mg | 0
    0.9% saline hydration | 0
    no longer combative | 45
    restraints removed | 45
    sodium 136 mEq/L | 0.5
    potassium 3.1 mEq/L | 0.5
    chloride 105 mEq/L | 0.5
    bicarbonate 9 mEq/L | 0.5
    BUN 2 mg/dL | 0.5
    creatinine 2.1 mg/dL | 0.5
    glucose 707 mg/dL | 0.5
    calcium 9.4 mg/dL | 0.5
    total protein 7.6 g/dL | 0.5
    AST 60 IU/L | 0.5
    ALT 53 IU/L | 0.5
    bilirubin 0.8 mg/dL | 0.5
    acetaminophen <5 μg/mL | 0.5
    salicylate <4 mg/dL | 0.5
    lactate >11.1 mmol/L | 0.5
    ethanol 214 mg/dL | 0.5
    osmolality 392 mOsm/kg | 0.5
    β-hydroxybutyrate 2.4 mg/dL | 0.5
    hyperglycemia | 0.5
    metabolic acidosis | 0.5
    arterial pH 7.10 | 0.5
    pCO2 18.8 mmHg | 0.5
    pO2 133.1 mmHg | 0.5
    elevated anion gap | 0.5
    osmolal gap >20 mOsm/kg | 0.5
    normal β-hydroxybutyrate | 0.5
    no ketonuria | 0.5
    glycosuria | 0.5
    moderate hemoglobinuria | 0.5
    no calcium oxalate crystalluria | 0.5
    no blood cells in urine | 0.5
    no infection in urine | 0.5
    negative urine drug screen | 0.5
    admitted to ICU | 0.5
    no ICU bed availability | 0.5
    remained in ED | 0.5
    nephrology consultation | 1
    bicarbonate 6 mEq/L | 4
    glucose 672 mg/dL | 4
    continued IV hydration | 4
    unresponsive | 5
    vomiting | 5
    aspiration | 5
    PEA | 5
    heart rate 29/min | 5
    chest compressions | 5
    endotracheal intubation | 5
    epinephrine 2 mg | 5
    atropine 1 mg | 5
    sodium bicarbonate 176 mEq | 5
    heart rate 110/min | 5
    blood pressure 121/88 mmHg | 5
    arterial pH 6.95 | 5
    pCO2 55.7 mmHg | 5
    pO2 88.1 mmHg | 5
    bicarbonate 12.4 mEq/L | 5
    bicarbonate drip | 5
    transferred to ICU | 5
    ventricular tachycardia | 6
    blood pressure 72/44 mmHg | 6
    dopamine drip | 6
    coagulopathy | 6
    INR 3.08 | 6
    fibrinogen 113 mg/dL | 6
    d-dimer >8.0 mcg/mL | 6
    fresh frozen plasma | 6
    platelet count 390 k/mm3 | 6
    hematocrit 47.7% | 6
    decreased left ventricular function | 6
    CK-MB elevation | 6
    troponin I elevation | 6
    hemodialysis | 12
    PEA | 15
    resuscitation | 15
    recurrent PEA | 15
    death | 19
    lactate >11.1 mmol/L | 19
    bicarbonate 12 mEq/L | 19
    glucose 327 mg/dL | 19
    insulin drip | 19
    hemodialysis | 19
    no serum lipase measurement | 19
    no serum amylase measurement | 19