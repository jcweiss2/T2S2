12 years old | 0
female | 0
admitted from the emergency department to the intensive care unit | 0
fever | -336
multiple asymmetrical joint swelling | -336
joint pain | -336
admission temperature 39.6°C | 0
heart rate 130 beats/min | 0
arterial blood pressure 127/57 mmHg | 0
respiratory rate 35 breaths/min | 0
oxygen saturation 93% on air | 0
hair lice | 0
multiple scratch marks on her scalp | 0
bilateral pleural effusion | 0
ejection systolic murmur grade 2/6 over the aortic area | 0
tender hepatomegaly | 0
liver span 10 cm | 0
multiple joint swelling | 0
redness | 0
tenderness | 0
right middle finger involvement | 0
right hip involvement | 0
both knees involvement | 0
ankles involvement | 0
white blood cell count 6000 cells/mm³ | 0
lymphocytes 0.9×10⁹ cells/l | 0
granulocytes 4.5×10⁹ cells/l | 0
monocytes 0.2×10⁹ cells/l | 0
reticulocytes 28×10⁹ cells/l | 0
platelets 156,000 cells/mm³ | 0
hemoglobin 107 g/l | 0
serum sodium 125 mmol/l | 0
serum potassium 4.8 mmol/l | 0
serum glucose 4.3 mmol/l | 0
serum urea 20.7 mmol/l | 0
serum creatinine 90 mmol/l | 0
lactate dehydrogenase 1427 IU/L | 0
aspartate aminotransferase 408 IU/L | 0
alanine transaminase 307 IU/L | 0
alkaline phosphatase 184 IU/L | 0
albumin 19 g/l | 0
gamma-glutamate transferase 110 IU/L | 0
creatine kinase 142 IU/L | 0
total bilirubin 145 mmol/l | 0
serum osmolality 289 mOsm/kg | 0
urine osmolality 647 mOsm/kg | 0
international normalized ratio 1.2 | 0
prothrombin time 14 | 0
activated partial thromboplastin time 36 | 0
sickle cell disease negative | 0
hepatitis A negative | 0
hepatitis C negative | 0
human immunodeficiency virus negative | 0
anti-HBs Ag antibodies positive | 0
chest X-ray bilateral pleural effusion | 0
widened mediastinum | 0
pear-shaped heart | 0
pericardial effusion | 0
sinus tachycardia | 0
diffuse ST-segment elevation | 0
generalized T-wave inversion | 0
transthoracic echocardiogram moderate size pericardial effusion | 0
no endocarditis | 0
no valvular heart disease |A|0
blood cultures obtained | 0
sputum cultures obtained | 0
urine cultures obtained | 0
ceftazidime started | 0
flucloxacillin started | 0
right chest tube thoracostomy inserted | 0
serous fluid drained 800 ml | 0
no air leak | 0
pleural fluid lactate dehydrogenase 5 IU/L | 0
pleural fluid albumin 19 g/L | 0
pleural fluid pH 7.37 | 0
Gram-positive cocci in clusters on pleural fluid Gram staining | 0
hair shaved | 0
anti-lice shampoo started | 0
sputum microscopy negative for acid-fast bacilli | 0
mycobacterium tuberculosis culture sample sent | 0
polymerase chain reaction test sent | 0
more tachypneic (RR 40 breaths/min) | 24
hypotensive (BP 90/40 mmHg) | 24
trachea intubated | 24
mechanical ventilation started | 24
antibiotics changed to meropenem | 24
dopamine infusion started | 24
norepinephrine infusion started | 24
air leak from right chest tube observed | 24
SpO2 maintained >95% on FiO2 0.4 | 24
bronchopleural fistula suspected | 24
echocardiography-guided pericardiocentesis performed | 24
pericardial pus aspirated 500 ml | 24
pig-tail catheter inserted into pericardium | 24
pericardial fluid proteins 42 g/l | 24
pericardial fluid albumin 27 g/l | 24
pericardial fluid Gram-positive cocci in clusters | 24
chest X-ray right minimal hydropneumothorax | 24
ultrasound abdomen perinephric collections | 24
subhepatic collections | 24
free fluid in abdomen | 24
free fluid in pelvis | 24
methicillin-sensitive Staphylococcus aureus cultured from sputum | 24
methicillin-sensitive Staphylococcus aureus cultured from blood | 24
methicillin-sensitive Staphylococcus aureus cultured from pleural fluid | 24
methicillin-sensitive Staphylococcus aureus cultured from pericardial aspirate | 24
urine cultures negative | 24
rheumatoid factor 48.8 IU/L | 24
cytomegalovirus IgM antibodies negative | 24
cytomegalovirus IgG titer 1/21,000 IU/L | 24
air leak through pericardial pig-tail catheter | 96
pus draining through pericardial pig-tail catheter | 96
air leak most marked during mechanical inspiration | 96
broncho-pericardial fistula suspected | 96
broncho-pleuropericardial fistula suspected | 96
pig-tail catheter clamped | 96
BP decreased to 80/50 mmHg | 96
HR increased to 120 beats/min | 96
BP and HR returned to baseline after de-clamping | 96
computed tomography pneumopericardium | 96
computed tomography hydropneumothorax | 96
radio-opaque contrast material injected into pericardial pig-tail catheter | 96
contrast spill into right pleural cavity | 96
CT fistulogram confirmed right pleural space and pericardium communication | 96
conservative management recommended | 96
abdominal collections aspirated laparoscopically | 120
disseminated intravascular coagulation developed | 264
bleeding from everywhere | 264
died of multi-organ failure | 312
parents refused autopsy | 312
