43 years old | 0
male | 0
smoker | 0
admitted to the hospital | 0
chest pain | 0
electrocardiogram changes | 0
postero-lateral myocardial infarction | 0
high serum troponin levels | 0
cardiac arrest | 0
ventricular fibrillation | 0
tMCS | 0
CentriMag Circulatory Support System | 0
cardiorespiratory collapse reversed | 12
coronary angiogram | 12
severe 3-vessel coronary artery disease | 12
stents placed | 12
intra-aortic balloon pump | 12
left ventricular ejection fraction 19% | 12
tMCS weaning | 120
tMCS explanted | 120
neurologically intact | 120
tMCS re-established | 128
tMCS explanted | 216
hemodynamic status deteriorated | 240
tMCS CentriMag instituted | 240
left groin sepsis | 240
arterial cannula re-sited | 240
sepsis cleared | 288
LVAD implantation | 288
bridge to transplantation | 288
ascending aortic intimal flap | 300
type A aortic dissection | 300
ECG-gated computerized tomographic aortogram | 300
intimal flap extended | 300
sino-tubular junction | 300
arch | 300
descending aorta | 300
abdominal aorta | 300
iliac arteries | 300
no communication between true and false lumens | 300
dissection repair | 312
LVAD insertion | 312
cardiopulmonary bypass | 312
left subclavian cannula | 312
right atrial cannula | 312
venous drainage | 312
ascending aorta clamped | 312
innominate artery | 312
aortic incision | 312
significant split | 312
sino-tubular junction | 312
distal ascending aorta | 312
tube graft | 312
Haemashield | 312
Teflon strips | 312
myocardial protection | 312
intermittent antegrade cold blood cardioplegia | 312
topical slush | 312
HeartMate 3 | 312
left ventricular apex | 312
inflow | 312
outflow graft | 312
aortic interposition graft | 312
cardiopulmonary bypass weaned | 312
intensive care unit | 336
ward | 504
discharged home | 672
functional status excellent | 4032
totally independent | 4032