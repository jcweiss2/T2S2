72 years old | 0
male | 0
Caucasian | 0
admitted to the hospital | 0
hypertension | -720
type-2 diabetes mellitus | -720
peripheral arterial disease of the lower limbs | -720
previous coronary artery bypass graft surgery | -720
dry cough | -720
fever | -720
anorexia | -720
loss of more than 10% of body weight | -720
dyspnea | -720
hypotensive | 0
tachycardic | 0
feverish | 0
jugular turgor at 45° | 0
bibasilar pulmonary rales | 0
new systolic mitral regurgitation murmur | 0
cardiorespiratory collapse | 0
mechanical ventilation | 0
continuous infusion of vasopressors | 0
oliguria | 0
poor peripheral perfusion | 0
cold extremities | 0
cyanosis | 0
capillary refill time >2 sec | 0
transferred to the intensive care unit | 0
pulmonary congestion | 0
cardiomegaly | 0
leukocytosis | 0
normocytic anemia | 0
elevated erythrocyte sedimentation rate | 0
elevated C-reactive protein plasma levels | 0
mitral valve thickening | 0
large flail of the anterior leaflet | 0
severe mitral regurgitant jet intensity | 0
severe mitral regurgitant jet area | 0
bilateral multiple B-lines in a diffuse pattern | 0
pulmonary edema | 0
definitive diagnosis of mitral native valve endocarditis | 0
cardiogenic shock | 0
severe acute mitral valve regurgitation | 0
empirical antimicrobial therapy | 0
ceftriaxone | 0
gentamicin | 0
norepinephrine | 0
intra-aortic balloon pump counterpulsation implant | 0
emergency mitral valve replacement surgery | 12
bioprosthetic mitral valve | 12
progressive improvement in cardiogenic shock | 12
gradual reduction of the vasopressor dose | 12
Gemella morbillorum isolated in blood cultures | 24
susceptibility testing | 24
sensitive to penicillin | 24
sensitive to ceftriaxone | 24
sensitive to vancomycin | 24
antibiotic regimen de-escalonated | 24
penicillin G | 24
gentamicin | 24
dependent on mechanical ventilation | 120
critical illness polyneuropathy | 120
refractory pulmonary congestion | 120
tracheostomy | 120
continuous ultrafiltration | 120
new episode of shock | 648
pulmonary edema | 648
lung compliance worsening | 648
need for mechanical ventilation with high pressures | 648
need for high fraction of inspired oxygen | 648
bioprosthetic mitral valve thickening | 648
severe stenosis | 648
emergency surgery for valve replacement | 648
died during the procedure | 648