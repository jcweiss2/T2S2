54 years old | 0
    female | 0
    farmer | 0
    no significant past medical history | 0
    admitted to the local hospital | -168
    fever | -168
    myalgia | -168
    fatigue | -168
    poor oral intake | -168
    lived in Jecheon-Si, Chungchung Province, South Korea | 0
    climbed a mountain | -672
    treated with antipyretics | -168
    fluid therapy | -168
    symptoms not relieved | -168
    somnolent | -72
    unable to follow commands | -72
    thrombocytopenia | -72
    leukopenia | -72
    elevated aspartate aminotransferase | -72
    elevated alanine aminotransferase | -72
    transferred to our hospital | -72
    temperature 37.2°C | 0
    blood pressure 125/81 mm/Hg | 0
    pulse 105 beats per minute | 0
    respiratory rate 22 breaths per minute | 0
    oxygen saturation 92% in ambient air | 0
    acutely ill | 0
    confused | 0
    Glasgow coma scale 13 | 0
    normal pupil light reflex | 0
    no meningeal irritation signs | 0
    clear conjunctivae | 0
    no palpable lymph nodes except both inguinal areas | 0
    no insect bite site | 0
    no eschar | 0
    no skin rash | 0
    no ecchymosis | 0
    mild leucopenia | 0
    thrombocytopenia | 0
    azotemia | 0
    hyperkalemia | 0
    elevated liver enzymes | 0
    increased creatine kinase | 0
    increased myoglobin | 0
    increased aldolase | 0
    negative blood cultures for bacteria | 0
    negative serum serology tests for Hantaan virus | 0
    negative serum serology tests for Leptospira interrogans | 0
    negative serum serology tests for Orientia tsutsugamushi | 0
    negative serum serology tests for Rickettsia typhi | 0
    reverse transcriptase polymerase chain reaction assay for SFTS virus | 0
    mild pulmonary congestion | 0
    bilateral pleural effusion | 0
    no evidence of structural lesions in the hepatobiliary system | 0
    no evidence of structural lesions in the kidney | 0
    no evidence of acute intracranial process | 0
    admitted to the medical intensive care unit | 0
    intravenous piperacillin/tazobactam | 0
    intravenous levofloxacin | 0
    emergent continuous renal replacement therapy | 0
    metabolic acidosis | 0
    hyperkalemia | 0
    died | 72
    rapidly progressive acute respiratory distress syndrome | 72
    multiple organ failure | 72
    SFTS virus demonstrated | 72
    no evidence of encephalitis | 0
    no evidence of hemorrhage | 0
    seizure-like motion | 0
    intermittent limb tremor | 0
    increased muscle enzymes after neuromuscular blocker use | 72
    fatal rhabdomyolysis | 72
    acute renal failure | 72
    myalgia | 0
    fever | 0
    thrombocytopenia | 0
    elevated creatine kinase | 72
    