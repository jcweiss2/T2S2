72 years old | 0
male | 0
cirrhosis | 0
hepatocellular carcinoma | 0
tocilizumab | 0
atezolizumab | 0
bevacizumab | 0
oral prednisone | 0
confusion | -312
lethargy | -312
bilateral lower extremity edema | -312
recurrent falls | -312
lacerations | -312
admitted to the emergency department | -312
admitted to the hospital | 0
feeling unwell | 0
temperature of 100.0°F | 0
blood pressure of 85/50 | 0
heart rate in the 80s | 0
increasing confusion | 0
red, hot, and painful leg ulceration | 0
elevated white blood cell count | 0
left shift | 0
sepsis protocol initiated | 0
admitted to the intensive care unit | 0
broad-spectrum antimicrobials | 0
vancomycin | 0
piperacillin/tazobactam | 0
changed to vancomycin, cefepime, and metronidazole | 24
acute kidney injury | 24
specimens for bacterial culture obtained | 0
blood cultures drawn | 0
M. canis positive | 0
Gram-stained photomicrographs | 0
subculture images | 0
antimicrobial susceptibility testing | 0
beta-lactamase production | 0
resistant to penicillin, ampicillin, and amoxicillin | 0
Staphylococcus aureus | 0
clinical improvement | 48
repeat blood cultures negative | 48
fever resolved | 48
leg wounds improved | 48
total white blood cell and neutrophil counts trended downwards | 48
IV cefepime continued | 48
oral cefdinir as outpatient therapy | 120
discharged | 120