6-year-old | 0  
    boy | 0  
    referred to our center | 0  
    evaluation of an adrenal mass | 0  
    visited the Emergency Department | prior to transfer (assumed several hours before transfer, timestamp -24)  
    generalized tonic-clonic type seizure | -24  
    posterior reversible encephalopathy syndrome | -24  
    hypertension | -24  
    brain computed tomography | -24  
    brain magnetic resonance imaging | -24  
    abdominal CT | -24  
    adrenal mass suggestive of pheochromocytoma | -24  
    treated with oral nifedipine | -24  
    treated with intravenous labetalol HCl | -24  
    treated with intravenous dexamethasone | -24  
    hypertensive encephalopathy | -24  
    transferred to our center | -24  
    born at 40 weeks of gestation | 0  
    no remarkable perinatal complications | 0  
    no medical history | 0  
    no treatment history | 0  
    family history of hyperthyroidism | 0  
    family history of thyroid cancer | 0  
    no headache | 0  
    no palpitation | 0  
    no diaphoresis | 0  
    weight gain 20 kg in past 10 months | -8760  
    pulse rate 110 beats/min | 0  
    blood pressure 170/110 mmHg | 0  
    respiratory rate 18 times/min | 0  
    body temperature 36.6℃ | 0  
    moon face | 0  
    central obesity | 0  
    Buffalo hump | 0  
    abdominal striae | 0  
    hirsutism | 0  
    height 125 cm | 0  
    weight 35 kg | 0  
    body mass index 23.04 kg/m² | 0  
    normal complete blood counts | 0  
    normal electrolytes | 0  
    normal liver function | 0  
    normal renal function tests | 0  
    fasting glucose 96 mg/dL | 0  
    hemoglobin A1c 5.7% | 0  
    proteinuria | 0  
    glycosuria | 0  
    urine calcium/creatinine ratio 0.23 | 0  
    normal electrocardiogram | 0  
    normal echocardiography | 0  
    normal kidney doppler ultrasonography | 0  
    abdominal CT showing 2.7 cm right adrenal mass | 0  
    tiny stone in right distal ureter | 0  
    abdominal MRI showing 3.3 cm right adrenal mass | 0  
    elevated 24-hour urinary free cortisol | 0  
    elevated midnight serum cortisol | 0  
    unsuppressed serum cortisol after low-dose DST | 0  
    undetectable plasma ACTH | 0  
    ruled out primary aldosteronism | 0  
    ruled out pheochromocytoma | 0  
    normal aldosterone/renin ratio | 0  
    normal plasma metanephrine | 0  
    normal plasma normetanephrine | 0  
    normal 24-hour urine metanephrine | 0  
    normal 24-hour urine normetanephrine | 0  
    complained of abdominal pain | after admission (assumed a few hours after admission, timestamp +24)  
    hematuria | +24  
    anuria | +24  
    abdominal CT showing bilateral distal ureter stones | +24  
    drowsy | +24  
    blood pressure not controlled | +24  
    oral losartan K | +24  
    spironolactone | +24  
    minoxidil | +24  
    intravenous nicardipine | +24  
    elevated blood urea nitrogen | +24  
    elevated creatinine | +24  
    transferred to ICU | +24  
    underwent CRRT | +24  
    preparation of ureteral stent indwelling | +24  
    fever developed | +24  
    elevated C-reactive protein | +24  
    broad-spectrum antibiotics administered | +24  
    started IV etomidate | +24  
    serum cortisol level monitored | +24  
    etomidate dose decreased | +24  
    IV hydrocortisone started | +24  
    serum cortisol maintained | +24  
    ureteral stent indwelling | +24  
    blood pressure improved | +24  
    discontinued losartan K | +24  
    discontinued minoxidil | +24  
    discontinued nicardipine | +24  
    improvement of oliguria | +24  
    renal function improved | +24  
    CRRT discontinued | +24  
    IV etomidate discontinued | +24  
    IV hydrocortisone increased | +24  
    underwent laparotomy | +24  
    resection of right adrenal mass | +24  
    adrenocortical adenoma confirmed | +24  
    surgery successful | +24  
    IV hydrocortisone changed to oral | +24  
    ureteral stones removed | +24  
    calcium carbonate apatite stones | +24  
    discharged | +24  
    replacement therapy with hydrocortisone | +24  
    <|eot_id|>
    
    6-year-old | 0
    boy | 0
    referred to our center | 0
    evaluation of an adrenal mass | 0
    visited the Emergency Department | -24
    generalized tonic-clonic type seizure | -24
    posterior reversible encephalopathy syndrome | -24
    hypertension | -24
    brain computed tomography | -24
    brain magnetic resonance imaging | -24
    abdominal CT | -24
    adrenal mass suggestive of pheochromocytoma | -24
    treated with oral nifedipine | -24
    treated with intravenous labetalol HCl | -24
    treated with intravenous dexamethasone | -24
    hypertensive encephalopathy | -24
    transferred to our center | -24
    born at 40 weeks of gestation | 0
    no remarkable perinatal complications | 0
    no medical history | 0
    no treatment history | 0
    family history of hyperthyroidism | 0
    family history of thyroid cancer | 0
    no headache | 0
    no palpitation | 0
    no diaphoresis |(concealed)
    weight gain 20 kg in past 10 months | -8760
    pulse rate 110 beats/min | 0
    blood pressure 170/110 mmHg | 0
    respiratory rate 18 times/min | 0
    body temperature 36.6℃ | 0
    moon face | 0
    central obesity | 0
    Buffalo hump | 0
    abdominal striae | 0
    hirsutism | 0
    height 125 cm | 0
    weight 35 kg | 0
    body mass index 23.04 kg/m² | 0
    normal complete blood counts | 0
    normal electrolytes | 0
    normal liver function | 0
    normal renal function tests | 0
    fasting glucose 96 mg/dL | 0
    hemoglobin A1c 5.7% | 0
    proteinuria | 0
    glycosuria | 0
    urine calcium/creatinine ratio 0.23 | 0
    normal electrocardiogram | 0
    normal echocardiography | 0
    normal kidney doppler ultrasonography | 0
    abdominal CT showing 2.7 cm right adrenal mass | 0
    tiny stone in right distal ureter | 0
    abdominal MRI showing 3.3 cm right adrenal mass | 0
    elevated 24-hour urinary free cortisol | 0
    elevated midnight serum cortisol | 0
    unsuppressed serum cortisol after low-dose DST | 0
    undetectable plasma ACTH | 0
    ruled out primary aldosteronism | 0
    ruled out pheochromocytoma | 0
    normal aldosterone/renin ratio | 0
    normal plasma metanephrine | 0
    normal plasma normetanephrine | 0
    normal 24-hour urine metanephrine | 0
    normal 24-hour urine normetanephrine | 0
    complained of abdominal pain | +24
    hematuria | +24
    anuria | +24
    abdominal CT showing bilateral distal ureter stones | +24
    drowsy | +24
    blood pressure not controlled | +24
    oral losartan K | +24
    spironolactone | +24
    minoxidil | +24
    intravenous nicardipine | +24
    elevated blood urea nitrogen | +24
    elevated creatinine | +24
    transferred to ICU | +24
    underwent CRRT | +24
    preparation of ureteral stent indwelling | +24
    fever developed | +24
    elevated C-reactive protein | +24
    broad-spectrum antibiotics administered | +24
    started IV etomidate | +24
    serum cortisol level monitored | +24
    etomidate dose decreased | +24
    IV hydrocortisone started | +24
    serum cortisol maintained | +24
    ureteral stent indwelling | +24
    blood pressure improved | +24
    discontinued losartan K | +24
    discontinued minoxidil | +24
    discontinued nicardipine | +24
    improvement of oliguria | +24
    renal function improved | +24
    CRRT discontinued | +24
    IV etomidate discontinued | +24
    IV hydrocortisone increased | +24
    underwent laparotomy | +24
    resection of right adrenal mass | +24
    adrenocortical adenoma confirmed | +24
    surgery successful | +24
    IV hydrocortisone changed to oral | +24
    ureteral stones removed | +24
    calcium carbonate apatite stones | +24
    discharged | +24
    replacement therapy with hydrocortisone | +24
    