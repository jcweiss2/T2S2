10 years old | 0
male | 0
pre-term | -4380
developmental delays | -4380
short stature | -2190
Russell–Silver syndrome | -2190
proteinuria | -2190
hypoalbuminemia | -2190
nephrotic syndrome | -2190
high-dose steroid | -2190
calcineurin inhibitor | -2190
renal function deteriorated | -2190
right renal vein thrombosis | -1096
pulmonary embolism | -1096
anticoagulants | -1096
persistent pulmonary hypertension | -1096
sildenafil | -1096
living donor kidney transplantation | 0
immunosuppression | 0
prednisolone | 0
mycophenolate mofetil (MMF) | 0
tacrolimus | 0
discontinued MMF | 70
steroid tapered | 70
tacrolimus continued | 70
pneumocystis pneumonia | 90
mechanical ventilation | 90
intravenous sulfamethoxazole/trimethoprim | 90
steroid increased | 90
dysuria | 135
gross hematuria | 135
blood urea nitrogen (BUN) 24 mg/dL | 135
creatinine (Cr) 0.56 mg/dL | 135
C-reactive protein (CRP) 0.42 mg/dL | 135
urinalysis | 135
red blood cell (RBC) count > 100/high power fields (HPF) | 135
white blood cell (WBC) count > 100/HPF | 135
urine culture for bacteria negative | 135
urine BK virus negative | 135
urine John Cunningham (JC) virus polymerase chain reaction (PCR) positive | 135
urine adenovirus culture positive | 135
hemorrhagic cystitis | 135
hydration | 135
pain control | 135
dysuria persisted | 142
hematuria persisted | 142
fever | 159
general weakness | 159
chest tightness | 159
mild cough | 159
persistent dysuria | 159
persistent hematuria | 159
BUN 175 mg/dL | 159
Cr 8.29 mg/dL | 159
CRP 30.23 mg/dL | 159
emergent hemodialysis | 159
piperacillin/tazobactam | 159
sputum culture negative | 159
blood culture negative | 159
urine culture negative | 159
adenovirus real-time PCR of sputum positive | 159
blood cytomegalovirus (CMV) antigen positive | 159
disseminated adenovirus infection | 159
immunosuppression reduction | 159
ganciclovir | 159
renal allograft biopsy | 159
diffuse necrotizing granulomatous tubulointerstitial nephritis | 159
infectious tubulointerstitial nephritis | 159
JC virus PCR positive | 159
serum CMV PCR positive | 159
coinfection | 159
ganciclovir targeting CMV | 159
antibiotic therapy | 159
granulocyte colony-stimulating factor | 159
immunoglobulin | 159
transfusion | 159
hemodialysis | 159
cidofovir | 167
nephrotoxicity | 167
renal impairment dose | 167
post-hematopoietic stem cell transplant adenovirus infection induction treatment | 167
on-going hemodialysis | 167
serum adenovirus PCR positive | 171
cerebrospinal fluid adenovirus PCR positive | 171
renal function not recovered | 171
generalized tonic-clonic seizure | 171
vancomycin | 171
meropenem | 171
acyclovir | 171
meningitis | 171
anemia | 171
leukopenia | 171
thrombocytopenia | 171
bone marrow suppression | 171
mechanical ventilation | 171
continuous renal replacement therapy | 171
deteriorated | 215
death | 215