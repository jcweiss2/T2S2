28 years old | 0
female | 0
admitted to the emergency department | 0
fever | -216
persistent cough | -216
fatigue | -216
progressive dyspnea | -216
end-stage kidney disease | 0
lupus nephritis Grade VI | 0
maintenance hemodialysis | 0
arteriovenous fistula | 0
hydroxychloroquine | 0
mycophenolic acid | 0
protected contact with sister | -168
wearing a surgical mask | -168
sister recovered from flu-like illness | -168
sister tested positive for COVID-19 | -168
sister asymptomatic | -168
decreased breath sounds | 0
crepitations at lung bases | 0
SpO2 88% on room air | 0
minor respiratory distress | 0
received 5L oxygen via nasal cannula | 0
desaturated further (SpO2 75%) | 0
septic shock | 0
intubated | 0
resuscitated with 500ml normal saline | 0
low dose noradrenaline | 0
mean arterial pressure 70 mm Hg | 0
electrocardiogram normal | 0
cardiac enzymes normal | 0
echocardiography normal | 0
lymphocytopenia | 0
increased C-reactive protein | 0
increased d-dimer | 0
increased lactate dehydrogenase | 0
increased ferritin | 0
blood urea nitrogen elevated | 0
creatinine elevated | 0
bilateral ground-glass opacities | 0
COVID-19 confirmed by RT-PCR | 0
admitted to ICU isolation chamber | 0
diagnostic work-up for infections | 0
evaluation for SLE flare | 0
no cutaneous manifestations of SLE | 0
no oral ulcers | 0
elevated anti-dsDNA | 0
decreased C3 complement | 0
decreased C4 complement | 0
no anti-cardiolipin antibodies | 0
no anti-β2GP1 antibodies | 0
no lupus anticoagulant | 0
no thrombocytopenia | 0
diagnostic dilemma between lupus pneumonitis and COVID-19 | 0
cultures derived for bacterial infections | 0
remained febrile | 0
bedside sonographic examination excluded deep vein thrombosis | 0
empiric therapy with lopinavir/ritonavir | 0
empiric therapy with ribavirin | 0
empiric therapy with piperacillin/tazobactam | 0
prophylactic anticoagulation | 0
hemodialysis every 48 hours | 0
supportive ICU care | 0
double lumen central line inserted for hemodialysis | 0
malfunctioning fistula | 0
SpO2/FiO2 ratio 150 | 72
ARDS-net ventilation | 72
prone positioning ventilation | 72
PEEP 10 cm H2O | 72
pulse methylprednisolone therapy initiated | 96
SpO2/FiO2 ratio increased to 300 | 96
vasopressors discontinued | 96
successfully extubated | 144
high flow nasal cannula | 144
SpO2 over 96% | 144
lymphocytes increased | 144
C-reactive protein decreased | 144
d-dimer decreased | 144
lactate dehydrogenase decreased | 144
ferritin decreased | 144
placed on 2L oxygen via nasal cannula | 192
no respiratory distress | 192
cultures negative for bacterial infections | 192
maintenance hemodialysis continued | 192
steroid therapy continued | 192
oxygen supportive care discontinued | 240
methylprednisolone tapered to 60mg/day | 240
RT-PCR test negative | 408
repeated microbiology tests negative | 408
discharged to home isolation | 456
maintenance oral steroid therapy | 456
followed-up by family physician | 456
