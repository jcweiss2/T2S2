16 years old | 0
male | 0
admitted to the hospital | 0
fever | 0
fatigue | 0
scleral icterus | 0
jaundice | 0
dark urine | 0
right abdominal pain | 0
right shoulder pain | 0
ulcerative colitis | -8760
corticosteroid-dependent course | -8760
acute exacerbations | -8760
aminosalicylates | -8760
immunomodulators | -8760
infliximab | -744
induction course of infliximab | -744
latest UC flare | -504
colonoscopy | -504
pancolitis | -504
IV corticosteroids | -504
infliximab | -504
alkaline phosphatase (ALP) | -504
leukocytosis | 0
anemia | 0
thrombocytopenia | 0
transaminitis | 0
aspartate aminotransferase (AST) | 0
alanine aminotransferase (ALT) | 0
hyperbilirubinemia | 0
C reactive protein (CRP) | 0
computed tomography (CT) | 0
multiple multi-loculated abscesses | 0
right hepatic lobe | 0
gas | 0
intrahepatic thrombosis | 0
right portal vein | 0
splenomegaly | 0
bilateral pleural effusions | 0
diffuse colonic wall thickening | 0
abscess drainage | 0
interventional radiology | 0
Peptostreptococci | 0
skin flora | 0
Escherichia coli | 0
acid-fast bacilli stain | 0
bacteremic | 0
Streptococcus viridans | 0
septic shock | 24
ICU management | 24
vancomycin | 24
meropenem | 24
ceftriaxone | 24
metronidazole | 24
repeat CT | 240
repeat CT | 480
amoxicillin-clavulanate | 720
discharged | 720
nasogastric tube | 720
exclusive enteral nutrition | 720
liver loculations improved | 4320
ultrasonography | 4320
normalization of liver enzymes | 4320
inflammatory markers | 4320
severe pancolitis | 7920
total colectomy | 7920
surgical gross pathology | 7920
moderately to severely active chronic pancolitis | 7920
mural abscesses | 7920
diffuse tan-red and hyperemic mucosa | 7920
scattered diffuse areas of ulceration | 7920
nodularity | 7920
pseudopolyps | 7920
ileum | 7920
appendix | 7920
ischemia | 7920
dysplasia | 7920
granulomas | 7920