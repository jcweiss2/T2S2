84 years old | 0
male | 0
admitted to the hospital | 0
right inguinal pain | -72
fever | -72
decreased appetite | -72
limited mobility | -72
obesity | 0
permanent atrial fibrillation | 0
apixaban | 0
chronic kidney disease stage IIIb | 0
distant repaired abdominal aortic aneurysm | 0
endovascular graft | 0
motor vehicle accident | -216
left knee hemarthrosis | -216
left lower limb cellulitis | -216
hypotensive | 0
blood pressure 95/61 mmHg | 0
borderline febrile to 37.8°C | 0
hypoxic | 0
oxygen saturation of 90% | 0
heart rate of 75/min | 0
weight on admission 114.4 kg | 0
alert and oriented | 0
cellulitis | 0
erythema | 0
previous hemarthrosis scar | 0
inoculation | 0
acute on chronic renal impairment | 0
creatinine 111 μmol/L | 0
albumin 32 g/L | 0
total bilirubin 18 μmol/L | 0
creatinine kinase 72 U/L | 0
aspartate aminotransferase 14 U/L | 0
alanine transferase 10 U/L | 0
white cell count 8.7 × 10^9/L | 0
neutrophil count 7.24 × 10^9/L | 0
lymphocytes 0.66 × 10^9/L | 0
pH 7.45 | 0
HCO3 22 mmol/L | 0
lactate 2.3 mmol/L | 0
C-reactive protein 95 mg/L | 0
C-reactive protein 150 mg/L | 48
Sequential Organ Failure Assessment score 3 | 24
intravenous flucloxacillin 2 g | 0
gentamicin 420 mg | 0
vancomycin 1 g | 0
IV crystalloid fluid resuscitation | 0
metaraminol infusion | 0
hypoxia improved | 72
blood cultures positive | 24
S. schleiferi ssp. coagulans identified | 24
urease and coagulase-positive testing | 24
piperacillin/tazobactam 4.5 g | 24
vancomycin 2 g loading dose | 24
vancomycin 1 g twice daily | 24
antimicrobials rationalized to IV flucloxacillin | 48
transthoracic and transesophageal echocardiography | 48
CT-position emission tomography | 72
moderate focal FDG uptake | 72
exposure to unwell pet Maltese terrier's otorrhea | -168
canine otitis externa | -168
topical 23 mg/mL miconazole nitrate | -168
5 mg/mL prednisolone acetate | -168
0.696 mg/mL polymyxin B | -168
ocular and lower limb exposure | -168
canine aural samples posttreatment tested positive | -168
Staphylococcus intermedius group | -168
vascular surgical opinion | 72
indefinite antimicrobial suppression | 72
oral flucloxacillin 1 g twice a day | 72
6-week course of IV flucloxacillin 2 g 4 h | 72
pulmonary edema | 120
diuresis with daily furosemide | 120
discharged | 168
outpatient parental antimicrobial therapy | 168
oral antimicrobial suppression | 168