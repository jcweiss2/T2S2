92 years old | 0
female | 0
hypertension | -672
atrial fibrillation | -672
dementia with Lewy bodies | -672
falls at home | -672
sick sinus syndrome | -672
bradycardia | -672
pacemaker implantation | -672
orthostatic hypotension | -672
admitted to acute geriatric unit | 0
transferred to geriatric rehabilitation care unit | 24
rabeprazole | 24
mianserin | 24
right leg wound | 24
no fever | 24
no inflammation | 24
local antiseptic dressings | 24
daily monitoring | 24
fever | 672
erythema | 672
edema of right leg | 672
lymphangitis | 672
dermohypodermitis diagnosis | 672
intravenous amoxicillin | 672
venous Doppler performed | 672
no thrombosis | 672
injury extension to entire lower limb | 672
purplish discoloration of skin | 672
bullae | 672
necrosis | 672
severe pain | 672
morphine administration | 672
limited leg movements | 672
necrotizing fasciitis | 672
blood cultures performed | 672
empiric broad-spectrum antibiotic therapy | 672
switched to piperacillin | 672
switched to tazobactam | 672
switched to gentamicin | 672
blood pressure 93/50 mmHg | 672
heart rate 91 bpm | 672
body temperature 34.3°C | 672
respiratory rate 32 bpm | 672
oxygen saturation 84% | 672
reduced consciousness | 672
distended abdomen | 672
dyspnea | 672
computed tomography scan | 672
no pneumoniae | 672
no abdominal infection | 672
no pelvic infection | 672
white cell count 4.6 cells/mm3 | 672
hemoglobin 13.0 g/dL | 672
platelet count 15.1×104 cells/mm3 | 672
C-reactive protein 70 mg/dL | 672
blood glucose 1.4 mmol/L | 672
procalcitonin 43 ng/mL | 672
troponin 3.73 μg/L | 672
pH 7.19 | 672
HCO3 14.4 mmol/L | 672
blood lactate 9.0 mmol/L | 672
urine analysis no infection | 672
septic shock | 672
fluid challenge | 672
extension of necrotic disease | 672
precarious medical condition | 672
transfer to La Pitié Salpêtrière Hospital | 672
surgical debridement | 672
mechanical ventilation | 672
inotropic support | 672
antibiotic administration | 672
death | 672
K. pneumoniae identified | 672
hypermucoviscous colonies | 672
positive string test | 672
resistance to amoxicillin | 672
resistance to piperacillin | 672
resistance to ticarcillin | 672
K2 serotype | 672
RmpA present | 672
aerobactin present | 672
yersiniabactin present | 672
ST86 sequence type | 672
