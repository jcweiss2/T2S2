81 years old | 0
male | 0
admitted to the hospital | 0
ischemic stroke | -8760
hypertension | -8760
stable stage 3 nephropathy | -8760
multiple myeloma type IgA lambda | -8760
symptomatic anemia | -730
monoclonal gammaglobulinemia | -730
treatment with melphalan | -730
treatment with prednisone | -730
treatment with bortezomib | -730
disease progression | -730
treatment with lenalidomide | -730
treatment with dexamethasone | -730
dyspnea | 0
general discomfort | 0
muscle weakness | 0
poor performance status | 0
tachypnea | 0
normal body temperature | 0
normal blood pressure | 0
no clinical signs of pneumonia | 0
no clinical signs of cardiac decompensation | 0
respiratory compensated metabolic acidosis | 0
increased anion gap | 0
elevated arterial lactate level | 0
lactic acidosis | 0
type B lactate acidosis | 0
metastatic prostate cancer | 0
elevated PSA level | 0
enlarged prostate | 0
hydronephrosis of the right kidney | 0
small nodules in the liver | 0
enlarged mediastinal and paratracheal lymph nodes | 0
sclerotic bone metastases | 0
treatment with cyproterone acetate | 24
treatment with prednisone | 24
treatment with thiamine | 24
clinically deteriorated | 24
increasing lactate levels | 24
lowering pH levels | 24
unconscious | 48
admitted to the ICU | 48
received NaHCO3 | 48
adrenaline-resistant cardiac arrest | 72
DNR will | 72
no resuscitation | 72
autopsy | 72
locally advanced and metastatic prostate cancer | 72
Gleason score 5 + 5 = 10 | 72
encasement of the right ureter | 72
metastases in the thoracic and lumbar spine | 72
metastases in the liver | 72
metastases in the lungs | 72
metastases in the peritoneum | 72
bilateral tumor thrombi | 72
no signs of activity of multiple myeloma | 72
no signs of cardiac ischemia | 72
frameshift mutation in exon 8 of the TP53 gene | 72
activating mutation in exon 10 of the PIK3CA gene | 72
no mutations in PTEN and IDH1 | 72