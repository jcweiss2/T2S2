55 years old | 0
male | 0
trivial fall | -720
severe back pain | -720
analgesics | -720
bed rest | -720
relieved pain | -720
increased back pain | -60
incapacitated | -60
persistent back pain | 0
restriction of movements | 0
gibbus at the thoracolumbar junction | 0
spasm of the para-spinal muscles | 0
restricted and painful movements of the spine | 0
normal motor power | 0
normal sensation | 0
intact reflexes | 0
normal bladder function | 0
normal bowel function | 0
anorexia | 0
loss of weight | 0
well-controlled type-2 diabetic | 0
oral medications for diabetes | 0
no other medication | 0
no allergy | 0
good cardiac status | 0
good pulmonary status | 0
no other constitutional symptoms | 0
surgical fixation of the fracture of humerus | -8760
uneventful postoperative recovery | -8760
no history of childhood illnesses | 0
slightly raised C-reactive protein | 0
raised erythrocyte sedimentation rate | 0
high normal white cell count | 0
normal bone profile | 0
normal renal function test | 0
normal liver function test | 0
compression fracture of the T12 vertebra | 0
marrow edema | 0
evidence suggestive of fluid in the fracture site | 0
normal cord | 0
normal signal intensity from the intervertebral discs | 0
prevertebral soft-tissue swelling | 0
epidural soft-tissue component indenting the anterior dural sac | 0
dual-energy X-ray absorptiometry scan | 0
osteopenic | 0
T-score of -2 | 0
computed tomography scan of the T12 vertebra | 0
intact posterior cortex | 0
transpedicular biopsy | 0
kyphoplasty | 0
general anaesthesia | 0
prone position | 0
Relton Hall frame | 0
transpedicular biopsy needles | 0
image control | 0
minimal resistance | 0
no material on aspiration | 0
saline injection | 0
aspiration | 0
sero-sanguineous material mixed with pus | 0
microbiology | 0
cytology | 0
fluid analysis | 0
deferred kyphoplasty | 0
supine position | 0
extubation | 0
severe bronchospasm | 0
decrease in saturation | 0
intubation | 0
arterial blood gas analysis | 0
severe respiratory acidosis | 0
pH 7.16 | 0
PaCO2 72 mm Hg | 0
PaO2 82 mm Hg | 0
bilateral multiple lung infiltrates | 0
mechanical ventilation | 0
intensive care unit | 0
intravenous vancomycin | 0
improved | 24
weaned off from the ventilator | 24
endo-tracheal tube detached | 24
high dependency unit | 24
clear chest | 72
resolution of infiltrates | 72
culture report | 72
Staphylococcus aureus | 72
sensitive to imipenum and linezolid | 72
intravenous linezolid | 72
oral administration | 120
thoracolumbar orthosis | 0
protected spine | 0
recovered uneventfully | 168
CRP and ESR returned to normal | 168
symptom free | 4320