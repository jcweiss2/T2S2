73 years old | 0
    woman | 0
    Ecuadorian indigenous ancestry | 0
    evaluated in the emergency department | 0
    intense and diffuse colicky abdominal pain | -48
    abdominal distension | -48
    inability to eliminate flatus | -48
    hypothyroidism | -175200
    conventional cholecystectomy | -175200
    no prior history of colitis | -175200
    no prior history of gastrointestinal disease | -175200
    increased polymerase chain reaction | 0
    no leukocytosis | 0
    no neutrophilia | 0
    no acidosis | 0
    mild hypokalemia | 0
    obstructive abdomen | 0
    simple tomography of abdomen and pelvis | 0
    contrast-enhanced tomography of abdomen and pelvis | 0
    no transition zone | 0
    no pneumoperitoneum | 0
    small amount of fluid in Douglas sac | 0
    stool studies did not show parasites | 0
    stool studies did not show blood | 0
    non-surgical medical treatment initiated | 0
    analgesia | 0
    bowel rest | 0
    hydration | 0
    clinical improvement | 72
    oral route restarted | 96
    gastrointestinal disturbances recurred | 96
    pain | 96
    distension | 96
    inability to eliminate flatus | 96
    colonoscopy performed | 168
    mucosal patches | 168
    erosions | 168
    edema localized at sigmoid | 168
    edema localized at descendant colon | 168
    edema localized at transverse colon | 168
    lesions biopsied | 168
    sent to pathology | 168
    sent to microbiology | 168
    ulceration of epithelium | 168
    lymphoplasmacytic infiltration | 168
    eosinophiles | 168
    congestion | 168
    hemorrhage | 168
    parasitic bodies with phagocyted red blood cells | 168
    serum antibodies against E. histolytica | 168
    negative | 168
    metronidazole started | 168
    gradual worsening abdominal distension | 336
    gradual worsening pain | 336
    feeding intolerance | 336
    persistent mild hypokalemia | 336
    normal renal function | 336
    normal liver function | 336
    down trending leukocytes | 336
    repeat abdominal tomography | 336
    pneumoperitoneum | 336
    colonic perforation | 336
    exploratory laparotomy conducted | 336
    fecal peritonitis | 336
    pneumoperitoneum | 336
    phlegmonous descending colon | 336
    massive colon dilation | 336
    multiple transmural perforations in sigma | 336
    multiple transmural perforations in descending colon | 336
    multiple transmural perforations in transverse colon | 336
    total colectomy | 336
    ileostomy | 336
    rectal stump closure | 336
    no surgical complications | 336
    hypotension | 360
    sepsis | 360
    managed in intensive care unit | 360
    fluids | 360
    vasoactive drugs | 360
    post-operative antimicrobial treatment | 360
    meropenem | 360
    metronidazole IV | 360
    metronidazole PO | 360
    tinidazole | 360
    superficial surgical site infection | 408
    multiresistant organisms | 408
    carbapenem-resistant Klebsiella pneumoniae | 408
    extended spectrum beta-lactamase producing Escherichia coli | 408
    treated with colistin | 408
    wound opened | 408
    heal by secondary intention | 408
    serial dressing changes | 408
    discharged | 720
    mucosal ulceration throughout entire colon | 336
    submucosa involvement | 336
    significant edema | 336
    congestion | 336
    inflammatory infiltrate | 336
    lymphocytes | 336
    plasmocytes | 336
    eosinophils | 336
    macrophages | 336
    necrotic areas | 336
    granulation tissue | 336
    E. histolytica trophozoites loaded with red blood cells | 336

