44 years old | 0
male | 0
admitted to the hospital | 0
rash | -72
vesicle on the left side of his forehead | -72
headache | -144
fever | -72
diagnosed with HZO | -72
treated with antiviral drugs | -72
treated with analgesics | -72
continuous fever | -72
worsening of left-sided frontal headache | -24
nausea | -24
blurred vision | -24
diplopia | -24
transferred to the hospital | 0
alert | 0
febrile | 0
crust on his forehead | 0
normal cardiopulmonary findings | 0
normal neurological findings | 0
heart rate 78 beats/min | 0
blood pressure 110/60 mmHg | 0
respiratory rate 20 breaths/min | 0
visual acuity 6/12 bilaterally | 0
no abnormalities in the ocular tissues | 0
no visual field defects | 0
horizontal diplopia | 0
lateral rectus muscle paresis in the left eye | 0
6th cranial nerve palsy | 0
no evidence of infection | 0
white blood cell count normal | 0
erythrocyte sedimentation rate elevated | 0
C-reactive protein level elevated | 0
blood culture performed | 0
brain MRI revealed lateral bulging and irregular marginal enhancement in the cavernous sinus | 0
admitted to the intensive care unit | 0
treated with second-generation cephalosporin | 0
Streptococcus constellatus subsp. constellatus detected in the blood culture | 24
switched to clindamycin | 24
echocardiography performed | 24
antithrombotic therapy with low molecular weight heparin | 24
symptoms improved | 168
discharged | 168
dental treatment | -216
pain in the left maxillary area | -96
follow-up for one year | 720