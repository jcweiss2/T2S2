35 years old | 0
    morbidly obese | 0
    woman | 0
    alcohol use disorder | 0
    admitted | 0
    decreased urine output | 0
    anasarca | 0
    presumed alcoholic cirrhosis | 0
    acute kidney injury | 0
    creatinine 2.9 | 0
    baseline creatinine 1.1 | 0
    normal creatinine 0.5-1.2 mg/dL | 0
    liver dysfunction | 0
    MELD score 32 | 0
    estimated 52.6% 3-month mortality rate | 0
    shock | 0
    transfer to medical intensive care unit | 0
    initiation of hemodialysis | 0
    initiation of vasopressors | 0
    initiation of broad-spectrum antibiotics | 0
    weaned off vasopressors | 504
    purpuric plaques on bilateral lower extremities | 504
    physical examination of bilateral, lateral, and medial thighs | 504
    greater than 20-cm retiform purpuric plaques | 504
    central necrotic eschar | 504
    surrounding indurated stellate red-brown plaques | 504
    hyperpigmented plaque on abdomen | 504
    peau d'orange on abdomen | 504
    normal calcium | 504
    hypo-albuminemia corrected calcium 10.0 | 504
    normal calcium 8.8-10.2 mg/dL | 504
    normal parathyroid hormone 61.1 | 504
    normal parathyroid hormone 10-69 pg/mL | 504
    low phosphorus 2.0 | 504
    normal phosphorus 2.5-4.5 mg/dL | 504
    excisional biopsy | 504
    calcification within small vessels | 504
    calcification between adipocytes | 504
    fat necrosis | 504
    consistent with calciphylaxis | 504
    treatment with intravenous sodium thiosulfate | 504
    titrated to 25 g/d | 504
    received vitamin K | 504
    received pentoxifylline | 504
    received 1 dose of zoledronic acid | 504
    persistence of necrotic eschars | 504
    medical maggot therapy initiated | 504
    maggot larvae applied to right lateral thigh | 504
    maggots enclosed with mesh | 504
    maggots began debriding necrotic tissue | 504
    debridement planned for 48 to 72 hours | 504
    serosanguinous oozing occurred | 504
    maggots removed after 24 hours | 504
    right thigh showed debridement | 504
    3-cm-deep concavity | 504
    palpably hollowed eschar | 504
    discontinued maggot therapy | 528
    massive hemorrhage from right lateral thigh | 576
    hemorrhage resolved with pressure and suture ligation | 576
    8 units of blood transfused | 576
    hemorrhagic shock | 576
    subcutaneous heparin discontinued | 576
    bled intermittently from deep wounds | 576
    bleeding controlled with pressure dressings | 576
    continued treatment with STS | 576
    continued treatment with vitamin K | 576
    continued treatment with pentoxifylline | 576
    skin improved clinically | 576
    no new lesions developed | 576
    existing indurated plaques softened | 576
    renal function recovered | 576
    hemodialysis discontinued | 576
    maggot therapy | 576
    placement of percutaneous gastrostomy tube | 672
    pneumoperitoneum | 672
    septic shock | 672
    patient died | 672
    