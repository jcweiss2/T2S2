33 years old | 0
female | 0
pregnant | 0
11th week of gestation | 0
admitted to the hospital | 0
high fever | 0
lower back pain | 0
intravenous antibiotic treatment | 0
pyelonephritis | 0
platelet count decreased | 0
disseminated intravascular coagulation | 48
sepsis | 48
body temperature 40°C | 48
tachycardia | 48
systolic murmur | 48
transthoracic echocardiography | 48
severe mitral valve regurgitation | 48
blood cultures grew MSSA | 48
intravenous gentamicin | 48
intravenous teicoplanin | 48
recombinant human soluble thrombomodulin not used | 48
inflammatory markers showed gradual improvement | 48
clinical condition worsened | 192
high-dose diuretic | 192
inotropic support | 192
noninvasive positive pressure ventilation | 192
mitral valve destruction | 192
minimally invasive thoracoscopic mitral valve repair | 240
fetal heart rate showed no abnormalities | 240
routine evaluation | 240
rapid sequence induction of anesthesia | 240
intravenous propofol | 240
rocuronium bromide | 240
fentanyl | 240
tracheal intubation | 240
general anesthesia | 240
target propofol concentration | 240
oxygen-air mixture | 240
remifentanil | 240
standard radial artery catheter | 240
Swan–Ganz catheter | 240
bispectral index | 240
cerebral oximetry monitoring | 240
intraoperative transesophageal echocardiography | 240
severe MR | 240
rupture of the chordae tendineae | 240
hypothermic CPB | 240
pump flow rate | 240
maternal uteroplacental perfusion | 240
fetal monitoring | 240
abdominal and transvaginal Doppler flow ultrasound | 240
successful repair | 240
weaned off the CPB | 348
inotropic support | 348
tracheal tube extubated | 348
postoperative condition favorable | 348
transvaginal ultrasound | 348
fetal heart rate | 348
hydrops fetalis | 432
dilation and curettage | 432
blood cultures did not detect bacterial growth | 480
antibiotics administered | 480
total of 8 weeks | 672