37 years old | 0
male | 0
admitted to the abdominal surgery department | 0
pain | 0
open postoperative wound in the left subcostal area | 0
multiple enterocutaneous fistulas | 0
daily output of up to 2000 ml of gastric and enteric contents | 0
high-degree obesity (BMI 48 kg/m²) | -120
many unsuccessful efforts of weight loss | -120
bariatric surgery—distal gastrectomy | -120
Roux-en-Y gastric bypass with Braun anastomosis | -120
Shalimov plug (staple line on proximal intestine) | -120
adhesive small bowel obstruction | -792
emergency surgery (relaparotomy, adhesiolysis, nasointestinal intubation) | -792
gastroenteroanastomosic leakage | -672
peritonitis | -672
surgical wound dehiscence | -672
total parenteral nutrition | -672
fistuloclysis | -672
daily fistula output about 2000 ml | -672
complex non-surgical treatment | -672
condition stabilized | -672
surgical fistula closure (suturing a fistula in a wound) | -504
fever of 38.7°C | -504
bowel content appeared in the wound | -504
surgical wound dehiscence | -504
fistula output increased to 2000 ml per day | -504
emergency relaparotomy in the left subcostal area | -480
bypass gastroenterostomy | -480
septic shock | -480
multiple enteroatmospheric fistulas | -480
output of bowel content up to 2500 ml per day | -480
abdominal wall phlegmon in the left subcostal area | -480
emergency relaparotomy | -432
collateral enteroenteric anastomosis | -432
fistula output did not decrease | -432
transferred to our clinic | -360
weight loss of 55 kg | -360
abdominal wall wound of irregular shape 15×10 cm | 0
rough edges in epigastrium | 0
wound edges covered with fresh granulation tissue | 0
wound bottom formed by small bowel loops | 0
enterocutaneous fistula 2.5 cm diameter | 0
enterocutaneous fistula 1 cm diameter with Kehr’s T-tube | 0
removed Kehr’s T-tube during wound revision | 0
gastroenteric anastomosis leakage with enteral feeding tube | 0
two small bowel lumens filled with enteric contents with bile | 0
recess anterior abdominal wall | 0
drainage tube through a counterincision | 0
skin inflamed, macerated, hyperemic | 0
small bowel contents actively aspirated | 0
total fistula output 1500 ml per day | 0
anemia (Hb 87 g/L) | 0
hypoproteinemia (total protein 55 g/L) | 0
hypoalbuminemia (albumin 32 g/L) | 0
hypokalemia (K 2.9 mmol/L) | 0
hyperlactatemia (lactate 2.3 mmol/L) | 0
elevated fibrinogen (5.1 g/L) | 0
CT chest, abdomen, pelvis: pulmonary embolism | 0
free fluid in left pleural cavity | 0
atelectasis of basal segment of left lung | 0
defect of abdominal wall with destruction of VIII-X ribs | 0
gastroatmospheric fistula | 0
thrombosis of left common femoral vein | 0
hepatomegaly | 0
liver steatosis | 0
free liquid in abdomen and pelvis | 0
fistulography with contrast | 0
gastroenteroanastomosis leakage identified | 0
intensive care management | 0
electrolyte imbalance correction | 0
sepsis control | 0
nutritional support (TPN, fistuloclysis) | 0
therapy of thromboembolic complications | 0
wound treatment | 0
active aspiration of gastric and bowel contents | 0
skin protection | 0
nasogastric tube aspiration | 0
complex non-operative management | 0
reconstructive surgery (laparotomy, distal gastrectomy, etc.) | 720
midline laparotomy | 720
adhesiolysis | 720
three entero-enteric anastomoses | 720
enterocutaneous fistulas resected | 720
Roux-gastrojejunostomy | 720
transversostomy | 720
resection of small bowel with fistulas | 720
colostomy closure | 720
transversodescendostomy | 720
total parenteral nutrition for 5 days | 720
infusion therapy | 720
secretion suppression | 720
thromboembolic prevention | 720
daily wound dressing | 720
wound healed | 720
sutures removed on day 15 | 720
discharged home on day 21 | 720
uneventful recovery | 720
laparotomy, adhesiolysis, colostomy closure | 8760
transversodescendostomy | 8760
discharged home on day 9 | 8760
satisfactory quality of life | 8760
pulmonary embolism | 0
no fresh infarct pneumonia | 0
gastroenteroanastomosis leakage identified via fistulogram | 0
active aspiration via drainage tube | 0
Foley tube for fistuloclysis | 0
postoperative wound dehiscence | -672
postoperative wound dehiscence | -504
postoperative wound dehiscence | -480
postoperative wound dehiscence | -432
postoperative wound dehiscence | 0
postoperative wound dehiscence | 720
postoperative wound dehiscence | 8760
