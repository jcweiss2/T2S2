66 years old | 0 | 0 
male | 0 | 0 
admitted to the hospital | 0 | 0 
intermittent high-grade fever | -216 | 0 
generalized dull-aching abdominal pain | -216 | 0 
passing turbid urine | -240 | -216 
decrease in urine output | -240 | -216 
swelling of both feet | -240 | -216 
treated with intravenous medications | -168 | -168 
type II diabetes mellitus | -2628 | 0 
on regular medication for diabetes | -2628 | 0 
conscious | 0 | 0 
afebrile | 0 | 0 
tachycardic | 0 | 0 
heart rate of 136/min | 0 | 0 
blood pressure was 110/70 mmHg | 0 | 0 
renal angle tenderness bilaterally | 0 | 0 
high total leukocyte counts | 0 | 0 
elevated urea and creatinine levels | 0 | 0 
pyuria with leukocyte esterase positivity | 0 | 0 
activated partial thromboplastin time was prolonged | 0 | 0 
sepsis-induced coagulopathy | 0 | 0 
enlarged kidneys with bilateral renal abscesses | 0 | 0 
emergency ultrasound-guided drainage of renal abscesses | 24 | 24 
transfusion of blood products | 24 | 24 
pus smear from renal abscesses showed septate fungal hyphae | 24 | 24 
intravenous meropenem | 0 | 24 
intravenous voriconazole | 24 | 24 
intravenous amphotericin B | 48 | 216 
cultures from both renal abscesses revealed growth of Aspergillus fumigatus | 48 | 48 
worsening renal function | 72 | 216 
acute pulmonary edema | 120 | 216 
hyperkalemia | 120 | 216 
metabolic acidosis | 120 | 216 
hemodialysis | 144 | 216 
noninvasive ventilation | 144 | 216 
sudden cardiac arrest | 216 | 216 
aspiration | 216 | 216 
succumbed to his illness | 216 | 216