42 years old | 0
female | 0
admitted to the hospital | 0
juvenile idiopathic arthritis | -37800
anakinra | -10950
hydroxychloroquine | -8760
chronic adrenal insufficiency | -37800
hydrocortisone | -37800
seizure disorder | -37800
culture negative infective endocarditis | -10080
cardioembolic stroke | -10080
mechanical fall | -24
C7 vertebral fracture | 0
acute on chronic hypoxic and hypercapnic respiratory failure | 0
rescue BiPAP support | 0
admission to the intensive care unit | 0
encephalopathic | 0
respiratory acidosis | 0
carbon dioxide retention | 0
intubated | 0
computed tomography thorax | 0
left-sided opacification | 0
left-sided pneumonia | 0
diaphragmatic weakness | 0
tracheotomy | 312
percutaneous endoscopic gastrostomy | 312
subarachnoid hemorrhage | -720
comminuted fracture of the distal left tibia | -720
progressive muscular weakness | -8760
elevated serum aldolase | 0
normalized serum aldolase | 96
elevated thyroid-stimulating hormone | 0
normal free thyroxine | 0
elevated alanine aminotransferase | 0
elevated aspartate aminotransferase | 0
normal bilirubin | 0
chronically low creatinine | 0
rheumatology consultation | 0
diaphragmatic weakness | 0
muscle biopsy | 0
myopathy | 0
electron microscopy | 0
abnormal autophagosomes | 0
curvilinear bodies | 0
hydroxychloroquine-induced myopathy | 0
discontinuation of hydroxychloroquine | 0
recovery | 576
steroid-induced myopathy | 0
type II fiber atrophy | 0
CIDP | 0
critical illness myopathy | 0
inflammatory myopathy | 0
discontinuing hydroxychloroquine | 0
reducing dose of steroids | 0