40 years old | 0
female | 0
admitted to the hospital | 0
high-grade fever | -48
myalgia | -48
nausea | -48
right hypochondriac pain | -48
diagnosed with COVID 19 | -336
hypertension in father | 0
no previous history of any chronic disease | 0
no medications | 0
no allergy | 0
no psychological illness | 0
fever | 0
generalized body aches | 0
mild tenderness on the right hypochondrium | 0
positive Murphy's sign | 0
no jaundice | 0
no scratch marks on the body | 0
high white cell count | 0
increased neutrophils | 0
elevated inflammatory markers | 0
C-reactive protein (CRP) | 0
D-dimers | 0
ferritin | 0
interleukins | 0
bilateral lower lung patchy pulmonary consolidations | 0
left-sided-pleural effusion | 0
thickened gall bladder wall | 0
surrounding pericholecystic fluid | 0
minimal free fluid in the abdomen and the pelvis | 0
acalculous cholecystitis | 0
broad spectrum antibiotics | 0
IV Piperacillin Tazobactum | 0
azithromycin | 0
hypotensive | 12
resuscitated with IV fluids | 12
ICU care | 12
no mechanical intubation | 12
inconclusive COVID real-time reverse transcriptase (Rrt-PCR) | 12
normotensive | 24
high-grade fever | 24
CT abdomen | 24
bilateral pleural effusion | 24
consolidation | 24
ground-glass opacities | 24
atelectasis | 24
no intra-abdominal collection | 24
IV meropenem | 24
fever settled | 48
stable | 216
discharged | 216
follow-up | 744
no symptoms | 744
stable throughout follow up period | 744