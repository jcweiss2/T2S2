40 years old | 0
male | 0
admitted to the hospital | 0
new-onset uncontrolled seizures | 0
unresponsive | 0
intubated | 0
sedated | 0
status epilepticus | 0
treated with anticonvulsants | 0
admitted to the neurological critical care unit | 0
no significant past medical history | 0
lived and worked in swimming pool maintenance | 0
had not traveled outside of the state | 0
experienced progressively worsening migraines | -720
migraines refractory to pharmacologic therapy | -720
nausea | -720
vomiting | -720
intermittent neck stiffness | -720
decreased appetite | -720
unintentional weight loss | -720
presented to an outside hospital | -192
complaining of severe headaches | -192
photophobia | -192
neck and back pain | -192
slurred speech | -192
tremors | -192
drooling | -192
left facial droop | -192
imaging returned negative | -192
symptoms attributed to migraine headache | -192
discharged home | -192
noncontrast computed tomography (CT) imaging of his head and spine | 0
unremarkable | 0
elevated white blood cell (WBC) count | 0
electroencephalogram | 0
moderate to severe diffuse slowing | 0
lumbar puncture (LP) | 0
mildly elevated opening pressure | 0
low glucose | 0
elevated protein | 0
elevated WBCs | 0
vancomycin and piperacillin-tazobactam administered | 0
Gram stain | 0
India Ink stain | 0
cerebrospinal fluid (CSF) demonstrated encapsulated, variably sized yeast cells | 0
BioFire FilmArray Meningitis/Encephalitis Panel | 0
positive for Cryptococcus neoformans/Cryptococcus gattii | 0
CrAg LFA cryptococcal antigen tests | 0
positive on both CSF and serum | 0
empiric antibiotics exchanged with intravenous amphotericin B | 24
flucytosine | 24
cerebrospinal fluid cultures grew C gattii | 24
identified by matrix-assisted laser desorption ionization time-of-flight mass spectrometry | 24
produced the characteristic blue color on l-canavanine, glycine, 2-bromothymol blue (CGB) agar | 24
multilocus sequence typing | 24
genotype was VGI | 24
remained unresponsive | 24
worsening fevers | 24
shivering | 24
neck stiffness | 24
thoracic CT | 48
left lung consolidation | 48
bronchoalveolar lavage | 48
infectious diseases consultants recommended continuation of antifungal therapy | 48
serial LP | 48
thorough evaluation of the patient’s immune status | 48
LP repeated 4 more times | 72
opening pressures of >55 cmH2O | 72
persistently elevated protein | 72
decreased glucose | 72
elevated leukocyte counts | 72
no evidence of immunocompromised state | 72
negative human immunodeficiency virus (HIV) 1/2 Ag-antibody (Ab) | 72
hepatitis A/B/C panel | 72
QuantiFERON-TB Gold | 72
alpha-1-antitrypsin | 72
antimitochondrial Ab | 72
antinuclear Ab assays | 72
immunoglobulin (Ig) panel | 72
normal IgA | 72
mildly decreased IgG | 72
mildly decreased IgM | 72
normal CD4/CD8 ratio | 72
mildly decreased absolute lymphocyte count | 72
absence of lymphoproliferation or leukemia | 72
normal CSF angiotensin-converting enzyme | 72
reduced absolute CD4 | 72
reduced absolute CD8 | 72
reduced IgG | 72
reduced IgM | 72
serial magnetic resonance imaging (MRI) | 96
symmetric cortical and subcortical diffusion restriction | 96
leptomeningeal enhancement | 96
hemorrhagic transformation of the left posterior parietal lobe | 96
focal areas of restricted diffusion in the right upper cervical spinal cord | 96
remained unable to follow commands | 120
neurological status decompensated | 120
eye-opening to purposeful withdrawal from pain | 120
abnormal decerebrate posturing | 120
compromise of brainstem reflexes | 120
discharged to inpatient hospice | 336
died | 336
autopsy performed | 336
extensive granulomatous meningitis | 336
numerous cryptococcal organisms | 336
diffuse bilateral cerebral cortical infarcts | 336
hemorrhage in the left posterior parieto-occipital region | 336
small infarct in the cervical spinal cord | 336
large cryptococcoma in the upper lobe of the left lung | 336
rare cryptococcal organisms diffusely present throughout bilateral lungs | 336
cause of death determined to be from complications of disseminated cryptococcosis | 336
cryptococcal meningitis | 336