63 years old | 0
male | 0
164 cm | 0
79 kg | 0
admitted to the hospital | 0
left hip fracture | -10
tibia fracture | -10
road traffic accident | -10
transsphenoidal approach operation | -4380
panhypopituitarism | -4380
diabetes mellitus | -4380
mild dyspnea | -10
arterial blood gas analysis | -10
pH 7.423 | -10
PaCO2 37.3 mmHg | -10
PaO2 50.1 mmHg | -10
SaO2 86.5% | -10
FiO2 0.2 | -10
alveolar-arterial oxygen gradient increased | -10
chest x-ray normal | -10
dyspnea worsened | -72
hypoxemia worsened | -72
chest computed tomography | -72
thromboembolism in the right interlobar pulmonary artery | -72
thromboembolism in the right lower lobe segmental artery | -72
thromboembolism in the subsegmental pulmonary artery | -72
heparin treatment initiated | -72
dyspnea improved | -72
hypoxemia improved | -72
transthoracic echocardiography | -96
no abnormality or thrombus | -96
left lower limb venography | -120
no venous thrombus | -120
inferior vena cava filter not inserted | -120
operation scheduled | -120
heparin stopped | -24
prothrombin time normal | 0
activated partial thromboplastin time normal | 0
BUN/Cr increased | 0
patient not premedicated | 0
standard monitoring devices applied | 0
Allen's test | 0
left radial artery cannulated | 0
initial blood pressure 120/70 mmHg | 0
5 L of 100% O2 applied | 0
initial arterial blood gas analysis | 0
pH 7.43 | 0
PaCO2 38.1 mmHg | 0
PaO2 102.9 mmHg | 0
SaO2 98% | 0
spinal anesthesia administered | 0
tetracaine administered | 0
epinephrine administered | 0
sensory block to T10 confirmed | 5
Hartmann's solution administered | 5
no significant changes in BP or heart rate | 5
pneumatic tourniquet inflated | 40
hypotension | 40
cardiac arrest | 40
cardiopulmonary resuscitation instituted | 40
transesophageal echocardiography | 40
multiple emboli in the right atrium | 40
interatrial septum bulging into the left atrium | 40
epinephrine administered | 40
atropine administered | 40
norepinephrine administered | 40
sodium bicarbonate administered | 40
vital signs improved | 55
operation resumed | 55
patient transferred to ICU | 135
mechanical ventilation continued | 135
heparin treatment initiated | 135
D-dimer 9467 ng/ml | 135
D-dimer increased to 52,796 ng/ml | 216
PaO2 improved | 216
patient extubated | 216
heparin treatment continued | 480
D-dimer decreased | 480
chest CT and echocardiography normal | 480
patient transferred to general ward | 720