47 years old | 0
woman | 0
presented to the emergency department | 0
weakness | 0
numbness of the limbs | 0
nausea | 0
fatigue | 0
dyspnea | 0
fever | -168
cough | -168
acute upper respiratory infection | -168
influenza virus A | -168
weakness | -120
numbness of the limbs | -120
history of GBS | -6048
clear consciousness | 0
blood pressure 84/58 mmHg | 0
heart rate 115 beats/minute | 0
peripheral oxygen saturation 99% | 0
respiratory rate 22 breaths/minute | 0
body temperature 35.7°C | 0
manual muscle testing strength 3/5 lower extremities | 0
manual muscle testing strength 4/5 upper extremities |. 0
electrocardiogram sinus tachycardia | 0
elevated ST segment V2-6 | 0
cardiothoracic ratio 53% | 0
pulmonary congestion | 0
high troponin I 1.3 ng/mL | 0
high brain natriuretic peptides 896 pg/mL | 0
creatine kinase 235 IU/L | 0
creatine kinase-myocardial band 15.5 IU/L | 0
polymerase chain reaction positive influenza virus A | 0
serology negative Campylobacter | 0
serology negative coxsackievirus | 0
serology negative adenovirus | 0
serology negative cytomegalovirus | 0
serology negative parvovirus B19 | 0
serology negative Epstein-Barr virus | 0
serology negative human herpesvirus 6 | 0
serology negative enterovirus | 0
serology negative hepatitis | 0
serology negative HIV | 0
transthoracic echocardiogram LV end-diastolic diameter 38 mm | 0
ejection fraction 25% | 0
LV wall thickened 14 mm | 0
myocardial edema | 0
cardiac computed tomography no coronary artery stenosis | 0
endomyocardial biopsy lymphocytes present | 0
endomyocardial biopsy eosinophils absent | 0
endomyocardial biopsy giant cells absent | 0
fulminant myocarditis | 0
VA-ECMO support | 0
intra-aortic balloon pumping support | 0
sedation | 0
shock state persisted | 0
large quantities norepinephrine administered | 0
severely reduced LV function | 6
ejection fraction 4% | 6
aortic valve hardly opened | 6
liver enzyme level increased | 72
myocardial injury | 72
shocked liver | 72
bilirubin increased | 72
bilirubin peaked 5.6 mg/dL | 72
aspartate aminotransferase increased 409 IU/dL | 72
alanine aminotransferase increased 120 IU/dL | 72
condition improved | 168
left ventricular ejection fraction 67% | 168
weaned from VA,ECMO | 168
weaned from IABP | 168
ventilator weaned | 264
cessation of sedation | 192
motor disorders in limbs remained | 192
sensory disorders in limbs remained | 192
manual muscle testing strength 0/5 lower extremities | 192
manual muscle testing strength 1/5 upper extremities | 192
absent deep tendon reflexes | 192
sensory disturbance glove-and-stocking type | 192
nerve conduction study decreased amplitude compound muscle action potential median nerve | 192
nerve conduction study decreased amplitude compound muscle action potential ulnar nerve | 192
nerve conduction study amplitude disappeared tibial nerve | 192
acute motor axonal neuropathy | 192
no albuminocytologic dissociation cerebrospinal fluid | 192
axonal GBS | 192
immunoadsorption rounds 5 | 216
motor disorders improved | 216
sensory disorders improved | 216
discharged | 648
no Conflict of Interest | 0
weakness | -48
numbness of the limbs | -48
manual muscle testing strength 4/5 upper extremities | 0
weaned from VA-ECMO | 168
