baby boy | 0
born by emergency cesarean section | 0
severe preeclampsia in the mother | -672
gestational week 25 6/7 | 0
birthweight 665 g | 0
intubated in the delivery room | 0
transferred to the neonatal intensive care unit | 0
mechanical ventilation | 0
total parenteral nutrition (TPN) | 24
minimal enteral nutrition with breast milk | 24
delayed meconium passage | 48
abdominal distension | 48
increased gastric residuals | 48
necrotizing enterocolitis (NEC) | 48
gastric free drainage | 144
broad-spectrum antibiotic therapy | 144
perforated NEC | 144
surgery | 144
short bowel syndrome | 144
stoma formation | 144
thyroid screening tests | 336
low serum levels of fT4 | 336
low TSH | 336
high cortisol | 336
high serum total bilirubin level | 336
high direct reacting bilirubin (DB) | 336
enteral levothyroxine 5 µg/kg/day | 336
no response to treatment | 432
enteral levothyroxine 10 µg/kg/day | 432
poor absorption of the drug | 432
rectal levothyroxine treatment | 504
increased fT4 levels | 576
decreased bilirubin levels | 576
death | 1848
severe bronchopulmonary dysplasia | 1848
surgical NEC | 1848
short bowel syndrome | 1848
sepsis | 1848