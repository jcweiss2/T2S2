83 years old | 0
female | 0
atrial fibrillation | -672
anticoagulation with apixaban | -672
hypertension | -672
hyperlipidemia | -672
type 2 diabetes mellitus | -672
small bowel obstruction | -24
exploratory laparotomy | -24
ventral hernia repair | -24
abdominal wound infections | -24
multiple debridements | -24
fever | -12
chills | -12
purulent drainage from abdominal wounds | -12
septic | -12
7.5 Fr triple lumen right internal jugular vein CVC placement | -12
possible arterial cannulation | -12
contrast computed tomography scan | -6
CVC penetration of right internal jugular vein | -6
CVC penetration of right subclavian artery | -6
CVC termination in aortic arch | -6
right-sided aortic arch anatomical variant | -6
separate origins of RSCA and RCCA | -6
tortuous course of arch vessels | -6
LCCA arising from aorta | -6
RCCA arising from aorta | -6
RSCA arising from aorta | -6
LSCA with Kommerel’s diverticulum | -6
transfer to facility | 0
planned endovascular intervention | 0
central arterial stent graft placement | 0
open brachial access | 0
right brachial artery cutdown | 0
systemic heparinization | 0
intravascular ultrasound | 0
angiography | 0
identification of vertebral artery origin | 0
stent graft deployment | 0
CVC removal | 0
balloon angioplasty | 0
completion angiogram | 0
extubation | 0
observation in surgical intensive care unit | 0
heparin infusion | 0
transition to apixaban | 48
transfer to floor | 24
discharge | 168
arterial duplex | 720
transition to apixaban monotherapy | 720
medication regimen adjustment | 720