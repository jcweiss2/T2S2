70 years old | 0
male | 0
admitted to the hospital | 0
jaundice | -504
vomiting | -504
total serum bilirubin 5.7 mg/dl | -504
direct bilirubin 4.7 mg/dl | -504
INR 1.2 | -504
normal ALT | -504
normal AST | -504
normal serum electrolyte | -504
normal serum creatinine | -504
mild hepatomegaly | -504
dilated intra and extra hepatic biliary channels | -504
no features of cirrhosis of liver | -504
no portal hypertension | -504
hypo-echoic lesion in the head of pancreas | -504
CECT scan | -504
soft tissue mass arising from head of pancreas | -504
gastric wall invasion | -504
decision for surgical intervention | -504
preoperative plan for pancreaticodudenctomy | -504
evaluated by cardiac physician | -504
evaluated by pulmonary physician | -504
evaluated by anesthesia physician | -504
found fit for surgery | -504
intraoperative finding similar to preoperative imaging | 0
common hepatic artery injury | 0
repair with Proline 8/0 | 0
intraoperative Doppler on hepatic artery shows normal flow | 0
RI 0.6 | 0
PSV 100 cm/s pre anastomotic | 0
PSV 125 cm/s post anastomotic | 0
SAT 71 ms | 0
pyloric preserving pancreaticodudenctomy | 0
admitted to Intensive care | 0
stable on POD 1 | 24
Doppler on hepatic artery revealed no detectable flow | 24
liver enzymes highly elevated | 24
ALT 1278 U/L | 24
AST 973 U/L | 24
CECT revealed completely thrombosed common hepatic artery | 24
intrahepatic small accessory left hepatic artery | 24
middle hepatic artery | 24
arised from Left gastric artery | 24
decision to follow the patient | 24
ALT start to decrease | 48
AST start to decrease | 48
bilirubin start to decrease | 48
shifted from ICU to word | 72
Doppler on hepatic artery did not detect any flow | 72
ALT 137 U/L | 240
AST 34 U/L | 240
total bilirubin 1.3 mg/dl | 240
discharged | 240
follow up two weeks later | 336
normal liver function tests | 336
non-detectable hepatic artery flow | 336
follow up six months later | 2160
normal lab parameters | 2160
CECT scan | 2160
completely thrombosed hepatic artery | 2160
small accessory left hepatic artery | 2160
middle hepatic artery | 2160