21 years old | 0
    male | 0
    obese | 0
    cough | -72
    fevers | -72
    shortness of breath | -72
    pleuritic chest pain | -72
    light-headedness | -24
    near syncope | -24
    acutely worsened dyspnoea | -24
    denies contact with sick persons | 0
    denies exertional chest pain | 0
    denies weight loss | 0
    denies night sweats | 0
    denies abdominal pain | 0
    denies changes in bladder or bowel habits | 0
    denies recent travel | 0
    denies surgery | 0
    denies prolonged immobilization | 0
    febrile (38.9°C) | 0
    tachycardic (121 beats per minute) | 0
    normotensive (104/66 mmHg) | 0
    hypoxic saturating 82% on room air | 0
    improved to 100% with non-rebreather mask at 15 L/min | 0
    COVID-19 diagnosed by PCR | 0
    acute sub-massive pulmonary embolism diagnosed by CTPA | 0
    unfractionated heparin (UFH) initiated | 0
    hypotensive | 12
    massive PE diagnosed | 12
    catheter-directed thrombolysis (CDT) of bilateral pulmonary arteries | 12
    patient improved clinically | 72
    plans made for discharge | 72
    acute respiratory failure | 96
    hypotension | 96
    intubated | 96
    cardiac arrest | 96
    return of spontaneous circulation (ROSC) obtained | 96
    vasopressors initiated | 96
    veno0arterial extracorporeal membrane oxygenation (ECMO) initiated | 96
    pulmonary artery angiogram demonstrated interval worsening of bilateral pulmonary emboli | 96
    recurrent massive PE confirmed | 96
    repeat CDT performed | 96
    ventilation parameters improved | 120
    vasopressors discontinued | 120
    weaning of ECMO began | 120
    venous duplex ultrasound demonstrated deep venous thrombus of right femoral vein | 120
    venous duplex ultrasound demonstrated deep venous thrombus of right popliteal vein | 120
    inferior vena cava (IVC) filter placed | 120
    UFH transitioned to low-molecular weight heparin | 120
    repeat pulmonary artery angiogram demonstrated improvement in emboli burden | 240
    successfully weaned from ECMO | 240
    decannulated | 240
    septic shock treated | 264
    development of right thigh haematoma | 960
    compartment syndrome requiring surgical debridement | 960
    transitioned to rivaroxaban | 960
    discharged to acute rehabilitation facility | 1248
    returned home | 1608
    able to perform activities of daily living independently | 1608
    remained anticoagulated on rivaroxaban | 1608
    no major adverse events 4 months following discharge | 1608
    <|eot_id|>
    