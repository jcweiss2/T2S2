77 years old | 0
male | 0
unstable angina | -2880
coronary stent insertion | -2880
Sigmart | -2880
aspirin | -2880
Almarl | -2880
Herben | -2880
admitted to the hospital | 0
TKA | 0
spinal anesthesia | 0
tourniquet application | 0
bupivacaine | 0
dexmedetomidine | 0
crystalloid administration | 0
estimated blood loss | 0
drowsy mental state | 24
severe pain on the right thigh | 24
overnight shivering | 24
Tridol Injection | 24
Glasgow coma scale score of 8/15 | 24
vital signs | 24
electrocardiogram | 24
stiff and dark brown right thigh | 24
oliguria | 24
dark colored urine | 24
elevated CK | 19
elevated CK-MB | 19
elevated AST | 19
elevated BUN/Cr | 19
normal troponin-I | 19
coagulation panel | 19
thrombocytopenia | 19
high levels of fibrinogen degradation product and D-dimer | 19
progressive deterioration of DIC | 19
elevated serum myoglobin | 25
myoglobinuria | 25
red blood cell count | 25
rhabdomyolysis diagnosis | 25
AKI diagnosis | 25
DIC diagnosis | 25
norepinephrine infusion | 25
arterial line placement | 25
central line placement | 25
fluid treatment | 25
dialysis | 25
Lasix administration | 25
sodium bicarbonate administration | 25
Denogan administration | 25
restored mental status | 27
elevated body temperature | 29
cardiac arrest | 32
CPR | 32
death | 33
discharge | -1