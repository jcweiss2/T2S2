25 years old | 0
male | 0
asymptomatic COVID-19 infection | -672
fever | -96
abdominal pain | -96
vomiting | -96
diarrhea | -96
elevated Erythrocyte Sedimentation Rate | -96
elevated C-Reactive Protein | -96
normal white blood cell count | -96
amoxicillin/clavulanic acid | -96
cefuroxime | -48
diffuse erythematous and maculopapular rash | -48
admitted to the hospital | 0
dyspnoea | 0
diffuse abdominal pain | 0
rash | 0
bilateral conjunctivitis | 0
neutrophilia | 0
thrombocytopenia | 0
lymphopenia | 0
high ferritin | 0
high D-dimer | 0
increased serum creatinine | 0
increased gamma-glutamyl transferase | 0
increased alkaline phosphatase | 0
increased total bilirubin | 0
thoraco-abdominal Computed Tomography | 0
uncomplicated ileocaecal inflammation | 0
mesenteric lymphadenopathy | 0
splenomegaly | 0
normal lung parenchyma | 0
discrete pericardial effusion | 0
transthoracic echocardiography | 0
normal cardiac morphology | 0
normal cardiac function | 0
intravenous ciprofloxacin | 0
metronidazole | 0
hypotension | 24
high anion gap metabolic acidosis | 24
lactic acid accumulation | 24
fluid resuscitation | 24
norepinephrine | 24
type 1 respiratory insufficiency | 24
High Flow Nasal Oxygen | 24
sedation | 24
intubation | 24
mechanical ventilation | 24
thoraco-abdominal CT | 48
terminal ileitis | 48
diffuse colitis | 48
increased lymphadenopathy | 48
hepatosplenomegaly | 48
new ascites | 48
bilateral pleural effusions | 48
meropenem | 48
vancomycin | 48
exploratory laparoscopy | 48
moderate clear ascites | 48
mildly dilated left ventricle | 72
moderately decreased ejection fraction | 72
anteroseptal akinesia | 72
hypokinesia | 72
circumferential pericardial effusion | 72
cardiomegaly | 72
pulmonary edema | 72
elevated high sensitive troponin T | 72
elevated NT-pro-BNP | 72
dobutamine | 72
levosimendan | 72
Cardiac MRI | 96
moderately dilated left ventricle | 96
moderately reduced systolic function | 96
non-ischemic myocardial injury | 96
focal myocardial edema | 96
pericardial inflammation | 96
MIS-A diagnosis | 96
intravenous immunoglobulins | 96
pulse corticosteroids | 96
improvement | 120
weaned off ventilatory support | 120
weaned off inotropic support | 120
weaned off vasopressor support | 120
antibiotics discontinued | 144
ECG showed regression of PR depression | 144
TTE showed improved anteroseptal contractility | 144
TTE showed increased LVEF | 144
TTE showed regressed pericardial effusion | 144
corticosteroids continued orally | 144
proton pump inhibitor | 144
calcium/vitamin D supplements | 144
heart failure therapy | 144
low-dose aspirin | 144
asymptomatic | 240
without inflammation | 240
resting ECG normal | 240
TTE showed normalisation of left ventricular diameters | 240
TTE showed normalisation of systolic function | 240
heart failure therapy discontinued | 240
low-dose aspirin discontinued | 240