64 years old | 0 | 0 
female | 0 | 0 
admitted to the hospital | 0 | 0 
severe headache | -24 | 0 
right periorbital and mid-facial swelling | -24 | 0 
fever | -336 | -168 
headache | -336 | -168 
light pain in the right ear | -336 | -168 
purulent secretion from the ear | -336 | -168 
swelling and redness of the skin behind the right ear | -336 | -168 
tinnitus | -336 | -168 
hearing disorder | -336 | -168 
Amoxicillin | -336 | -168 
painkillers | -336 | -168 
anti-inflammatory drugs | -336 | -168 
arterial hypertension | 0 | 0 
angiotensin-converting enzyme inhibitors | 0 | 0 
right facial and periorbital swelling | 0 | 0 
right blepharoptosis | 0 | 0 
chemosis | 0 | 0 
proptosis | 0 | 0 
visual acuity of 7/12 on her right eye | 0 | 0 
no visual fields abnormalities | 0 | 0 
normal intraocular pressures | 0 | 0 
no relative afferent pupillary defect | 0 | 0 
normal color vision | 0 | 0 
no signs of optic disc swelling | 0 | 0 
febrile | 0 | 0 
conscious | 0 | 0 
somnolent | 0 | 0 
no neurological deficits | 0 | 0 
normal cardiovascular examination | 0 | 0 
normal respiratory examination | 0 | 0 
elevated white blood cells count | 0 | 0 
elevated erythrocyte sedimentation rate | 0 | 0 
elevated C-reactive protein | 0 | 0 
normal renal function | 0 | 0 
normal liver function | 0 | 0 
prothrombin G20210A mutation | 0 | 0 
normal coagulation profile | 0 | 0 
normal urinalysis | 0 | 0 
non-opacification of the right cavernous sinus | 0 | 0 
Ceftriaxone | 0 | 48 
Enoxaparin | 0 | 48 
shortness of breath | 96 | 96 
reduced oxygen saturation | 96 | 96 
unilateral homogeneous opacification on right lobar lung | 96 | 96 
air bronchograms | 96 | 96 
non-invasive mechanical ventilation | 96 | 168 
Amikacin | 96 | 168 
Piperacillin–Tazobactam | 96 | 168 
improvement of symptoms | 168 | 168 
transfer back to the Service | 168 | 168 
control contrast-enhanced magnetic resonance angiography | 168 | 168 
persistence of the lacunar image in the right cavernous sinus | 168 | 168 
diminished periorbital swelling | 168 | 168 
discharged | 336 | 336 
oral anticoagulant – Acenocoumarol | 336 | 0 
follow-up CT venogram | 720 | 720 
full recovery | 720 | 720