67 years old | 0
    male | 0
    small cell lung cancer | 0
    coronary artery disease | 0
    chronic obstructive pulmonary disease | 0
    type 2 diabetes | 0
    admitted to the intensive care unit | 0
    weakness | 0
    pancytopenia | 0
    sepsis | 0
    urinary tract infection | 0
    bed-bound | -72
    chemotherapy with etoposide | -4320
    chemotherapy with carboplatin | -4320
    radiation therapy | -4320
    one dose of atezolizumab | -4320
    broad-spectrum antibiotics | 0
    neuopogen | 0
    supportive therapy | 0
    hematemesis | 24
    blood-loss anemia | 24
    blood counts stabilized posttransfusion | 24
    peripheral smear | 24
    no schistocytes | 24
    no abnormal platelet morphology | 24
    pancytopenia confirmed | 24
    spherocytes confirmed | 24
    computed tomography of abdomen/pelvis | 24
    computed tomography angiography of abdomen/pelvis | 24
    no splenomegaly | 24
    hypertriglyceridemia (385) | 24
    elevated ferritin (32100) | 24
    MRSA bacteremia | 24
    suspicion for endocarditis | 24
    transthoracic echocardiogram | 24
    no vegetation | 24
    HLH diagnosis | 24
    fever | 24
    hyperferritinemia | 24
    hypertriglyceridemia | 24
    high-dose steroids | 24
    etoposide discussed | 24
    etoposide withheld | 24
    worsening sepsis | 24
    exacerbating immunosuppression | 24
    decline | 24
    resuscitation | 48
    intubation | 48
    pressors | 48
    no improvement | 48
    comfort care only | 48
    expired | 48
    elevated soluble IL2 receptor (22268 U/mL) | 48
    MRSA-related infective endocarditis | 48
    secondary HLH | 48
    chemotherapy treatment | -2880
    radiation therapy treatment | -2880
    no recurrence of disease | -672
    HLH triggered by MRSA-septicemia | 48
    MAHS excluded | 48
    elevated ferritin >500 | 24
    elevated soluble CD25 | 24
    no splenomegaly | 24
    persistent fever | 24
    pancytopenia | 24
    hypertriglyceridemia | 24
    hyperferritinemia | 24
    blood cultures positive for MRSA | 24
    no vegetation on echocardiogram | 24
    HLH criteria met | 24
    low or absent NK cell activity | 24
    hemophagocytosis in bone marrow | 24
    hemophagocytosis in spleen | 24
    hemophagocytosis in lymph node | 24
    hemophagocytosis in cerebrospinal fluid | 24
    hypofibrinogenemia | 24
    HLH diagnosis confirmed | 48
    HLH treatment initiated | 24
    HLH prognosis | 48
    patient death | 48
    postmortem findings | 48
    Southern Regional Meeting presentation | 0
    written informed consent | 0
    ethical approval not required | 0
    no conflicts of interest | 0
    no financial support | 0
    
