14 years old | 0  
    female | 0  
    nausea | -72  
    vomiting | -72  
    abdominal pain | -72  
    admitted to the local clinic | 0  
    acute viral gastroenteritis | 0  
    hyperglycemia (glucose, 500 mg/dL) | 0  
    ketonuria | 0  
    transferred to emergency unit | 0  
    worsening mental status | 0  
    intravenous fluid | 0  
    short-acting insulin | 0  
    mother has type 2 diabetes mellitus | 0  
    lethargic | 0  
    severely dehydrated | 0  
    drowsy (GCS=14) | 0  
    tachycardia (124 beats/min) | 0  
    tachypnea (40 breaths/min) | 0  
    hypothermia (35℃) | 0  
    blood pressure 106/56 mmHg | 0  
    weight decreased by 1.7 kg in previous month | -720  
    weight 48 kg | 0  
    body mass index 20 kg/m² | 0  
    chest x-ray no abnormalities | 0  
    abdominal x-ray no abnormalities | 0  
    metabolic acidosis (pH 6.92) | 0  
    glucose 569 mg/dL | 0  
    corrected sodium 133 mmol/L | 0  
    potassium 3.2 mmol/L | 0  
    corrected calcium 8.5 mg/dL | 0  
    phosphate 2.1 mg/dL | 0  
    blood urea nitrogen 25.9 mg/dL | 0  
    creatinine 0.57 mg/dL | 0  
    lactate 0.6 mmol/L | 0  
    urinalysis ketones present | 0  
    urinalysis glucose present | 0  
    C-peptide 0.26 ng/mL | 0  
    glycosylated hemoglobin 15.7% | 0  
    antiglutamic acid decarboxylase positive (1.72 U/mL) | 0  
    anti-islet cell antibody negative | 0  
    anti-insulin antibody negative | 0  
    type 1 diabetes | 0  
    severe DKA | 0  
    fluid therapy (0.45% saline) | 0  
    continuous intravenous insulin infusion | 0  
    hourly neurological evaluations | 0  
    remained drowsy | 0  
    no signs of cerebral edema | 0  
    generalized tonic seizure | 4  
    bradycardia | 4  
    cardiopulmonary arrest | 4  
    external cardiac massage | 4  
    epinephrine injection | 4  
    spontaneous circulation resumed | 4  
    metabolic acidosis after resuscitation (pH 7.05) | 4  
    hypophosphatemia (1.2 mg/dL) | 4  
    K2HPO4 administered | 4  
    KCl administered | 4  
    phosphorus replacement 1.9 mEq/kg/day | 4  
    brain CT scan no brain edema | 4  
    dexamethasone prescribed | 4  
    mannitol prescribed | 4  
    admitted to ICU | 4  
    remained drowsy (GCS=14) | 4  
    vital signs stable | 4  
    stuporous (GCS=9) | 16  
    shallow respiration | 16  
    weak respiration | 16  
    slow respiration | 16  
    endotracheal intubation | 16  
    respiratory acidosis (pH 6.80) | 16  
    severe hypophosphatemia (0.4 mg/dL) | 16  
    phosphate replacement increased to 3.8 mEq/kg/day | 16  
    repeat brain CT no abnormalities | 16  
    electrolyte normalization started | 48  
    pH normalization started | 48  
    mechanical ventilation required | 48  
    phosphate 1.4 mg/dL | 48  
    phosphate replacement increased to 5.7 mEq/kg/day | 48  
    fluid replacement continued | 48  
    potassium replacement continued | 48  
    insulin administration continued | 48  
    vital signs stable on day 3 | 72  
    self-respiration recovered | 72  
    arterial blood gas normal (pH 7.39) | 72  
    phosphate 3.5 mg/dL | 72  
    weaning from inotropic support | 72  
    weaning from ventilator support | 72  
    transferred to general ward | 96  
    oral feeding started | 96  
    multiple subcutaneous insulin injections started | 96  
    phosphate supplementation stopped | 96  
    electroencephalogram no epileptiform discharges | 96  
    electroencephalogram no slow waves | 96  
    discharged on day 10 | 240  
    no neurologic complications | 240  
    follow-up no neurologic complications | 240  
    follow-up no respiratory problems | 240  
    no further phosphate supplementation required | 240  

