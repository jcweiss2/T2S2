2 years old | 0
male | 0
Caucasian | 0
admitted to the Emergency Room | 0
high fever | 0
not relieved by antipyretic treatment | 0
febrile | 0
body temperature 39.2°C | 0
severely ill | 0
extremely irritable | 0
heart rate 170/min | 0
blood pressure 98/51 mmHg | 0
petechial lesions | 0
disseminated on the torso and limbs | 0
suspecting meningococcemia | 0
intravenous fluids | 0
ceftriaxone | 0
hypotension | 0
inotropic support | 0
intubation | 0
mechanical ventilation | 0
transferred to the pediatric Intensive Care Unit | 0
Neisseria meningitidis serogroup B isolated | 0
cerebrospinal fluid sample normal | 0
antibiotic therapy continued | 0
inflammatory markers levels decreased | 48
C-reactive protein decreased | 48
inotropic agents stopped | 120
extubated | 168
general improvement | 168
spikes of fever | 168
broader antibiotic therapy | 168
ceftriaxone | 168
gentamicin | 168
teicoplanin | 168
blood and urine cultures negative | 168
lumbar puncture negative | 168
chest X-ray normal | 168
brain magnetic resonance imaging normal | 168
transferred to the General Pediatrics Unit | 312
stable but still febrile | 312
physical examination unremarkable | 312
cutaneous ulcers | 312
hemoglobin 8.1 g/L | 312
red blood cells 3,050,000/mm3 | 312
mean corpuscular volume 80.6 fl | 312
white blood cell count 25,830/mm3 | 312
polymorphonuclear leucocytes 16,140/mm3 | 312
Platelets count 1,090,000/mm3 | 312
C-reactive protein 44.80 mg/L | 312
febrile | 312
fever spikes | 312
broad-spectrum antibiotic treatment | 312
conditions worsened | 504
extremely irritable | 504
more frequent fever spikes | 504
higher temperatures | 504
C-reactive protein 89.70 mg/L | 504
erythrocyte sedimentation rate 36 mm/h | 504
Ferritin 173 ug/L | 504
neopterine 31.0 nmol/L | 504
TNF 29.8 ng/L | 504
antibiotic therapy broadened | 504
meropenem | 504
teicoplanin | 504
cultures collected negative | 504
erythematous-papular rash | 528
hepatomegaly | 528
bilateral cervical lymphadenopathy | 528
suspecting viral infection | 528
serological tests | 528
Adenovirus | 528
EBV | 528
CMV | 528
Parvovirus B19 | 528
negative results | 600
neck ultrasound | 600
reactive lymph nodes | 600
suspecting vasculitis | 600
atypical Kawasaki | 600
electrocardiogram | 600
echocardiography | 600
no atrial shunt | 600
no mitral or tricuspid regurgitation | 600
good biventricular contractility | 600
hyper echogenicity of mitral papillary muscles | 600
outflows free | 600
normal coronaries | 600
IVIG administered | 624
no effect on fever spikes | 624
IVIG administration repeated | 672
poor clinical improvement | 672
hemoglobin 7.4 g/dL | 696
red blood cells 3,050,000/mm3 | 696
mean corpuscular volume 76.4 fl | 696
white blood cell count 23,470/mm3 | 696
polymorphonuclear leucocytes 11,050/mm3 | 696
Platelets count 98,000/mm3 | 696
LDH 1091 U/L | 696
normal renal function | 696
albumin 31 g/L | 696
AST 86 IU/L | 696
ALT 117 IU/L | 696
GGT 300 U/L | 696
sodium 135 mmol/L | 696
triglycerides 361 mg/dL | 696
coagulation pattern compatible with severe discoagulopathy | 696
prothrombin 15% | 696
activated partial thromboplastin time 45 sec | 696
fibrinogen 1 g/L | 696
Vitamin K administered | 696
fresh frozen plasma administered | 696
coagulation pattern normalized | 696
bone marrow aspirate | 696
no signs of hemophagocytic lymphohistiocytosis | 696
conjunctival injection | 720
fissured dry lips | 720
facial and feet edema | 720
KD diagnosis | 720
MAS suspected | 720
IVMP administered | 768
inflammatory markers decreased | 840
fever spikes reduced | 840
afebrile | 888
follow-up echocardiogram | 888
no cardiac worsening | 888
follow-up at 3 months | 2160
healthy child | 2160
normal physical examination | 2160
normal laboratory tests | 2160
normal inflammatory markers | 2160
normal ECG | 2160
follow-up echocardiogram confirmed no cardiac worsening | 2160