41 years old | 0
premenopausal woman | 0
admitted to the hospital | 0
worsening abdominal pain | 0
vomiting | 0
non-bloody diarrhoea | 0
fever | 0
intermittent abdominal pain | -504
returned from overseas travel to Indonesia | -504
Stage 4 endometriosis | -0
bilateral endometriomas | -0
rectal nodule | -0
obliterated pouch of Douglas | -0
fixed anterior uterus | -0
previous caesarean section | -0
well controlled asthma | -0
no recent sexual intercourse | 0
no uterine instrumentation | 0
no history of PID | 0
no history of sexually transmitted infections | 0
not taking any regular medication | 0
not on any contraceptives | 0
regular menstrual cycles | 0
tachycardic | 0
hypotensive | 0
febrile | 0
right renal angle tenderness | 0
generalised lower abdominal tenderness | 0
rebound | 0
guarding | 0
right adnexal tenderness | 0
no palpable masses | 0
no cervical motion tenderness | 0
normal cervix | 0
no abnormal vaginal discharge | 0
elevated lactate | 0
leucocytosis | 0
neutrophilia | 0
elevated C-reactive protein | 0
acute kidney injury | 0
elevated creatinine | 0
reduced estimated glomerular filtration rate | 0
negative quantitative beta hCG | 0
negative urinalysis | 0
negative microscopy | 0
negative culture | 0
negative endocervical swabs | 0
negative blood cultures | 0
positive stool culture | 0
Campylobacter jejuni | 0
bilateral enlarged ovaries | 0
septated cysts | 0
low-density mass | 0
fat stranding | 0
multiple endometriomas | 0
right ovarian cyst | 0
left ovarian cysts | 0
fixed ovaries | 0
kissing ovaries sign | 0
negative sliding sign | 0
bowel adherent to posterior wall of uterus | 0
bowel nodules | 0
colitis | 0
urosepsis | 0
appendicitis | 0
tubo-ovarian abscesses | 0
empirically managed for sepsis | 0
fluid resuscitation | 0
broad-spectrum intravenous antibiotics | 0
ceftriaxone | 0
metronidazole | 0
condition deteriorated | 24
ongoing fever | 24
tachycardia | 24
hypotension | 24
inotropic support | 24
intravenous amoxicillin | 24
clavulanic acid | 24
azithromycin | 24
Campylobacteriosis | 24
repeat CT abdomen pelvis | 120
interval increase in left multiloculated adnexal mass | 120
increased surrounding fat stranding | 120
free fluid in pelvis | 120
bowel wall thickening | 120
exploratory laparoscopy | 120
urgent laparoscopic washout | 120
drainage of tubo-ovarian abscesses | 120
sterile abscess culture fluid | 120
Escherichia coli | 120
right adnexal tissue histopathology | 120
abscess formation | 120
no evidence of endometriosis | 120
intravenous antibiotics | 120
intravenous fluids | 120
condition improved | 120
discharged from hospital | 168
outpatient follow-up | 168
repeat pelvic scan | 168