43 years old | 0
male | 0
admitted to the hospital | 0
jaundice | -168
nausea | -168
vomiting | -168
abdominal pain | -168
flu-like syndrome | -168
fever | -168
chills | -168
headache | -168
myalgia | -168
arthralgia | -168
tea-colored urine | -96
decreased urine output | -96
asymptomatic chronic HBV infection | -7920
asymptomatic chronic HBV infection diagnosis | -7920
abdominal upper quadrant tenderness | 0
profound jaundice | 0
no hepatosplenomegaly | 0
no ascites | 0
normal neurological examination | 0
acute kidney injury | 0
elevated total bilirubin | 0
elevated indirect bilirubin | 0
elevated liver transaminases | 0
anemia | 0
thrombocytopenia | 0
hypoalbuminemia | 0
positive bilirubin in urine | 0
positive urobilinogen in urine | 0
no hemoglobin in urine | 0
negative Covid-19 PCR | 0
positive HBsAg | 0
positive IgM anti-HBc | 0
positive anti-HBe | 0
negative HBeAg | 0
negative hepatitis C | 0
negative hepatitis D | 0
negative HIV | 0
normal liver size and parenchyma on ultrasound | 0
severe liver fibrosis on hepatic elastography | 0
altered consciousness | 48
metabolic acidosis | 48
oliguria | 48
severe malaria diagnosis | 48
intravenous artesunate treatment | 48
oral primaquine treatment | 48
continuous renal replacement therapy | 48
intubation | 48
transferred to intensive care unit | 48
pulmonary edema | 120
septic shock | 120
multiorgan dysfunction | 120
death | 168
cardiopulmonary resuscitation | 168