74 years old | 0
male | 0
hypertension | 0
insulin-dependent diabetes mellitus type 2 | 0
diabetic retinopathy | 0
weight loss | -672
iron deficiency anemia | -672
tumor in the colon ascendens | -672
liver metastases | -672
right hemicolectomy | -672
low-grade pT3cN0 adenocarcinoma | -672
absence of metastases in 24 excised lymph nodes | -672
lymphovascular growth | -672
no vascular or perineural growth | -672
activated BRAF mutation | -672
loss of expression of MLH1 and PMS2 | -672
mismatch repair-deficient (MMR-D)/microsatellite-instable (MSI) tumor | -672
initiated therapy with pembrolizumab | 0
symptoms of a cold | -168
leukocytosis | -168
increase in C-reactive protein | -168
dry coughing | -504
no fever | -504
increase in AST and ALT | -504
ICI-induced hepatitis grade 2 | -504
initiated prednisolone therapy | -504
decrease in C-reactive protein and AST | -504
increase in white blood cells and neutrophils | -504
dyspnea | -408
myocardial infarction suspected | -408
elevation of troponin T | -408
septal hypokinesia | -408
no dynamic change in troponin T | -408
somnolence | -408
difficulty walking | -408
dysarthria | -384
hoarseness | -384
pain in neck and right leg | -384
difficulty raising right leg | -384
increased dose of prednisolone | -384
no signs of stroke | -384
increased creatine kinase and myoglobin levels | -384
ICI-induced myositis suspected | -384
gradual decrease in creatinine levels | -384
antibodies against acetylcholine receptor and titin present | -384
albumin present in cerebrospinal fluid | -384
unable to sit up | -336
severe dysarthria and dysphagia | -336
absent reflexes | -336
intubated | -336
given methylprednisolone | -336
given intravenous immunoglobulins | -336
given infliximab | -312
felt better | -312
better muscle strength in hands | -312
carbon dioxide retention | -288
noninvasive ventilation | -288
sinus bradycardia | -288
died | -288
autopsy showed significant stenosis of right coronary artery | -288
no fibrosis or signs of recent myocardial infarction | -288
tongue softened | -288
no surgical complication after hemicolectomy | -288
metastasis in right liver lobe | -288
inflammatory infiltration of lymphocytes in intercostal musculature, diaphragm, cervical musculature, and tongue | -288
fibrosis in one area of heart | -288
inflammatory infiltrate in small area of heart | -288
hepatocellular cancer (HCC) in liver | -288
HCC positive for hepatocytes and negative for glypican, CDX2, CK20, and CK7 | -288
fibrosis stage 2-3 in porta field | -288
cause of death determined as respiratory insufficiency due to polymyositis | -288