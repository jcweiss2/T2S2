61 years old | 0
male | 0
admitted to the hospital | 0
diarrhea | -24
nausea | -24
foul-smelling belching | -24
vomiting | -24
stabbing epigastric pain | -24
intermittent chills | -24
dizziness | -24
denied fever | -24
denied headache | -24
no recent travel | -24
no sick contacts | -24
no unusual food intake | -24
20-year history of ulcerative colitis | -6720
total procto-colectomy with ileal–anal anastomosis | -5040
ulcerative colitis in remission | -5040
diabetes mellitus | 0
hypercholesterolemia | 0
hypertension | 0
sitagliptin–metformin | 0
atorvastatin | 0
enalapril | 0
metoprolol tartrate | 0
no excessive consumption of NSAIDs | 0
no smoking | 0
no alcohol abuse | 0
hypotensive | 0
blood pressure 80/56 mmHg | 0
pulse 60 | 0
respiratory rate 16 | 0
temperature 36°C | 0
abdomen soft | 0
abdomen non-distended | 0
abdomen mildly tender | 0
leukocytosis | 0
elevated lactate | 0
anion gap metabolic acidosis | 0
acute kidney injury | 0
creatinine 299 µmol/L | 0
non-contrast CT of the chest, abdomen, and pelvis | 0
emphysema in the wall of the stomach | 0
air in peri-gastric veins | 0
portal venous gas | 0
left adrenal nodule | 0
intravenous fluids | 0
piperacillin/tazobactam | 0
pantoprazole | 0
admitted to the intensive care unit | 0
rapid resolution of symptoms | 24
admission stool studies negative | 24
diet advanced gradually | 24
renal function improved | 24
follow-up CT of the abdomen and pelvis | 72
resolution of the EG | 72
discharged home | 72
oral pantoprazole | 72
ciprofloxacin | 72
metronidazole | 72
follow-up with gastroenterology | 168
follow-up CT abdomen | 432
gastric intramural air | 0
pneumatosis intestinalis | 0
gastric emphysema | 0
Enterobacter spp. | 0
Staphylococcus aureus | 0
Pseudomonas aeruginosa | 0
Candida albicans | 0
alcohol abuse | 0
gastric surgery | 0
recent gastroenteritis | 0
corrosive ingestion | 0
chronic consumption of NSAIDs/steroids | 0
COPD | 0
immunosuppression | 0
raised intra-gastric pressures | 0
dissection of air from the mediastinum | 0
trauma | 0
malignancy | 0
inflammation | 0
ischemia | 0
low-grade fever | 0
chills | 0
mild-to-severe abdominal pain | 0
diarrhea | 0
hematochezia | 0
shock | 0
abdominal distension | 0
epigastric tenderness | 0
decreased bowel sounds | 0
metabolic acidosis | 0
sepsis | 0
plain radiography | 0
CT | 0
irregular, mottled appearance of the air | 0
thickened gastric wall | 0
portal vein | 0
gastric ischemia | 0
acute abdomen | 0
perforation | 0
necrosis | 0
IV fluids | 0
nasogastric tube placement | 0
nutritional support | 0
broad-spectrum antibiotics | 0
anti-fungal medications | 0
esophagogastroduodenoscopy | 0
gastric strictures | 0
gastric contractures | 0