37 years old | 0
male | 0
admitted to the hospital | 0
fever | -96
headache | -96
myalgia | -96
epigastralgia | -96
nausea | -96
diarrhoea | -96
active smoking | 0
no splenic disorders | 0
no alcohol excess | 0
not immunocompromised | 0
no cardiac symptoms | 0
dog bite | -72
temperature 38.2°C | 0
heart rate 130 b.p.m. | 0
blood pressure 118/72 mmHg | 0
pulse oxygen saturation 100% | 0
bite wound on right hand | 0
no rash | 0
no sign of cellulitis | 0
no soft tissue necrosis | 0
C-reactive protein 417 mg/L | 0
white blood cell count 9.45 G/L | 0
procalcitonin 8.42 μg/L | 0
thrombocytopaenia | 0
acute kidney injury | 0
abnormal liver enzymes | 0
high sensitivity-troponin T elevated | 0
N-terminal brain natriuretic peptide elevated | 0
mild diffuse ST-segment elevation | 0
micro-Q waves in inferior and lateral leads | 0
mild global left ventricular hypokinesia | 0
decrease in LV ejection fraction | 0
preserved right ventricular function | 0
no pericardial effusion | 0
blood cultures drawn | 0
parenteral cefotaxime | 0
Capnocytophaga canimorsus identified | 45
cefotaxime changed to amoxicillin | 47
favourable clinical course | 47
recovery of biological markers | 47
coronary computed tomography angiography | 48
normal coronary arteries | 48
cardiovascular magnetic resonance | 120
non-dilated LV | 120
normal global systolic function | 120
focal areas of subepicardial oedema | 120
early hyper-enhancement in LV inferolateral wall | 120
late gadolinium-enhancement imaging | 120
diagnosis of acute myocarditis | 120
increased T2 time | 120
increased extracellular volume | 120
discharged | 168
no further symptoms at 1 year | 8760