8 years old | 0
male | 0
admitted to the hospital | 0
high fever | -168
constitutional symptoms: malaise | -168
constitutional symptoms: fatigue | -168
constitutional symptoms: anorexia | -168
constitutional symptoms: myalgias | -168
reddish maculopapular skin rashes forearms | -168
reddish maculopapular skin rashes ankles | -168
grotesque pitting edema (anasarca) involving the face | -168
grotesque pitting edema (anasarca) involving the trunk | -168
grotesque pitting edema (anasarca) involving the extremities | -168
pure motor symmetrical progressive weakness, pelvifemoral region | -168
muscles excruciatingly painful | -168
flaccid weakness | -168
bedbound | -168
generalized pitting anasarca | 0
no family history of relevant autoimmune disorders | 0
negative history of Raynaud's phenomenon | 0
negative history of polyarthralgias | 0
negative history of polyarthritis | 0
negative history of bulbar symptomatology: dysphonia | 0
negative history of bulbar symptomatology: pharyngeal dysphagia | 0
negative history of bulbar symptomatology: respiratory muscle weakness | 0
negative history of soft-tissue calcifications | 0
negative history of oral ulceration | 0
no positive history of preceding vaccination | 0
no endocrine disorders | 0
no nutritional disorders | 0
no metabolic disorders | 0
no exposure to drugs | 0
no exposure to toxic substances | 0
conscious | 0
oriented | 0
sick looking | 0
distraught | 0
flaccid quadriparesis | 0
Grade 1 deep tendon reflexes | 0
diffuse Grade 1/5 Medical Research Council muscular weakness | 0
exquisite pain | 0
muscles diffusely tender to palpation | 0
symmetric proximal and axial weakness | 0
grotesque pitting swelling of the face | 0
grotesque pitting swelling of the neck | 0
grotesque pitting swelling of the abdomen | 0
grotesque pitting swelling of the extremities | 0
grotesque pitting swelling of the scrotum | 0
multiple erythematous maculopapular rashes extensor surfaces of the elbows | 0
multiple erythematous maculopapular rashes medial malleoli of the ankles | 0
no evidence of calcinosis | 0
no focal neurological signs | 0
hypoalbuminemia (1.8 mg/dl) | 0
hypotension (90/60 mmHg) | 0
tachycardia (140/min) | 0
normal echocardiogram | 0
normal renal functions | 0
no albuminuria | 0
serum procalcitonin negative | 0
sepsis work up negative | 0
viral serologies negative | 0
complete blood counts normal | 0
serologic tests for antinuclear antibodies (ANA) normal | 0
rheumatoid factor normal | 0
ANA profile normal | 0
perinuclear ANCA normal | 0
cytoplasmic-ANCA normal | 0
antistreptolysin-O titers normal | 0
thyroid functions normal | 0
hepatitis serologies normal | 0
electrocardiography normal | 0
cardiac injury enzymes normal | 0
chest radiography unremarkable | 0
abdominal ultrasonography unremarkable | 0
creatine phosphokinase elevated (12000U/L) | 0
lactate dehydrogenase elevated (6980U/L) | 0
nerve conduction studies normal | 0
electromyography (EMG): increased muscle membrane irritability | 0
EMG: increased insertional activity | 0
EMG: spontaneous fibrillations | 0
EMG: low amplitude short duration polyphasic myopathic MUPs | 0
left vastus lateralis muscle biopsy | 0
diagnosis of JDM | 0
Jo-1 IgG antibody positive | 0
anti-Mi2 antibody positive | 0
reduced C3 complement levels | 0
reduced C4 complement levels | 0
diagnosis of acute JDM | 0
baffling clinical syndromic constellation: hypotension | 0
baffling clinical syndromic constellation: hemoconcentration (high hematocrit of 56%) | 0
baffling clinical syndromic constellation: “shock”-like syndrome | 0
baffling clinical syndromic constellation: hypoalbuminemia | 0
baffling clinical syndromic constellation: massive generalized pitting edema | 0
fulminant SCLS | 0
intense pain | 0
myalgias | 0
incessant crying | 0
parenteral Tramadol (50 mg IV Q8H) | 0
paracetamol around the clock | 0
hemodynamic instability | 0
cardiovascular monitoring | 0
central venous pressure monitoring | 0
aggressive fluid resuscitation | 0
high-dose catecholamine therapy | 0
blood pressure below systolic BP (SBP) of 90 mmHg | 0
volume infusion | 0
moderate dose dopamine | 0
norepinephrine infusion | 0
SBP supported at 90 mm Hg | 0
pulse methylprednisolone (30 mg/kg/day) | 0
high-dose IVIg (2 g/kg/day) | 0
theophylline 200 mg BD | 0
salbutamol 2 mg BD | 0
leukotriene inhibitors (montelukast) | 0
fresh frozen plasma | 0
20% albumin | 0
hemodynamic indices improvement | 72
immunomodulatory therapy: Prednisolone 1.5 mg/kg | 72
immunomodulatory therapy: Azathioprine 2.5 mg/kg/day | 72
motoric recovery | 336
amelioration of edema (50% from baseline) | 336
ambulating | 336
discharged | 672
normal motoric power | 2016
switched to alternate-day glucocorticoid schedule | 2016
cautious reduction of maintenance dose | 2016
gradual taper of prednisolone | 2016
gradual taper of azathioprine | 2016
clinical remission | 17520
immunomodulatory therapy tapered off | 8760
