49 years old | 0
    male | 0
    hospitalized | 0
    fever | -96
    pyrexia | -96
    cough | -96
    shortness of breath | -96
    diabetes | 0
    sliding-scale insulin | 0
    HbA1c 12.3% | 0
    fasting blood sugar 250 mg/dL | 0
    post prandial blood sugar 350 mg/dL | 0
    interleukin 637.93 pg/mL | 0
    C-reactive protein 17.84 mg/L | 0
    D-Dimer 460 ng/mL | 0
    creatinine 0.8 mg/dl |;0
    lymphocyte 9.5% | 0
    neutrophil 84% | 0
    intensive care unit admission | 0
    Remdesivir IV | 0
    methylprednisolone IV | 0
    bilateral pneumonia | 0
    swelling | 0
    discomfort in left eye | 0
    malaise | 0
    proptosis | 0
    chemosis | 0
    periorbital cellulitis | 0
    partial ophthalmoplegia | 0
    visual acuity 6/6 | 0
    MRI findings | 0
    mucormycosis | 0
    rhino-orbital-cerebral extension | 0
    bone erosion | 0
    FESS | 0
    debridement of necrotic tissue | 0
    post-Covid pneumonia | 0
    sepsis | 0
    difficult airway | 0
    restricted mouth opening | 0
    facial nerve palsy | 0
    general anesthesia | 0
    ASA III | 0
    glycopyrrolate 0.2 mg | 0
    fentanyl 150 mg | 0
    propofol 100 mg | 0
    rapid sequence induction | 0
    scoline 2 mg/kg | 0
    endotracheal tube placement | 0
    xylocard 1.5 mg/kg | 0
    vecuronium 0.1 mg/kg | 0
    oxygen | 0
    nitrous | 0
    sevoflurane 1% | 0
    elective ventilation | 0
    uncontrolled diabetes | 0
    active mucormycosis | 0
    surgery executed | 0
    complications managed | 0
    discharged | 0