32 years old | 0
female | 0
referred because of pain localized in the mid-dorsal region | -8760
pain onset several months earlier | -8760
progressive worsening of pain | -8760
pain aggravated with local palpation | -8760
pain aggravated with trunk movement | -8760
weakness in the lower limbs | -8760
radiographic study identified expansive lesion in T8 | -8760
local kyphosis | -8760
imminent instability | -8760
CT scan performed | -8760
MRI performed | -8760
bone involvement | -8760
invasion of the medullary canal | -8760
percutaneous CT-guided core-needle biopsy | -8760
histologic report confirmed giant-cell tumor | -8760
total en bloc spondylectomy of T8 | 0
anterior-column reconstruction with titanium mesh | 0
structural allograft | 0
pedicle screw instrumentation from T6 to T10 | 0
eighth dorsal nerve routes sacrificed | 0
surgery duration 5 hours | 0
immediate postoperative period favorable | 0
no reported neurologic deficits | 0
pulmonary rehabilitation started by second postoperative day | 48
progressive dyspnea initiated by third postoperative day | 72
impaired gas exchange | 72
CT scan confirmed bilateral hemothorax | 72
bilateral thoracentesis | 72
recovery from symptoms | 72
worsening of general status by 19th postoperative day | 456
fever | 456
dyspnea | 456
decreased gas exchange | 456
increase in inflammatory markers | 456
CT scan revealed moderate fluid collection in both lungs | 456
empyema | 456
septic state | 456
transfer to intensive care unit | 456
surgical debridement of infected tissues | 456
allograft extraction | 456
titanium mesh extraction | 456
iliac crest tricortical autograft for anterior support | 456
posterior pedicle instrumentation kept | 456
copious irrigation of surgical wound | 456
drains placed in thoracic cavity | 456
drains placed in paravertebral spaces | 456
blood cultures identified Enterobacter aerogenes | 456
pus samples identified Enterobacter aerogenes | 456
explanted mesh samples identified Enterobacter aerogenes | 456
allograft samples identified Enterobacter aerogenes | 456
pathogen-directed i.v. antibiotic therapy initiated | 456
lower respiratory tract infection diagnosed 10 days after revision | 624
Acinetobacter baumannii identified in sputum samples | 624
septated empyema resurged in paravertebral space | 624
combined anterior and posterior approach for drainage | 624
posterior open drainage 12 days later | 960
subcutaneous abscess | 960
methicillin-resistant Staphylococcus aureus isolated | 960
Pseudomonas aeruginosa isolated | 960
discharge from hospital 79 days after initial admission | 1896
custom-molded thoracolumbar brace prescribed | 1896
physical therapy maintenance | 1896
asymptomatic after 9 months | 6552
no evidence of infection | 6552
no evidence of tumor relapse | 6552
follow-up imaging shows encouraging evolution | 6552
no bone graft resorption | 6552
no failure of instrumentation | 6552
