80 years old | 0
female | 0
admitted to the hospital | 0
abdominal pain | 0
vomiting | 0
barium meal examination | -24
peritoneal irritation signs | 0
tenderness | 0
guarding in the abdomen | 0
reduced white blood cell count | 0
increased serum C-reactive protein level | 0
sepsis | 0
abdominal X-ray | 0
barium leakage from the sigmoid colon | 0
abdominal computed tomography | 0
free air in the intraperitoneal cavity | 0
barium peritonitis with sigmoid colon perforation | 0
emergency surgery | 0
Hartmann’s procedure | 0
intraperitoneal drainage | 0
imipenem/cilastatin sodium | 0
doripenem | 0
serum CRP level decreased | 240
serum CRP level increased | 240
WBC count increased | 312
systemic CT examination | 312
methylprednisolone | 312
persistent inflammatory reaction | 312
WBC count improved | 315
serum CRP level improved | 315
discharged | 840