72 years old | 0
    female | 0
    nonalcoholic steatohepatitis | -1464
    duodenal varices | -1464
    portosystemic encephalopathy | -1464
    incomplete retrograde obliteration | -1464
    grade II encephalopathy | -1464
    plasma ammonia level 147 µg/dL | -1464
    ICG15 41% | -1464
    Hepatitis B surface antigen negative | -1464
    Hepatitis C virus antibody negative | -1464
    antinuclear antibody negative | -1464
    antimitochondrial antibody negative | -1464
    endoscopy revealed huge tortuous duodenal varices | -1464
    3D-CT showed duodenal varices supplied by right colic vein and pancreatoduodenal vein | -1464
    spleen volume 189 mL | -1464
    liver volume 595 mL | -1464
    spleen/liver volume ratio 0.32 | -1464
    portal vein diameter 7.0 mm | -1464
    splenic vein diameter 6.0 mm | -1464
    retrograde obliteration via internal jugular vein | -1464
    occlusive balloon catheter insertion into right ovarian vein | -1464
    obliteration attempt with microcoils, glucose, ethanol, ethanolamine oleate | -1464
    3D-CT post-obliteration showed incomplete obliteration | -1464
    encephalopathy improved to grade 0 | -1464
    plasma ammonia level reduced to 39 µg/dL | -1464
    febrile | 0
    drowsy | 0
    urinary incontinence | 0
    emergency admission | 0
    diagnosis of recurrence of hepatic encephalopathy | 0
    body temperature 39.7°C | 0
    disoriented | 0
    neck rigidity not evident | 0
    Kernig's sign negative | 0
    hemoglobin 9.7 g/dL | 0
    total leukocyte count 14500/µL | 0
    total platelet count 13.1 × 10^4/µL | 0
    total bilirubin 1.3 mg/dL | 0
    albumin 3.5 g/dL | 0
    aspartate transaminase 37 U/L | 0
    alanine transaminase 28 U/L | 0
    prothrombin time 91.6% | 0
    C-reactive protein 16.4 mg/dL | 0
    procalcitonin 30.8 ng/mL | 0
    serum ammonia 34 µg/dL | 0
    Child-Pugh score 9 (class B) | 0
    radiological investigation showed mild ascites | 0
    cerebral CT normal | 0
    endoscopy showed reduced duodenal varices | 0
    embolized coil partially migrated into duodenal lumen | 0
    lumbar puncture revealed purulent cerebrospinal fluid | 0
    cerebrospinal fluid cell count 1542/µL | 0
    cerebrospinal fluid sugar 31 mg/dL | 0
    cerebrospinal fluid proteins 540 mg/dL | 0
    bacterial meningitis diagnosis | 0
    bacteremia due to coil migration | 0
    admitted to intensive care unit | 0
    intravenous antibiotics (meropenem hydrate) | 0
    culture results positive for klebsiella aerogenes | 120
    antibiotics changed to cefepim | 120
    cefepim administered for 14 days | 120
    repeat blood and CSF cultures positive on day 5 | 120
    subsequent cultures negative on days 7, 9, 12 | 168, 216, 288
    anemia due to precursory bleeding from coil migration | 0
    risk of re-bleeding | 0
    trans-ileocolic vein obliteration attempted | 120
    right pararectal mini-laparotomy | 120
    sheath insertion into superior mesenteric vein | 120
    balloon catheter insertion into right colic vein | 120
    duodenal varices completely obliterated | 120
    portal venous pressure increased to 25.5 cmH2O | 120
    ascites increased | 120
    partial splenic embolization with 60% infarction | 288
    wedged hepatic venous pressure 23.0 cmH2O | 288
    3D-CT showed completed embolization of duodenal varices | 360
    spleen volume decreased to 85 mL | 360
    liver volume increased to 889 mL | 360
    corrected spleen/liver volume ratio 0.10 | 360
    portal vein diameter 9.0 mm | 360
    splenic vein diameter 5.0 mm | 360
    body temperature rose to 39.2°C | 600
    blood culture positive for klebsiella aerogenes | 600
    cefepim re-administered for 14 days | 600
    blood cultures negative on days 34 and 41 | 816, 984
    neurological status recovered by day 34 | 816
    ICG15 improved to 19% | 816
    discharged | 1008
    