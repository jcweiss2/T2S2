36 years old| 0
woman| 0
admitted to Hospital das Clínicas, University of São Paulo, Brazil | 0
pregnancy | 0
in vitro fertilization (IVF) performed | -840
attempted IVF three times without success | -840
IVF procedure complicated with mild OHSS | -840
mild OHSS did not require hospitalization or treatment | -840
unknown protocols for ovarian stimulation and ovulation induction | -840
abdominal enlargement | -840
oocyte retrieval (25 oocytes collected) | -840
two embryos transferred | -826
human albumin administered intravenously | -826
admitted to our service | -672
abdominal discomfort | -672
hyperemesis | -672
low urine output | -672
weight gain (7 kg in previous seven days) | -672
core temperature normal | -672
blood pressure normal | -672
abdomen distended | -672
ascites detectable during physical examination | -672
breathing normal | -672
oxygen saturation in room air normal | -672
small bilateral pleural effusions observed on thoracic radiographs | -672
transabdominal ultrasonographic examination at admission | 0
viable intrauterine twin pregnancy | 0
bilateral multiloculated cystic ovaries | 0
ascites | 0
hemoglobin 15 g/dL | 0
hematocrit 42.7% | 0
leukocyte count 18,540/mm3 | 0
platelet count 450,000/μL | 0
serum sodium 133 mmol/L | 0
potassium 4.7 mmol/L | 0
creatinine 0.6 mg/dL | 0
albumin 3.5 g/dL | 0
AST 45 IU/L | 0
ALT 27 IU/L | 0
bilirubin levels normal | 0
thyroid function normal | 0
serum E2 level 6,204 pg/mL | 0
human chorionic gonadotropin level 14,765 mIU/mL | 0
serology for viral hepatitis negative | 0
OHSS suspected | 0
supportive care in ICU initiated | 0
intravenous crystalloid hydration | 0
20% albumin (150 mL/day) started | 0
heparin (5,000 IU three times a day) administered | 0
thromboembolic prophylaxis | 0
patient responded well | 0
maintained adequate urine output | 0
hemoconcentration resolved | 0
discharged to obstetric ward | 168
developed fever | 168
shivering | 168
renal failure (creatinine 1.68 mg/dL) | 168
C-reactive protein increased from 42.7 to 116 mg/L | 168
respiratory compromise | 168
transvaginal paracentesis performed | 168
4 L of ascites aspirated | 168
fluid analysis revealed 520 cells/mm3 | 168
400 polymorphonuclear (PMN) cells/mm3 | 168
total protein concentration 5.0 g/dL | 168
Escherichia coli recovered from ascitic fluid culture | 168
ceftriaxone initiated | 168
human albumin administered at 1.5 g/kg on first day | 168
human albumin administered at 1.0 g/kg on third day | 168
general condition improved | 168
renal function improved | 168
no other source of infection discovered | 168
another transvaginal paracentesis | 216
discomfort from tense ascites alleviated | 216
fluid cell count improved (520/mm3 to 280/mm3) | 216
ceftriaxone discontinued | 264
remained in hospital for another month | 672
two further episodes of bacteremia | 672
blood cultures positive for Escherichia coli ESBL | 672
blood cultures positive for Acinetobacter baumannii | 672
E. coli treated with piperacillin/tazobactam | 672
A. baumannii treated with meropenem | 672
transvaginal paracentesis (5 L of ascites aspirated) | 672
albumin infusion for alleviation of abdominal hypertension and discomfort | 672
discharged from hospital | 1440
readmitted at 31 weeks of gestation | 1440
assessment of fetal vitality | 1440
premature rupture of membranes at 34 weeks | 1680
Caesarean section performed | 1680
mother and both babies discharged in good condition | 1728
