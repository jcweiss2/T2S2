65 years old | 0
male | 0
height: 165.2 cm | 0
body weight: 55 kg | 0
admitted to the hospital | 0
presumptive cholangiocarcinoma | 0
previously healthy | 0
unremarkable medical history | 0
elevated C-reactive protein | 0
total bilirubin 0.6 mg/dl | 0
direct bilirubin 0.3 mg/dl | 0
MELD score 6 | 0
axillary body temperature 36.7°C | 0
normal vital signs | 0
normal preoperative chest radiography | 0
normal transthoracic echocardiography | 0
tumor involving both the right and left intrahepatic bile duct and common bile duct | 0
enlarged lymph node around the common hepatic artery | 0
probable metastasis | 0
bilateral invasion of the bile duct | 0
tumor unresectable | 0
LDLT planned | 0
anesthesia induced | 0
intravenous thiopental sodium 350 mg | 0
atracurium 30 mg | 0
sevoflurane | 0
endotracheal intubation | 0
sevoflurane for anesthetic maintenance | 0
BIS monitored | 0
right radial artery cannulated | 0
right femoral artery cannulated | 0
right femoral vein cannulated | 0
warming blanket applied | 0
ambient temperature set at 25°C | 0
warming blanket temperature set at 40°C | 0
fluid warming system prepared | 0
body temperature monitored | 0
initial body temperature 36.7°C | 0
inhalant anesthetic changed to isoflurane | -30
anesthesia maintained with remifentanil | -30
anesthesia maintained with atracurium | -30
lymph node excised for frozen biopsy | -120
common bile duct clamped | -120
bile duct clamping | -120
common bile duct resected | -120
frozen biopsy negative for cancer cells | -60
LDLT continued | -60
donor hepatectomy started | -60
nasogastric tube placed | -60
AVA catheter inserted | -60
pulmonary artery catheter inserted | -30
body temperature not measured for half an hour | -30
last recorded skin temperature 36.9°C | -30
CBT measured with pulmonary artery catheter | 0
initial CBT 37.6°C | 0
fluid warming system turned off | 0
warming blanket set to cooling mode | 0
room temperature adjusted to 22°C | 0
donor hepatectomy converted to open hepatectomy | 30
massive bleeding from inferior vena cava | 30
CBT continuously rose to 39.5°C | 120
mild reactive tachycardia | 120
ETCO2 within normal range | 120
arterial blood gas analysis showed no acidosis | 120
no signs of malignant hyperthermia | 120
no signs of infection | 120
thyroid function tests normal | 120
BIS monitored | 120
hyperthermia discussed with surgeon | 120
surgeon suggested clamping of common bile duct as cause of hyperthermia | 120
bile drained | 210
CBT rapidly declined | 210
total duration of bile duct clamping 5 hours | 210
anhepatic phase started | 270
CBT 37.5°C | 270
CBT decreased to 36.9°C | 300
warming blanket turned on | 300
fluid warming system turned on | 300
room temperature set at 25°C | 300
CBT maintained at 36.7-37.3°C | 360
anesthesia time 14 hours | 840
patient received crystalloid | 840
patient received colloid solution | 840
patient received 5% albumin | 840
patient received cell saver blood | 840
urine output 2165 ml | 840
patient transferred to ICU | 840
body temperature at tympanic membrane 37.6°C | 840
WBC count slightly increased | 840
CRP 2.12 mg/dl | 840
total bilirubin 1.3 mg/dl | 840
direct bilirubin 0.9 mg/dl | 840
postoperative chest radiographs showed no remarkable interval change | 840
all cultures showed no growth of bacteria or fungus | 840
patient transferred to general ward on fifth postoperative day | 1200
no postoperative complications | 1200