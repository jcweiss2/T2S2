2 years old | 0
girl | 0
chromosomal abnormality of 1p36 deletion syndrome | 0
developmental delay | 0
intellectual disability | 0
seizures | 0
vision problems | 0
hearing problems | 0
distinctive facial features | 0
brain anomalies | 0
orofacial clefting | 0
congenital heart disease | 0
cardiomyopathy | 0
renal anomalies | 0
admitted to clinic for evaluation of gastroesophageal reflux | 0
pulmonary arterial banding at 4 weeks of age for ventricular septal defect | 0
Ebstein anomaly | 0
lip alveolus | 0
palate cleft | 0
laryngomalacia | 0
hypothyroidism | 0
psychomotor retardation | 0
gastroesophageal reflux | 0
home oxygen therapy | 0
tube feeding | 0
upper-gastrointestinal series on day 2 of admission | 0
fever | 48
diarrhea | 48
use of high-flow nasal cannula | 48
respiratory distress | 48
respiration stabilized | 48
circulation stabilized | 48
diarrhea resolved | 48
fever persisted | 48
higher fever (>39°C) between days 16 and 22 | 384
tachycardia (140–180 bpm) between days 16 and 22 | 384
mild lactate level elevation (2–4 mmol/L) between days 16 and 22 | 384
mild decrease of SpO2 to high 70% range between days 16 and 22 | 384
elevated blood urea nitrogen (39–54 mg/dL) between days 16 and 22 | 384
fever unexplained by mild dehydration | 384
tachycardia unexplained by mild dehydration | 384
preserved general condition | 384
preserved peripheral circulation | 384
marginal elevation of C-reactive protein level | 384
negative cultures | 384
no bacterial infection | 384
antibiotics not administered | 384
abrupt presentation of further higher fever (40–41°C) on day 23 | 552
respiratory distress on day 23 | 552
abdominal distention on day 23 | 552
hypotensive shock | 552
thrombocytopenia | 552
renal dysfunction | 552
liver dysfunction | 552
coagulation disorder | 552
mixed acidosis | 552
multiple-organ failure (MOF) | 552
disseminated intravascular coagulation (DIC) | 552
initiation of intensive care | 552
mechanical ventilation | 552
inotropes | 552
antibiotics | 552
decompression of stomach gas using nasogastric tube | 552
decompression of intestinal gas using Nélaton’s catheter | 552
accumulation of intestinal gas | 552
rapid extreme stiffening of abdomen | 552
complete loss of elasticity | 552
skin reddening on lower extremities | 552
skin reddening on lower abdomen | 552
circulatory failure in lower extremities | 552
circulatory failure in lower abdomen | 552
progression of MOF | 552
progression of DIC | 552
no urine produced after shock onset | 552
urine output 1.7 mL/kg/h prior to shock | 552
urine output more than 3.0 mL/kg/h previous 3 days | 552
assessment for open decompressive laparotomy | 552
advanced bleeding tendency | 552
inability to perform laparotomy | 552
death | 566
autopsy performed 23.5 h after death | 566
severe abdominal distention at autopsy | 566
extreme skin reddening on lower abdomen | 566
extreme skin reddening on lower extremities | 566
small amount of ascites | 566
intestinal dilation due to gas retention | 566
no organic intestinal tract obstruction | 566
intestinal mucosa macroscopically unremarkable | 566
localized dot hemorrhage in colonic mucosa | 566
congestion in intestinal wall | 566
no edema in intestinal wall | 566
no inflammation in intestinal wall | 566
extensive pneumonia | 566
accumulation of extensive intestinal gas unclarified | 566
secondary ACS induced by intestinal gas accumulation | 566
septic shock | 566
progression of pneumonia | 566
systemic inflammation induced by pneumonia | 566
triggering septic shock | 566
triggering DIC | 566
MOF progression | 566
DIC progression | 566
skin reddening on lower abdomen and extremities half a day before death | 566
abdominal distension progression | 566
severe abdominal distention contributing to circulatory failure | 566
IAP not measured | 566
no impeded blood flow on lower extremities prior to shock | 566
lack of apparent edema | 566
no muscle relaxant effect on abdomen stiffness | 566
diagnosis of secondary ACS | 566
accumulation of excessive intestinal gas | 566
no organic occlusive intestinal lesion | 566
no intestinal edema | 566
no bacterial pathogen identified | 566
no association with chromosomal abnormality | 566
sudden unexplained death | 566
lack of high-quality evidence for decision making | 566
IAP monitoring not performed | 566
fatal secondary ACS due to intestinal gas | 566
