18 years old | 0
female | 0
admitted to the emergency room | 0
alleged history of attempted suicide | -24
consumed paraquat | -24
difficulty in opening mouth | 0
decreased urine output | 0
no history of vomiting | 0
no history of loose stools | 0
no history of abdominal pain | 0
no history of seizures | 0
no history of fever | 0
conscious and oriented | 0
neck edema | 0
mucosal erosion of tongue | 0
mucosal erosion of palate | 0
mucosal erosion of lips | 0
oral bleeding | 0
pulse rate 98 beats per min | 0
blood pressure 130/80 mmHg | 0
respiratory rate 22 per min | 0
difficulty in breathing | 0
laryngeal edema | 0
intubated | 0
gastric lavage | 0
charcoal given | 0
elective ventilation | 0
IV fluids | 0
antiemetic | 0
high serum urea | 0
high serum creatinine | 0
dialysis | 24
normal thyroid function | 0
normal liver function | 0
normal urine examination | 0
bilateral grade I changes in kidneys | 0
normal 2D echo | 0
normal ECG | 0
corrosive injury to esophagus | 0
corrosive injury to proximal stomach | 0
Klebsiella pneumoniae | 48
intravenous methylprednisolone | 0
IV cyclophosphomide | 0
IV dexamethasone | 48
injection N-acetylcysteine | 0
vitamin C | 0
vitamin E | 0
expired | 288
septicemia | 288
respiratory failure | 288