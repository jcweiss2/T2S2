26 years old | 0
female | 0
Vietnamese descent | 0
admitted to the hospital | 0
widespread symmetric erythematous pustular eruption | 0
diffuse burning sensation | 0
facial swelling | 0
subjective fevers | 0
malaise | 0
mifepristone consumption | -48
tachycardia | 0
elevated temperature | 0
total lymphocyte count 18,000/mm3 | 0
absolute neutrophils 17,800/mm3 | 0
albumin 2.3 g/dL | 0
calcium 6.5 mg/dL | 0
alkaline phosphatase 31 U/L | 0
sodium 131 mmol/L | 0
potassium 3.2 mmol/L | 0
bicarbonate 19 mmol/L | 0
phosphorus 1.8 mg/dL | 0
glucose 179 mg/dL | 0
skin swab cultures negative | 0
blood cultures negative | 0
skin swab polymerase chain reaction negative | 0
quantitative human chorionic gonadotropin 1982.0 mIU/mL | 0
last reported menstrual period 5 weeks prior | -840
methylprednisolone treatment | 0
ceftriaxone treatment | 0
clindamycin treatment | 0
punch biopsy | 0
subcorneal pustules with neutrophil spongiosis | 0
papillary dermal edema with hemorrhage | 0
brisk perivascular mixed inflammatory infiltrate | 0
focal small-vessel vasculitis | 0
diagnosis of acute generalized exanthematous pustulosis | 0
diphenhydramine treatment | 0
triamcinolone treatment | 0
hypotension | 24
tachycardia | 24
admitted to critical care service | 24
central and arterial lines placement | 24
fluid resuscitation | 24
blood pressure recovery | 48
tachycardia resolution | 48
lines removal | 48
transferred to family medicine | 48
discharge | 72
pregnancy termination | 72 
no shortness of breath | 0
no mucous membrane involvement | 0
no target lesions | 0
no blisters | 0
no eosinophilia | 0
no visceral involvement | 0 
no hepatitis | 0
no nephritis | 0
no myocarditis | 0
no pneumonitis | 0