62 years old | 0
male | 0
HIV positive | 0
bioprosthetic aortic valve replacement | -12000
admitted to the hospital | 0
sepsis | 0
blood cultures positive for Staphylococcus aureus | 0
septic shock | 0
respiratory insufficiency | 0
renal failure | 0
CT-scan of the chest and abdomen | 0
transesophageal echocardiography (TEE) | 0
no endocarditis | 0
treatment with broad-spectrum antibiotics | 0
clinical condition improved | 168
discharged from ICU | 168
symptoms of a stroke | 168
CT detected a thromboembolism | 168
vegetation on the right coronary cusp of the aortic valve bioprothesis | 168
aortic root abscess | 168
neurological symptoms declined | 240
acute deterioration of the patient's hemodynamic conditions | 288
admitted to the intensive care unit | 288
high dose vasopressor therapy | 288
transthoracic echocardiography (TTE) | 288
shunting from the aortic root to the right atrium | 288
contrast enhanced computed tomography | 288
cardiac surgery | 288
removal of the bioprosthesis | 288
periannular abscess opening into the right atrium | 288
pericardial patch plasty | 288
new bioprosthesis implanted | 288
clinical status improved | 312
left the ICU | 456
discharged | 1344