20 years old | 0  
    woman | 0  
    primigravida | 0  
    transferred to our hospital | 0  
    breathing difficulty | -96  
    delivering a dead fetus | -96  
    intubated in emergency department | 0  
    respiratory distress | 0  
    shifted to critical care department | 0  
    no significant past medical history | 0  
    no significant genetic history | 0  
    no history of preeclampsia | 0  
    no history of gestational diabetes | 0  
    no history of infections during pregnancy | 0  
    Glasgow coma scale (GCS) E4M6Vt | 0  
    temperature 101°F | 0  
    pulse 122 beats/minute | 0  
    blood pressure 118/78 mm Hg | 0  
    no rash | 0  
    bilateral crepitations | 0  
    chest X-ray PA view bilateral infiltrates | 0  
    echo assessment poor LV systolic function | 0  
    echo assessment no RA/RV dilatation | 0  
    treated for pneumonia | 0  
    treated for sepsis | 0  
    treated for acute kidney injury (AKI) | 0  
    treated for peripartum cardiomyopathy | 0  
    hemodynamics improved | 0  
    cardiopulmonary-renal functions improved | 0  
    persistent high-grade fever | 0  
    gross muscle weakness | 120  
    all four limbs weakness | 120  
    predominantly proximal muscles weakness | 120  
    dark colored urine | 120  
    positive urine myoglobin | 120  
    raised ESR 47 mm/hour | 120  
    raised CPK 109,200 U/L | 120  
    raised LDH 460 U/L | 120  
    normal thyroid function tests | 120  
    SLE ruled out | 120  
    negative ANA | 120  
    negative anti-dsDNA antibody | 120  
    rhabdomyolysis differential diagnosis | 120  
    no major recovery with hemodialysis | 120  
    no major recovery with supportive measures | 120  
    proximal muscle weakness | 120  
    inflammatory myopathy suspected | 120  
    MRI cervical spine diffuse edema | 120  
    EMG myopathic pattern | 120  
    muscle biopsy inflammatory reaction | 120  
    endomysial infiltration with lymphocytes | 120  
    few necrotic muscle fibers | 120  
    polymyositis diagnosed | 120  
    IV steroids (methylprednisolone 1 g/day) | 120  
    prednisolone 60 mg/day | 120  
    tracheostomy performed | 240  
    responded well to steroids | 168  
    limbs power recovered progressively | 168  
    CPK levels decreased | 168  
    liberated from mechanical ventilator | 456  
    decannulated | 456  
    bulbar weakness persisted | 456  
    intermittent cough | 456  
    intolerance to oral feeds | 456  
    retained secretions | 456  
    videolaryngoscopy confirmed dysphagia | 456  
    cricopharyngeal muscle discordance | 456  
    feed through Ryles tube | 456  
    CPK levels decreased to 1066 U/L | 456  
    able to walk without support | 456  
    started oral feeds | 456  
    discharged | 456  
    tapering dose of oral steroids | 456  
    followed up after 2 weeks | 456  
    monthly follow-up | 456  
    prednisone 60 mg/day for 6 weeks | 456  
    steroid dose tapered every week by 5 mg for 8 weeks | 456  
    steroid dose tapered off by 2.5 mg every week | 456  
    counseled to avoid conception for a year | 456  
    fetal loss | 456  
    pregnancy as a trigger factor | 456  
    postpartum PM | 456  
    new onset PM | 456  
    differential diagnosis of puerperal fever | 456  
    pregnancy trigger new onset PM | 456  
    consent acquired | 456