33 years old | 0
female | 0
admitted for higher level of care | 0
acute respiratory failure | 0
mechanical ventilation | 0
methicillin sensitive Staphylococcus aureus bacteremia | 0
tricuspid valve endocarditis | 0
spontaneous right sided pneumothorax | -240
chest tube placement | -240
temperature 100.9 F | 0
pulse 113/min | 0
respiratory rate 18/min |
