85 years old | 0
female | 0
homemaker | 0
rheumatoid arthritis | -6720
hyperlipidemia | -6720
asthma | -6720
cerebrovascular accident | -144
received first dose of MODERNA COVID-19 vaccine | -720
minor pain at injection site | -720
received second dose of MODERNA COVID-19 vaccine | 0
generalized weakness | 12
muscle cramps | 12
loss of appetite | 12
nausea | 12
dark brown to black urine | 12
admitted to ER | 48
exhausted | 48
hypoactive bowel sounds | 48
mild abdominal tenderness | 48
elevated serum creatinine | 48
elevated BUN | 48
decreased GFR | 48
elevated AST | 48
elevated ALT | 48
elevated alkaline phosphatase | 48
elevated CPK | 48
elevated troponin | 48
myoglobin in urine | 48
started on bicarbonate-rich intravenous fluids | 48
heart failure with preserved ejection fraction | 48
started on broad-spectrum intravenous antibiotics | 72
temporary dialysis catheter inserted | 72
received hemodialysis | 72
started on empiric glucocorticoids | 96
cerebrospinal fluid analysis | 96
transferred to intensive care unit | 120
intubated on ventilator support | 120
cardiac arrest | 168
palliative care consultation | 168
terminally extubated | 168
died | 168
clopidogrel | -144
metoprolol | -144
nifedipine | -6720
rosuvastatin | -6720
telmisartan | -6720
tofacitinib | -144
trazodone | -144
physiotherapy | -144
non-weight bearing exercises | -144
family history of autoimmune disease | 0 
no previous history of tobacco or alcohol abuse | 0
no previous COVID-19 infection | 0
no recent history of trauma or surgery | 0
no recent over-the-counter medications | 0