87 years old | 0
female | 0
admitted to the emergency unit | 0
abdominal pain | -24
diarrhea | -24
hypertension | 0
third-degree atrioventricular block | 0
pacemaker | 0
fall | -24
dizziness | -24
lower abdominal pain | -24
watery stool | -24
right-sided pelvic pain | -24
blood pressure 122/50 mmHg | 0
pulse 63/min | 0
respiratory rate 20/min | 0
saturation 90% on room air | 0
temperature 35.5°C | 0
tenderness over the pubic bone | 0
tenderness over the lower abdomen | 0
no peritoneal reaction | 0
right hip region swelling | 0
right hip region tenderness | 0
normal rectal examination | 0
hemoglobin 6.5 mmol/l | 0
white blood cell count 10.6 × 109/l | 0
platelets 102 × 109/l |:0
creatinine 196 µmol/l | 0
C-reactive protein 29 mg/l | 0
pH 7.16 | 0
lactate 13.6 mmol/l | 0
X-ray of the pelvic region | 0
right-sided nondisplaced pubic ramus fracture | 0
arterial blood gas repeated after 9 hours | 9
pH 7.42 | 9
lactate 2.7 | 9
near normalization of blood gas parameters | 9
i.v. fluid administration | 9
pelvic fracture caused by fall due to severe dehydration and diarrhea | 9
condition worsened after 21 hours | 21
severe abdominal pain | 21
C-reactive protein increased to 123 mmol/l | 21
suspicion of intestinal ischemia | 21
exploratory laparotomy | 21
intra-operative detection of necrosis of sigmoid colon | 21
intra-operative detection of necrosis of proximal part of rectum | 21
flexible sigmoidoscopy | 21
non-vital mucosa 10–25 cm from anus | 21
non-vital ileum 20 cm from ileocecal region | 21
adherent non-vital ileum to rectosigmoid junction | 21
retroperitoneal hematomas in pelvic region | 21
no hematoma near inferior mesenteric artery | 21
resection of non-vital intestinal segments | 21
ileostomy performed | 21
sigmoideostomy performed | 21
minor bleeding during procedure | 21
postoperative severe sepsis | 21
intensive care unit admission | 21
recovery | 21
discharged | 240
histopathology showing necrosis due to ischemia | 21
no sign of vasculitis | 21
no sign of thrombosis | 21
