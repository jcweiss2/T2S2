37 years old | 0
male | 0
psychiatric history | 0
harmful use of alcohol | 0
harmful use of cocaine | 0
admitted to emergency services | 0
fell from the third floor of a building | -1
hemodynamically unstable | 0
aggressive fluid therapy | 0
X-rays of the pelvis | 0
X-rays of the thorax | 0
chest tube inserted | 0
pleural effusion | 0
serosanguineous fluid discharge | 0
Echo-FAST | 0
abundant free fluid | 0
transferred to the operating room | 0
emergency laparotomy | 0
4-liter hemoperitoneum | 0
active arterial bleeding | 0
complete avulsion of the hepatic artery | 0
multiple hepatic lacerations | 0
ligate the proper hepatic artery | 0
temporary abdominal closure | 0
vacuum pack technique | 0
admitted to the Resuscitation Unit | 0
hemodynamic recovery | 12
CT scan | 12
no neurological lesions | 12
absence of blood flow in the hepatic artery | 12
hepatic dysfunction | 12
ALT 3800 | 12
TBil 6 | 12
74000 platelets/μl | 12
IP 40% | 12
ischemic hepatitis | 12
abdomen closed definitively | 72
discharge of bile contents | 168
abdominal drainages | 168
suspicion of ischemic cholangiopathy | 168
transparietohepatic cholangiography | 168
destructuring of the intra- and extrahepatic bile duct | 168
ischemic cholangiopathy | 168
internal–external transhepatic drainage | 168
clinical improvement | 216
MRI | 216
multiple hepatic infarctions | 216
diffuse IC | 216
septic shock | 960
cholangitis | 960
multiple bilomas | 960
CT scan | 960
irreversible IC | 960
sepsis control | 960
waiting list for liver transplantation | 960
liver transplantation | 1680
biliary reconstruction | 1680
hepaticojejunostomy | 1680
re-operations | 1704
arteriographies | 1704
hemoperitoneum | 1704
bilateral mydriasis | 1816
decreased level of consciousness | 1816
brain CT scan | 1816
multiple bilateral ischemic lesions | 1816
right occipital hemorrhage | 1816
limit the therapeutic effort | 1816
died | 1816