70 years old | 0
male | 0
non-hypertensive | 0
non-smoker | 0
well-controlled diabetic | 0
HbA1c 6.83% | 0
presented for unresolving back pain | 0
COVID-19-induced pneumonia | -1440
slightly elevated white blood cell (WBC) 15,200/mm3 | 0
no abnormal monoclonal gammopathy | 0
contrast-enhanced chest-abdomen-pelvis computed tomography (CT) | 0
mediastinal calcified lymph nodes | 0
dense infiltrative retroesophageal prevertebral lesion | 0
retractile subpleural fibrous bands | 0
stepwise increase in WBC | 0
stepwise increase in C-reactive protein (CRP) | 0
broad spectrum antibiotherapy initiated | 0
dorsal MR conducted | 72
expanding prevertebral lesion from T2 till T9 | 72
tuberculosis testing negative | 0
HIV testing negative | 0
brucellosis testing negative | 0
blood culture negative | 0
serum galactomannan assay negative | 0
RT-PCR COVID-19 negative | 0
first percutaneous CT-guided biopsy inconclusive | 0
rising WBC count | 0
rising CRP | 0
control dorsal MR carried out | 240
slight progression of the lesion | 240
empirical antifungal therapy with fluconazole and amphotericin B initiated | 336
second CT-guided biopsy performed | 408
necrotic lesions observed | 408
fungal organisms with acute-angle-branching hyphae observed | 408
culture showed growth of Aspergillus fumigatus | 408
antifungal therapy switched to voriconazole | 432
dosage 400 mg b.i.d. for the first day | 432
dosage reduced to 200 mg b.i.d. | 456
surgical thoracotomy not executed | 432
CRP levels decreased | 432
increasing levels of creatinine | 432
progressive oliguria | 432
hemodialysis sessions | 432
acutely developed paraplegia | 552
altered mental state | 552
ICU transfer | 552
head CT performed | 552
no focal abnormality in the brain parenchyma | 552
adequate gray matter-white matter differentiation | 552
lumbar puncture | 552
sterile cultures | 552
dorsal MR performed | 552
recent spinal cord compression at T6 to T8 | 552
antifungal treatment insufficient | 552
renal function deteriorating | 552
neurological function deteriorating | 552
comatose | 672
intubated | 672
passing away | 672
