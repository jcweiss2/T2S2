intermittent high-grade fever | -72
generalized dull-aching abdominal pain | -72
passing turbid urine | -240
decrease in urine output | -240
swelling of both feet | -240
treated with intravenous medications | -168
type II diabetes mellitus | 0
conscious | 0
afebrile | 0
tachycardic with heart rate of 136/min | 0
renal angle tenderness bilaterally | 0
high total leukocyte counts with left shift | 0
elevated urea and creatinine levels | 0
pyuria with leukocyte esterase positivity | 0
activated partial thromboplastin time was prolonged | 0
sepsis-induced coagulopathy | 0
enlarged kidneys with bilateral renal abscesses | 0
emergency ultrasound-guided drainage of renal abscesses | 12
transfusion of blood products | 12
coagulopathy | 12
pus smear from renal abscesses from both sides showed septate fungal hyphae | 24
initiated on intravenous meropenem | 0
initiated on intravenous voriconazole | 24
initiated on intravenous amphotericin B | 24
cultures from both renal abscesses revealed growth of Aspergillus fumigatus | 48
worsening renal function | 72
acute pulmonary edema | 72
hyperkalemia | 72
metabolic acidosis | 72
initiated on hemodialysis | 72
initiated on noninvasive ventilation | 72
sudden cardiac arrest | 216
aspiration | 216
death | 216