47 years old | 0
    obese | 0
    woman | 0
    BMI of 42 | 0
    large incisional hernia at midline laparotomy | 0
    referred for laparoscopic correction | 0
    hypertension | 0
    transabdominal gynecologic surgery | 0
    peripheral vascular disease | 0
    multiple angioplasties of the iliac arteries | 0
    carbon dioxide used to create pneumoperitoneum | 0
    intraabdominal pressure maintained at 12mm Hg | 0
    laparoscopic correction | 0
    extensive adhesiolysis | 0
    15-minute break | 120
    decompression of the abdomen | 120
    total duration of the pneumoperitoneum 215 minutes | 0
    blood pressure remained stable | 0
    hernia defect measured 20 cm × 16 cm | 0
    application of two 30cm×20cm expanded polytetrafluoroethylene meshes | 0
    meshes fixed with tackers | 0
    meshes fixed with transabdominal sutures | 0
    recovery was uneventful | 0
    postoperative day 3 | 72
    paralytic ileus | 72
    no localized tenderness | 72
    plain abdominal x-ray | 72
    ultrasound showed distended bowel | 72
    C-reactive protein significantly raised | 72
    relaparoscopy | 72
    intraabdominal pressure maintained at 12 mm Hg | 72
    procedure took not more than 12 minutes | 72
    bowel distension | 72
    no signs of contamination | 72
    no perforation | 72
    no ischemia | 72
    no action undertaken | 72
    systemic inflammatory response syndrome | 72
    respiratory insufficiency | 72
    transfer to intensive care unit | 72
    stabilized | 72
    required less support | 72
    no apparent infection | 72
    postoperative day 9 | 216
    bloody diarrhea | 216
    colonoscopy | 216
    severe ischemic colitis in the transverse colon | 216
    mesenteric angiography | 216
    occluded superior mesenteric artery | 216
    compensatory distended inferior mesenteric artery | 216
    pinpoint stenosis at origin | 216
    balloon angioplasty | 216
    anticoagulants | 216
    steadily improved | 216
    5 days later | 288
    situation deteriorated | 288
    another colonoscopy | 288
    multiple perforations of the ischemic transverse colon | 288
    laparotomy | 288
    fecal peritonitis | 288
    multiple perforations of the ischemic ascending and transverse colon | 288
    resection of the ischemic colon | 288
    removal of contaminated meshes | 288
    postoperative deterioration | 288
    death | 384
    histological examination of resected bowel | 384
    extensive ischemia | 384
    multiple transmural ulcerations | 384
    multiple perforations | 384
    no autopsy | 384
    <|eot_id|>