89 years old | 0
    male | 0
    vomiting | -96
    epigastric distension | -96
    no bowel movements | -96
    no flatus | -96
    gallstones | -87600
    right upper quadrant pain | -87600
    hypertension | -87600
    diabetes | -87600
    pulmonary tuberculosis | -420000
    schistosomiasis | -420000
    moderate drinking | 0
    no smoking | 0
    no allergies | 0
    unremarkable family history | 0
    temperature 36.2 °C | 0
    heart rate 77 beats per min | 0
    respiratory rate 20 breaths per min | 0
    blood pressure 137/74 mmHg | 0
    abdominal tenderness | 0
    no rebound tenderness | 0
    hyperactive bowel sounds | 0
    normal lung examination | 0
    normal heart examination | 0
    normal routine blood examination | 0
    normal liver function | 0
    normal renal function | 0
    normal coagulation function | 0
    normal troponin | 0
    normal procalcitonin | 0
    high-sensitivity C-reactive protein increased (26.1 mg/L) | 0
    abdominal CT showed cholecystoduodenal fistula | 0
    abdominal CT showed jejunal gallstone ileus | 0
    abdominal CT showed pneumobilia | 0
    cholecystitis | 0
    Rigler’s triad | 0
    ceftriaxone sodium and sulbactam sodium administered | 0
    octreotide acetate administered | 0
    esomeprazole administered | 0
    nasogastric tube inserted | 0
    gastrointestinal decompression | 0
    nutrition support | 0
    amino acid administered | 0
    lipid emulsion administered | 0
    no indication for emergency surgery | 0
    propulsive enteroscopy performed (first time) | 0
    deep ulcer in duodenal bulb | 0
    yellow purulent secretion | 0
    mucosal edema | 0
    stone incarceration in upper jejunum | 0
    food residue proximal to gallstone | 0
    basket and snare used to remove food residue | 0
    failed to remove stone | 0
    laser lithotripsy performed (first time) | 0
    sodium bicarbonate injected (first time) | 0
    propulsive enteroscopy performed (second time) | 24
    stone smaller than before | 24
    laser lithotripsy performed (second time) | 24
    sodium bicarbonate injected (second time) | 24
    no passage of gas | 168
    gastrointestinal decompression drainage 800-1000 mL per day | 168
    transferred to Department of Biliary-pancreatic Surgery | 168
    laparoscopic duodenoplasty | 408
    cholecystectomy | 408
    enterolithotomy | 408
    repair | 408
    severe inflammation and edema around gallbladder | 408
    jejunal gallstone ileus confirmed | 408
    gallbladder removed | 408
    cauliflower drainage tube placed | 408
    purse-string suturing performed | 408
    jejunum cut | 408
    gallstone removed | 408
    intestine wall sutured | 408
    drainage tubes placed | 408
    tachycardia (170 beats per min) | 432
    normal white blood cell count | 432
    mild anemia (hemoglobin 117.0 g/L) | 432
    hypoproteinemia (32.5 g/L) | 432
    urea elevated (14.74 mmol/L) | 432
    creatinine elevated (149 µmol/L) | 432
    NT-proBNP elevated (5458 pg/mL) | 432
    normal troponin | 432
    atrial fibrillation | 432
    pulmonary arterial hypertension (44 mmHg) | 432
    enlargement of right heart | 432
    tricuspid insufficiency | 432
    deslanoside administered | 432
    amiodarone hydrochloride administered | 432
    sinus rhythm restored | 432
    hypourocrinia | 432
    anuric | 432
    transferred to intensive care unit | 432
    hyperpyrexia (39 °C) | 432
    disturbance of consciousness | 432
    white blood cell count increased (10.11 × 109 cells/L) | 432
    neutrophilic granulocyte percentage 90.5% | 432
    prothrombin time prolonged (57.9 s) | 432
    international normalized ratio elevated (6.02) | 432
    troponin elevated (5476.8 pg/mL) | 432
    NT-proBNP elevated (31194 pg/mL) | 432
    creatinine elevated (347 µmol/L) | 432
    procalcitonin elevated (31.01 ng/mL) | 432
    high-sensitivity C-reactive protein increased (220.0 mg/L) | 432
    Enterococcus faecium cultured | 432
    meropenem administered | 432
    tigecycline administered | 432
    linezolid administered | 432
    teicoplanin administered | 432
    continuous renal replacement therapy | 432
    plasma transfusion | 432
    coronary dilating drugs | 432
    abdominal tenderness | 432
    rebound tenderness | 432
    exudate around drainage tube | 432
    hypotension | 432
    drainage tube replaced | 432
    noradrenaline administered | 432
    pituitrin administered | 432
    platelet count decreased | 432
    teicoplanin administered | 432
    urine volume recovered | 432
    vital signs stable | 432
    white blood cell count decreased (2.48 × 109 cells/L) | 456
    moderate anemia (hemoglobin 61.0 g/L) | 456
    creatinine elevated (225 µmol/L) | 456
    troponin elevated (44.7 pg/mL) | 456
    NT-proBNP elevated (3229 pg/mL) | 456
    procalcitonin elevated (1.74 ng/mL) | 456
    transferred to Department of Biliary-pancreatic Surgery | 456
    cefoperzone sodium and tazobactam sodium administered | 456
    lethargy | 504
    mouth breathing | 504
    coma | 528
    pupils unresponsive to light | 528
    abdominal CT postoperative changes | 528
    exudative effusion around operative region | 528
    chest CT infection in right lung | 528
    head CT cerebral infarction | 528
    transferred to intensive care unit | 528
    anti-infective therapy | 528
    enteral nutrition | 528
    electrolytes maintenance | 528
    oxygen therapy | 528
    blood pressure decreased | 576
    oxyhemoglobin saturation decreased | 576
    death | 576