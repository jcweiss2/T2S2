38 years old | 0
Afro-Caribbean female | 0
admitted to the hospital | 0
bleeding from an ulcerating left fungating parotid tumour | 0
pea-sized mass | -8760
fine-needle aspiration cytology | -8760
ACC | -8760
refused surgery | -8760
lost to follow-up | -8760
tumour slowly increased in size | -8760
rapid growth | -168
malnourished | 0
14 by 12 cm fungating parotid mass | 0
areas of necrosis | 0
haemorrhage | 0
hemoglobin 9.3 g/L | 0
albumin level <10 g/L | 0
electrolytes normal | 0
liver function tests normal | 0
coagulation profile normal | 0
nutritional support | 0
hemostasis | 0
acute confusion | 48
agitated | 48
thrombosis of the contralateral transverse sinus | 48
thrombosis of the distal part of the right common femoral vein | 48
warfarin | 48
inferior vena caval filter | 48
INR 8.0 | 288
bleeding from the tumour site | 288
warfarin stopped | 288
Vitamin K | 288
fresh-frozen plasma | 288
INR 2.0 | 336
warfarin switched to low-molecular-weight heparin | 336
platelet count dropped | 432
heparin-induced thrombocytopenia | 432
lepirudin | 432
platelets returned to normal | 444
septicemia | 456
broad-spectrum antibiotics | 456
radical left-sided parotidectomy | 672
type-1 modified radical neck dissection | 672
latissimus dorsi pedicled muscle flap reconstruction | 672
facial nerve sacrificed | 672
accessory nerve preserved | 672
internal jugular vein preserved | 672
zygomatic arch removed | 672
tumour herniating into the oral cavity | 672
oral mucosa excised | 672
split skin graft | 672
histology confirmed moderately differentiated ACC | 672
vascular invasion | 672
lymph nodes harvested | 672
disease staged as pT4pN0M0 | 672
hematoma formation | 720
septicemia due to infected central venous catheter | 720
antibiotics | 720
split skin graft re-grafted | 720
discharged | 1560
normalized serum albumin level | 1560
adjuvant postoperative radiotherapy | 1560
no signs of local or regional disease | 1560
lung metastasis | 4560
died | 4560