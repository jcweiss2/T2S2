67 years old | 0
female | 0
resident of Goiânia, Goiás (Brazil) | 0
rheumatoid arthritis | 0
hydroxychloroquine use (400 mg daily for 4 years) | 0
denies history of diabetes mellitus | 0
denies history of high blood pressure | 0
denies smoking | 0
denies alcohol consumption | 0
traveled to Italy | -1344
returned to Brazil | -1320
unverified fever | -1320
dry cough | -1320
malaise | -1320
RT-qPCR test for COVID-19 (Biopur®) | -1296
presented to emergency room | -1224
hospitalized | -1224
fever | -1224
chills | -1224
nausea | -1224
diagnosis of COVID-19 confirmed by RT-qPCR | -1200
chest computed tomography (CT) | -1200
ground-glass opacities | -1200
consolidations involving more than 75% of lung volume | -1200
oseltamivir started | -1224
enoxaparin started | -1176
transferred to ICU | -1152
respiratory failure | -1152
SARS diagnosis | -1152
azithromycin started | -1152
piperacycline with tazobactam started | -1152
mechanical ventilation | -1152
septic shock with pulmonary focus | -1152
meropenem started | -1056
chest CT scan on April 14 | 432
radiological improvement | 432
extubated | 576
regained consciousness | 576
noticed hearing loss in right ear | 576
discharged from ICU | 648
discharged from hospital | 816
audiometry on August 27, 2019 | -6720
hearing loss at 6 and 8 kHz in right ear | -6720
normal thresholds in left ear | -6720
evaluated by otorhinolaryngologist | 1296
normal otoscopic findings | 1296
disabling tinnitus | 1296
severe sensorineural hearing loss in right ear | 1296
isolated hearing loss at 4 and 8 kHz in left ear | 1296
impedance testing (type A curve) | 1296
no bilateral contralateral stapedial acoustic reflexes | 1296
combined corticosteroid therapy (oral and intratympanic) | 1296
prednisolone (60 mg for 7 days) | 1296
prednisolone (40 mg for 7 days) | 1296
prednisolone (20 mg for 5 days) | 1296
prednisolone (10 mg for 5 days) | 1296
intratympanic dexamethasone applications | 1296
topical anesthesia with 2% tetracaine spray | 1296
44% phenol on eardrum | 1296
increased blood pressure during corticosteroid therapy | 1296
blood pressure normalized after oral corticosteroid | 1296
no other adverse effects | 1296
brain MRI on May 20, 2020 | 1344
multiple microhemorrhagic lesions | 1344
splenium of corpus callosum | 1344
cerebellum | 1344
medium cerebellar peduncles | 1344
subcortical white matter | 1344
no ischemic injuries | 1344
no changes in auditory canal | 1344
magnetic resonance angiography of brain and neck | 1344
no changes | 1344
audiometry on June 23, 2020 | 1728
improvement in 250 kHz in right ear | 1728
improvement in 4, 6, and 8 kHz in left ear | 1728
persistent tinnitus | 1728
