18 years old | 0
female | 0
born at 24 weeks + 3 days | -720
via emergent cesarean delivery | -720
breech presentation | -720
cord prolapse | -720
birth weight of 645 g | -720
HIV negative | -720
mother 36 years old | -720
Apgar score of 4 | -720
Apgar score of 8 | -720
mechanical ventilation | -720
central umbilical catheters | -720
total parenteral nutrition | -720
empiric antibiotics | -720
skin sensors for monitoring | -720
late-onset sepsis | -720
Escherichia coli bacteremia | -720
cefepime | -720
day of life 9 | -720
day of life 20 | -720
skin abrasion | -720
erythema | -720
induration | -720
plaque with a necrotic center | -720
ulcer | -720
extension to subcutaneous cell tissue | -720
necrotic area | -720
thermic instability | -720
metabolic acidosis | -720
hyperglycemia | -720
hypotension | -720
suspected mucormicosis | -720
liposomal amphotericin B (L-AmB) | -720
fungal biomarkers | -720
serum galactomannan | -720
1,3 beta-D-glucan | -720
skin biopsy | -720
microbiological and pathological studies | -720
refractory shock | -720
metabolic acidosis | -720
renal failure | -720
died | 36
Rhizopus spp. | -720
broad aseptate hyphae | -720
right angle branching | -720
MALDI-TOF MS | -720
polymerase chain reaction (PCR) | -720
sequencing region D1/ D2 -24S RNA long subunit- | -720
internal transcribed spacer region | -720
Rhizopus arrhizus | -720
fungal blood cultures | -720
negative | -720
superficial infection | -720
vesicle or pustule | -720
erythematous plaque | -720
ulcerate | -720
gangrenous form | -720
painful papule | -720
necrotizing cellulitis | -720
necrotic plaque | -720
necrotic eschar | -720
skin abscesses | -720
premature infant | -720
immunocompromised hosts | -720
diabetes | -720
invasive and fatal infections | -720
inmate and adaptative immune systems | -720
immaturity | -720
parenteral nutrition use | -720
antibiotic use | -720
orogastric tubes | -720
venous catheters | -720
skin sensors | -720
cutaneous aspergillosis | -720
hyalohyphomycosis | -720
Fusarium | -720
necrotizing fasciitis | -720
clostridial gas gangrene | -720
sepsis-associated purpura fulminans | -720
bacterial cellulitis | -720
pyoderma gangrenosum | -720
culture and histopathology | -720
tissue biopsy | -720
laboratory processing | -720
routine culture media | -720
broad, hyaline and aseptate hyphae | -720
vascular invasion | -720
necrotic tissue | -720
PCR assays | -720
mass spectrometry tests | -720
MALDI-TOF MS | -720
identification of the fungus | -720
species level | -720
surgical debridement | -720
anti-fungal treatment | -720
L-AmB | -720
associated or not with another agent | -720
ischemic necrosis | -720
infected tissue | -720
arrival of leukocytes | -720
anti-fungal agents | -720
site of infection | -720
pediatric patients | -720
pooled data | -720
antifungal therapy | -720
surgical debridement | -720
lower risk of death | -720
death | -720
aggressive approach | -720
infection control | -720
traditional diagnostic methods | -720
microbiology and histopathology | -720
modern tests | -720
mass spectrometry | -720
molecular studies | -720
rapid and accurate etiological diagnosis | -720