31 years old | 0
pregnant | 0
no family history of congenital heart disease | 0
referred to centre | 0
foetal aortic valve stenosis | -112
detected at 18 + 0 weeks of gestation | -112
maternal transabdominal foetal ultrasound imaging | -56
severe foetal aortic valve stenosis | -56
poorly contracting dilated left ventricle | -56
severe mitral valve regurgitation | -56
local endocardial fibroelastosis | -56
mitral valve inflow biphasic | -56
regurgitant velocity exceeded 4 m | -56
maximum systolic flow velocity across aortic valve 2 m/s | -56
flow across oval foramen left to right | -56
flow inside aortic arch retrogradely | -56
percutaneous ultrasound-guided foetal balloon valvuloplasty attempted | -24
general maternofoetal anaesthesia | -24
function of left ventricle deteriorated | -24
mitral valve flow integral exhibited mostly a-wave filling | -24
foetus lying in dorsoanterior cephalic position | -24
left ventricle pointed posteriorly | -24
foetoscopic assistance employed | -24
three 11 Fr catheter sheaths placed | -24
amniotic cavity insufflated with carbon dioxide | -24
foetus rotated in dorsoposterior position | -24
upper extremities postured along foetal sides | -24
insufflation gas removed | 0
18 gauge needle advanced into foetal left ventricle | 0
needle placed underneath obstructed aortic valve | 0
successful foetal balloon valvuloplasty achieved | 0
mother and foetus tolerated procedure well | 0
no complications observed | 0
interventional materials removed | 0
maternal skin incisions closed | 0
marked improvement of flow across aortic valve | 24
increase in flow velocity from 1.75 m/s to more than 3 m/s | 24
foetus delivered in third week after prenatal intervention | 504
scheduled for postnatal re-valvuloplasty on second day of life | 504
stent insertions in ductus arteriosus and atrial septum | 504
insertion of flow occluders into both pulmonary branches | 504
left ventricular function improved over time | 504
baby died at 6 months of age | 1008
Escherichia coli septicaemia | 1008
long-standing central venous line | 1008
cardiac surgery addressing mitral valve regurgitation and branch pulmonary artery obstruction | 1008
parental informed consent obtained | -24
procedure performed in accordance with Declaration of Helsinki | -24