45 years old | 0
male | 0
Asian | 0
admitted to the hospital | 0
fever | -144
cough | -144
dyspnoea | -144
diarrhoea | -144
vomiting | -144
abdominal pain | -144
bilateral crackles on lung bases | 0
severe pain located in the epigastrium | 0
rigidity and guarding of the abdominal wall | 0
SpO2 82% on room air | 0
heart rate 109 beats per minute | 0
blood pressure 89/47 mm Hg | 0
intubated | 0
mechanically ventilated | 0
resuscitated with low-dose noradrenaline and crystalloid fluids | 0
SARS-CoV-2 infection | 0
leukocytosis | 0
lymphocytopenia | 0
increased C-reactive protein | 0
increased lactate dehydrogenase | 0
increased lactate | 0
increased d-dimers | 0
blood urea nitrogen 6.1 mmol/L | 0
creatinine 119 μmol/L | 0
chest CT scans revealed bilateral peripheral ground-glass opacities | 0
pulmonary embolism | 0
abdominal CT scans depicted thickened bowel wall | 0
portal vein thrombosis | 0
emergency exploratory laparotomy | 12
contained small intestinal perforation | 12
peritonitis | 12
resection of an ischaemic area of the jejunum | 12
histopathologic examination revealed epithelial necrosis | 12
haemorrhagic infarction changes | 12
neutrophilic inflammation | 12
fibrin deposition | 12
admitted to ICU | 12
administered empiric therapy with ribavirin | 12
meropenem | 12
vancomycin | 12
therapeutic anticoagulation with enoxaparin | 12
ARDS-net ventilation | 12
administration of hydrocortisone | 12
vasopressors | 12
supportive ICU care | 12
developed acute kidney injury | 24
blood urea nitrogen 7.9 mmol/L | 24
creatinine 309 μmol/L | 24
mild metabolic acidosis | 24
hyperkalaemia | 24
anuric | 24
state of shock | 24
administered CRRT | 24
extracorporeal blood purification therapy with CytoSorb filter | 24
transfused with two packs of red blood cells | 24
initiated diuresis | 72
weaned off vasopressors | 72
lactate level normalized | 72
inflammatory biomarkers normalized | 72
CRRT discontinued | 72
extubated | 168
renal function normalized | 336
RT-PCR for COVID-19 negative | 456
discharged from hospital | 816
prescribed oral rivaroxaban | 816