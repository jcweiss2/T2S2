preterm baby boy | 0
born by vaginal delivery | 0
32 weeks of gestation | 0
antenatal steroids | -168
premature rupture of membranes | -168
spontaneous labour | -168
Apgar 9-10 | 0
examination normal at birth | 0
birth weight 1800 g | 0
head circumference 30.5 cm | 0
admitted to neonatal intensive care unit | 0
orally fed | 0
elevated procalcitonin | 0
received antibiotics | 0
fever | 24
screeches | 24
C-reactive protein 77 mg/L | 24
white blood cell 4.81 x 10^9/l | 24
lumbar puncture normal | 24
haemoculture positive for Gram-negative bacillus | 24
intubated | 48
severe apnoea | 48
altered hemodynamic status | 48
painful distended and contractured abdomen | 48
large gastric residual | 48
clear gastric residual appearance | 48
regular stools | 48
normal stools | 48
abdominal X-ray non-abnormal | 48
ultrasound non-abnormal | 48
C-reactive protein 155 mg/L | 48
normal white blood cell | 48
thrombocytopenia | 48
exploratory laparotomy | 48
perforated appendicitis | 48
peritonitis | 48
appendectomy | 48
peritoneal lavage with warm saline | 48
favourable outcome | 72
histopathology confirmed diagnosis | 72
no signs of Hirschprung's disease | 72
follow-up at 5 months of age | 2160
reassuring follow-up | 2160