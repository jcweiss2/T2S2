43 years old | 0
male | 0
schizophrenia | 0
asthma | 0
polysubstance use disorder | 0
ongoing IVDU | 0
presented to the institution | 0
fever | 0
chills | 0
left-sided pleuritic chest pain | 0
admission for methicillin-sensitive Staphylococcus aureus TV endocarditis | -25920
paraspinal abscess | -25920
percutaneous drainage | -25920
6 weeks of intravenous antibiotic therapy | -25920
arrival | 0
febrile | 0
tachycardic | 0
normotensive | 0
adequate oxygen saturation on room air | 0
started on intravenous antimicrobial therapy | 0
transthoracic echocardiography | 0
30-mm mobile mass on the TV | 0
vegetation | 0
evaluated by a multidisciplinary heart valve team | 0
management of schizophrenia | 0
management of substance use disorder | 0
7 days of appropriate antimicrobial therapy | 0
continued febrile | 168
positive blood cultures | 168
repeat computed tomography scans | 168
ongoing septic pulmonary emboli | 168
tricuspid valve replacement offered | 168
refused open surgical procedure | 168
decision to debulk the TV vegetation | 168
consent obtained | 168
taken to a hybrid operating room | 168
general anesthesia | 168
endotracheal tube | 168
left-sided central venous catheter | 168
TEE guidance | 168
intraoperative preprocedural TEE imaging | 168
vegetation measuring 32 × 26 mm | 168
attached to the septal and anterior leaflets | 168
mild TR | 168
normal right ventricular systolic function | 168
TV annulus measured at 37 mm | 168
no vegetations on other cardiac valves | 168
AngioVac vacuum-assisted thrombectomy system | 168
right internal jugular and femoral venous access | 168
fluoroscopy | 168
inflow cannula advanced to TV vegetation | 168
extracorporeal circulation | 168
flows of 2-3 L/min | 168
real-time debulking observed | 168
additional manipulations of the inflow cannula | 168
satisfactory debulking | 168
flow stopped | 168
largest components removed | 168
small residual components | 168
moderate TR postprocedure | 168
no structural damage noted | 168
vegetation retrieved for culture | 168
hemodynamically stable | 168
vegetation cultures positive for methicillin-sensitive Staphylococcus aureus | 168
6 weeks of antibiotic therapy | 168
started on suboxone | 168
discharged to a family member’s home | 168
represented with methicillin-resistant Staphylococcus aureus bacteremia | 3024
transesophageal echocardiography | 3024
no abscess | 3024
no worsening vegetation | 3024
6 weeks of antimicrobial therapy | 3024
discharged home | 3024
stable condition | 3024
no further interventions | 3024
