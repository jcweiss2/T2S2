57 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
lepromatous leprosy | -720 | -720 | Factual
treatment with rifampicin/clofazimine/dapsone | -720 | 0 | Factual
abdominal distension | 0 | 0 | Factual
constipation | 0 | 0 | Factual
vomiting | 0 | 0 | Factual
10-kg weight loss | -720 | 0 | Factual
peripheral lymphadenopathy | 0 | 0 | Factual
distended abdomen | 0 | 0 | Factual
positive shifting dullness | 0 | 0 | Factual
mural thickening of the terminal ileum | 0 | 0 | Factual
enlarged mesenteric lymph nodes | 0 | 0 | Factual
mesenteric fat stranding | 0 | 0 | Factual
intra-abdominal free fluid | 0 | 0 | Factual
abdominal granulomatous infection | 0 | 0 | Possible
neoplastic process | 0 | 0 | Possible
abdominal paracentesis | 0 | 0 | Factual
atypically large lymphocytes | 0 | 0 | Factual
high-grade lymphoma | 0 | 0 | Factual
flow cytometry | 0 | 0 | Factual
abnormal CD4/CD8 double-negative T-cell population | 0 | 0 | Factual
cervical lymph node biopsy | 0 | 0 | Factual
high-grade peripheral T-cell lymphoma | 0 | 0 | Factual
bone marrow examination | 0 | 0 | Factual
no involvement of T-cell NHL | 0 | 0 | Factual
stage IV lymphoma | 0 | 0 | Factual
dexamethasone | 0 | 0 | Factual
tumor-lysis syndrome precautions | 0 | 0 | Factual
severe sepsis | 24 | 24 | Factual
transfer to medical ICU | 24 | 24 | Factual
antibiotics | 24 | 168 | Factual
antifungals | 24 | 168 | Factual
ICU care | 24 | 168 | Factual
EPOCH chemotherapy protocol | 168 | 1008 | Factual
CNS prophylaxis | 168 | 1008 | Factual
intrathecal methotrexate | 168 | 1008 | Factual
complete metabolic remission | 1008 | 1008 | Factual
febrile neutropenia episodes | 1008 | 1200 | Factual
recurrent bacteremia | 1008 | 1200 | Factual
generalized weakness | 1008 | 1008 | Factual
no sensory changes | 1008 | 1008 | Factual
no clear fatigability | 1008 | 1008 | Factual
decreased power in proximal and distal muscles | 1008 | 1008 | Factual
normal distal latencies | 1008 | 1008 | Factual
normal compound muscle action potential | 1008 | 1008 | Factual
normal conduction velocities | 1008 | 1008 | Factual
normal F waves | 1008 | 1008 | Factual
normal sensory nerve studies | 1008 | 1008 | Factual
needle electromyogram | 1008 | 1008 | Factual
poor recruitment effects | 1008 | 1008 | Factual
repetitive nerve stimulation | 1008 | 1008 | Factual
significant incremental response | 1008 | 1008 | Factual
presynaptic neuromuscular junction disorder | 1008 | 1008 | Possible
LEMS | 1008 | 1008 | Possible
intravenous immunoglobulins | 1008 | 1012 | Factual
improvement of motor function | 1012 | 1012 | Factual
ambulation | 1012 | 1012 | Factual
consolidation by autologous bone marrow transplant | 1200 | 1200 | Factual
recurrent bacteremia and sepsis | 1200 | 1200 | Factual
multiorgan failure | 1200 | 1200 | Factual
death | 1200 | 1200 | Factual