28 years old | 0
female | 0
8 weeks pregnant | 0
admitted to the hospital | 0
acute severe asthma | -1
short non-infective prodrome | -1
hypoxic cardiac arrest | -1
ventricular fibrillation | -1
resuscitation to sinus tachycardia | -1
endotracheal intubation | -1
therapeutically cooled to 33°C | 0
salbutamol | 0
ipratropium | 0
aminophylline | 0
hydrocortisone | 0
magnesium | 0
ketamine | 0
inhalation anesthesia with 1 MAC isoflurane | 0
severe hypercapnic acidosis | 0
neuromuscular blockade | 0
intravenous sedatives stopped | 48
neuromuscular blockers stopped | 48
generalised status myoclonus | 48
isoflurane stopped | 96
comatose | 96
absent motor response to painful stimulus | 96
preserved pupillary reflexes | 96
preserved corneal reflexes | 96
preserved cough reflexes | 96
preserved gag reflexes | 96
spontaneously breathing | 96
severe generalised status myoclonus | 96
refractory to three antiepileptic medications | 96
electroencephalography showed generalised periodic discharges | 96
no discernable background rhythm | 96
reversible causes of coma eliminated | 96
plasma neuron-specific enolase | 240
NSE 51 mcg/L | 240
somatosensory-evoked potential | 240
unhelpful due to myoclonus motion artefacts | 240
brain magnetic resonance imaging | 240
bilateral basal ganglia and frontoparietal cortex infarction | 240
severe hypoxic encephalopathy | 240
medical consensus regarding poor prognosis | 240
extubated | 240
died | 264