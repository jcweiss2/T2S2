newborn female | 0
born at 24 weeks + 3 days | 0
breech presentation | 0
cord prolapse | 0
birth weight of 645 g | 0
HIV negative mother | 0
Apgar score of 4 | 0
Apgar score of 8 | 5
mechanical ventilation | 0
central umbilical catheters | 0
total parenteral nutrition | 0
empiric antibiotics | 0
skin sensors | 0
late-onset sepsis | 216
Escherichia coli bacteremia | 216
antimicrobial therapy with cefepime | 216
adhesive patch removal | 480
skin abrasion | 480
erythema | 480
induration | 480
plaque with necrotic center | 480
ulcer | 528
subcutaneous cell tissue | 528
necrotic area | 528
intensive treatment | 528
wound care team | 528
healings | 528
hydrating dermal wound dressings | 528
sodium alginate | 528
carboxymethylcellulose | 528
hydrocolloids | 528
thermic instability | 528
metabolic acidosis | 528
hyperglycemia | 528
hypotension | 528
clinical deterioration | 528
cutaneous mucormicosis | 528
skin biopsy | 528
empiric antifungal treatment | 528
liposomal amphotericin B | 528
fungal biomarkers | 528
serum galactomannan | 528
1,3 beta-D-glucan | 528
refractory shock | 552
renal failure | 552
death | 564
fungal cultures | 528
Rhizopus spp. | 528
histopathology | 528
broad aseptate hyphae | 528
right angle branching | 528
Mucorales | 528
mass spectroscopy | 528
MALDI-TOF MS | 528
polymerase chain reaction | 528
PCR | 528
Rhizopus arrhizus | 528
fungal blood cultures | 528 
R. oryzae | 528 
necrotic eschar | 528 
skin abscesses | 528 
gangrenous form | 528 
superficial infection | 528 
vesicle | 528 
pustule | 528 
erythematous plaque | 528 
ulcerate | 528 
necrotizing cellulitis | 528 
necrotic plaque | 528 
distant tissues | 528 
infection control | 528 
surgical debridement | 528 
anti-fungal treatment | 528 
ischemic necrosis | 528 
leukocytes | 528 
anti-fungal agents | 528 
infection site | 528 
gastrointestinal tract | 528 
skin | 528 
lungs | 528 
rhinocerebral spaces | 528 
primary cutaneous mucormycosis | 528 
secondary cutaneous mucormycosis | 528 
disseminated infection | 528 
rhinocerebral mucormycosis | 528 
minor local skin trauma | 480 
vascular invasion | 528 
thrombosis | 528 
infarctions | 528 
necrotic surrounding tissue | 528 
autopsy | 564 
tissue biopsy | 528 
laboratory processing | 528 
routine culture media | 528 
broad hyaline | 528 
aseptate hyphae | 528 
vascular invasion | 528 
necrotic tissue | 528 
PCR assays | 528 
mass spectrometry tests | 528 
MALDI-TOF MS | 528 
faster diagnosis | 528 
accurate diagnosis | 528 
species level | 528 
traditional methods | 528 
microbiological | 528 
histopathological | 528 
necrotizing cellulitis | 528 
Mucorales | 528 
underlying disease | 528 
predisposing factors | 528 
disease severity | 528 
surgical debridement | 528 
anti-fungal treatment | 528 
L-AmB | 528 
another agent | 528 
ischemic necrosis | 528 
infected tissue | 528 
leukocytes | 528 
anti-fungal agents | 528 
efficacy | 528 
pediatric patients | 528 
mucormycosis | 528 
antifungal therapy | 528 
surgical debridement | 528 
lower risk | 528 
death | 564 
high suspicion | 0 
prompt recognition | 0 
aggressive approach | 0 
infection control | 0 
traditional diagnostic methods | 528 
microbiology | 528 
histopathology | 528 
modern tests | 528 
mass spectrometry | 528 
molecular studies | 528 
rapid diagnosis | 528 
accurate diagnosis | 528 
etiological diagnosis | 528 
extremely premature infant | 0 
necrotizing cellulitis | 528 
Mucorales | 528 
facility | 0 
informed consent | 0 
Institutional Ethics Committee | 0 
Clínica Universitaria Bolivariana | 0 
Universidad Pontificia Bolivariana | 0 
Álvaro Hoyos | 0 
María Adelaida Mejía | 0 
Verónica Herrera | 0 
Andrés Soto | 0 
Clara Rico | 0 
Alejandro Díaz-Díaz | 0 
critical review | 0 
conflicting interests | 0 
declaration | 0 
acknowledgements | 0