43 years old | 0
male | 0
admitted to the hospital | 0
shortness of breath | -336
non-productive cough | -720
subjective fevers | -720
chills | -720
weakness | -720
malaise | -720
azithromycin | -336
presumed diagnosis of pneumonia | -336
no past medical history of autoimmune | 0
no past medical history of systemic | 0
no past medical history of immune-compromising conditions | 0
no sick contacts | 0
no recent travel | 0
no tuberculosis | 0
no chemical exposure | 0
no nausea | 0
no vomiting | 0
no diarrhea | 0
no muscular weakness | 0
no neurological symptoms | 0
no orthopnea | 0
no paroxysmal nocturnal dyspnea | 0
able to walk approximately five blocks without getting dyspneic | 0
20 pack year smoking history | 0
no known drug allergies | 0
no other medications | 0
negative social history | 0
unremarkable family history | 0
desk job | 0
negative occupational history | 0
afebrile | 0
respiratory rate of 26 breaths/min | 0
heart rate of 115 beats/min | 0
room air saturation of 75% | 0
blood pressure of 90/60 mm Hg | 0
hyperkeratosis over the index fingers | 0
hyperkeratosis over the thumbs | 0
thickening over the metacarpophalangeal joints | 0
thickening over the proximal interphalangeal joints | 0
early resuscitation | 0
6 L of oxygen via nasal cannula | 0
30 cc/kg of normal saline | 0
normalization of blood pressure | 0
normalization of heart rate | 0
white blood cell count of 25,000 units/L | 0
hemoglobin level of 13.5 g/dL | 0
platelet count of 385 × 10^9/L | 0
sodium level of 133 mg/dL | 0
BUN of 13 mg/dL | 0
creatinine of 0.69 mg/dL | 0
troponin of 0.09 μg/L | 0
B-type natriuretic peptide of 79 pg/mL | 0
normal alkaline phosphatase | 0
normal bilirubin level | 0
aspartate transaminase of 259 units/L | 0
alanine transaminase of 266 units/L | 0
CPK of 7,500 International Units/L | 0
albumin of 2.4 g/dL | 0
globulin level of 4.2 g/dL | 0
arterial blood gas values of 7.37/43/52 | 0
lactic acid of 2.4 mg/dL | 0
ESR of 35 mm/h | 0
CRP of 24 mg/L | 0
procalcitonin level of 34 ng/mL | 0
ANA with speckled pattern and 1:320 titers | 0
anti-Jo-1 antibody positive | 0
anti-CCP antibody positive | 0
pericardial effusion | 0
non-confluent areas of ill-defined opacities | 0
denser consolidations | 0
air bronchograms | 0
infiltrates | 0
atelectasis | 0
small right-sided pleural effusion | 0
patchy right-sided opacity | 0
moderate to large pericardial effusion | 0
intensive care unit transfer | 48
worsening hypoxia | 48
worsening hypotension | 48
non-invasive positive pressure ventilation | 48
mechanical ventilation | 48
pulmonary artery catheterization | 48
optimal fluid management | 48
veno-venous ECMO | 96
severe acute respiratory distress syndrome | 96
broad spectrum antibiotics | 0
vancomycin | 0
zosyn | 0
azithromycin | 0
high dose methylprednisolone | 0
minimal vasopressor requirements | 0
worsening pericardial effusion | 0
diagnostic pericardial window | 0
therapeutic pericardial window | 0
non-oliguric renal failure | 0
acute tubular necrosis | 0
hypotension | 0
sepsis | 0
rhabdomyolysis | 0
upper gastrointestinal bleed | 0
erosive gastritis | 0
proton pump inhibitors | 0
improvement in respiratory status | 120
improvement in cardiovascular status | 120
improvement in renal status | 120
decannulation from ECMO | 120
transition to mechanical ventilation | 120
extubation | 120
discharged home | 240
physical therapy assistance | 240
wean off steroid | 240
taper regimen | 240
follow-up with rheumatology | 240