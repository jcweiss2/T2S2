40 years old| 0
    male | 0
    admitted to the hospital | 0
    hypertension | -8760
    atrial fibrillation | -8760
    severe uncontrolled hyperthyroidism | -8760
    thyroid storm | -8760
    medical intensive care unit admission | -8760
    intubation | -8760
    noncompliance with medications | -1416
    central chest pain | -2
    palpitation | -2
    agitation | -2
    nausea | -2
    blood pressure 181/112 mmHg | -2
    irregularly irregular pulse | -2
    heart rate 140 beats/min | -2
    tachypneic | -2
    respiratory rate 38/min | -2
    temperature 37.6°C | -2
    oxygen saturation 85% on room air | -2
    oxygen saturation 96% on 5 L oxygen | -2
    anxious | 0
    agitated | 0
    diffuse goiter | 0
    clammy skin | 0
    warm skin | 0
    bibasilar crackles | 0
    no lower limb edema | 0
    fast atrial fibrillation | 0
    ST-segment elevation V3-V6 | 0
    mild leukocytosis | 0
    normal hemoglobin | 0
    normal platelets | 0
    normal renal function tests | 0
    normal liver function tests | 0
    proBNP 1100 pg/mL | 0
    undetectable thyroid-stimulating hormone | 0
    serum thyroxin >100 pmol/L | 0
    Burch-Wartofsky score 60 | 0
    serum troponin T 1200 ng/L | 0
    acute anterior wall myocardial infarction | 0
    thyroid storm diagnosis | 0
    dual antiplatelet therapy started | 0
    aspirin | 0
    clopidogrel | 0
    unfractionated heparin infusion | 0
    propylthiouracil 200 mg every 4 hours | 0
    hydrocortisone 200 mg stat | 0
    hydrocortisone 100 mg every 8 hours | 0
    cholestyramine 4 mg every 6 hours | 0
    Lugol's solution 10 drops every 8 hours | 0
    isosorbide dinitrate infusion 25 mcg/min | 0
    intravenous furosemide 40 mg | 0
    chest pain progression | 2
    increased tachypnea | 2
    additional intravenous furosemide | 2
    isosorbide dinitrate infusion increased to 50 mcg/min | 2
    high-risk coronary angiography consent | 4
    anesthesia standby | 4
    femoral access procedure | 4
    diluted contrast solution 50:50 | 4
    15 ml contrast used | 4
    single vessel disease | 4
    distal LAD 100% embolic occlusion | 4
    TIMI 3 | 4
    blood flow restored | 4
    chest pain settled | 4
    ECG improvement | 4
    ejection fraction 35% | 4
    anterior wall hypokinesia | 4
    grade 2 diastolic dysfunction | 4
    moderately dilated left atrium | 4
    BP improved to 130/80 | 48
    heart rate 70%u201380 beats/min | 48
    respiratory rate <20/min | 48
    oxygen saturation >96% | 48
    bisoprolol started | 48
    intravenous furosemide switched to oral | 48
    ECG atrial fibrillation controlled | 168
    T wave inversion anterior leads | 168
    T4 improved to 67 pmol/L | 168
    hydrocortisone tapered | 168
    cholestyramine stopped | 168
    Lugol's solution stopped | 168
    PTU switched to carbimazole | 168
    discharge medications initiated | 168
    DAPT | 168
    rivaroxaban for 1 month | 168
    clopidogrel and rivaroxaban for 1 year | 168
    rosuvastatin 20 mg | 168
    furosemide 40 mg daily | 168
    bisoprolol 10 mg | 168
    spironolactone 25 mg | 168
    valsartan 160 mg | 168
    medication compliance | 168
    ECG atrial fibrillation controlled after 1 month | 744
    T4 dropped to 23 pmol/L | 1008
    ejection fraction improved to 49% | 2160
