65 years old | 0
male | 0
autoimmune hepatitis | 0
hypertension | 0
hyperlipidemia | 0
benign prostatic hypertrophy | 0
admitted to intensive care unit | 0
severe symptomatic hypotonic hyponatremia | -720
diffuse large B-cell lymphoma of the liver | -720
furosemide | 0
allopurinol | 0
prazosin | 0
folic acid | 0
ursodiol | 0
pantoprazole | 0
prednisolone | 0
transferred to oncology service | 24
cyclophosphamide | 24
rituximab | 24
dexamethasone | 24
tumor lysis syndrome | 72
renal failure | 72
hemodialysis | 72
volume overload | 72
respiratory failure | 72
intubation | 72
mechanical ventilation | 72
extubated | 168
transferred back to oncology service | 168
chest CT on hospital day 18 | 432
PEA arrest | 432
central airway obstruction | 432
blood clots | 432
emergent intubation | 432
return of spontaneous circulation | 432
cachectic | 432
temperature 38.2°C | 432
pulse 72/min | 432
blood pressure 107/61 mmHg | 432
respiratory rate 21 | 432
oxygen saturation 97% | 432
FiO2 50% | 432
pupils equally round and reactive | 432
nonresponsive to verbal or physical stimuli | 432
dried blood in oropharynx | 432
bloody secretions from endotracheal tube | 432
significant anasarca | 432
unremarkable cardiovascular exam | 432
unremarkable pulmonary exam | 432
unremarkable abdominal exam | 432
WBC 3.8 103/uL | 432
hemoglobin 9.5 g/dL | 432
BUN 56 mg/dL | 432
creatinine 1.69 mg/dL | 432
CT abdomen and pelvis | 408
thick-walled cavitary lesion in left lower lobe | 408
non-contrast chest CT | 432
air fluid level in cavitary lesion | 432
bronchoscopy | 576
blood clots admixed with thick mucus | 576
CT pulmonary angiography | 576
1.9 × 1.5 cm saccular contrast-enhancing lesion | 576
bronchoalveolar lavage consistent with Mucor | 576
pulmonary artery pseudoaneurysm | 576
pulmonary mucormycosis | 576
isavuconazonium | 576
embolization of PAP | 576
no further hemoptysis | 576
irreversible anoxic brain injury | 576
renal failure worsened | 576
family elected to forgo hemodialysis | 576
forgo cardiopulmonary resuscitation | 576
passed away | 864
