near-drowning incident | -1
bystander CPR | -1
abdominal pain | 0
diffuse abrasions on torso | 0
pneumoperitoneum | 0
pneumomediastinum | 0
intraabdominal free fluid | 0
hollow viscus perforation | 0
laparotomy | 1
gross contamination with food debris | 1
total gastroesophageal junction disruption | 1
hemodynamically labile | 1
damage control procedure | 1
distal esophagus stapled closed | 1
proximal stomach stapled closed | 1
mediastinal drain placed | 1
gastrostomy tube placed | 1
nasogastric tube placed | 1
septic shock | 24
respiratory failure | 24
prolonged intubation | 24
deep venous thrombosis | 24
pulmonary embolism | 24
bilateral pleural effusions | 24
general deconditioning | 24
parenteral nutrition started | 24
extubated | 432
leak in esophagus | 432
enteral nutrition initiated | 432
discharged | 1200
Ivor-Lewis distal esophagectomy | 2160
gastric pull-up | 2160
esophagogastric anastomosis | 2160
extubated | 2163
jejunostomy tube placed | 2163
esophagram showed no leak | 2170
initiated on liquid diet | 2170
discharged | 2170
tolerate regular diet | 2600
gaining weight | 2600 
recovering well | 2600