88 years old | 0
female | 0
admitted to the hospital | 0
right hip pain | -432
fell while walking | -432
transferred to our hospital | -18
history of hypertension | 0
history of dementia | 0
intertrochanteric fracture | -96
COVID-19 | -96
sepsis | -18
ischemic colitis | -18
urinary tract infection | -18
hypotension | -18
transferred to ICU | -18
transferred to isolation ward | -19
blood pressure dropped | -19
hip pain | -18
conservative observation | -432
visited another hospital | -96
planned surgical treatment | -96
diagnosed with COVID-19 | -96
postponed surgery | -96
treated for sepsis | -18
treated for ischemic colitis | -18
transferred to our hospital for surgery | -18
preoperative laboratory findings | 0
hemoglobin | 0
platelet | 0
serum albumin | 0
C-reactive protein | 0
sodium | 0
arterial blood gas analysis | 0
prothrombin time | 0
international normalized ratio | 0
activated partial thromboplastin Time | 0
D-dimer | 0
chest computed tomography | 0
diffuse PTE | 0
consolidation in the right lower lobe | 0
ground glass opacity | 0
pleural effusion | 0
rib fractures | 0
abdominopelvic CT scan | 0
deep vein thrombus | 0
transthoracic echocardiography | 0
ejection fraction | 0
aortic stenosis | 0
mitral regurgitation | 0
echogenic material in the left atrium | 0
electrocardiography | 0
cardiology consultation | 0
heparinization | 0
insertion of IVC filter | 0
admitted to the operating room | 0
preoperative vital signs | 0
induction of anesthesia | 0
tracheal intubation | 0
maintenance of anesthesia | 0
intraoperative monitoring | 0
intraoperative transesophageal echocardiography | 0
mean arterial pressure | 0
fluid administration | 0
bleeding | 0
urine output | 0
anesthetic time | 0
operating time | 0
reversal of anesthesia | 0
tracheal extubation | 0
transferred to ICU | 0
postoperative day 2 | 48
removal of ECMO sheaths | 48
transferred to general ward | 48
postoperative day 8 | 192
removal of IVC filter | 192
discharged | 192