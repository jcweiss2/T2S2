59 years old | 0
male | 0
admitted to the hospital | 0
ascending aortic aneurysm | -720
atrial fibrillation | -720
congestive heart failure | -720
bilateral lower extremity venous stasis ulcers | -720
stage 3 chronic kidney disease | -720
multinodular goiter | -720
ground-level fall | -1
felt heart racing | -1
denies dyspnea | -1
denies chest pain | -1
denies loss of consciousness | -1
deterioration of health | -720
unable to properly care for bilateral lower extremity wounds | -720
cleaning wounds with water and washcloth | -720
septic shock | 0
blood pressure 84/53 mm Hg | 0
heart rate 124 beats per minute | 0
lactate 3 mg/dL | 0
3 lower extremity ulcers | 0
necrotic skin and subcutaneous tissue | 0
maggots | 0
C-reactive protein 6.97 mg/L | 0
creatinine 3.54 mg/dL | 0
elevated troponin 0.06 ng/mL | 0
elevated white blood cell count 14.8 × 103 cells per mL | 0
electrocardiogram showed atrial fibrillation | 0
chest X-ray showed enlarged heart | 0
X-ray imaging showed bilateral areas of subcutaneous gas formation | 0
admitted to ICU | 0
sepsis bundle initiated | 0
fluid resuscitation | 0
vasopressor support with norepinephrine | 0
blood cultures obtained | 0
broad-spectrum antibiotics started | 0
vancomycin started | 0
piperacillin/tazobactam started | 0
acute coronary syndrome protocol initiated | 0
amiodarone started | 0
debridement of bilateral lower extremity necrotic skin and soft tissue | 24
gram negative rods and gram positive cocci grew in blood cultures | 24
S fonticola and MSSA identified | 48
S fonticola resistant to amoxicillin/clavulanate | 48
vancomycin discontinued | 96
piperacillin/tazobactam de-escalated to ceftriaxone | 96
cardiac echocardiogram showed dilation of all cardiac chambers | 120
left ventricular systolic function severely depressed | 120
transesophageal echocardiogram showed severe left ventricular systolic dysfunction | 168
mitral valve vegetation | 168
mobile echo density consistent with thrombus | 168
cardiac catheterization showed severe 2 vessel coronary artery disease | 168
ceftriaxone changed to cefepime | 168
discharged to skilled nursing facility | 240
completed 6 weeks of antibiotic therapy | 1008
uneventful recovery | 1008