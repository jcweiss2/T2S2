30 years old | 0
    housewife | 0
    presented to hospital emergency | 0
    ingestion of 15 g of KMnO4 powder | -15
    suicidal attempt | -15
    no other drugs ingested | -15
    arrived at hospital within 15 minutes | -15
    drowsy | 0
    hypoxia | 0
    stridor | 0
    oxygen saturation 85% | 0
    ABG pH 7.32 | 0
    pO2 52.1 | 0
    pCO2 46 | 0
    HCO3 22 | 0
    SpO2 86.1% | 0
    tachycardia | 0
    heart rate 116/min | 0
    blood pressure 110/70 mmHg | 0
    temperature 98.2°F | 0
    multiple patches of blackish-brown stain on face and hands | 0
    shifted to medical ICU | 0
    oral cavity examination: brownish black staining | 0
    copious secretions | 0
    vocal cords swollen | 0
    almost complete airway obstruction | 0
    planned percutaneous tracheostomy | 0
    attempted intubation | 0
    difficult intubation | 0
    stained and edematous pharyngeal structures | 0
    stained and edematous laryngeal structures | 0
    sloughed debris in posterior pharynx | 0
    placed 6.5 mm endotracheal tube | 0
    fiber optic bronchoscopic guidance | 0
    intermittent positive pressure ventilation | 0
    invasive ventilatory support | 0
    broad-spectrum antibiotics | 0
    steroids | 0
    proton-pump inhibitor | 0
    intravenous fluids | 0
    improved oxygenation | 24
    ABG pH 7.37 | 24
    pO2 113 | 24
    pCO2 33.9 | 24
    HCO3 19.2 | 24
    SpO2 98.1% | 24
    improved sensorium | 24
    upper GI endoscopy on day 1 | 24
    diffuse ulceration in esophagus | 24
    necrotic areas in esophagus | 24
    diffuse ulceration in fundus of stomach | 24
    necrotic areas in fundus of stomach | 24
    bronchoscopy | 24
    edematous and inflamed mucosa in tracheo-bronchial tree | 24
    hemorrhagic patches in tracheo-bronchial tree | 24
    normal renal parameters | 0
    normal hepatic parameters | 0
    normal electrolytes | 0
    normal complete hemogram | 0
    normal methemoglobin level | 0
    deranged liver function tests on day 2 | 48
    rising serum bilirubin | 48
    total serum bilirubin 4.5 mg/dl | 72
    serum glutamic pyruvic transaminase 354 IU | 72
    deranged coagulation profile | 72
    INR 2.06 | 72
    decreased platelet counts 80,000/cumm | 72
    clinical picture of acute hepatic necrosis | 72
    improved coagulation profile on day 4 | 96
    elevated serum transaminase levels | 96
    reduced oral cavity staining | 96
    reduced upper airway edema | 96
    reduced vocal cord swelling | 96
    extubation attempted | 96
    cuff leak check | 96
    copious oral secretions post-extubation | 96
    difficulty swallowing | 96
    difficulty breathing | 96
    reintubation | 96
    percutaneous tracheostomy | 96
    weaned off ventilator next day | 120
    shifted to ward | 120
    tracheostomy tube in situ | 120
    total parenteral nutrition started on day 5 | 120
    started clear liquids on day 8 | 192
    improved liver functions | 192
    improved coagulation profile | 192
    decannulated on day 9 | 216
    discharged | 216
    follow-up after 3 months normal | 216
    no psychiatric illness in the past | -672
    happily married | -672
    no pyloric stenosis | 216
    no esophageal strictures | 216
    no kidney involvement | 216
    no pancreas involvement | 216
    no cardiovascular depression | 216
    no heart block | 216
    no hypotension | 216
    no shock | 216
    no cardiac arrest | 216
    no GI hemorrhage | 216
    no methemoglobinemia | 216
    no disseminated intravascular coagulation | 216
    no acute respiratory distress syndrome | 216
    no pancreatitis | 216
    no subcortical hemorrhages | 216
    no papillary hemorrhages | 216
    no lung consolidation | 216
    no severe fatty liver changes | 216
    no peritonitis | 216
    no perforation | 216
    no difficulty intubation initially | 0
    no failed intubation | 0
    no requirement for emergency tracheostomy initially | 0
    no requirement for crico-thyroidotomy | 0
    no nebulized epinephrine | 0
    no inhalational induction with sevoflurane | 0
    no gastric lavage | 0
    no activated charcoal | 0
    no methylene blue | 0
    no vitamin C | 0
    no argon plasma coagulation | 0
    no parenteral nutrition delay | 0