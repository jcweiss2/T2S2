65 years old | 0
male | 0
admitted to emergency room | 0
fever | 0
chills | 0
loss of consciousness | 0
no response to physical stimulation | 0
muscle strength of right limb grade 0 | 0
muscle strength of left limb grade 2 | 0
Babinski’s sign positive on the right lower limb | 0
leukocyte count of 17.5×10^9/L | 0
neutrophil count of 16.28×10^9/L | 0
C-reactive protein count of 84.29 mg/L | 0
blood cultures grew Streptococcus viridans | 0
no abnormalities in electrocardiogram | 0
no abnormalities in myocardial infarction markers | 0
catheter ablation | -336
refractory AF | -336
computed tomography scan of the brain | 0
large area of left craniocerebral infarction | 0
air emboli in the right lobe | 0
chest CT | 0
air between the left atrium and esophagus | 0
pericardial effusions | 0
diagnosed with AEF | 0
diagnosed with sepsis | 0
diagnosed with cerebral infarction | 0
urgent surgical operation | 0
intraoperative gastroscopy | 0
esophageal fistula | 0
fresh blood | 0
standard posterolateral thoracotomy | 0
dense adhesions between the lower esophagus and the pericardium | 0
necrotic tissues dropped | 0
massive bleeding | 0
1 cm-diameter defect in the posterior wall of the left atrium | 0
4-0 Prolene suture | 0
autologous pericardial tissue | 0
closure of the bleeding point and fistula | 0
3-incision esophagectomy | 0
simultaneous anastomosis | 0
intensive care unit monitoring | 0
anti-infection administration | 0
nutritional support | 0
anticoagulation | 0
supportive treatments | 0
died of sepsis and multiple organ failure | 576
esophagectomy | 0
simultaneous reconstruction | 0 
atrial-esophageal fistula | -336