44 years old | 0
female | 0
obese | 0
admitted to the hospital | 0
inhalation injury | 0
burn injury | 0
second-to-third degree burn injury | 0
32% total body surface area burn | 0
intubated with endotracheal tube | 0
ETT no 6.5 | 0
depth of placement 22 cm | 0
fixed with thread on the right lip corner | 0
spontaneous breathing | 0
symmetrical breathing | 0
respiratory rate 20x/minute | 0
SpO2 100% | 0
T-piece 10 lpm | 0
blood pressure 128/79 mmHg | 0
heart rate 98x/minute | 0
warm extremities | 0
capillary refill time <2 seconds | 0
no spontaneous bleeding | 0
head and neck edema | 0
burn injury on the mucous membranes of the lips, mouth, and eyes | 0
full of edema | 0
nasogastric tube insertion | 0
brownish fluid obtained | 0
high value of leucocytes 28880 103/µl | 0
rise in blood glucose value to 242 mg/dL | 0
low albumin value of 2.5 gr/dL | 0
sputum obtained from the tracheal secretions | 0
Acinetobacter baumanii bacteria | 0
treated with tigecycline | 0
grade II-III burn injury | 0
stress ulcer | 0
leucocytosis | 0
percutaneous dilatational tracheostomy | 18
early tracheostomy | 18
PDT performed | 18
ventilator set to PSV/CPAP | 18
PS 10 Peep 5 trig 3 FiO2 50% | 18
intubated successfully | 18
treated in the ICU | 18
tangential excision | 24
debridement | 24
25% plasbumin transfusion | 24
100 ml for 2 days | 24
discharged from the ICU | 168
moved to a normal ward | 168
still canulated | 168
able to breathe spontaneously | 168
discharged from the hospital | 336
referred back to the first hospital | 336
no follow-up for Pseudomonas infection at the PDT site | 336