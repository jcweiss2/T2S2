19 years old | 0
    male | 0
    ALL | 0
    Philadelphia positive | 0
    fever | 0
    anemia | 0
    thrombocytopenia | 0
    hypercalcemia | 0
    normal white cell count | 0
    intravenous fluids | 0
    clodronate | 0
    prednisolone | 0
    vincristine | 0
    idarubicin | 0
    Lasparaginase | 0
    intrathecal methotrexate | 0
    fever | 240
    diarrhea | 240
    E.coli | 240
    Klebsiella pneumoniae | 240
    ceftazidime | 240
    amikacin | 240
    responded well to treatment | 240
    clinically stable | 240
    small painful nodule over left thigh | 504
    Pseudomonas aeruginosa | 504
    ciprofloxacin | 504
    imipenem | 504
    MRSA | 504
    nasal swab | 504
    E.coli | 504
    urine sample | 504
    change ceftazidime to imipenem | 504
    change amikacin to ciprofloxacin | 504
    vancomycin | 504
    continuously febrile | 504
    central venous catheter removed | 504
    induction chemotherapy on hold | 504
    G-CSF initiated | 504
    pyrexial | 504
    thigh nodule developed into cellulitis | 504
    fluid collection | 504
    surgical incision and drainage | 504
    continued deterioration | 504
    cellulitis extending toward perineum | 504
    febrile | 504
    hypotensive | 504
    transferred to ICU | 504
    hemodynamically unstable | 720
    ventilatory support | 720
    inotropic support | 720
    central blood cultures | 720
    peripheral blood cultures | 720
    A. xylosoxidans | 720
    gram negative bacillus | 720
    oxidase and nitrate positive | 720
    negative reaction for urea | 720
    negative reaction for mannitol | 720
    negative reaction for sucrose | 720
    negative reaction for maltose | 720
    sensitive to colistin | 720
    sensitive to imipenem | 720
    sensitive to ceftazidime | 720
    sensitive to piperacillin/tazobactam | 720
    intravenous colistin | 720
    removal of central venous catheter | 720
    further deterioration | 720
    cardiac arrest | 720
    death | 720
    septic shock | 720
    multiorgan failure | 720
    