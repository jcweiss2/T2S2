25 years old | 0
male | 0
congenital macrocephaly | 0
hydrocephalus | 0
presented to the emergency department | 0
behavioral changes | -72
insomnia | -72
language impairment | -72
head CT scan | 0
discharged | 0
benzodiazepine | 0
antipsychotic drug | 0
returned the same day | 0
worsening symptoms | 0
decreased level of consciousness | 0
high fever | 0
non-collaborative | 0
eyes closed | 0
miotic pupils | 0
no conjugated eye deviation | 0
dysarthria | 0
low production of speech | 0
no focal signs of neurological dysfunction | 0
auricular temperature 39.9 ºC | 0
blood pressure 103/54 mmHg | 0
HR 127 bpm | 0
blood gas analysis | 0
blood workup | 0
mild leukocytosis | 0
neutrophilia | 0
slight lymphopenia | 0
normal C-reactive protein | 0
normal procalcitonin | 0
lumbar puncture | 0
ceftriaxone | 0
ampicillin | 0
acyclovir | 0
CSF total proteins 66.5 mg/dl | 0
CSF 38 cells/mm3 | 0
no mononuclear cell predominance | 0
viral encephalitis | 0
focal onset impaired awareness seizures | 24
levetiracetam | 24
sodium valproate | 24
acyclovir treatment | 0
CSF PCR panel negative | 120
autoimmune encephalitis suspected | 120
lumbar puncture repeated | 120
antibody testing | 120
methylprednisolone | 120
EEG bi@hemispherical cerebral activity disorganization | 120
EEG polymorphic continuous bilateral theta@delta activity | 120
brain MRI no signal changes | 120
Anti-NMDAR antibodies confirmed | 120
anti-NMDAR encephalitis diagnosis | 120
ICU admission | 144
respiratory distress | 144
decreased level of consciousness | 144
fluctuating heart rate | 144
low arterial blood pressure | 144
vasopressors | 144
severe bradycardia | 144
pauses up to 5 seconds | 144
severe dystonia | 144
dyskinesia | 144
sialorrhea | 144
IVIg | 480
rituximab | 480
infectious complications | 720
discharge to rehabilitation facility | 2160
decreased level of consciousness at discharge | 2160
no verbal response | 2160
no collaboration | 2160
bilateral stereotypical movements | 2160
oro@mandibular dyskinesia | 2160
memory lapses | 2160
25 years old|0
male|0
congenital macrocephaly|0
hydrocephalus|0
presented to the emergency department|0
behavioral changes|-72
insomnia|-72
language impairment|-72
head CT scan|0
discharged|0
benzodiazepine|0
antipsychotic drug|0
returned the same day|0
worsening symptoms|0
decreased level of consciousness|0
high fever|0
non-collaborative|0
eyes closed|0
miotic pupils|0
no conjugated eye deviation|0
dysarthria|0
low production of speech|0
no focal signs of neurological dysfunction|0
auricular temperature 39.9 ºC|0
blood pressure 103/54 mmHg|0
HR 127 bpm|0
blood gas analysis|0
blood workup|0
mild leukocytosis|0
neutrophilia|0
slight lymphopenia|0
normal C-reactive protein|0
normal procalcitonin|0
lumbar puncture|0
ceftriaxone|0
ampicillin|0
acyclovir|0
CSF total proteins 66.5 mg/dl|0
CSF 38 cells/mm3|0
no mononuclear cell predominance|0
viral encephalitis|0
focal onset impaired awareness seizures|24
levetiracetam|24
sodium valproate|24
acyclovir treatment|0
CSF PCR panel negative|120
autoimmune encephalitis suspected|120
lumbar puncture repeated|120
antibody testing|120
methylprednisolone|120
EEG bi-hemispherical cerebral activity disorganization|120
EEG polymorphic continuous bilateral theta-delta activity|120
brain MRI no signal changes|120
Anti-NMDAR antibodies confirmed|120
anti-NMDAR encephalitis diagnosis|120
ICU admission|144
respiratory distress|144
decreased level of consciousness|144
fluctuating heart rate|144
low arterial blood pressure|144
vasopressors|144
severe bradycardia|144
pauses up to 5 seconds|144
severe dystonia|144
dyskinesia|144
sialorrhea|144
IVIg|480
rituximab|480
infectious complications|720
discharge to rehabilitation facility|2160
decreased level of consciousness at discharge|2160
no verbal response|2160
no collaboration|2160
bilateral stereotypical movements|2160
oro-mandibular dyskinesia|2160
memory lapses|2160
