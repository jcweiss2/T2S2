44 years old | 0
male | 0
hepatitis B | -672
primary hepatocellular carcinoma | 0
chronic viral hepatitis B | -672
no cirrhosis | -672
multiphasic contrast-enhanced Magnetic Resonance Imaging (MRI) | 0
mass in the right hepatic lobe | 0
small lesions | 0
arterial hypervascularity | 0
Alpha-fetoprotein (AFP) greater than 3,630 ng/mL | 0
Barcelona Clinic Liver Cancer (BCLC) stage B | 0
transarterial chemoembolization | 0
first TACE | 0
30 mg THP loaded by 100–300 µm drug micro-ball | 0
8 mL iodized oil | 0
350 µm gelfoam sponge particles | 0
fever | 24
severe liver damage | 24
white blood cell (WBC) 8.5×10^9/L | 24
neutrophil granulocyte (GRAN) 91.4% | 24
alanine aminotransferase (ALT) 2.6 upper limit of normal value (ULN) | 24
aspartate aminotransferase (AST) 7.9 ULN | 24
total bilirubin (TBIL) 1.9 ULN | 24
treatment for liver preservation | 24
other treatments | 24
ALT returned to normal range | 720
AST returned to normal range | 720
TBIL returned to normal range | 720
WBC 9.2×10^9/L | 720
GRAN 82.7% | 720
abdominal enhancement MRI showed significant necrosis of the lesions | 720
AFP dropped to 1,708 ng/mL | 720
repeated fever | 912
cough | 912
anti-infection treatment | 912
body temperature reached a maximum of 39 °C | 912
Chest computed tomography (CT) showed pneumonia | 912
pneumorachis with iodine oil deposition | 912
hepatic abscess | 912
anti-infection treatment (Tazobactam Sodium/Piperacillin Sodium for Injectio) | 912
pigtail catheter drainage | 912
bacteria culture was negative | 912
significant reduction in the original lesion | 1092
new lesions in the liver increased | 1092
AFP rose to more than 3,630 ng/mL | 1092
second TACE | 1344
60 mg THP plus 20 mL iodized oil | 1344
third TACE | 1560
60 mg THP plus 8 mL iodized oil | 1560
fourth TACE | 1776
60 mg THP plus 7mL iodized oil | 1776
fifth TACE | 1992
60 mg THP plus 4 mL iodized oil plus 350 µm gelatin sponge particles | 1992
fever began | 1996
WBC 14.1×10^9/L | 1996
GRAN 98.5% | 1996
ALT 163 U/L | 1996
AST 249 U/L | 1996
TBIL 73 µmol/L | 1996
anti-infection and liver protection treatment | 1996
fainted | 2008
difficulty breathing | 2008
enhancing CT showed a large amount of gas in the lesions and in the portal veins | 2008
hepatic portal venous gas (HPVG) | 2008
bacteria cultured showed that Streptococcus anginosus from hepatic puncture tube drainage was positive | 2008
died | 2010