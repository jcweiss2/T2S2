49 years old | 0
female | 0
presented to the hospital | 0
fatigue | -72
dizziness | -72
intermittent fever | -72
minor scratch on her left foot | -72
trauma at her left foot | -168
computed tomography (CT) | 0
large vegetation at the aortic valve cusp | 0
pericardial effusion | 0
antibiotic therapy | 0
referred to the department of cardiology | 0
referred to the center for emergency surgery | 0
standard sternotomy | 0
pericardium opened | 0
hemorrhagic pericardial effusion | 0
cardiopulmonary bypass (CPB) | 0
aortotomy | 0
large vegetation identified | 0
septic perforations of the aortic wall | 0
Prolene 4–0 sutures | 0
aortic valve replaced | 0
SJM mechanical valve | 0
uneventful weaning of CPB | 0
chest closed | 0
transferred to the intensive care unit (ICU) | 0
large quantities of blood in the thoracic drainage | 1
hemodynamic unstable | 1
reoperation initiated | 1
resuscitation | 1
sternum reopened | 1
CPB | 1
rupture of the left ventricular lateral wall | 1
Dor plasty not feasible | 1
myocardial phlegmon excised | 1
histopathological examination | 1
myocardial infarction | 1
multiple bacteria in coronary capillary vessels | 1
bacterial imbibition of myocardial tissue | 1
Dacron patch | 1
myocardial reconstruction | 1
venous bypass graft | 1
BioGlue | 1
cardiac activity reestablished | 1
no bleeding | 1
extracorporeal life support (ECLS) | 1
CPB weaned | 1
chest closure | 1
abscess at the left foot lanced | 72
antibiotics administered | 0
Staphylococcus aureus infection | 0
clindamycin and flucloxacillin | 0
echocardiography | 120
left ventricular ejection fraction | 120
mild pericardial effusion | 120
pseudoaneurysm detected | 8760
reoperation | 8760
aneurysm resection | 8760
rehabilitation | 9072
patient recovered | 9072