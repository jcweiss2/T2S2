60 years old | 0 | 0 
male | 0 | 0 
admitted to the hospital | 0 | 0 
biopsy proven PAN | -8760 | 0 
paroxysmal atrial fibrillation | -8760 | 0 
hypertension | -8760 | 0 
dyslipidemia | -8760 | 0 
non-insulin dependent diabetes mellitus | -8760 | 0 
prior admissions for PAN flares | -8760 | 0 
admission for septic shock | -17520 | -17520 
scrotal pain | 0 | 0 
fever of 103°F | 0 | 0 
fatigue | 0 | 0 
tachycardic to 130 beats per minute | 0 | 0 
hypotensive to 103/40 mm Hg | 0 | 0 
broad-spectrum antibiotics | 0 | 24 
vancomycin | 0 | 24 
Zosyn | 0 | 24 
kidney function worsened | 24 | 48 
switch in antibiotics to meropenem | 48 | 48 
creatinine level continued to rise | 48 | 72 
fevers without a specific source of an infection | 48 | 168 
no focus was found on the CT chest, abdomen, and pelvis | 72 | 72 
stopping all antibiotics | 72 | 72 
macular rash | 168 | 168 
rash progressed slowly to involve his axillary area | 168 | 192 
rash progressed to involve his chest, head, neck, and abdomen | 192 | 216 
decline of his mental status | 192 | 216 
worsening of skin lesions | 216 | 216 
element of bullae and vesicles | 216 | 216 
dermatology team was involved | 216 | 216 
biopsy was obtained | 216 | 216 
initiating local steroid cream | 216 | 216 
rash became pustular | 264 | 264 
high grade fever of 109°F | 264 | 264 
transfer to the intensive care unit | 264 | 264 
pulse steroids | 264 | 312 
fever subsided | 312 | 312 
improvement of the initial rash | 312 | 312 
decreased progression of sloughing | 312 | 312 
complete resolution of acute kidney injury | 312 | 312 
taper in steroids | 312 | 336 
skin biopsy | 216 | 216 
urine analysis | 0 | 0 
CT chest/abdomen/pelvis | 72 | 72 
CBC/BMP/coagulation | 0 | 0 
DRESS | 0 | 0 
GPP | 0 | 0 
PAN typical rash | 0 | 0 
Steven Johnson syndrome | 0 | 0 
leukocytoclastic vasculitis | 0 | 0 
subcorneal pustular dermatosis | 0 | 0 
cutaneous candidiasis | 0 | 0 
AGEP | 168 | 312 
intra- and subcorneal spongiform | 216 | 216 
superficial, interstitial, mid-dermal infiltrate rich in neutrophils | 216 | 216 
dermal edema | 216 | 216 
tender erythematous nodules | 0 | 0 
purpura | 0 | 0 
livedo reticularis | 0 | 0 
ulcers | 0 | 0 
bullous or vesicular eruption | 0 | 0 
systemic corticosteroids | 264 | 312 
withdrawal of the offending drug | 72 | 72 
supportive care | 0 | 336 
symptomatic treatment of pruritus and skin inflammation | 216 | 336 
immunosuppressive management | 336 | 336 
discharged | 336 | 336