26 years old | 0
female | 0
primigravida | 0
ulcerative colitis | -672
abdominal pain | -504
fever | -504
bloody diarrhoea | -504
generalised weakness | -504
mesalazine | -504
6-mercaptopurine | -504
prednisolone | -504
analgesia | -504
intravenous fluids | -504
intravenous steroids | -504
discharged | -312
readmitted | 0
systemic signs of sepsis | 0
tachycardia | 0
hypotension | 0
pyrexia | 0
distended abdomen | 0
exquisitely tender on palpation | 0
positive rebound tenderness | 0
peritonitis | 0
severe colonic distension | 0
emergent caesarean section | 0
infra-umbilical midline incision | 0
fetus delivered | 0
apgar scores 9 at one minute | 0
apgar scores 9 at five minutes | 0
weight 1.474 kg | 0
height 36.2 cm | 0
total abdominal colectomy | 0
end ileostomy | 0
total operative time 96 min | 0
estimated blood loss 250 ml | 0
discharged | 216
ventilator support | 0
weaned off ventilator | 168
transitioned to neonatal progressive care unit | 168
discharged home | 336
pathologic examination | 0
toxic megacolon | 0
transmural inflammation | 0
erosion of the bowel wall | 0
completion proctectomy | 672
ileal reservoir | 672
ileoanal anastomosis | 672
diverting ileostomy | 672
operative time 177 min | 672
estimated blood loss 200 ml | 672
loop ileostomy reversed | 1200
2-3 bowel movements a day | 1200
constitutionally well | 1200
optimal healing of surgical wounds | 1200
reduced fertility | 1200
ileal pouch-anal anastomosis | 1200
neonate measured between 40 and 50th centile | 1200
satisfactory recovery | 1200