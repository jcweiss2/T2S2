46 years old | 0
female | 0
obesity | -7200
psoriatic arthritis | -7200
hypoparathyroidism | -7200
hypothyroidism | -7200
total thyroidectomy | -7200
multinodular goitre | -7200
elective sleeve gastrectomy | 0
gastric perforations | 0
friable mucosa | 0
abdominal sepsis | 4
transfer to intensive care | 4
critically low calcium level | 4
ionised calcium 0.78 mmol/L | 4
continuous intravenous calcium gluconate infusion | 4
normocalcaemia | 4
prolonged ICU admission | 4
abdominal operations | 4
weight loss 14 kg | 192
endocrinology advice | 336
hypothyroidism management | 336
TSH 5.83 mU/L | 336
intravenous triiodothyronine | 336
euthyroidism | 672
high dose intravenous calcium | 672
ionised calcium measured daily | 672
serum phosphate level 1.07 | 672
intravenous calcitriol | 1008
intravenous calcitriol ceased | 1013
intramuscular cholecalciferol | 1344
low 1,25(OH)vitamin D3 level | 1344
renal function normal | 1344
eGFR > 90 mL/min/1.73 m2 | 1344
intravenous calcitriol recommenced | 2016
reduced calcium gluconate requirements | 2016
intramuscular thyroxine | 2016
intravenous thyroxine | 2020
maintenance schedule established | 2020
discharge | 5760
normocalcaemia on review | 6048
weight 71.8 kg | 6048
BMI 29 kg/m2 | 6048