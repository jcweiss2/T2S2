42 years old | 0
male | 0
generalized weakness | -2160
fever | -2160
cough | -2160
weight loss | -2160
HIV-antibody test positive | -2160
sputum AFB smear positive | -2160
isoniazid | -40
rifampin | -40
ethambutol | -40
pyrazinamide | -40
fluconazole | -40
trimethoprim/sulfamethoxazole | -40
HIV-1 Western blot test positive | -40
CD4 cell count 10/µL | -40
HIV RNA titer 18,000 copies/mL | -40
oral thrush | 0
hepatosplenomegaly | 0
ascites | 0
hemoglobin 10.6g/dL | 0
white blood cell 2,700/µL | 0
platelet 58,000/µL | 0
total bilirubin 2.4mg/dL | 0
AST/ALT 131/48IU/L | 0
ALP 114IU/L | 0
GGT133 IU/L | 0
costophrenic angle blunting | 0
fluid shifting in the right hemithorax | 0
mild pneumonic infiltration in left lung | 0
anti-retroviral agents | 0
zidovudine | 0
lamivudine | 0
efavirenz | 0
hemoglobin 7.4g/dL | 3
white blood cell 1,070/µL | 3
platelet 13,000/µL | 3
rifampin discontinued | 3
zidovudine discontinued | 3
trimethoprim/sulfamethoxazole discontinued | 3
new pulmonary infiltrates | 5
septic shock | 5
piperacillin/tazobactam | 5
mechanical ventilator support | 6
Gram stain negative | 6
ordinary culture negative | 6
bone marrow aspiration | 9
bone marrow biopsy | 9
Histoplasma capsulatum | 9
death | 10