65 years old | 0
female | 0
end-stage osteoarthritis of the right knee | 0
joint pain | 0
hypertension | 0
gastroesophageal reflux disease | 0
history of DVT | -672
right total knee arthroplasty | 0
enoxaparin | 24
vague epigastric pain | 192
lethargy | 192
febrile episodes | 192
decreased appetite | 192
somnolence | 192
anxiety | 192
nausea | 192
temperature 101.7 F | 192
heart rate 111 | 192
respiration 20 | 192
blood pressure 123/87 | 192
oxygen saturation 92% | 192
hyponatremia | 192
hypokalemia | 192
glucose 60 | 192
hematocrit 25.3 | 192
creatinine 0.8 | 192
WBC count 14,900 | 192
platelet count 161,000 | 192
pulmonary embolism | 192
sepsis | 192
metabolic encephalopathy | 192
adrenal insufficiency | 192
chest CT scan | 192
MRI of the brain | 192
empirical intravenous antibiotics | 192
ceftriaxone | 192
vancomycin | 192
acyclovir | 192
CSF cultures | 192
urine cultures | 192
blood cultures | 192
aggressive intravenous volume support | 192
pressors | 192
basal cortisol levels | 192
cosyntropin stimulation | 192
abdominal CT | 192
bilateral adrenal hemorrhages | 192
enoxaparin discontinued | 192
high dose hydrocortisone | 192
glucocorticoid tapered | 192
discharged | 240
follow-up | 8760
excellent range of motion | 8760
X-rays demonstrate well-placed components | 8760
no evidence of loosening | 8760
returned to previous activity level | 8760
bowling | 8760