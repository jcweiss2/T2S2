18 years old|0
male|0
admitted to the hospital|0
unrestrained driver in a rollover motor vehicle accident|-unknown
prolonged extrication|-unknown
positive blood alcohol screen|-unknown
intubated at the scene|-unknown
taken to a Level-1 trauma center|-unknown
open book pelvic fracture|0
complete disruption of the posterior sacroiliac complex|0
vertical and rotational instability of the left hemipelvis|0
pubic symphysis diastasis|0
left greater than right sacroiliac joint disruption|0
left open comminuted femoral shaft fracture|0
left distal tibia shaft fracture|0
systolic blood pressure in the 80s|0
tachycardic|0
positive focused assessment with sonography for trauma scan in pelvic windows|0
pelvis bound with a sheet|0
secured using hemostats|0
pulses detected with Doppler ultrasound in bilateral lower extremities|0
poor response to initial fluid bolus|0
sustained tachycardia|0
taken to the angiography suite|0
significant slowing of flow within the left superior gluteal artery|0
significant slowing of flow within the left internal pudendal artery|0
radiographic blush|0
thought due to vasospasm|0
thought due to distal arterial injury|0
empiric Gelfoam embolization of the left internal iliac artery|0
hypotension stabilized|0
tachycardia stabilized|0
hemodynamic instability began to respond appropriately to resuscitation|0
pelvic fractures temporarily stabilized post-embolization through an external fixator|0
left femoral shaft fracture stabilized on PID 0|0
definitive fixation of the pelvis|48
definitive fixation of both sacroiliac joints through sacroiliac screws|48
left tibia intramedullary nailing|48
definitive fixation of the left femur through intramedullary nailing|96
remained intubated post-operatively until PID 6|144
transferred out of the Intensive Care Unit on PID 8|192
wounds followed throughout hospital course|0
incisions remained clean and dry throughout hospital stay|0
intermittently febrile throughout admission|0
increasing lymphocyte count on routine daily collection|0
computed tomography (CT) of the pelvis on PID 10|240
evidence of 15cm diameter simple-appearing fluid collection|240
scant gas collection lateral to the left hip|240
near area of surgical fixation|240
considered appropriate post-operative changes|240
no clinical evidence of infection on PID 10|240
elevated white blood cell count of 22.9|240
white blood cell count trending upward from 14.4 on PID 8|240
managed with observation|240
general surgery trauma team advised by orthopedics|240
cause of leukocytosis likely not related to fluid collection|240
progressed as expected over next few days|0
first evidence of minimal serous drainage from left hip/buttock wound|360
scant amount of drainage noted|360
minimal soiling of sheets|360
no foul smell|360
no evidence of purulence|360
no fluid could be expressed from the wound|360
managed expectantly with local wound care|360
wound without erythema|360
wound without induration|360
discharged to rehabilitation center|360
continued drainage from left buttock area|360
developed early signs of wound margin epidermolysis|360
readmitted to the hospital|528
evidence of increasing drainage|528
marginal erythema|528
induration|528
epidermolysis adjacent to the wound edge|528
clinical evidence of early sepsis|528
started on intravenous vancomycin|528
underwent local debridement of left hip/buttock wound|528
evidence of cavitation extending posterior to the greater trochanter|528
significant fat necrosis|528
epidermolysis|528
monitored closely|528
scheduled for repeat debridement|528
repeat CT scan noted questionable intramuscular abscess formation|528
ill-defined collection of fluid and gas in left gluteal musculature|528
aggressive repeat surgical debridement of left hip|576
massive gluteal muscle necrosis identified|576
wound cultures from left hip obtained on PID 22|528
tissue cultures from left hip obtained on PID 24|576
positive for Proteus mirabilis|528
positive for Serratiamarcescens|528
positive for Klebsiella pneumoniae|528
third surgical debridement of left hip wound|600
drain placed|600
continued on vancomycin for 8 days|0
piperacillin/tazobactam added for 10 days|0
wound noted on PID29 to have no erythema|696
wound noted on PID29 to have no drainage|696
significant decrease in swelling|696
continued induration of the abductor compartment|696
progressed with physical therapy|0
recovered as anticipated from traumatic injuries|0
significant gluteal fold asymmetry on left side|2928
necrosis|2928
atrophy|2928
significant gains in strength of left hip and buttock area|2928
continued to ambulate with Trendelenburg gait|2928
orthopedic fractures healed|2928
unable to return to competitive football|2928
sustained weakness of left hip and buttock area|2928
