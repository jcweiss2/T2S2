45 years old | 0
    male | 0
    presented to Accident and Emergency Department | 0
    fever | -48
    chills | -48
    productive cough | -48
    runny nose | -48
    gradual onset headache | -48
    temperature of 39.8°C | 0
    heart rate of 115 bpm | 0
    blood pressure of 130/70 mmHg | 0
    respiratory rate of 18/min | 0
    throat was injected | 0
    unremarkable ear examination | 0
    unremarkable oral cavity examination | 0
    slightly raised WBC count (15.45 × 10^9/L) | 0
    normal chest radiograph | 0
    symptomatic treatment for presumed upper respiratory tract infection | 0
    discharged from A and E | 0
    eight episodes of witnessed seizures | 6
    febrile | 6
    status epilepticus | 6
    heart rate of 173 bpm | 6
    blood pressure of 94/57 mmHg | 6
    normal cardiac auscultation | 6
    confused | 6
    impaired consciousness | 6
    preserved reflexes | 6
    equal and reactive pupils | 6
    no papilledema | 6
    WBC count increased to 31 × 10^9/L | 6
    predominant neutrophils (84%) | 6
    CRP levels elevated (245.6 ml/L) | 6
    intubated | 6
    urgent noncontrast CT of the brain | 6
    subtle fullness in right frontal region | 6
    mild sulcal effacement | 6
    diffuse mucosal thickening in paranasal sinuses | 6
    lumbar puncture performed | 6
    CSF leukocytosis | 6
    increased CSF protein levels | 6
    GCS dropped from 10 to 7 | 6
    contrast-enhanced MRI of the brain | 8
    large right frontotemporoparietal subdural collection | 8
    smaller left frontal subdural collections | 8
    severe mass effect in right cerebral hemisphere | 8
    midline shift | 8
    fluid-filled paranasal sinuses with mucosal hyperenhancement | 8
    small bony defect in posterior wall of left frontal sinus | 8
    adjacent meningeal enhancement | 8
    right frontal parenchymal edema | 8
    diagnosis of sinogenic meningoencephalitis | 8
    diagnosis of multiple subdural empyemas | 8
    retrospective confirmation of bone defect on initial CT | 8
    intravenous vancomycin | 8
    intravenous ceftriaxone | 8
    right decompressive craniectomy | 8
    evacuation of subdural empyema | 8
    FESS to address sinusitis | 8
    Streptococcus intermedius in pus | 8
    intravenous meropenem | 8
    intravenous vancomycin for 2 weeks | 8
    intensive care unit stay for 5 days | 8
    GCS improved to 10 | 8
    vital signs normalized | 8
    extubated on fourth postoperative day | 12
    follow-up CT showing improved mass effect | 12
    follow-up CT showing improved cerebral edema | 12
    discharged after 20 days | 480
    CRP 51.4 mg/L at discharge | 480
    no change in personality | 480
    no change in cognitive functions | 480
    no motor deficits | 480
    no sensory deficits | 480
    developed scar epilepsy | 480
    follow-up CTs showing parenchymal loss | 480
    follow-up CTs showing gliosis | 480
    oral sodium valproate | 480
    oral levetiracetam | 480

    