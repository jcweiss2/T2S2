42 years old | 0
female | 0
Caucasian | 0
admitted to the hospital | 0
diagnosed with acetylcholine receptor antibody positive oculo-bulbar myasthenia gravis | -2160
drooping eyelids | -2160
double vision | -2160
difficulty swallowing | -2160
diurnal variation | -2160
characteristic fluctuation of symptoms | -2160
failed bedside swallow evaluation | -2160
notable aspiration to thin liquids on modified barium swallow | -2160
underwent plasmapheresis | -2160
complete resolution of symptoms | -2160
IVIG | -2160
repetitive nerve stimulation study | -2160
antibody titers confirmed the diagnosis of postsynaptic neuromuscular junction disorder | -2160
started on pyridostigmine | -2160
prednisone | -2160
mycophenolate | -2160
generalized anxiety disorder | -2160
allergic rhinitis | -2160
recurrence of drooping eyelids | -672
change in voice | -672
concerns of impending myasthenia exacerbation | -672
started on regular plasma exchange | -672
CT chest showed 6.7 cm lobulated soft tissue mass in anterior mediastinum | -672
referred to cardiothoracic surgery for possible thymectomy | -672
fever | -120
chills | -120
cough | -120
minimal clear sputum production | -120
exertional shortness of breath | -120
decreased sense of taste | -120
decreased sense of smell | -120
decreased appetite | -120
traveled to nearby city | -168
chest x-ray showed patchy infiltrates in left lower lobe | -120
elevated white count | -120
lymphopenia | -120
respiratory pathogen panel came back negative | -120
tested for COVID-19 RT-PCR | -120
COVID-19 RT-PCR came back positive | -120
bedside negative inspiratory force obtained was 65 cm H2O | -120
discharged from emergency department | -120
self-quarantine for next fourteen days | -120
follow CDC guidelines | -120
immunomodulatory therapy continued | -120
plasmapheresis deferred | -120
recovered from COVID-19 infection | 168
no complications | 168
no myasthenic crisis | 168
no myasthenia exacerbation | 168
no changes to immunosuppressive medications | 168