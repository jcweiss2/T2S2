47 years old | 0
    male | 0
    kidney transplant | -61368
    diarrhea | -336
    nausea | -336
    vomiting | -336
    acute kidney injury | -336
    nausea | -336
    vomiting | -336
    diarrhea | -336
    inability to drink or eat | -336
    nausea | 0
    abdominal discomfort | 0
    vomiting | 0
    no shortness of breath | 0
    no cough | 0
    no fever | 0
    no chills | 0
    type two diabetes | 0
    hypertension | 0
    hyperlipidemia | 0
    endocarditis | 0
    coronary artery disease | 0
    heart failure with reduced ejection fraction | 0
    coronary artery bypass surgery | -78840
    mitral valve replacement | -78840
    tacrolimus | 0
    mycophenolic acid | 0
    no known allergies to medications | 0
    past tobacco smoker | 0
    alcohol rarely drank | 0
    no illicit drug use | 0
    family history of hypertension | 0
    family history of heart disease | 0
    family history of throat cancer | 0
    temperature 36.6°C | 0
    blood pressure 90/58 mmHg | 0
    heart rate 103 beats per minute | 0
    respiratory rate 16 breaths per minute | 0
    oxygen saturation 98% | 0
    BMI 42.2 | 0
    normal heart sounds | 0
    clear lung sounds | 0
    creatinine 6.7 mg/dL | 0
    potassium 5.7 mMol/L | 0
    blood urea nitrogen 175 mg/dL | 0
    bicarbonate 14 mMol/L | 0
    white-cell count 2.9 K/CUMM | 0
    lymphocytes 0.2 K/CUMM | 0
    INR 2.75 | 0
    chest radiograph prominent pulmonary vascular markings | 0
    chest radiograph enlarged cardiac silhouette | 0
    no pulmonary infiltrates | 0
    SARS-CoV-2 RNA positive | 0
    hypotension resolved after 1L normal saline | 0
    insulin | 0
    beta-agonists | 0
    calcium | 0
    polystyrene sulfonates | 0
    admitted to the hospital | 0
    vital signs stable | 72
    oxygen saturation 96% | 72
    diarrhea resolved | 72
    nausea resolved | 72
    vomiting resolved | 72
    tolerate soft diet | 72
    unresolved acute kidney injury | 72
    hyperkalemia | 72
    metabolic acidosis | 72
    leukopenia | 72
    mild thrombocytopenia | 72
    oliguria | 0
    renal ultrasonography normal | 72
    urinary sediment no cellular casts | 72
    intravenous fluid | 0
    5L normal saline administered | 0
    immunosuppressive therapy discontinued | 0
    warfarin 5 mg | 0
    warfarin 2 mg | 24
    INR continued to rise | 0
    productive cough | 96
    shortness of breath | 96
    oxygen saturation 85% | 96
    oxygen saturation 95% with nasal cannula | 96
    filgrastim 480 mcg administered | 96
    shortness of breath progressed | 102
    oxygen saturation decreased | 102
    HFNC 40 L/min | 102
    transferred to ICU | 102
    blood culture | 102
    sputum culture | 102
    chest radiograph multifocal air-space opacities | 102
    furosemide | 102
    vancomycin | 102
    cefepime | 102
    intubation | 120
    mechanical ventilation | 120
    blood pressure 75/46 mmHg | 120
    norepinephrine | 120
    vasopressin | 120
    worsening kidney function | 120
    anuria | 120
    CRRT initiated | 120
    white blood cell count increased to 35 K/CUMM | 120
    increased C-reactive protein | 120
    increased ferritin | 120
    increased lactate dehydrogenase | 120
    increased creatine phosphokinase | 120
    worsening bilateral opacities | 120
    echocardiography LVEF 20% | 120
    prosthetic mitral valve normal | 120
    mechanical ventilation continued | 120
    oxygen saturation decreased | 120
    atrial fibrillation | 120
    amiodarone | 120
    hypotension worsened | 120
    CRRT held | 120
    death | 216
    
    
    47 years old | 0
    male | 0
    kidney transplant | -61368
    diarrhea | -336
    nausea | -336
    vomiting | -336
    acute kidney injury | -336
    nausea | -336
    vomiting | -336
    diarrhea | -336
    inability to drink or eat | -336
    nausea | 0
    abdominal discomfort | 0
    vomiting | 0
    no shortness of breath | 0
    no cough | 0
    no fever | 0
    no chills | 0
    type two diabetes | 0
    hypertension |4 0
    hyperlipidemia | 0
    endocarditis | 0
    coronary artery disease | 0
    heart failure with reduced ejection fraction | 0
    coronary artery bypass surgery | -78840
    mitral valve replacement | -78840
    tacrolimus | 0
    mycophenolic acid | 0
    no known allergies to medications | 0
    past tobacco smoker | 0
    alcohol rarely drank | 0
    no illicit drug use | 0
    family history of hypertension | 0
    family history of heart disease | 0
    family history of throat cancer | 0
    temperature 36.6°C | 0
    blood pressure 90/58 mmHg | 0
    heart rate 103 beats per minute | 0
    respiratory rate 16 breaths per minute | 0
    oxygen saturation 98% | 0
    BMI 42.2 | 0
    normal heart sounds | 0
    clear lung sounds | 0
    creatinine 6.7 mg/dL | 0
    potassium 5.7 mMol/L | 0
    blood urea nitrogen 175 mg/dL | 0
    bicarbonate 14 mMol/L | 0
    white-cell count 2.9 K/CUMM | 0
    lymphocytes 0.2 K/CUMM | 0
    INR 2.75 | 0
    chest radiograph prominent pulmonary vascular markings | 0
    chest radiograph enlarged cardiac silhouette | 0
    no pulmonary infiltrates | 0
    SARS-CoV-2 RNA positive | 0
    hypotension resolved after 1L normal saline | 0
    insulin | 0
    beta-agonists | 0
    calcium | 0
    polystyrene sulfonates | 0
    admitted to the hospital | 0
    vital signs stable | 72
    oxygen saturation 96% | 72
    diarrhea resolved | 72
    nausea resolved | 72
    vomiting resolved | 72
    tolerate soft diet | 72
    unresolved acute kidney injury | 72
    hyperkalemia | 72
    metabolic acidosis | 72
    leukopenia | 72
    mild thrombocytopenia | 72
    oliguria | 0
    renal ultrasonography normal | 72
    urinary sediment no cellular casts | 72
    intravenous fluid | 0
    5L normal saline administered | 0
    immunosuppressive therapy discontinued | 0
    warfarin 5 mg | 0
    warfarin 2 mg | 24
    INR continued to rise | 0
    productive cough | 96
    shortness of breath | 96
    oxygen saturation 85% | 96
    oxygen saturation 95% with nasal cannula | 96
    filgrastim 480 mcg administered | 96
    shortness of breath progressed | 102
    oxygen saturation decreased | 102
    HFNC 40 L/min | 102
    transferred to ICU | 102
    blood culture | 102
    sputum culture | 102
    chest radiograph multifocal air-space opacities | 102
    furosemide | 102
    vancomycin | 102
    cefepime | 102
    intubation | 120
    mechanical ventilation | 120
    blood pressure 75/46 mmHg | 120
    norepinephrine | 120
    vasopressin | 120
    worsening kidney function | 120
    anuria | 120
    CRRT initiated | 120
    white blood cell count increased to 35 K/CUMM | 120
    increased C-reactive protein | 120
    increased ferritin | 120
    increased lactate dehydrogenase | 120
    increased creatine phosphokinase | 120
    worsening bilateral opacities | 120
    echocardiography LVEF 20% | 120
    prosthetic mitral valve normal | 120
    mechanical ventilation continued | 120
    oxygen saturation decreased | 120
    atrial fibrillation | 120
    amiodarone | 120
    hypotension worsened | 120
    CRRT held | 120
    death | 216