60 years old | 0
    male | 0
    anxiety disorder | 0
    presented to a community hospital | 0
    four-day history of increasing fatigue | -96
    increasing fatigue | -96
    weakness | -96
    cough | -96
    shortness of breath | -96
    sharp right-sided pleuritic chest pain | -96
    right upper quadrant abdominal pain | -96
    deep breathing | -96
    denied nausea | -96
    denied vomiting | -96
    review of systems was otherwise negative | -96
    heavy smoker | 0
    occasional alcohol consumption | 0
    denied intravenous recreational drugs use | 0
    febrile | 0
    oral temperature of 39.2°C | 0
    hemodynamically stable | 0
    edentulous | 0
    decreased air entry in right lower and middle lobes | 0
    bronchial breath sounds at right lung base | 0
    crepitations over rest of right lung | 0
    abdomen tender in right upper quadrant | 0
    elevated total leukocyte count (17.8×10^9 cells/L) | 0
    neutrophil predominance (16.12×10^9 cells/L) | 0
    blood cultures (aerobic and anaerobic) negative | 0
    chest radiography right-sided pneumothorax | 0
    right lower lobe consolidation | 0
    pleural fluid | 0
    noncontrast CT scan of abdomen | 0
    right-sided hydropneumothorax | 0
    areas of pulmonary consolidation | 0
    loculated pleural fluid | 0
    admitted to hospital | 0
    chest tube placed | 0
    empirical antimicrobial therapy with levofloxacin | 0
    empirical antimicrobial therapy with metronidazole | 0
    pleural fluid sample submitted | 0
    no polymorphonuclear cells on Gram stain | 0
    no bacteria observed on Gram stain | 0
    aerobic culture no bacterial growth after 72h | 72
    Gram-positive spore-forming bacillus recovered on anaerobic culture after 48h | 48
    identified as Clostridium bifermentans | 48
    antimicrobial susceptibility testing performed | 48
    susceptible to amoxicillin-clavulanate | 48
    susceptible to cefoxitin | 48
    susceptible to clindamycin | 48
    susceptible to meropenem | 48
    susceptible to metronidazole | 48
    susceptible to penicillin | 48
    significant dyspnea | 72
    chest pain | 72
    CT scan of chest with contrast | 72
    right main pulmonary artery embolus | 72
    clinically deteriorated | 72
    admission to intensive care unit | 72
    antimicrobial therapy changed to piperacillin-tazobactam | 72
    antimicrobial therapy changed to levofloxacin | 72
    heparin initiated | 72
    thoracotomy | 360
    decortication of right lung | 360
    empyema fluid obtained | 360
    C bifermentans recovered again | 360
    postoperative antimicrobial therapy with piperacillin-tazobactam | 360
    intermittent low-grade fevers (~38°C) | 360
    ongoing hypoxia requiring 2L oxygen | 360
    repeat chest radiography loculated right-sided pneumothorax | 360
    small amount of fluid in empyema cavity | 360
    second thoracotomy | 1056
    right rib resection | 1056
    empyema drainage | 1056
    lung tissue obtained | 1056
    aerobic culture sterile | 1056
    anaerobic culture sterile | 1056
    antimicrobial therapy changed to ceftriaxone | 1056
    antimicrobial therapy changed to metronidazole | 1056
    echocardiogram performed | 1056
    no evidence of endocarditis | 1056
    no valvular pathology | 1056
    gradually improved | 1056
    discharged home | 1824
    prescription for oral metronidazole | 1824
    additional 10 days of therapy as outpatient | 1824
    arbitrary treatment duration of six weeks | 1824
    chest radiography right-sided pneumothorax | 0
    right lower lobe consolidation | 0
    pleural fluid | 0
    CT scan demonstrated pulmonary embolus | 72
    pneumothorax with empyema | 0
    no intra-abdominal abnormality | 0
    negative blood cultures | 0
    Gram-positive bacillus identified | 48
    patient required ICU admission | 72
    postoperative fevers | 360
    postoperative hypoxia | 360
    repeat surgery | 1056
    sterile cultures after second surgery | 1056
    echocardiogram negative for endocarditis | 1056
    oral metronidazole prescribed at discharge | 1824
    