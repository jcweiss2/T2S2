19 years old | 0
male | 0
admitted to the hospital | 0
severe pain in the nuchal area | -48
mild occipital headache | -48
mild sore throat | -72
fever | -48
chills | -48
nuchal rigidity | 0
opposition to passive anteflexion and rotation of the head | 0
mild redness and enlargement of tonsils | 0
limited straight leg raise maneuver | 0
leucocytosis | 0
neutrophilia | 0
elevated C-reactive protein | 0
elevated procalcitonin | 0
CT examination of the head | 0
chest radiogram | 0
lumbar puncture | 12
cerebrospinal fluid examination | 12
borderline pleocytosis | 12
normal proteinorhachia | 12
empiric antimicrobial therapy | 0
ceftriaxone | 0
vancomycin | 0
parenteral rehydration | 0
analgesic therapy | 0
headache disappeared | 24
pain in the nuchal area worsened | 24
erythema and tenderness of the skin | 24
generalised urticarial allergic exanthema | 24
antimicrobial therapy changed | 24
piperacillin–tazobactam | 24
clindamycin | 24
erythema and edema of the left lateral part of the neck | 48
palpable mass in the left lateral part of the neck | 48
CT of the neck | 48
collection of liquid | 48
thrombosis of the left internal jugular vein | 48
hypodense collection of fluid | 48
magnetic resonance imagining of the cervical spinal column | 48
epidural effusion | 48
cultivation of the oropharyngeal swab | 48
blood cultures | 48
Klebsiella pneumoniae | 48
antimicrobial therapy changed | 120
ceftriaxone | 120
clindamycin | 120
decline of C-reactive protein | 120
decline of procalcitonin | 120
pain in the neck area improved | 120
local erythema of the skin improved | 120
surgical revision and drainage of the abscess | 168
cultivation of pus | 168
Klebsiella pneumoniae | 168
antimicrobial therapy continued | 168
postsurgical course unremarkable | 192
patient transferred back to the intensive care unit | 192
patient afebrile | 192
minor pain near the surgical wound | 192
no pain in the cervical area | 192
no limitations of movement in the neck | 192
C-reactive protein level | 192
clindamycin stopped | 192
piperacillin–tazobactam continued | 192
follow-up CT scan | 240
complete regression of the cervical abscess | 240
partial recanalization of the left internal jugular vein | 240
complete regression of the epidural effusion | 240
C-reactive protein level | 240
antimicrobial regime changed | 240
moxifloxacin | 240
patient discharged | 360
asymptomatic | 432
CRP below 5 mg/L | 432
moxifloxacin treatment discontinued | 432