92 years old | 0
    woman | 0
    presented to the emergency department | 0
    fever | -48
    myalgia | -48
    anorexia | -48
    general weakness | -48
    hypertension | 0
    lived in a rural region | 0
    frequently in contact with grass | 0
    frequently in contact with domestic animals | 0
    alert | 0
    insect bite on left shoulder | 0
    blood pressure 94/54 mmHg | 0
    pulse rate 85 beats per minute | 0
    temperature 37.5°C | 0
    respiratory rate 20 breaths per minute | 0
    oxygen saturation 95% on room air | 0
    leukopenia | 0
    thrombocytopenia | 0
    white blood cell count 1,300 cells/μL | 0
    platelet count 100 × 10³/μL | 0
    elevated aspartate aminotransferase 88 IU/L | 0
    elevated alanine aminotransferase 40 IU/L | 0
    ceftriaxone administration | 0
    SFTSV detected | 24
    SFTSV viral load 186,606 copies/mL | 24
    conservative treatment | 24
    stable until day 4 | 24
    sudden-onset pneumonia | 120
    chest X-ray confirmed pneumonia | 120
    respiratory failure | 120
    high-resolution CT subtle bronchiolitis in upper lobes | 120
    high-resolution CT bronchial wall thickening in lower lobes | 120
    cefepime administration | 120
    vancomycin administration | 120
    voriconazole loading dose 6 mg/kg | 120
    voriconazole maintenance dose 4 mg/kg | 120
    serum Aspergillus galactomannan antigen level 6.1 | 120
    mechanical ventilation started | 144
    intensive care unit admission | 144
    bronchoalveolar fluid gram stain | 144
    bronchoalveolar fluid culture | 144
    fungus culture | 144
    septic shock | 144
    multifocal consolidations on chest X-ray | 144
    intravenous immunoglobulin administration | 168
    serum Aspergillus galactomannan antigen level 3.7 | 168
    serum Aspergillus galactomannan antigen level 1.6 | 216
    died | 264
    respiratory failure | 264
    refractory hypotension | 264
    metabolic acidosis | 264
    leukopenia persisted | 0
    thrombocytopenia persisted | 0
    CD4+ lymphocyte count remained low | 0
    neutropenia | 0
    bilateral lung infiltration | 120
    no corticosteroid administration | 0
    no other pathogens identified | 264
    low CD4 T+-cell count | 0
    high SFTSV viral load | 24
    no follow-up chest CT scan | 264
    no post-mortem examination | 264
    