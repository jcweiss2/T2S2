41 years old | 0 | 0 
female | 0 | 0 
admitted to the hospital | 0 | 0 
history of untreated hypertension | 0 | 0 
morbid obesity | 0 | 0 
chronic back pain | 0 | 0 
IVDU | 0 | 0 
low back pain | -336 | 0 
diffuse abdominal pain | -336 | 0 
lower extremity weakness | -336 | 0 
anorexia | -336 | 0 
fever | -336 | 0 
chills | -336 | 0 
shortness of breath | -336 | 0 
dizziness | -336 | 0 
constipation | -336 | 0 
acetaminophen use | -336 | 0 
gabapentin use | -336 | 0 
hydrocodone use | -336 | 0 
methamphetamines use | -336 | 0 
marijuana use | -336 | 0 
blood pressure of 79/53 mmHg | 0 | 0 
heart rate of 149 bpm | 0 | 0 
lactic acid of 4.2 mg dl-1 | 0 | 0 
WBC 37 500 u l-1 | 0 | 0 
erythrocyte sedimentation rate 75 mm h-1 | 0 | 0 
urine toxicology positive for cannabis | 0 | 0 
urine toxicology positive for amphetamines | 0 | 0 
midline tenderness of the lumbar spine | 0 | 0 
3/5 strength in bilateral lower extremities | 0 | 0 
bilateral shoulder warmth | 0 | 0 
bilateral shoulder erythema | 0 | 0 
bilateral shoulder tenderness | 0 | 0 
limited range of motion | 0 | 0 
multiple needle puncture sites | 0 | 0 
puncture wounds on the right foot | 0 | 0 
blood cultures collected | 0 | 0 
vancomycin started | 0 | 0 
metronidazole started | 0 | 0 
aztreonam started | 0 | 0 
IV fluids started | 0 | 0 
MRSA in blood cultures | 24 | 24 
sensitivities to vancomycin | 24 | 24 
sensitivities to rifampin | 24 | 24 
sensitivities to levofloxacin | 24 | 24 
sensitivities to clindamycin | 24 | 24 
sensitivities to daptomycin | 24 | 24 
sensitivities to linezolid | 24 | 24 
bilateral shoulder plain radiographs | 24 | 24 
arthrocentesis of the AC joints | 24 | 24 
WBC of 93 137 u l-1 in one shoulder | 24 | 24 
WBC of 32 043 u l-1 in the other shoulder | 24 | 24 
MRSA in aspirates | 24 | 24 
emergent surgical debridement of the shoulders | 48 | 48 
intubation | 48 | 48 
MRI of the lumbar spine | 48 | 48 
L3-L5 osteomyelitis | 48 | 48 
facet septic arthritis | 48 | 48 
dorsal paraspinous myositis | 48 | 48 
L2-L5 epidural abscess | 48 | 48 
bilateral psoas myositis | 48 | 48 
bilateral psoas abscesses | 48 | 48 
MRI of the bilateral shoulders | 48 | 48 
septic arthritis of the AC joints | 48 | 48 
right distal trapezius abscess | 48 | 48 
left supraclavicular abscess | 48 | 48 
MRI of the brain | 48 | 48 
TTE | 48 | 48 
no valvular vegetations | 48 | 48 
repeat surgical debridement of the shoulders | 120 | 120 
neurosurgery evaluation | 120 | 120 
leukocytosis | 120 | 168 
peak WBC of 52 100 u l-1 | 168 | 168 
trough levels of vancomycin monitored | 120 | 168 
repeat blood cultures positive for MRSA | 120 | 168 
antibiotics escalated to daptomycin | 240 | 240 
antibiotics escalated to ceftaroline | 240 | 240 
blood cultures became negative | 336 | 336 
rifampin added | 336 | 336 
repeat MRI of the lumbar spine | 336 | 336 
worsening epidural abscess | 336 | 336 
surgical drainage with drain placement | 432 | 432 
intraoperative wound cultures positive for MRSA | 432 | 432 
intraoperative wound cultures positive for Proteus mirabilis | 432 | 432 
drains removed | 672 | 672 
discharged | 672 | 672 
oral levofloxacin prescribed | 672 | 724 
oral rifampin prescribed | 672 | 724 
lost to follow-up | 724 | 724