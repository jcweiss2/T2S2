47 years old | 0
female | 0
admitted to the hospital | 0
headache | -48
blurred vision | -48
Glasgow coma scale (GCS) 15 | 0
afebrile | 0
no neurological alterations | 0
visual field intact | 0
body mass index (BMI) 28.2 | 0
mild psoriasis | 0
gastroesophageal reflux disease (GERD) | 0
cholelithiasis | 0
no relevant infections | 0
no previous surgeries | 0
no routine medications | 0
mother of two children | 0
regular menses | 0
blood pressure within normal limits | 0
heart rate within normal limits | 0
microcromic microcytic anemia | 0
reticulocytosis | 0
hemoglobin (Hb) 8.6g/dL | 0
hematocrit (HCT) 27.8% | 0
mean cell volume (MCV) 64.5 | 0
mean corpuscular hemoglobin (MCH) 20 pg | 0
mean corpuscular hemoglobin concentration (MCHC) 30.9 g/dL | 0
red blood cell distribution width (RDW) 20.2 % | 0
leucocytes count within normal limits | 0
inflammatory indexes within normal limits | 0
hormone blood concentrations normal | 0
thyroid-stimulating hormone (TSH) 0.238 μU/mL | 0
follicle-stimulating hormone (FSH) 0.6 mU/mL | 0
β-17-estradiol 35.8 pg/mL | 0
urine osmolality normal | 0
CT scan of the skull | -48
large mass arising from the sella | -48
eroding the bony structures | -48
invading the nasal cavity | -48
MRI confirmed solid-cystic lesion | 0
abutting both cavernous sinuses | 0
wrapping both carotid siphons | 0
diagnosed with pituitary adenoma | 0
scheduled for surgery | 0
headache treated with pain medications | 0
no vision problems | 0
sudden worsening of headache | 24
gaze palsy | 24
nuchal rigidity | 24
GCS fell to 6 | 24
emergency CT scan | 24
no parenchymal infarction | 24
no extra-axial bleeding | 24
no fluid collection | 24
no ischemia | 24
urgent craniotomy | 24
right frontotemporal approach | 24
brain swelling | 24
dense pus covering the brain surface | 24
purulent material within the tumor | 24
drained | 24
taken to intensive care unit (ICU) | 24
died a few days later | 72
pathological analysis confirmed nonfunctioning pituitary adenoma | 72
chronic inflammation | 72
necrosis | 72
cultures of intraoperative material negative | 72
spontaneous rupture of secondary pituitary abscess | 24
acute purulent meningoencephalitis | 24