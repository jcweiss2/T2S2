30 years old | 0
male | 0
gunshot injury to the chest | -936
two gunshot wounds | -936
damage control laparotomy | -936
right nephrectomy | -936
liver packing | -936
re-look laparotomies | -936
acute kidney injury | -936
haemodialysis | -936
bile leak | -936
endoscopic retrograde cholangiogram | -936
common bile duct stent | -936
sepsis | -936
pulmonary embolism | -936
anticoagulation with warfarin | -672
discharged | -672
colicky abdominal pain | -8
non-productive cough | -8
Grade III dyspnoea | -8
pyrexia | -8
International Normalized Ratio (INR) >10 | -8
bilateral pleural effusions | -8
blood products given | -8
empiric broad-spectrum antibiotics started | -8
warfarin stopped | -8
respiratory distress | 0
signs of cardiac tamponade | 0
X-ray showed bilateral pleural effusions and cardiomegaly | 0
emergency echocardiogram | 0
pericardial effusion | 0
2 cm defect/aneurysm in the lateral right ventricular wall | 0
surgical repair of the right ventricular aneurysm | 24
ventricular function was moderate | 24
ejection fraction 45% | 24
femoro-femoral bypass | 24
full sternotomy incision | 24
pericardial adhesions | 24
bypass perfusion time was 132 min | 24
aortic cross-clamp was applied | 24
heart arrested with antegrade cold blood cardioplegia | 24
cross-clamp time was 41 min | 24
significant bloody pericardial effusion | 24
RVA detected on the lateral wall | 24
bile collection in the sub-diaphragmatic area | 24
closed suction drain placed in the subdiaphragmatic position | 24
diaphragmatic defect closed | 24
RVA excised | 24
bovine pericardial patch used to close the defect | 24
sternal closure | 24
pericardial and mediastinal drain placement | 24
transferred to the intensive care unit | 24
post-operative stay in the intensive care unit | 48
post-operative stay in the general ward | 48
discharged home | 168
therapeutic anticoagulation | 168
follow-up ECHO scheduled | 168
histology revealed a true aneurysm | 168
fibrosis | 168
haemorrhage with organization | 168
haemosiderin deposition | 168
fibrin | 168
dystrophic calcification | 168
focal endarteritis obliterans | 168