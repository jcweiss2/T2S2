77 years old | 0 | 0 
female | 0 | 0 
breast cancer | -10080 | -10080 
chemotherapy | -10080 | -10080 
radiation to the chest | -10080 | -10080 
severe aortic stenosis | -10080 | 0 
coronary artery disease | -10080 | 0 
90% occlusion of the left anterior descending artery | -10080 | 0 
admitted to the hospital | 0 | 0 
tissue aortic valve replacement | 0 | 5 
saphenous vein graft bypass | 0 | 5 
left internal mammary artery dissected | 0 | 5 
induction of anesthesia | 0 | 0 
intubation | 0 | 2 
discontinuation of cardiopulmonary bypass | 5 | 5 
decline in cerebral head saturations | 5 | 5 
use of vasopressors | 5 | 24 
taken to the intensive care unit | 5 | 5 
extubated | 2 | 2 
persistent lactic acidosis | 5 | 48 
high-dose vasopressor support | 5 | 48 
mixed cardiogenic and vasoplegic shock | 5 | 48 
lethargic | 15 | 15 
leftward gaze | 15 | 15 
right upper extremity weakness | 15 | 15 
symptoms resolved | 15 | 15 
bilateral tongue ecchymoses | 15 | 15 
tongue numbness | 15 | 720 
dysgeusia | 15 | 720 
CT scan of her head | 15 | 15 
CT angiogram of her brain and neck | 15 | 15 
mild calcification at the bifurcation of the right common carotid artery | 15 | 15 
50% focal stenosis of the distal left common carotid artery | 15 | 15 
right lingual artery completely occluded | 15 | 15 
mild distal collateral flow | 15 | 15 
left lingual artery with multifocal irregularities | 15 | 15 
postoperative platelet count | 5 | 5 
prothrombin time (PT) | 5 | 5 
international normalized ratio (INR) | 5 | 5 
fibrinogen | 5 | 5 
ADAMTS13 inhibitor screen | 24 | 24 
volume resuscitation | 24 | 48 
low-dose epinephrine | 24 | 24 
high-dose norepinephrine | 24 | 48 
vasopressin | 24 | 48 
systemic vascular resistance improved | 48 | 48 
otolaryngology service consulted | 24 | 24 
serial examinations of the patient’s tongue | 24 | 720 
flexible bronchoscopes | 24 | 720 
persistent tongue numbness | 24 | 720 
dysgeusia | 24 | 720 
supportive therapy | 24 | 720 
tongue sensation and taste returned to baseline | 1440 | 1440 
discharged | 720 | 720