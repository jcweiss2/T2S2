64 years old | 0
male | 0
admitted with worsening skin lesions | 0
concerns for sepsis | 0
lesions suspicious for abscesses | 0
appeared rapidly over a few weeks | -672
diabetes | -672
not visited primary care physician’s office prior to presentation | -672
hemodynamically stable | 0
tachycardia to 130 beats per minute | 0
scattered pustules on scalp | 0
crusted papules on scalp | 0
atrophic cribriform plaques on thigh | 0
atrophic cribriform plaques on chest | 0
slit-like ulcerations with irregular borders in axilla bilaterally | 0
no tracts | 0
no subcutaneous nodulations | 0
axillary lymphadenopathy | 0
jagged red to purplish ulcerations on right third phalanx | 0
overhanging borders | 0
overlying peripheral erythema | 0
tenderness | 0
empirically treated with vancomycin | 0
empirically treated with piperacillin-tazobactam | 0
intravenous fluids | 0
leukocytosis of 15,000/μL | 0
neutrophilic predominance | 0
elevated inflammatory markers | 0
high sensitivity C-reactive protein (hsCRP) of 31.56 mg/L | 0
lactate dehydrogenase (LDH) of 546IU/mL | 0
mild transaminitis | 0
blood cultures with no growth | 0
normal electrolytes | 0
punch biopsy from border of ulcers on finger | 0
punch biopsy from scalp | 0
punch biopsy from upper thigh | 0
bacterial cultures showed no growth | 0
mycobacterial cultures showed no growth | 0
fungal cultures showed no growth | 0
viral cultures showed no growth | 0
biopsy from finger showed ulcerative dermatitis | 0
sub-adjacent neutrophilic infiltrate | 0
concerning for early stages of pyoderma gangrenosum | 0
discharged with close follow-ups | 24
prednisone taper | 24
clobetasol | 24
doxycycline | 24
satisfied Delphi consensus criteria for PG | 24
biopsy-proven neutrophilic infiltrate of the ulcer edge | 24
rapid progression of skin lesions | 24
peripheral erythema | 24
undermined borders | 24
tenderness at ulceration site | 24
multiple ulcerations | 24
cribriform scars at sites of healed ulcers | 24
biopsy results from thigh showed intraepidermal vesicular dermatitis | 24
biopsy results from scalp showed intraepidermal vesicular dermatitis | 24
atypical lymphoid infiltrate | 24
lymphocytes had atypia | 24
CD25 positivity | 24
immunostaining showed positivity for CD2 | 24
immunostaining showed positivity for CD3 | 24
immunostaining showed positivity for CD5 | 24
immunostaining showed positivity for CD25 | 24
immunostaining showed negative ALK1 | 24
immunostaining showed negative CD8 | 24
immunostaining showed negative CD20 | 24
immunostaining showed negative CD34 | 24
flow-cytometry | 24
HTLV1/2 levels | 24
suspicion of T-cell lymphoma | 24
negative autoimmune panel | 24
negative human immunodeficiency virus (HIV) | 24
negative rapid plasma reagin (RPR) | 24
negative hepatitis serologies | 24
negative Quantiferon assay | 24
urine protein electrophoresis showing polyclonal gammopathy | 24
no monoclonal band on fixation | 24
HTLV1/2 serology positive | 24
elevated interleukin-2 (IL2) receptor levels | 24
flow cytometry consistent with ATLL | 24
CD4+/CD25+/CD7- cells | 24
developed altered mental status | 48
severe hypercalcemia | 48
corrected calcium was 17.8 mg/dL | 48
unresponsive to aggressive hydration | 48
unresponsive to multiple doses of calcitonin | 48
upgraded to critical care | 48
hypercalcemia non-parathyroid hormone dependent | 48
given zoledronic acid | 48
eventual improvement | 48
developed hypoxic respiratory failure | 72
disseminated intravascular coagulopathy | 72
requiring emergent intubation | 72
PET/CT scan showed extensive organ-system lymphomatous involvement | 72
lymphomatous involvement in lungs | 72
lymphomatous involvement in spleen | 72
lymphomatous involvement in kidneys | 72
lymphomatous involvement in diaphragm | 72
lymphomatous involvement in scalp | 72
multi-level lymphadenopathy | 72
axillary/chest wall lymphadenopathy | 72
retroperitoneal lymphadenopathy | 72
pelvic lymphadenopathy | 72
cervical chains lymphadenopathy | 72
rapid decompensation | 72
goals of care discussed | 72
made full comfort care | 72
eventually passed away | 72
