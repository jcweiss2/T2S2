66 years old | 0
male | 0
admitted to the hospital | 0
fever | -240
cough | -240
sputum production | -240
progressive jaundice | -240
chronic alcoholic | 0
diabetes mellitus | 0
liver cirrhosis | 0
cerebral infarction | -3456
dysphagia | -240
plain chest X-ray | -72
bilateral lower lung field haziness | -72
abdominal CT scan | -72
27-mm liver mass | -72
aspiration pneumonia | -72
hepatocellular carcinoma | -72
intravenous antibiotics | -72
ceftriaxone | -72
azithromycin | -72
difficulty swallowing food | 0
reflexive cough | 0
intact gag reflexes | 0
decreased pharyngeal elevation | 0
swollen bilateral anterior neck area | -336
lower left quadrant of the anterior neck swollen | -336
mild tenderness | -336
follow-up plain radiograph of the chest | 0
leukocytosis | 0
neutrophilia | 0
increased C-reactive protein | 0
VFSS | 24
puree-like diet | 24
boiled rice | 24
semi-blended diet | 24
curd-type yogurt | 24
small and large amounts of fluid | 24
soft tissue posterior to the upper esophagus severely swollen | 24
retropharyngeal mass | 24
mechanical obstruction | 24
aspiration | 24
high risk of suffocation | 24
moderate-to-severe grade residues | 24
valleculae | 24
pyriform sinuses | 24
tube feeding | 24
unsuccessful insertion of nasogastric tube | 24
urgent contrast-enhanced CT scan of the neck | 24
loculated fluid collection | 24
retropharyngeal | 24
anterior cervical | 24
pericarotid | 24
prevertebral spaces | 24
upper mediastinum | 24
airway severely narrowed | 24
subglottic region | 24
reactive intraparotid or superficial cervical lymph nodes | 24
left side of the neck | 24
retropharyngeal abscess | 24
mediastinitis | 24
emergency tracheostomy | 48
incision to drain the abscess | 48
intravenous administration of ampicillin-sulbactam | 48
afebrile | 72
culture of the purulent discharge | 72
methicillin-resistant Staphylococcus aureus | 72
Klebsiella pneumoniae | 72
ceftriaxone-vancomycin | 72
CRP decreased | 120
intensive care | 240
general ward | 240
follow-up VFSS | 432
supraglottic penetration | 432
pharyngeal residue | 432
oral feeding training | 432
nasogastric tube feeding | 432
tracheostomy tube removed | 504
third VFSS | 576
silent aspiration | 576
full oral feeding | 576
follow-up chest CT | 576
improvement in the mediastinal extension | 576
WBC count normalized | 576
CRP normalized | 576
discharged | 1104