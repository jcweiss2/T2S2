79 years old | 0
white | 0
female | 0
IgG/λ MM | -144
hypertension | 0
type 2 diabetes mellitus | 0
dyslipidemia | 0
hyperuricemia | 0
increase in total serum proteins | -144
increase in γ-globulins | -144
increase in heavy IgG chains | -144
increase in free λ light chains | -144
IgG/λ monoclonal gammopathy | -144
anemia | -144
lytic bone lesions | -144
medullary aspirate | -144
plasmocytes with abnormal phenotypic characteristics | -144
oral melphalan | -144
prednisolone | -144
ECOG Performance Status 1 | -144
admitted to the emergency department | 0
fatigue | 0
severe bone pain | 0
diarrhea | 0
hemodynamic instability | 0
oliguric | 0
requiring oxygen | 0
decrease in breath sounds | 0
anemia | 0
leukocytosis | 0
neutrophilia | 0
thrombocytopenia | 0
C-reactive protein | 0
renal failure | 0
hypoalbuminemia | 0
arterial blood gas analysis | 0
type 1 respiratory insufficiency | 0
hyperlactacidemia | 0
bilateral pleural effusion | 0
diagnostic thoracentesis | 0
pleural fluid compatible with an exudate | 0
septic shock | 24
multiorgan failure | 24
renal failure | 24
hematological failure | 24
neurological failure | 24
cardiovascular failure | 24
respiratory failure | 24
broad-spectrum antibiotics | 24
sustained low-efficiency daily diafiltration | 24
deterioration | 48
dyspnea | 48
tachypnea | 48
desaturation | 48
aggravated pleural effusion | 48
therapeutic thoracentesis | 72
serosanguineous fluid | 72
pleural fluid analysis | 72
monoclonal γ-globulin spike | 72
flow cytometry | 72
abnormal PCs | 72
cytological exam | 72
immunocytochemical study | 72
bacteriological exam | 72
multi-resistant Escherichia coli | 72
myelomatous pleural effusion | 72
bacterial overinfection | 72
respiratory insufficiency | 96
poor prognosis | 96
extramedullary disease | 96
MPE | 96
palliative care | 120
death | 240