73 years old | 0
    man | 0
    presented to the emergency department | 0
    painless jaundice | -168
    elevated liver function tests | -168
    obstructive cholestatic pattern | -168
    intrahepatic duct dilatation | 0
    hypodense metastatic lesions | 0
    mass effect on the common hepatic duct | 0
    presumed primary cholangiocarcinoma | 0
    subjective heaviness to his eyes | 0
    cranial nerve deficit | 0
    admitted | 0
    ERCP | 24
    stent insertion | 24
    clinically improved the biliary obstruction | 24
    cytology brushing | 24
    undiagnostic | 24
    partial ptosis of the left eyelid | 48
    complete ptosis of the right eyelid | 48
    binocular diplopia | 48
    retro-orbital pain | 48
    partial left CNIII palsy | 48
    complete right CNIII palsy | 48
    CT scan | 48
    MRI of the brain and orbits | 48
    bilateral nodular lesions involving the cavernous sinus | 48
    maximum intensity projection 18F-FDG PET/CT | 48
    diffuse extensive nodal disease | 48
    extranodal disease | 48
    multiple abdominal organs involvement | 48
    bone involvement | 48
    soft tissues involvement | 48
    bilateral intense avidity of the cavernous sinus | 48
    targeted fine needle aspiration biopsies | 72
    left level III cervical node | 72
    hepatic lesion | 72
    B cells | 72
    CD10 expression | 72
    CD19 expression | 72
    CD20 expression | 72
    CD23 expression | 72
    Ki67 proliferation index 90% | 72
    rearrangement of c-MYC gene | 72
    confirmed Burkitt's lymphoma | 72
    CSF analysis | 72
    flow cytometry | 72
    negative for malignant cells | 72
    commenced on hyper-CVAD chemotherapy | 96
    neutropenic sepsis | 168
    admission to intensive care unit | 168
    de-escalation to mini R-CHOP | 168
    escalated to R-CHOP | 168
    intrathecal methotrexate | 168
    restaging 18F-FDG PET/CT | 672
    complete resolution of generalized Burkitt's lymphoma deposits | 672
    return to normal metabolic activity | 672
    full function of bilateral oculomotor nerves | 672
    clinical remission | 672
    