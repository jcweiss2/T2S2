43 years old | 0
    woman | 0
    abdominal pain | -720
    lumbar pain | -720
    nausea | -720
    nonproductive retching | -720
    denied fever | 0
    cesarean sections | unknown
    cholecystectomy | unknown
    hiatoplasty for hiatal hernia | -52560
    thoracic kyphosis | 0
    painful abdominal palpation | 0
    negative rebound tenderness test | 0
    normal bowel sounds | 0
    hemoglobin 15.8 g% | 0
    creatinine 1.09 mg/dL | 0
    hematocrit 48.9% | 0
    potassium 3.8 mEq/L | 0
    leucocytes 18.4 × 103/mm3 | 0
    sodium 140 mEq/L | 0
    bands 0% | 0
    ALT 20 U/L |# hello-world
Just another repository

This is a test readme.
