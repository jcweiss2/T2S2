18 years old | 0  
    male | 0  
    admitted to the hospital | 0  
    RSV infection | -2160  
    failure to thrive | -2160  
    prominent bulging of the anterior fontanel | -2160  
    severe intracranial hypertension | -2160  
    hydrocephalus | -2160  
    ventriculoperitoneal shunt placement | -2160  
    deflection of the growth curve | -2160  
    generalized sclerosis of the bone | -2160  
    osteoclast-poor osteopetrosis | -2160  
    TCIRG1 mutation | -2160  
    allogeneic HSCT | -1344  
    impaired vision of the right eye | -1344  
    acute otitis media | -1200  
    otitis media with effusion | -1200  
    placement of tympanostomy tubes | -840  
    dehiscent jugular bulb | -840  
    conductive hearing loss | -840  
    small tympanic cavity | -840  
    thickened superstructures and footplates of the stapes | -840  
    upward and medial angulation of the petrous bone apex | -840  
    inclined and verticalized tegmen | -840  
    rehabilitation with hearing aid | -840  
    monocular blindness | -840  
    stable blood values | -840  
    favorable development | -840  
    recurrence of otitis media | 0  
    good general health | 0  
    stable audiometric thresholds | 0  

<|eot_id|>
