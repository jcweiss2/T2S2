32 years old | 0
male | 0
bipolar disorder | -152
lithium | -152
weight gain | -61
olanzapine | -61
nausea | -61
vomiting | -61
severe epigastric pain | -61
no haematemesis | -61
no melaena | -61
no jaundice | -61
no previous history of pancreatitis | -61
no gall stone disease | -61
family history for diabetes negative | -61
heart rate 105-115/min | 0
blood pressure 110/56 mm Hg | 0
respiratory rate 24-28/min | 0
febrile | 0
epigastric tenderness | 0
guarding | 0
normal liver dullness on percussion | 0
absent bowel sound | 0
bulky pancreas | 0
pancreatic oedema | 0
no peripancreatic collection | 0
no abnormality on upper GI endoscopy | 0
increasing pain intensity | 0
referred to back | 0
breathlessness | 240
admitted to intensive care unit | 240
low arterial O2 saturation | 240
dyspnoea | 240
all drugs stopped | 240
serum lipase 900 U/L | 240
serum triglyceride 560 mg/dL | 240
blood sugar 230 and 478 mg/dL | 240
normal serum calcium level | 240
mild derangement in liver function tests | 240
HIV serology status nonreactive | 240
mask oxygen | 240
intubated | 240
mechanical ventilation | 240
lung protective strategy | 240
left sided pleural effusion | 240
contrast enhanced computed tomography scan abdomen | 312
pancreatic necrosis | 312
oedema | 312
peripancreatic collection | 312
no cholelithiasis | 312
no choledocholithiasis | 312
large pelvic fluid collection | 312
left sided percutaneous drain | 312
USG guided percutaneous drainage | 312
inotropic and vasopressor support | 312
repeat CECT | 504
pancreatic necrosis | 504
gas formation in pancreas | 504
peripancreatic areas | 504
CT severity index 6-7/10 | 504
diagnosis of EP | 504
sepsis | 504
appropriate antibiotics | 504
peripancreatic drain | 504
culture report from drained fluid | 504
anaerobic enteric organisms | 504
intravenous imipenem and clindamycin | 504
peripancreatic region irrigated with metronidazole | 504
sustained low efficiency dialysis | 504
acute kidney injury | 504
hyperglycaemia controlled with regular insulin infusion | 504
extubated | 624
enteral feeding | 624
nasojejunal | 624
discharged from the hospital | 1152
drug and life style advice | 1152
correcting dysglycaemia | 1152
dyslipidaemia | 1152
increased body weight | 1152
olanzapine replaced | 1152
lost about 15 kg body weight | 1152
no symptoms/signs of pancreatitis | 1152