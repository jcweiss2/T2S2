66 years old | 0\
male | 0\
dual-chamber pacemaker implanted | -10584\
sick sinus syndrome | -10584\
paroxysmal atrial fibrillation | -10584\
severe lumbar back pain | 0\
mental status changes | 0\
hypotension | 0\
acute renal failure | 0\
hypoxemic respiratory failure | 0\
intubation | 0\
severe sepsis | 0\
hemodynamic support with 2 vasoactive agents | 0\
blood cultures yielded methicillin-sensitive Staphylococcus aureus | 0\
vancomycin | 0\
nafcillin | 0\
transthoracic echocardiogram | 0\
left ventricular ejection fraction of 55% | 0\
positive bubble study | 0\
patent foramen ovale | 0\
computed tomography scan of the chest, abdomen, and pelvis | 0\
osteomyelitis of the lower spine | 0\
magnetic resonance imaging of the brain | 0\
multiple small, 2- to 3-mm, acute infarctions | 0\
septic emboli to the distal extremities | 0\
transesophageal echocardiogram | 0\
vegetation within the right atrium | 0\
vegetation attached to the pacemaker lead | 0\
mobile structure attached to the pacemaker lead within the right ventricle | 0\
cardiothoracic surgery consulted | 0\
laser lead extraction procedure | 0\
bilateral femoral veins accessed | 0\
16F GORE DrySeal Flex introducer sheath | 0\
8F sheath | 0\
9F sheath | 0\
8F catheter | 0\
91.4-cm 12F 45-degree curved sheath | 0\
115-cm Indigo CAT8 XTORQ | 0\
intracardiac echocardiography | 0\
aspiration | 0\
vegetation removed | 0\
laser lead extraction | 0\
pocket inspected | 0\
pocket closed | 0\
Penumbra and ICE systems removed | 0\
hemostasis achieved | 0\
vegetations sent to pathology | 0\
pathology of the vegetation specimens | 0\
gram-positive cocci in chains | 0\
culture-positive for methicillin-sensitive Staphylococcus aureus | 0\
condition improved | 48\
condition deteriorated | 72\
tissue necrosis of the distal upper and lower extremities | 72\
lactic acidosis | 72\
worsening renal failure | 72\
care withdrawn | 72\
extubated to comfort care | 72\
died | 72