66 years old | 0
female | 0
admitted to hospital | 0
fever | -192
close contact with confirmed COVID-19 case | -192
SARS-CoV-2 RNA detected | -192
nasopharyngeal and throat swab | -192
RT-PCR method | -192
E-gene Ct 22.04 | -192
RdRp Ct 35.09 | -192
Roche LightCycler 480 | -192
initial supportive treatment for COVID-19 | -192
hypertension | 0
osteopenia | 0
Perindopril/Amlodipine | 0
Cholecalciferol (vitamin D3) | 0
ex-smoker | 0
20 pack years | 0
no history of immunosuppression | 0
no chronic organ dysfunction | 0
no history of fungal colonisation | 0
independent in activities of daily living | 0
fever | 0
respiratory rate 26/min | 0
pulse 80/min | 0
blood pressure 120/70 mmHg | 0
low oxygen saturation (SpO2 89% on room air) | 0
increase in work of breathing | 0
bibasal coarse crepitations | 0
arterial blood gas sampling | 0
pH 7.44 | 0
PaO2 70 mmHg | 0
PaO2/FiO2 = 334 | 0
PaCO2 34 mmHg | 0
lactate 0.9 mmol/L | 0
white blood cell count (WCC) 5.3 × 10^9/L | 0
neutrophil differential count 3.9 × 10^9/L | 0
lymphocyte count 1.2 × 10^9/L | 0
liver function tests | 0
AST 52U/L | 0
ALT 32 U/L | 0
GGT 61U/L | 0
LDH 429 U/L | 0
renal function normal | 0
blood cultures | 0
Facklamia hominis | 0
urine culture | 0
Escherichia coli | 0
Ceftriaxone | 0
Ceftriaxone 1g daily | 0
Azithromycin | 0
Azithromycin 500mg daily | 0
supplemental oxygen | 0
subcutaneous enoxaparin sodium | 0
venous thromboembolism prophylaxis | 0
no specific therapy targeting COVID-19 infection | 0
deteriorated rapidly | 48
progressive dyspnoea | 48
increasing oxygen requirement | 48
admitted to ICU | 48
temperature 39.5°C | 48
respiratory rate 40/min | 48
oxygen saturation 91% on high flow nasal prongs (HFNP) | 48
FiO2 40% | 48
40 L/m of airflow | 48
moderate increase in work of breathing | 48
trans-thoracic echocardiogram | 48
normal biventricular function | 48
mild right ventricular dilatation | 48
arterial blood gas | 48
pH 7.46 | 48
PaO2 59 mmHg | 48
PaO2/FiO2 = 148 | 48
PaCO2 31 mmHg | 48
awake prone positioning | 48
elective endotracheal intubation | 48
mechanical ventilation | 48
lung-protective ventilation | 48
Tidal volume 4–6 ml/kg | 48
PEEP 12 cmH2O | 48
Plateau pressure <30 cmH2O | 48
PaO2 >60 mmHg | 48
pH > 7.2 | 48
ARDS net protocol | 48
further deterioration in ventilatory parameters | 96
severe ARDS criteria | 96
PaO2/FiO2 = 82 mmHg | 96
PEEP = 12 cmH2O | 96
worsening respiratory function | 192
hypercapnoea | 192
fever absent | 192
increased inflammatory markers | 192
C reactive protein 351mg/L | 192
deranged LFTs | 192
ALT = 125 U/L | 192
AST = 154 U/L | 192
GGT = 611 U/L | 192
ALP = 229 U/L | 192
raised ferritin | 192
raised D-dimer | 192
fibrinogen 5.8g/L | 192
chest radiology | 192
significant progression of bilateral consolidative opacities | 192
respiratory tract specimens | 192
non-bronchoscopic endotracheal aspirate (ETT) | 192
persistent SARS-CoV-2 RNA | 192
Piperacillin/Tazobactam | 192
prone ventilation | 192
improvement in ventilatory parameters | 192
fungal elements | 192
Gram staining | 192
Aspergillus fumigatus complex | 192
Horse blood agar | 192
Chocolate agar | 192
uniseriate conidial heads | 192
phialides limited to the upper two thirds of the vesicle | 192
culture mount stained with lactophenol cotton blue | 192
new onset of fever | 240
progressive bilateral consolidation | 240
Voriconazole | 240
6 mg/kg loading | 240
3mg/kg twice daily | 240
rapid clinical and radiological progress | 288
fevers settled | 288
inflammatory markers improved | 288
liver function normalized | 288
steady-state Voriconazole trough levels | 288
2.72mg/L | 288
extubated | 372
treatment de-escalated | 372
oral Voriconazole | 372
300mg twice daily | 372
ward rehabilitation | 432
two negative SARS-CoV-2 RT-PCR clearance swabs | 432
discharged home | 456
contrast-enhanced computed tomography (CECT) | 540
bilateral organising pneumonia | 540
fibrosis | 540
probable small segmental pulmonary embolism | 540
left upper lobe | 540
Voriconazole ceased | 540
total duration of treatment one month | 540
risk of drug-drug interaction | 540
Apixaban | 540
abnormal liver function testing | 540
Voriconazole trough level 3.6mg/L | 540
mild dry cough | 540
improved effort tolerance | 540
no systemic features | 540