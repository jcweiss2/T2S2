22 years old | 0
male | 0
admitted to ICU | 0
fever | -240
cough | -192
sputum production | -192
respiratory distress | -24
altered sensorium | -24
tachycardia | 0
tachypnea | 0
hypotension | 0
hypoxemia | 0
right lower lobe consolidation | 0
intubation | 0
mechanical ventilation | 0
bronchoalveolar lavage | 0
blood samples sent for culture | 0
provisional diagnosis of acute febrile illness | 0
provisional diagnosis of pneumonia | 0
provisional diagnosis of septic shock | 0
piperacillin-tazobactum started | 0
vancomycin started | 0
antimalarials started | 0
tests for malaria done | 0
tests for leptospirosis done | 0
tests for dengue done | 0
tests for typhoid done | 0
all tests negative | 0
prone ventilation | 0
ARDS net protocol | 0
PaO2/FiO2 ratio 100 | 0
MRSA positive in blood culture | 24
MRSA positive in BAL culture | 24
i.v. vancomycin added | 24
PaO2/FiO2 ratio improved | 120
extubation | 168
post-extubation hypoxia | 168
respiratory rate 28-30/min | 168
computed tomography pulmonary angiogram | 168
high resolution computed tomography chest | 168
patchy consolidation | 168
cavity in lateral basal segment of right lower lobe | 168
pulmonary angiogram normal | 168
vancomycin continued | 168
respiratory rate settled | 672
discharged | 672