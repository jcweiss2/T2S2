three years old | 0
female | 0
complex congenital heart disease | -672
previous cardiac surgeries | -672
admitted to the pediatric intensive care unit | 0
shock | 0
cardiopulmonary arrest | 0
resuscitation | 0
thrombosis in her right ventricle-to-pulmonary artery conduit | 0
severe hypoxic-ischemic encephalopathy | 0
acute kidney injury | 0
neurological rehabilitation | 0
transition to home ventilation | 0
treatment for dystonia | 0
treatment for heart failure | 0
treatment for endocarditis | 0
treatment for pulmonary embolism | 0
stem cell therapy for neurological dysfunction | 0
metformin therapy initiated | -408
metformin dose increased | -144
new wide complex bradycardia | 0
peaked T waves | 0
blood pressure = 90/40 mmHg | 0
respiratory rate = 26 breaths per minute | 0
temperature = 37.2 °C | 0
oxygen saturation = 87% | 0
poorly perfused | 0
prolonged capillary refill time | 0
lethargic | 0
severe lactic acidosis | 0
hyperkalemia | 0
managed for hyperkalemia | 0
propranolol discontinued | 0
hypotensive | 0
dopamine infusion | 0
norepinephrine infusion | 0
higher ventilator support | 0
clinical status improved | 3
support therapies weaned | 3
similar episode recurred | 12
rise in serum lactate | 12
hyperkalemia | 12
metformin discontinued | 12
no further episodes | 12
clinical status returned to baseline | 12
creatinine levels doubled | -120
metformin dose increased | -144
renal insufficiency | -120
intravascular depletion | -120
metformin levels not collected | 0 
sepsis ruled out | 0
rhabdomyolysis ruled out | 0
creatinine kinase levels normal | 0
blood cultures sterile | 0