39 years old | 0
female | 0
gestational age 32 weeks | 0
presented to the emergency room | 0
shortness of breath | 0
progressive limb weakness | 0
history of worsening neck pain | -17520
weakness in right arm | -1440
weakness in left arm | -1440
weakness in both legs | -1440
no complaints of anosmia | 0
no complaints of seizure | 0
no complaints of blurred vision | 0
no complaints of slurred speech | 0
no complaints of dysphagia | 0
no complaints of hoarseness | 0
no complaints of skewed face | 0
numbness from neck down | 0
no urination disturbances | 0
no defecation disturbances | 0
fever | -72
no medical history of cancer | 0
no family history of cancer | 0
history of contraceptive injection for 15 years | -131400
consumption of ibuprofen | -17520
consumption of paracetamol | -17520
intact mental status | 0
no meningeal signs | 0
cranial nerve palsy | 0
tetraplegia | 0
hypoesthesia below C3-C4 spinal cord segments | 0
abnormal proprioception in all extremities | 0
increased tendon reflexes in both arms | 0
positive Babinski reflex | 0
positive Chaddock reflex | 0
PCR positive for COVID-19 | 0
chest radiography paracardial infiltrates | 0
respiratory failure | 0
increased D-dimer (2000 mg/dL) | 0
hypokalemia | 0
admitted to intensive care unit | 0
intubation | 0
treatment with high-dose n-acetylcysteine | 0
treatment with remdesivir | 0
treatment with zinc | 0
treatment with vitamin D | 0
treatment with vitamin C | 0
fetal distress | 0
emergency cesarean section | 0
successful surgery | 0
baby did not survive | 0
brain MRI mass in foramen magnum | 0
cervical MRI mass with homogenous contrast enhancement | 0
spinal cord edema | 0
administered steroids | 0
rapid deterioration | 0
tumor excision by craniotomy | 0
histopathological examination transitional type WHO grade 1 meningioma | 0
histopathological examination angiomatous type WHO grade 1 meningioma | 0
whorl pattern | 0
proliferating meningothelial cells with oval to spindle nuclei | 0
psammoma bodies | 0
proliferation of blood vessels with hyalinization | 0
brief increased awareness after surgery | 0
continued deterioration | 0
close monitoring | 0
blood pressure decreased to 60/30 mmHg | 0
administered norepinephrine | 0
suspected sepsis | 0
death due to septic shock | 0
death due to respiratory failure | 0
