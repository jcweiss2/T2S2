36 years old | 0
male | 0
police officer | 0
admitted to the hospital | 0
snakebite | -2
anti-snake venom | -2
IV fluids | -2
antibiotics | -2
supportive care | -2
decreased urine output | 24
deranged renal functions | 24
hemodialysis | 24
dull drowsy state | 72
stable hemodynamic | 72
bilateral decreased air entry | 72
swelling at the site of bite | 72
cellulitis | 72
blister formation | 72
hemoglobin 7.6 g/dL | 72
total leucocyte count 15,000 | 72
platelets 50,000 | 72
normal coagulation profile | 72
activated partial thromboplastin time 15 seconds | 72
International Normalized Ratio 1.19 | 72
bedside clotting time 5 minutes | 72
bleeding time 32 seconds | 72
deranged kidney function tests | 72
urea 167 mg/dL | 72
creatinine 6.17 mg/dL | 72
total creatine phosphokinase 52,168 | 72
transaminitis | 72
serum glutamic-oxaloacetic transaminase/pyruvic transminase 1,985/252 | 72
total bilirubin 4.56 | 72
direct bilirubin 0.64 | 72
indirect bilirubin 3.92 | 72
sepsis | 72
procalcitonin 4.79 | 72
oxygen support | 72
intravenous antibiotics | 72
antivenom | 72
acute kidney shutdown | 72
anuric status | 72
hemodialysis | 72
heparin free | 72
ultrafiltration | 72
persistent fall in hemoglobin | 120
multiple blood transfusions | 120
hemolysis | 120
fragmented cells | 120
spherocytes | 120
lactate dehydrogenase 4,128 | 120
worsening of hypoxemia | 168
bilateral infiltrates on chest X-ray | 168
pleural effusion | 168
high-flow nasal cannula oxygen support | 168
hemoptysis | 168
CT chest | 168
multifocal peribronchial air space opacification | 168
ground-glass opacification | 168
moderate pleural effusion | 168
lung collapse | 168
probable diagnosis of diffuse alveolar hemorrhage | 168
steroids | 168
methylprednisolone 80 mg/day | 168
coagulation profile | 168
thrombocytopenia | 168
bilateral pleural drain | 168
transudative picture | 168
sterile | 168
two-dimensional echocardiography | 168
good biventricular systolic functioning | 168
ejection fraction 55% | 168
ultrasound abdomen | 168
bulky hypoechoic bilateral kidneys | 168
reduced corticomedullary differentiation | 168
autoimmune pathology | 168
antinuclear antibodies negative | 168
antineutrophil cytoplasmic antibodies negative | 168
perinuclear antineutrophil cytoplasmic antibodies negative | 168
sputum culture | 168
E. coli | 168
antibiotics upgraded to meropenem | 168
no signs of improvement | 240
hemoptysis continued | 240
progressive fall in hemoglobin | 240
persistent AKI | 240
plasma exchange therapy | 480
first plasma exchange | 480
centrifugation technology | 480
internal jugular venous access | 480
5% Hum albumin | 480
replacement fluid | 480
monitoring for electrolytes/fluid balance | 480
proteins | 480
coagulation profile | 480
renal parameters improved | 480
urine output 25 to >50 mL/hour | 480
secondary sepsis | 504
leukocytosis | 504
procalcitonin 21 | 504
polymyxin B | 504
electively intubated | 504
worsening type I respiratory failure | 504
five sessions of consecutive plasma exchange | 504
intermittent hemodialysis | 504
renal support | 504
clinical signs of recovery | 528
improving oxygen requirement | 528
settling leukocytosis | 528
renal function improved | 528
creatinine 3.5 mg/dL | 528
urine output improved | 528
from 500 mL/24 hour to 2,100 mL/24 hour | 528
pulmonary hemorrhage settled | 528
minimal tracheal bleed | 528
static hemoglobin | 528
bronchoscopy | 528
clear airways | 528
repeat high resolution computed tomography chest | 528
multifocal peribronchial consolidations | 528
bilateral effusion | 528
antibiotics | 528
supportive care | 528
successful weaning trials | 552
extubated | 552
low-flow oxygen | 552
hemodynamically stable | 552
serial X-rays | 552
clearing out infiltrates | 552
residual right basal collapse consolidation | 552
discharged | 720
stable condition | 720
creatinine 1.2 | 720
good urine output | 720
cleared out chest X-ray | 720
follow-up in outpatient department | 720
healthy | 720
no sequelae | 720
fully recovered AKI | 720
creatinine 0.96 | 720
chest X-ray clear | 720