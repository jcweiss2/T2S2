21 years old | 0
female | 0
pregnant | 0
admitted to the obstetric department | 0
pre-term labor | 0
nifedipine administration | 0
pulmonary edema | 1
hypoxemia | 1
transfer to ICU | 1
blood pressure 101/61 mm Hg | 1
sinus tachycardia | 1
oxygen saturation 98% | 1
loud first heart sound | 1
diastolic murmur | 1
bilateral wheezing | 1
jugular venous distension | 1
systolic blood pressure fall | 2
desaturation | 2
metabolic acidosis | 2
hyperlactatemia | 2
intubation | 2
ventilation | 2
pulmonary edema confirmed by chest X-ray | 2
severe mitral stenosis | 2
normal left ventricular function | 2
enlargement and pressure overload of the left atrium | 2
severe pulmonary hypertension | 2
loop diuretics administration | 4
full-dose heparin administration | 4
no fetal distress | 4
severe rheumatic mitral stenosis | 4
spontaneous vaginal delivery | 12
baby alive | 12
baby transferred to intensive neonatal care unit | 12
mother in critical state | 12
hypotension | 12
endometritis | 12
sepsis | 12
ceftriaxone administration | 12
ampicillin administration | 12
valvuloplasty postponed | 12
infection resolution | 192
percutaneous double balloon mitral valvuloplasty | 192
mitral mean gradient reduced | 192
mitral area increased | 192
pulmonary pressure normalized | 192
extubation | 216
recovery | 216