9 years old | 0
    female | 0
    fever | 0
    jaundice | 0
    right upper quadrant abdominal pain | 0
    rhabdomyosarcoma of the right deltoid and triceps muscles | -1440
    VAC chemotherapy (vincristine, 1.5 mg/m2/day; actinomycin-D, 1.35 mg/m2/day; cyclophosphamide, 1.2 g/m2/day for 3 days) | -1440
    wide excision of the tumor | -1440
    postoperative VAC chemotherapy | -1440
    mild abdominal pain | -192
    neutropenic fever | -192
    white blood cell 0.78×103/μL | -192
    hemoglobin 6.9 g/dL | -192
    platelets 4×103/μL | -192
    intravenous broad-spectrum antibiotics (piperacillin and tazobactam) | -192
    transfusion (red blood cells, platelets) | -192
    granulocyte colony stimulating factor | -192
    mild elevation of liver enzymes (AST, 103 U/L; ALT, 77 U/L) | -192
    total bilirubin 1.5 mg/dL | -192
    abdominal pain aggravated | -168
    persistent fever | -168
    pancytopenia (WBC, 0.42×103/μL; Hb, 8.1 g/dL; platelet, 6×103/μL) | -168
    marked increase in liver enzymes (AST, 519 U/L; ALT, 370 U/L) | -168
    hyperbilirubinemia (total bilirubin, 4.8 mg/dL) | -168
    prolonged prothrombin time (1.17 international normalized ratio) | -168
    active partial thromboplastin time (55.2 seconds) | -168
    hepatomegaly, 3.5 cm distal from the right costal margin | -168
    sepsis | -168
    antibiotics changed to vancomycin and meropenem | -168
    addition of intravenous immunoglobulin | -168
    fever peaked to 38.9°C | -144
    severe abdominal pain | -144
    icteric sclerae | -144
    aggravated hepatomegaly | -144
    abdominal distension | -144
    body weight increased by 6.1% (2.5 kg) | -144
    AST/ALT 1,172/810 U/L | -144
    total/direct bilirubin 6.1/3.1 mg/dL | -144
    abdominal Doppler ultrasonography showed reversed blood flow of the right portal vein | -144
    SOS diagnosis | -144
    treatment with defibrotide (32 mg/kg/day in four divided doses) | -144
    transferred to the intensive care unit | -144
    condition became unstable | -144
    chest radiography showing diffuse pleural effusion | -144
    irritable | -144
    did not recognize her mother and medical personnel | -144
    liver enzyme levels peaked (AST 2,110 U/L; ALT 1,908 U/L) | -144
    total bilirubin 15.1 mg/dL | -144
    direct bilirubin 8.6 mg/dL | -144
    ammonia level increased (135 μg/dL) | -144
    hepatic encephalopathy | -144
    vasopressor infusion | -144
    paracentesis of the ascites | -144
    glycerin enema | -144
    rifaximin | -144
    lactulose (through an L-tube) | -144
    mechanical ventilation started | -96
    defibrotide treatment continued for 10 days | -144
    body weight began to decrease | -72
    fever gradually subsided | -72
    laboratory results showed improvement | -72
    weaned from mechanical ventilator | 408
    abdominal US normalized blood flow of the right portal vein | 528
    discharged | 744
    bilirubin level normalized | -
    parents refused further chemotherapy | -
    subsequent surveillance imaging studies showed no evidence of recurrence of cancer | -
    no sequelae to the liver | -
    
