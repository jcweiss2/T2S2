61 years old | 0
    male | 0
    non-Hodgkin’s lymphoma | 0
    prior radiation therapy | 0
    coronary artery disease | 0
    coronary artery bypass graft | 0
    mechanical aortic valve replacement | 0
    severe bicuspid aortic valve stenosis | 0
    presented to outside hospital | 0
    fever | 0
    malaise | 0
    respiratory distress | 0
    treated with broad-spectrum intravenous antibiotics | 0
    sepsis | 0
    intubated | 0
    respiratory failure | 0
    methicillin-sensitive Staphylococcus aureus in blood cultures | 0
    transesophageal echocardiogram | 0
    vegetation on mechanical aortic valve | 0
    prosthetic endocarditis | 0
    antibiotic therapy narrowed to intravenous oxacillin, gentamicin, rifampin | 0
    pulseless electrical activity cardiac arrest | -144
    complete heart block | -144
    placement of external MRI-compatible pacemaker | -144
    placement of right ventricle MRI-compatible active-fixation lead | -144
    left subclavian approach | -144
    stenosis of internal jugular veins | -144
    computed tomography of head | -144
    multifocal bilateral infarcts | -144
    small areas of adjacent parenchymal hemorrhage | -144
    subarachnoid hemorrhage | -144
    persistent ventilator requirement | -144
    left pneumothorax | -144
    chest tube placement | -144
    progressive renal injury | -144
    acute tubular necrosis | -144
    transferred to our institution | -144
    intubated | -144
    sedated | -144
    corneal reflexes present | -144
    gag reflexes present | -144
    grimaced in response to upper extremity noxious stimuli | -144
    no response to lower extremity noxious stimuli | -144
    white blood count 22,700/μL | -144
    hemoglobin 9.4 g/dL | -144
    platelets 402,000/μL | -144
    creatinine 3.2 mg/dL | -144
    limited transthoracic echocardiogram | -144
    aortic valve vegetation | -144
    trace aortic regurgitation | -144
    brain MRI requested | -24
    repeat contrast CT contraindicated | -24
    noncontrast CT insufficiently sensitive | -24
    MRI approved | 0
    MRI-compatible temporary active-fixation right ventricular pacing lead | 0
    externalized pacemaker generator | 0
    use of transmit-receive head coil | 0
    imaging in normal mode | 0
    repositioning of generator to upper left chest | 0
    insulating generator from direct skin contact | 0
    gauze pads inserted | 0
    transparent film dressing | 0
    pre-MRI impedance 773 ohms | 0
    pre-MRI thresholds 0.3 V at 0.4 ms | 0
    pacing mode VOO at 80 bpm | 0
    transcutaneous pacing pads placed | 0
    monitored by intensive care nurse | 0
    MRI completed uneventfully | 0
    post-MRI impedance unchanged | 0
    post-MRI thresholds unchanged | 0
    post-MRI battery capacity unchanged | 0
    chest roentgenograph no lead migration | 0
    bilateral multifocal infarcts | 0
    septic emboli | 0
    no brain abscess | 0
    cardiac CT requested | 24
    over-breathing ventilator | 24
    administered benzodiazepine bolus | 24
    neuromuscular blockade | 24
    device reprogrammed to VOO at 70 bpm | 24
    hypoattenuated mass associated with mechanical aortic valve | 24
    vegetation | 24
    thickening of mitral-aortic intervalvular fibrosa | 24
    perivalvular involvement | 24
    no abscess | 24
    lead tip within right ventricular apex | 24
    operative mortality risk 40% | 24
    surgical intervention not offered | 24
    transition to comfort-oriented care | 24
    death | 48