59 years old | 0\
female | 0\
blood type O | 0\
Rh positive | 0\
liver cancer | -672\
transarterial embolization | -672\
sorafenib | -672\
dizziness | -672\
skin ulcers | -672\
radiation therapy | -24\
Piggyback LT | 0\
hepatitis B | 0\
entecavir | 0\
HBsAg 113.23 IU/mL | 0\
anti-HBs 0 mIU/mL | 0\
HBeAg 0.08 PEI µ/mL | 0\
anti-HBe >4.4 PEI µ/mL | 0\
anti-HBc 8.26 PEI µ/mL | 0\
human immunodeficiency virus negative | 0\
hepatitis A negative | 0\
hepatitis C negative | 0\
donor 21 years old | 0\
donor male | 0\
donor blood type O | 0\
donor Rh positive | 0\
donor HLA class-I A11, A30 | 0\
donor HLA class-II B13 | 0\
donor HLA class-III DR11, DR15 | 0\
donor HLA class-IV DQ6, DQ7 | 0\
recipient HLA class-I A2, A11 | 0\
recipient HLA class-II B13, B46 | 0\
recipient HLA class-III DR14, DR15 | 0\
recipient HLA class-IV DQ5, DQ6 | 0\
acute renal failure | 0\
hematoma around the liver | 0\
intravenous administration of hepatitis B immunoglobulin | 24\
immunosuppressive drugs | 24\
steroids | 24\
tacrolimus | 24\
continuous hemodialysis | 24\
intermittent infusion of fresh frozen plasma | 24\
leukocyte-depleted red blood cells | 24\
other blood products | 24\
active bleeding in the abdominal cavity ceased | 24\
renal function gradually recovered | 24\
massive tumor necrosis | 24\
necrosis accounted for ~90% | 24\
surviving tumor accounted for ~10% | 24\
fever | 240\
fever 37–39°C | 240\
fever peaking at 23:00 h daily | 240\
PCT levels rose to 10.3 ng/mL | 240\
PCT levels dropped to 3 ng/mL | 312\
blood cultures negative | 312\
cytomegalovirus negative | 312\
Epstein–Barr virus negative | 312\
obscure red spots on the patient’s chest | 312\
no symptoms such as itching | 312\
Nikolsky sign negative | 312\
tacrolimus administration changed to sirolimus | 408\
mycophenolate mofetil added | 408\
sputum culture suggested the presence of Acinetobacter baumannii | 432\
sputum culture suggested the presence of methicillin-resistant Staphylococcus aureus | 432\
rash advanced into erythematous macules and papules | 456\
rash spread to the limbs, palms, neck, and face | 456\
oral examination revealed white ulcers on both sides of the buccal mucosa and lips | 456\
severe bone marrow suppression | 456\
WBC count 0.86 × 10^9/L | 456\
PLT count 35 × 10^9/L | 456\
HGB level 70 g/L | 456\
transferred to the intensive care unit | 456\
gamma globulin administration | 456\
skin biopsy | 456\
fluorescence in situ hybridization of the peripheral blood | 456\
abdominal incision split | 696\
sutured again | 696\
bone marrow aspiration | 768\
bone marrow pathology report revealed no special lesions | 768\
bone marrow cell morphology examination revealed that the bone marrow cells were proliferating and active | 768\
megakaryocyte production was reduced | 768\
platelet levels decreased | 768\
FISH analysis of the peripheral blood followed by flow cytometry detected 3% donor lymphocytes | 792\
skin biopsy specimens exhibited epidermal dyskeratosis | 792\
basic vacuolization | 792\
lymphocytic infiltrates | 792\
consistent with grade-1 acute lt-GVHD | 792\
differential diagnoses include bacterial, fungal, and viral infections | 792\
drug reactions | 792\
toxic epidermal necrolysis | 792\
hemophagocytic syndrome | 792\
blood culture was negative at the onset of the rash | 792\
no history of allergies to drugs | 792\
no drugs were suspected of causing allergy | 792\
serological tests of the virus were negative | 792\
no macrophages phagocytosing neutrophils or platelets were observed in the bone marrow biopsy | 792\
collective findings, together with the clinical course, were consistent with the diagnosis of lt-GVHD | 792\
analysis of serum T-lymphocyte subsets revealed that the ratio of CD4:CD8 was reversed | 792\
concentration of serum immunoglobin M was reduced to 0.3 g/L | 792\
continuous platelet transfusion | 792\
use of thrombopoietin | 792\
PLT count dropped to 3.2 × 10^9/L | 792\
rash was significantly reduced | 912\
general condition continued to deteriorate | 912\
serum ferritin levels increased to 11,276.55 ng/mL | 912\
esophageal and oral ulcers continued to worsen | 912\
prevented the patient from eating | 912\
temperature rose to 39.4°C | 1128\
hallucinations | 1128\
destruction of the patient’s skin, bone marrow, and mucosal epithelium further increased her immunodeficiency | 1128\
resulting in her course of disease being accompanied by multiple infections | 1128\
MRSA | 1128\
Acinetobacter baumannii | 1128\
Enterococcus faecalis | 1128\
despite intensive treatments | 1128\
serum immunoglobin M level was reduced to 0 g/L | 1128\
succumbed to septic shock and multiple organ dysfunction syndrome | 1656