66 years old | 0
female | 0
advanced diffuse large B-cell lymphoma | -2190
diagnosed with DLBCL | -2190
R-CHOP | -2190
rituximab | -2190
cyclophosphamide | -2190
doxorubicin | -2190
vincristine | -2190
prednisone | -2190
autologous hematopoietic stem cell transplant | -1560
DLBCL recurred | -780
R-CHOP | -780
transthoracic echocardiogram | -720
left ventricular ejection fraction 55% to 60% | -720
global longitudinal strain -12% | -720
admitted to the hospital with acute decompensated heart failure | 0
left ventricular ejection fraction 25% | 0
global left ventricular dysfunction | 0
positron emission tomography scan | 0
progression of DLBCL | 0
new pulmonary nodules | 0
referred to CAR T cell therapy | 0
coronary computed tomography | 0
mild coronary artery disease | 0
cardiac magnetic resonance imaging | 0
no evidence of infiltrative or inflammatory disease | 0
anthracycline-induced cardiomyopathy | 0
furosemide | 0
guideline-directed medical therapy | 0
lisinopril | 0
metoprolol succinate | 0
referred to cardio-oncologist | 0
good exercise tolerance | 0
right heart catheterization | 0
mildly elevated biventricular filling pressures | 0
normal cardiac output | 0
CAR T cell therapy | 0
cytokine release syndrome | 0
fevers | 48
derangements in blood pressure | 48
oxygenation | 48
hypotension | 48
hypoxemia | 48
vasodilatory shock | 48
atrial or ventricular arrhythmias | 48
ventricular dysfunction | 48
invasive pulmonary artery catheter monitoring | 0
CardioMEMS device | 0
implanted | 0
three months of GDMT | 2160
repeat right heart catheterization | 2160
normal filling pressures | 2160
preserved cardiac output | 2160
successful placement of CardioMEMS device | 2160
repeat TTE | 2160
no improvement in LVEF | 2160
right ventricular performance improved | 2160
admitted for pre-treatment | 2160
lympho-depleting chemotherapy | 2160
fludarabine | 2160
cyclophosphamide | 2160
neutropenic fever | 2160
hypotension | 2160
intravenous antibiotics | 2160
GDMT held | 2160
axicabtagene ciloleucel | 2160
CAR T cells | 2160
infusion | 2160
mild CRS | 72
fevers | 72
sinus tachycardia | 72
systolic blood pressures in the 90s | 72
elevated pulmonary artery diastolic pressure | 72
intravenous furosemide | 72
tocilizumab | 72
worsening tachypnea | 120
new oxygen requirement | 120
second dose of tocilizumab | 120
diffuse pulmonary opacities | 120
noncardiogenic pulmonary edema | 120
atrial flutter | 288
rapid ventricular rates | 288
acute hypoxic respiratory failure | 288
cardiogenic pulmonary edema | 288
intubation | 288
low-dose norepinephrine | 288
amiodarone | 288
converted to sinus rhythm | 288
weaned off vasopressors | 432
extubated | 432
discharged to acute rehabilitation | 720
unable to restart GDMT | 720
hypotension | 720
pulmonary artery diastolic pressure 6 mmHg | 720
furosemide 20 mg daily | 1008
nausea | 1344
acute shortness of breath | 1440
oxygen saturation 88% | 1440
pulmonary edema | 1440
possible left lower lobe infiltrate | 1440
intubated | 1440
progressive hypoxic respiratory failure | 1440
multiple vasopressors | 1440
mixed septic and cardiogenic shock | 1440
cardiac arrest | 1440
ventricular tachycardia | 1440
expired | 1440