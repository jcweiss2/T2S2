45 years old | 0
female | 0
fall from 18 feet height | -504
difficulty in breathing | -48
completely treated pulmonary tuberculosis | -87600
reduced air entry on left chest | 0
epigastric tenderness | 0
bowel sounds present | 0
X-ray chest PA view showing hydropneumothorax | 0
CT scan chest showing hydropneumothorax | 0
ultrasonography abdomen 7 days before admission | -168
provisional diagnosis of traumatic hydropneumothorax | 0
intercostal drain tube insertion | 0
seropurulent fluid drainage | 0
gastric contents in drain | 0
nasogastric tube insertion | 0
Ryle's tube in left hydropneumothorax | 0
revised diagnosis as TDH with iatrogenic perforation | 0
surgical repair planned | 0
tachypnoeic (RR 36/min) | 0
SpO2 92% on O2 | 0
heart rate 118/min | 0
BP 130/78 mm Hg | 0
ABG: PaO2 64, PaCO2 39, pH 7.38 | 0
rapid sequence induction | 0
tracheal intubation | 0
IPPV initiated | 0
thoracic epidural catheter placement | 0
bupivacaine administered | 0
diaphragmatic rent (6x5 cm) discovered | 0
stomach and spleen herniated | 0
viscera reduced | 0
tear repaired | 0
fresh ICT inserted | 0
feeding gastrostomy performed | 0
mechanical ventilation in ICU | 0
reduced left chest air entry | 0
chest X-ray showing infiltrates | 0
ABG: PaCO2 58 | 0
pleural fluid culture: enterobacter | 0
ventilator dependency | 0
ABG: PaO2 55, PaCO2 58 | 0
tracheostomy performed | 336
enteral feeds via gastrostomy | 0
minimal ventilatory support | 0
high grade fever | 0
leucocytosis | 0
tachycardia | 0
SIRS | 0
infection controlled | 0
left lung expansion | 0
improved gas exchange | 0
haemodynamic stability | 0
ICT removed | 672
transfer to surgical department | 720
