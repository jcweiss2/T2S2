56 years old | 0
male | 0
admitted to the hospital | 0
chronic left leg ulcer | 0
liver cirrhosis | 0
congestive heart failure | 0
substance use disorder | 0
bacteremia | 0
fever | -72
chills | -72
leg pain | -72
non-healing wound | -72
alcohol use | -72
opioid use | -72
hypertension | -8760
hyperlipidemia | -8760
stroke | -8760
hepatitis C | -8760
heart failure | -8760
polysubstance use | -8760
aspirin | -72
atorvastatin | -72
ferrous sulfate | -72
folic acid | -72
gabapentin | -72
metoprolol | -72
mirtazapine | -72
sacubitril | -72
valsartan | -72
thiamine | -72
methadone | -72
emergency room visit | -336
admission for leg ulcer | -336
blood culture | -336
vancomycin | -336
discharge | -336
readmission | -168
blood culture | -168
no growth | -168
discharge | -168
admission to hospital | 0
fever | 0
chills | 0
leg pain | 0
non-healing wound | 0
alcohol use | 0
opioid use | 0
normocytic anemia | 0
chronic thrombocytopenia | 0
elevated C-reactive protein | 0
normal lactic acid | 0
vancomycin | 0
ampicillin-sulbactam | 0
piperacillin-tazobactam | 0
urology consultation | 0
wound care consultation | 0
orthopedic consultation | 0
blood culture | 0
Empedobacter falsenii | 96
multidrug resistance | 96
urine culture | 96
no growth | 96
swab culture | 96
vancomycin-resistant Enterococcus faecalis | 96
cefepime | 96
fever resolution | 48
discharge | 168
trimethoprim-sulfamethoxazole | 168
follow-up appointment | 720
missed appointment | 720
readmission | 720
cellulitis | 720
urinary tract infection | 720
Klebsiella pneumoniae | 720
levofloxacin | 720
discharge | 720
readmission | 1440
acute hypoxemic respiratory failure | 1440
pneumonia | 1440
septic shock | 1440
encephalopathy | 1440
Klebsiella pneumoniae | 1440
Staphylococcus aureus | 1440