37 years old | 0
    male | 0
    admitted to the hospital | 0
    pain in left hemithorax | -168
    pain in left upper abdomen | -168
    fever | -168
    body temperature of 39.1°C | -168
    severe cough | -168
    purulent greenish sputum | -168
    mild pain in left hypochondrium | -168
    cough | -120
    shortness of breath | -120
    alcohol abuser | -131400
    tobacco smoker | -131400
    periodic upper abdominal pain | -17520
    inability to remain in a prone position due to dyspnea and cough | 0
    increased dyspnea | 0
    increased sputum volume | 0
    blood pressure 140/90 mmHg | 0
    heart rate 98 beats per minute | 0
    temperature 38.2°C | 0
    respiratory rate 23 breaths per minute | 0
    absent breath sound in lower half of left hemithorax | 0
    reduced breath sounds with wheezing under upper half of left hemithorax | 0
    hemoglobin 12.5 g/dL | 0
    white blood cells 16,800/mm³ | 0
    platelets 590,000/mm³ |2
    