44 years old | 0
female | 0
arterial hypertension | 0
dyslipidemia |&nbsp;
obesity | 0
sought the emergency department | -48
acute onset of rapidly progressive erythematous rash | -48
rash emerged on thighs | -48
rash emerged on armpits | -48
rash emerged on inframammary fold | -48
rash progressed to whole body | -48
aspirin | 0
losartan | 0
atorvastatin | 0
application of dexamethasone | -48
used tampons (menstruation) | -72
hypotensive | 0
blood pressure 65/42 mmHg | 0
heart rate 113 bpm | 0
febrile (39.4 °C) | 0
somnolent | 0
morbilliform rash | 0
pustular lesions | 0
diagnosis of septic shock | 0
Sequential Organ Failure Score 8 | 0
considered toxic shock syndrome | 0
considered DRESS | 0
considered AGEP | 0
started on vancomycin | 0
started on piperacillin/tazobactam | 0
started on clindamycin | 0
received norepinephrine | 0
received vasopressin | 0
intravenous fluid resuscitation | 0
leukocytosis | 0
neutrophilia | 0
white blood cell 15.70 × 109/L | 0
acute kidney failure | 0
serum creatinine 2.3 mg/dL | 0
blood urea nitrogen 46 mg/dL | 0
estimated glomerular filtration rate 40.8 mL/min | 0
increased total bilirubin | 0
increased serum transaminases | 0
metabolic acidosis | 0
hyperlactatemia | 0
chest x-ray parahiliar bilateral reticular infiltrates | 0
nasopharyngeal swab RT-PCR positive for SARS-CoV-2 | 0
acute kidney failure worsened | 24
vancomycin discontinued | 24
substituted for daptomycin | 24
elevated creatine phosphokinase | 24
concern on rhabdomyolysis | 24
concern on deep tissue involvement | 24
skin biopsy performed | 24
diffuse spongiosis | 24
intradermic subcorneal micro pustules | 24
neutrophilic content | 24
reactive changes of microvascular endothelium | 24
diagnosis of AGEP | 24
considered toxic shock syndrome | 24
considered DRESS | 24
considered septic shock | 24
considered pustular psoriasis | 24
required vasopressors | 0
required corticosteroids (fludrocortisone and hydrocortisone) | 0
completed 10-day course of antibiotics | 240
local management with hyperoxygenated fatty acids | 0
progressive improvement in haemodynamics | 24
progressive improvement in skin lesions | 24
no longer required vasopressors | 120
extubated | 120
complete recovery of kidney function | 120
complete recovery of liver function | 120
chest CT no typical COVID-19 pneumonia | 120
developed critical polyneuropathy | 120
proximal limb weakness | 120
resolved with physical rehabilitation | 336
discharged | 336
