40 years old | 0
    male | 0
    admitted to the hospital | 0
    sudden chest pain | -5
    back pain | -5
    acute type A aortic dissection | 0
    hypertension | -87600
    heavy smoking | -175200
    creatinine elevation (237.6 mmol/L) | 0
    aortic false lumen formation | 0
    ascending aortic and total aortic arch replacement | 0
    stented elephant trunk implantation | 0
    cardiopulmonary bypass | 0
    transferred to ICU | 0
    red blood cells transfusion (4 U) | 0
    plasma transfusion (850 mL) | 0
    cryoprecipitate transfusion (20 U) | 0
    platelets transfusion (2 U) | 0
    lung protective ventilation | 0
    fluid management | 0
    continuous renal replacement therapy | 0
    airway secretion clearance | 0
    severe ARDS | 0
    oxygenation index (OI) drop to 51 | 0
    prone positioning (PP) | 0
    ECMO consideration | 0
    chest radiography (diffuse exudation of both lungs) | 0
    prone position ventilation | 0
    drain patency assessment every hour | 0
    circulatory changes monitoring | 0
    blood gas analysis | 0
    chest X-ray (reduced diffuse exudation) | 96
    oxygenation index improvement | 96
    acute kidney injury (AKI) grade II | 0
    coagulation dysfunction | 0
    acute myocardial injury | 0
    hypoproteinemia | 0
    high-risk stage 3 hypertension | 0
    PaO2/FiO2 ≤ 100 mmHg with PEEP ≥ 5 cmH2O | 0
    bilateral lung opacities | 0
    hypoxemia | 0
    hypercapnia | 0
    acute cardiac tamponade | 0
    mediastinal pericardial drainage | 0
    thoracic drainage | 0
    sternotomy | 0
    obesity | 0
    prolonged CPB | 0
    ischemic reperfusion injury | 0
    inflammatory mediators release | 0
    ventilator-induced lung injury | 0
    hemodynamic instability | 0
    brachial plexus injury | 0
    facial pressure ulcers | 0
    facial edema | 0
    vascular catheter kinking | 0
    elevated intraabdominal pressure | 0
    acute severe pancreatitis | 0
    pulmonary contusion | 0
    pulmonary embolism | 0
    sepsis | 0
    severe trauma | 0
    burns | 0
    transfusion-related acute lung injury (TRALI) | 0
    fluid overload | 0
    cardiac failure | 0
    bilateral shadows (on CXR or CT scan) | 0
    new/worsening respiratory symptoms | 0
    PaO2/FiO2 ≤ 100 mmHg with PEEP ≥ 5 cmH2O | 0
    acute onset | 0
    lung protective mechanical ventilation | 0
    oxygen therapy | 0
    intubation/mechanical ventilation | 0
    noninvasive ventilation | 0
    central venous pressure < 4 mmHg | 0
    PAOP < 8 mmHg | 0
    antipyretics | 0
    sedatives | 0
    analgesics | 0
    paralysis agents | 0
    inotropics | 0
    inhaled vasodilators | 0
    nitric oxide | 0
    prostacyclin | 0
    prostaglandin E1 | 0
    hemoglobin 7–9 g/dL | 0
    chest and back pain (tearing-like) | 0
    thoracic and abdominal aorta CTA | -5
    acute myocardial injury | 0
    hypoproteinemia | 0
    high-risk stage 3 hypertension | 0
    preoperative examination | 0
    general anesthesia | 0
    postoperative complications | 0
    ICU stay | 0
    ventilator use | 0
    postoperative mortality | 0
    postoperative severe ARDS | 0
    prone position ventilation treatment | 0
    intermittent short-term PP | 0
    improved oxygenation | 0
    reduced mortality rate | 0
    reduced ventilator duration | 0
    reduced ICU length of stay | 0
    improved respiratory mechanics | 0
    increased functional residual volume | 0
    reduced lung shunt | 0
    promoted pulmonary secretion discharge | 0
    improved ventilation flow ratio | 0
    OI upward trend | 0
    drainage tube compression risk | 0
    fatal bleeding risk (ECMO) | 0
    abnormal coagulation function | 0
    individualized treatment plan | 0
    sternotomy contraindication | 0
    PP time ≥ 12 hours | 0
    PP time < 6 hours | 0
    supine position | 0
    assessment of lung condition | 0
    hourly drain patency assessment | 0
    real-time circulatory monitoring | 0
    dynamic blood gas analysis follow-up | 0
    significant reduction in diffuse exudation | 96
    improved OI | 96
    written informed consent | 0
    no competing interests | 0
    CARE Checklist compliance | 0
    single blind peer review | 0
    informed consent statement | 0
    conflict-of-interest statement | 0
    CARE Checklist (2016) statement | 0
    provenance and peer review | 0
    peer-review model | 0
    specialty type | 0
    country/territory of origin | 0
    peer-review report’s scientific quality classification | 0