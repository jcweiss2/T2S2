11 years old | 0
female | 0
admitted to the hospital | 0
high fever | 0
nausea | 0
severe weakness | 0
myalgia | 0
main body ache | 0
conscious | 0
pale | 0
ill | 0
body temperature 39.5 °C | 0
pulse 120 bpm | 0
blood pressure 110/75 mmHg | 0
no rash | 0
no spontaneous bleeding | 0
no jaundice | 0
hemoglobin 14.8 g/dl | 0
hematocrit 40% | 0
platelet count 140000/mm3 | 0
Dengue IgM antibodies positive | 0
SARS-COV2 antigen nasopharynx test negative | 0
clinical diagnosis suspect of Dengue fever | 0
standard diet | 0
feverish | 24
looked ill | 24
short of breath | 24
nausea | 24
abdominal bloating | 24
platelet count 78000/mm3 | 24
platelet count 15000/mm3 | 48
blood pressure 110/90 mmHg | 48
pulse 90 bpm | 48
pleura effusion | 48
pleural effusion index 38.13% | 48
managed in the intensive care unit | 48
sharp acute abdominal pain | 72
abdominal ultrasonography | 72
liver function test elevated | 96
AST 151 IU/L | 96
ALT 59 IU/L | 96
C-reactive protein level 14.4 mg/L | 96
conservative treatment | 96
intravenous antibiotics | 120
abdominal pain lasted for 3 days | 120
abdominal bloating sensation lasted for 3 days | 120
patient's condition improved | 120
discharged from the hospital | 168
liver function enzyme restored | 168
follow-up post-treatment | 168