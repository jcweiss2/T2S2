14 years old | 0
African-American | 0
male | 0
right thigh pain | 0
painful ambulation | 0
no fever | 0
otherwise healthy | 0
no significant past medical history | 0
no trauma | 0
developed pain upon doing butterfly stretches | -24
football conditioning routine | -24
pulling sensation on active and passive movement | 0
full range of motion | 0
mild leukocytosis | 0
14,500/µL white blood cell count | 0
59% polymorphonuclear cells | 0
ESR 10 mm/h | 0
CRP 5.7 mg/dL | 0
CT pelvis with and without contrast | 0
concerning area of pelvic bone | 0
MRI pelvis with contrast | 0
intramuscular tears | 0
edema involving right obturator internus and externus muscles | 0
mild widening of right pubic bone apophysis | 0
edema at superior ramus | 0
thought to have osteitis pubis | 0
discharged | 0
crutches | 0
600 mg ibuprofen | 0
instructions to avoid sports | 0
follow-up with sports medicine in 1 week | 0
readmitted to the hospital | 0
worsening symptoms | 0
abdominal pain | 0
thigh pain | 0
inability to walk | 0
worsening pain in both shoulders | 0
generalized myalgias | 0
malaise | 0
emesis | 0
diarrhea | 0
tachycardia | 0
tachypnea | 0
afebrile | 0
normotensive | 0
limited range of motion at right hip | 0
diffuse tenderness to palpation in all quadrants of abdomen | 0
no distension | 0
no rebound | 0
no focal neurologic deficits | 0
white blood cell count 12,100/µL | 0
ESR 59 mm/h | 0
CRP 20.7 mg/dL | 0
CT abdomen and pelvis with contrast | 0
right obturator internus muscle fluid collection | 0
enhancement at site of muscle tear | 0
empirically given 1 gram ceftriaxone | 0
started on intravenous vancomycin | 0
admitted to intensive care unit | 0
oxacillin added to antibiotic regimen | 0
clindamycin added to antibiotic regimen | 0
blood cultures ordered | 0
urine cultures ordered | 0
urine cultures no growth | 0
blood cultures yielded MSSA | 48
vancomycin discontinued | 48
MRI left shoulder | 48
repeat MRI pelvis | 48
myositis in left shoulder | 48
enlarging fluid mass in right obturator internus muscle | 48
osteomyelitis of right pubic bone | 48
continued on IV oxacillin | 48
continued on IV clindamycin | 48
daily blood cultures positive for three consecutive days | 48
blood cultures negative for 2 days | 120
discontinuation of blood cultures | 120
underwent abscess drainage | 120
placed in prone position | 120
preprocedural CT redemonstrated hypodense region | 120
15-cm One-Step needle advanced into abscess | 120
5 cc cloudy tan-colored fluid collected | 120
sheath extended | 120
guide wire coiled within abscess | 120
sheath removed | 120
entrance route gauge increased | 120
8 French all-purpose drainage catheter inserted | 120
15 cc fluid aspirated | 120
total sedation time 21 minutes | 120
technically successful | 120
no immediate complications | 120
catheter maintained to external bulb suction | 120
no follow-up imaging | 120
febrile until postprocedure day 2 | 168
downward-trending white blood cells | 168
downward-trending ESR | 168
downward-trending CRP | 168
PICC placed | 216
continuation of IV antibiotics at home | 216
Ancef 2 grams every 8 hours for 6 weeks | 216
discharged | 336
denied pain during ambulation | 336
white blood cells 8900/µL | 336
ESR 79 mm/h | 336
scheduled for outpatient follow-up | 336
initial PT assessment | 384
limitation in ROM | 384
limitation in strength | 384
pressure bilaterally at anterior hips | 384
predominantly right sided hip rotation pain | 384
physical therapy for 6 weeks | 384
gradual improvement in ROM | 384
gradual improvement in strength | 384
ESR normalization | 672
CRP normalization | 672
completion of 6 weeks antibiotics | 1176
PICC removed | 1176
denied pain with ambulation | 1176
denied pain climbing stairs | 1176
full ROM | 1176
full strength | 1176
no further follow-up needed | 1176
