47 years old | 0  
    female | 0  
    hypothyroidism | -432  
    Hashimoto’s thyroiditis | -432  
    iron deficiency anemia | -432  
    lymphadenopathy | -432  
    ITP | -432  
    received first dose of Pfizer-BioNTech mRNA vaccine | 0  
    mild arm soreness | 48  
    no other adverse effects | 0  
    ITP diagnosed in 2002 | -432  
    pregnancy | -432  
    platelets decreased to 4000/mcL | -432  
    prednisone treatment | -432  
    complete remission | -432  
    ITP flare-up 6 years later | -432  
    platelets decreased to 3000/mcL | -432  
    IVIG and dexamethasone treatment | -432  
    complete remission | -432  
    direct platelet antibody level 1962 | -432  
    elevated rheumatoid factor 20.7 IU/mL | -432  
    negative ANA | -432  
    negative dsDNA | -432  
    negative anticardiolipin IgM and IgG | -432  
    negative lupus anticoagulant | -432  
    bone marrow biopsy: no lymphoproliferative disorder | -432  
    no increased blasts | -432  
    no clonal blast cells | -432  
    normal karyotype 46XX | -432  
    platelet counts 164000-36000 | -432  
    no maintenance therapy for ITP | -432  
    enlarged left axillary lymph node in 2018 | -432  
    left axillary adenopathy on CT 12/2018 | -432  
    retroperitoneal adenopathy on CT 6/2019 | -432  
    biopsy of left axillary lymph node: no malignancy | -432  
    excisional biopsy 3/2019: follicular hyperplasia | -432  
    flow cytometry negative for lymphocytic malignancy in 2018 | -432  
    fine needle aspirate negative for malignancy in 2019 | -432  
    presented to ER 18 days postvaccination | 432  
    easy bruising | 432  
    gum bleeding | 432  
    epistaxis | 432  
    denied trauma | 432  
    denied headache | 432  
    denied visual changes | 432  
    denied rectal bleeding | 432  
    denied gastrointestinal symptoms | 432  
    ecchymosis | 432  
    petechiae | 432  
    dried blood in oropharynx | 432  
    no splenomegaly | 432  
    no hepatomegaly | 432  
    CT head: negative for hemorrhage | 432  
    chest radiograph clear | 432  
    platelet count 1000/mcL | 432  
    previous platelet count 62000/mcL | 432  
    peripheral smear confirmed thrombocytopenia | 432  
    normal RBC morphology | 432  
    prothrombin time 16.2 seconds | 432  
    INR 1.5 | 432  
    reticulocyte count 2.2% | 432  
    LDH 310 U/L | 432  
    manual WBC differential: 13 atypical lymphocytes | 432  
    elevated alkaline phosphatase 109 U/L | 432  
    ANA negative | 432  
    normal WBC count and differential | 432  
    normal hemoglobin | 432  
    normal RDW | 432  
    normal aPPT | 432  
    normal haptoglobin | 432  
    normal basic metabolic panel | 432  
    negative SARS-CoV-2 test | 432  
    negative flu A and B | 432  
    fibrinogen 280 | 432  
    denied headaches | 432  
    received dexamethasone | 432  
    admitted to ICU | 432  
    platelet transfusion | 432  
    IVIG (Privigen) | 432  
    platelets improved to 61000/mcL | 432  
    platelets fell to 19000/mcL | 432  
    second platelet transfusion | 432  
    second IVIG | 432  
    platelets rose to 72000/mcL | 432  
    CT chest, abdomen, pelvis: resolution of adenopathy | 432  
    Sjogren’s SS-A antibody (RO) 2.8 AI | 432  
    repeat ANA positive 1:80 | 432  
    EBV DNA PCR positive 429 IU/mL | 432  
    negative hepatitis C | 432  
    negative hepatitis B | 432  
    negative HIV | 432  
    negative thyroid-stimulating hormone | 432  
    discharged | 432  
    received only first dose of vaccine | 432  

<|eot_id|>
