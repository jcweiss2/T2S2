65 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
no history of smoking | 0 | 0 | Factual
no underlying pulmonary diseases | 0 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
shortness of breath | -96 | 0 | Factual
fever | -96 | 0 | Factual
dry cough | -96 | 0 | Factual
fatigue | -96 | 0 | Factual
breath sounds reduced | 0 | 0 | Factual
oxygen saturation 93% | 0 | 0 | Factual
bilateral peripheral ground-glass attenuation | 0 | 0 | Factual
patchy consolidation | 0 | 0 | Factual
lung involvement 60%-70% | 0 | 0 | Factual
nasopharyngeal SARS-CoV-2 RT-PCR test positive | 0 | 0 | Factual
symptoms worsened | 0 | 504 | Factual
increased temperature | 0 | 504 | Factual
saturation with free breathing decreased | 0 | 504 | Factual
white cell count 7.93 х 109/ L | 0 | 504 | Factual
hemoglobin 159 g/l | 0 | 504 | Factual
platelet count 468 х 109/l | 0 | 504 | Factual
Westergren ESR 41 mm/h | 0 | 504 | Factual
interleukine 6 102 pg/ml | 0 | 504 | Factual
С-reactive protein 142 mg/l | 0 | 504 | Factual
ferritin 939.92 μg/ml | 0 | 504 | Factual
D-dimer 609 ng/ml | 0 | 504 | Factual
procalcitonin 0,11 ng/ml | 0 | 504 | Factual
treatment with dexamethason | 0 | 504 | Factual
treatment with heparin | 0 | 504 | Factual
treatment with tocilizumab | 0 | 504 | Factual
treatment with acetylcysteine | 0 | 504 | Factual
treatment with pantoprazole | 0 | 504 | Factual
treatment with nadroparin calcium | 0 | 504 | Factual
oxygen supplementation | 0 | 504 | Factual
air and pleural effusion in the right pleural cavity | 360 | 360 | Factual
collapse of the right lung | 360 | 360 | Factual
thoracentesis | 360 | 360 | Factual
thoracostomy | 360 | 360 | Factual
1400 ml of yellowish opaque liquid evacuated | 360 | 360 | Factual
linezolid therapy | 360 | 504 | Factual
imipenem/cilastatin therapy | 360 | 504 | Factual
oxygen supplementation with flow rate 8-10 l/min | 360 | 504 | Factual
daily drainage volume 300-1000 ml | 360 | 504 | Factual
pleural effusion with gas bubbles | 432 | 432 | Factual
focal area of subpleural infiltration | 432 | 432 | Factual
central cavity of destruction | 432 | 432 | Factual
air layer up to 47 mm | 432 | 432 | Factual
left side hydropneumothorax | 432 | 432 | Factual
pleural fluid analysis | 432 | 432 | Factual
exudative lymphocytic-rich effusion | 432 | 432 | Factual
Acinetobacter baumannii | 432 | 432 | Factual
Pseudomonas aeruginosa | 432 | 432 | Factual
Klebsiella pneumonia | 432 | 432 | Factual
needle thoracocentesis | 504 | 504 | Factual
new pleural drainage | 504 | 504 | Factual
air and creamy purulent mass aspirated | 504 | 504 | Factual
serofibrinous hemorrhagic fluid drawn | 504 | 504 | Factual
pleural empyema | 504 | 504 | Factual
transfer to the Surgical Department | 504 | 504 | Factual
right pleural space irrigated with antiseptic solutions | 504 | 1008 | Factual
lung expansion by continuous vacuum aspiration | 504 | 1008 | Factual
encapsulated pleural effusion | 736 | 736 | Factual
ultrasound-guided puncture | 736 | 736 | Factual
new drainage of the pleural cavity | 736 | 736 | Factual
antibiotic therapy | 504 | 1008 | Factual
colistimethatum natrium | 504 | 1008 | Factual
imipenem/cilastatin | 504 | 1008 | Factual
discharged from the hospital | 1008 | 1008 | Factual
oxygen saturation 97% | 1008 | 1008 | Factual
small amount of fluid in the right pleural cavity | 1008 | 1008 | Factual
lab test scores normal | 1008 | 1008 | Factual
С-reactive protein 11.7 mg/l | 1008 | 1008 | Factual
procalcitonin < 0,1 ng/ml | 1008 | 1008 | Factual