44 years old | 0  
    male | 0  
    admitted to the hospital | 0  
    progressive left facial necrosis | -240  
    blurred vision of the left eye | -240  
    left periorbital pain | -240  
    swelling | -240  
    fever | -240  
    general malaise | -240  
    crepitus | 0  
    fluctuation | 0  
    local heat over entire face and scalp | 0  
    decayed left upper second molar | -336  
    self-extracted left upper second molar | -336  
    intermittent sharp pain | -672  
    poor oral hygiene | -672  
    loss of appetite | -672  
    hyperglycemic (576 mg/dL plasma glucose) | 0  
    diffuse subcutaneous emphysematous changes of the neck and left upper thorax | 0  
    bilateral facial, periorbital, and scalp regions involvement | 0  
    leukocytosis (44400/uL) | 0  
    high CRP level (335 mg/L) | 0  
    metabolic acidosis (pH = 7.277, pCO2 = 12.8 mmHg) |# hello-world
just another repository
I am a student
