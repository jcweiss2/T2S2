Here is the table of events and timestamps:

18 years old | 0
male | 0
history of primary refractory acute myeloblastic leukemia | -1095
multiple relapses | -1095
allogeneic bone marrow transplant from cord blood | -27
delayed engraftment | -27
prolonged severe neutropenia | -27
vancomycin-resistant Enterococcus | -27
Streptococcus viridans | -27
Streptococcus mitis | -27
tedizolid | -27
cefepime | -27
Flagyl | -27
daptomycin | -27
filgrastim | 0
acyclovir | 0
Bactrim | 0
caspofungin | 0
fever | 0
tachycardia | 0
hypotension | 0
tachypnea | 0
distended abdomen | 0
localized peritonitis | 0
white cell count 0.2 x 10^9 /L | 0
absolute neutrophil count (ANC) of zero | 0
anemic | 0
hemoglobin of 7 g/L | 0
thrombocytopenic | 0
platelet count of 10 x 10^9 /L | 0
lactic acid of 3.1 mmol/L | 0
CT scan | 0
segmental ischemia of the small bowel | 0
fever to 38.2°C | 0
explore the operating room for an exploratory laparotomy | 0
15 cm ischemic bowel segment | 0
50 cm of small bowel resection | 0
primary anastomosis | 0
norepinephrine and vasopressin for blood pressure support | 0
transesophageal echo | 0
admitted to the intensive care unit | 0
pressors were weaned | 0
extubated | 0
transferred to the floor | 0
diet advanced on postoperative day (POD) 3 | 72
passed flatus | 72
new fevers | 96
increased abdominal pain | 96
lactic acidosis | 96
respiratory decompensation | 96
amphotericin B (AmBisome) started | 96
repeat CT scan | 96
area of necrotic small bowel remote from the initial anastomosis | 96
invasive fungal forms in both the omental and small intestinal resection specimens | 96
invasive fungal forms in both the omental and small intestinal resection specimens, invading through blood vessel walls, with associated hemorrhage and transmural ischemic necrosis, consistent with mucormycosis | 96
died | 120