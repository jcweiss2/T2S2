62 years old | 0
male | 0
diabetes mellitus | 0
hypertension | 0
fever | -48
dyspnea | -48
productive cough | -48
yellow purulent sputum | -48
smoked 20 cigarettes a day for approximately 40 years | 0
visited a hot spring | -240
no history of immunosuppression | 0
no history of recurrent infection | 0
no history of chemotherapy | 0
no history of steroid use | 0
blood pressure 118/60 mmHg | 0
heart rate 130 beats/min | 0
respiratory rate 28/min | 0
percutaneous oxygen saturation 95% | 0
body temperature 37.5℃ | 0
holoinspiratory coarse crackles in the right lung | 0
high anion gap metabolic acidosis | 0
increased lactate | 0
leukopenia | 0
thrombocytopenia | 0
renal dysfunction | 0
elevated transaminase | 0
infiltration of the right upper and middle lobes | 0
consolidation with air bronchogram in the right upper and middle lobes | 0
admitted to hospital | 0
consulted infectious disease specialist | 0
Gram-negative cocci and coccobacilli on sputum Gram staining | 0
initiated treatment with meropenem | 0
administered azithromycin | 0
intubated | 12
noradrenaline administered | 12
recuperated from shock | 24
respiratory condition gradually improved | 24
A. baumannii identified in sputum culture | 72
changed antibiotic regimen from meropenem to ampicillin/sulbactam | 72
extubated | 96
set up for nasal high-flow therapy | 96
transferred out of intensive care unit | 168
Serratia marcescens identified from sputum culture | 288
diagnosed HAP | 288
changed ampicillin/sulbactam to cefepime | 288
treated with intravenous antibiotics for 42 days | 1008
treated with oral ciprofloxacin for 14 days | 1008