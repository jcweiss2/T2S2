71 years old | 0
female | 0
hypertension | -720
dyspnea on exertion | 0
malaise | -2160
anorexia | -2160
fatigue | -2160
progressive unintentional weight loss | -2160
atrial fibrillation | 0
heart failure | 0
admission to hospital | 0
abdominal and pelvic ultrasound | 0
bilateral adnexal masses | 0
solid and cystic changes | 0
abdominal CT scan | 0
solid peritoneal deposits | 0
moderate to large volume ascites | 0
ovarian malignancy | 0
CA-125 level | 0
discharge from hospital | 120
outpatient clinic visit | 120
paracentesis | 120
malignant cells | 120
poorly differentiated carcinoma or sarcoma | 120
epithelioid morphology | 120
planned chemotherapy | 120
Paclitaxel | 131
Carboplatin | 131
interval debulking | 131
first dose of chemotherapy | 131
no allopurinol for TLS prophylaxis | 131
re-admission to hospital | 135
diarrhea | 135
fatigue | 135
generalized weakness | 135
afebrile | 135
clinically dehydrated | 135
blood work | 135
CBC | 135
Leukocytes | 135
Neutrophils | 135
Lymphocytes | 135
Monocytes | 135
Hemoglobin | 135
Platelets | 135
Potassium | 135
Phosphate | 135
Calcium | 135
Albumin | 135
BUN | 135
Creatinine | 135
Uric acid | 135
LDH | 135
temperature | 135
irregular heart rate | 135
blood pressure | 135
oxygen saturation | 135
respiratory rate | 135
volume resuscitation | 135
hypotension | 135
pre-renal acute kidney injury | 135
pancytopenic | 135
PRBC | 135
GCSF | 135
prophylactic antibiotics | 135
diagnosis of tumour lysis syndrome | 135
uric acid level | 135
Cairo-Bishop criteria | 135
Rasburicase | 135
maintenance dose | 135
ICU stay | 139
intubation | 139
progressive hypoxic respiratory failure | 139
volume overload | 139
vasopressor support | 139
septic shock | 139
CRRT | 139
blood cultures | 139
Group B streptococcus | 139
urine | 139
E. coli | 139
broad spectrum antibiotic therapy | 139
piperacillin-tazobactam | 139
fungemia | 143
clinical deterioration | 143
comfort care | 143
life support withdrawn | 143
death | 143
autopsy | 143
intramural uterine malignant neoplasm | 143
extensive necrosis | 143
undifferentiated endometrial stromal sarcoma | 143
metastatic involvement | 143
omentum | 143
bowel | 143
gastric mucosa | 143
pancreas | 143
kidneys | 143
marked autolytic changes | 143
granular casts | 143
proximal distal tubules | 143