57 years old | 0
female | 0
diabetes | -116 months
vitamin D deficiency | -116 months
CML in AP | -116 months
hepatosplenomegaly | -116 months
spleen size 25-cm | -116 months
liver size 22-cm | -116 months
imatinib treatment | -116 months
imatinib dose increased to 600 mg/day | -38 months
intolerant to imatinib | -38 months
pallor | -24 months
hepatosplenomegaly | -24 months
hemoglobin concentration 7 g/dL | -24 months
platelet count 194 000/μL | -24 months
WBC count 26 000/μL | -24 months
basophils 0% | -24 months
eosinophils 1% | -24 months
blasts 10% | -24 months
referred to tertiary care hospital | -24 months
BM test | -20 months
hypercellular BM | -20 months
blasts 11% | -20 months
CD45 positive | -20 months
CD34 positive | -20 months
CD33 positive | -20 months
CD117 positive | -20 months
CD56 negative | -20 months
karyotype 47,XX,+7,t(9,22)(q34,q11.2) | -20 months
FISH analysis | -20 months
BCR/ABL fusion signals 5% | -20 months
switched to dasatinib | 0
dasatinib 100 mg/day | 0
minimal interruption of treatment | 0
GCSF | 0
blood product transfusions | 0
shortness of breath | 3 months
lung infiltrates | 3 months
abdominal pain | 3 months
CT scan | 3 months
mild hepatosplenomegaly | 3 months
portal venous hypertension | 3 months
splenic lesion | 3 months
no lymphadenopathy | 3 months
complete cytogenetic remission | 6 months
disappearance of Philadelphia chromosome | 6 months
trisomy 7 | 6 months
FISH negative | 6 months
molecular analysis | 6 months
BCRABL p210 not detectable | 6 months
JAK-2 V617F mutation negative | 6 months
first isolated CNS relapse | 6 months
severe headache | 6 months
nausea | 6 months
generalized tonic-clonic seizures | 6 months
brain MRI | 6 months
abnormal signal intensity | 6 months
leptomeningeal infiltration | 6 months
CSF examination | 6 months
WBCs 130/μL | 6 months
blasts 51% | 6 months
immature cells | 6 months
flow cytometry | 6 months
myeloblasts 43% | 6 months
CD34 positive | 6 months
CD117 positive | 6 months
CD33 positive | 6 months
HLA-DR negative | 6 months
CD3 negative | 6 months
CD13 negative | 6 months
treated with dasatinib and TIT chemotherapy | 6 months
CSF clear | 11 months
refused further TIT chemotherapies | 11 months
refused allo-SCT | 11 months
second isolated CNS relapse | 14 months
severe headache | 14 months
brain MRI | 14 months
interval improvement | 14 months
new leukemic infiltrations | 14 months
CSF | 14 months
blast population 52% | 14 months
CD34 positive | 14 months
CD117 positive | 14 months
CD33 positive | 14 months
CD13 positive | 14 months
CD7 positive | 14 months
treated with whole-brain radiation therapy | 14 months
dasatinib 100 mg/day | 14 months
deep molecular remission | 14 months
hepatosplenomegaly | 24 months
CT scan | 24 months
spleen size 18 cm | 24 months
BM biopsy | 26 months
BM cellularity 50% | 26 months
trilineage hematopoiesis | 26 months
blasts <1% | 26 months
cytogenetic analysis normal | 26 months
karyotype 46,XX | 26 months
hypothyroidism | 38 months
levothyroxine | 38 months
minimal pleural effusion | 38 months
diuretics | 38 months
GCSF support | 38 months
dasatinib decreased to 70 mg/day | 38 months
dasatinib increased to 100 mg/day | 46 months
dasatinib halted | 52 months
diarrhea | 52 months
edema | 52 months
PegINF-α2a | 52 months
hepatosplenomegaly resolved | 52 months
PegINF-α2a discontinued | 64 months
spleen growth | 64 months
joint pains | 64 months
minimal left-sided pleural effusion | 64 months
chronic diarrhea | 64 months
lupus anticoagulant positive | 64 months
anticardiolipin IgG and IgM antibodies positive | 64 months
B2GP1 positive | 64 months
anti-dsDNA antibodies positive | 64 months
refused prophylactic anticoagulation | 64 months
referred to rheumatology department | 64 months
compliance/logistic issues | 64 months
ultrasonography | 70 months
spleen size 17.1 cm | 70 months
CML therapy on hold | 70 months
deep molecular remission | 70 months
BCR-ABL transcripts undetectable | 70 months
bloody diarrhea | 90 months
endoscopic biopsy | 90 months
adenocarcinoma of the rectum | 90 months
invasion of the uterus | 90 months
septic shock | 96 months
admitted to intensive care unit | 96 months
CT imaging | 96 months
splenic infarct | 96 months
massive ascites | 96 months
omental thickening | 96 months
peritoneal deposits | 96 months
adnexal mass | 96 months
rectal mass | 96 months
infiltration into the anal canal | 96 months
surrounding soft tissue | 96 months
bilateral inguinal lymph nodes | 96 months
pulmonary embolism | 96 months
bilateral pulmonary nodules | 96 months
palliative supportive care | 96 months
died | 96 months