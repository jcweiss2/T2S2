68 years old | 0
male | 0
admitted to the hospital | 0
chest pain | -72
acute dyspnea | -72
type 2 diabetes mellitus | 0
hypertension | 0
oral metformin hydrochloride | 0
valsartan | 0
hemoglobin A1c of 7.7% | 0
history of similar diseases in close relatives denied | 0
heart sounds normal | 0
coarse crackles in both lungs | 0
no other abnormalities detected | 0
white blood cell count high | 0
C-reactive protein levels high | 0
myocardial enzymes lactate dehydrogenase elevated | 0
aspartate aminotransferase elevated | 0
troponin-T positive | 0
anti-HIV antibody test negative | 0
chest radiography consolidation in right upper lobe | 0
bilateral congestion | 0
cardiac infarction | 0
bacterial pneumonia | 0
percutaneous coronary intervention | 0
admitted to intensive care unit | 0
oxygen saturation 92% | 0
respiratory rate 30 breaths/min | 0
intubated | 0
invasive mechanical ventilation | 0
progressive respiratory failure | 0
intravenous antibiotics | 0
levofloxacin 500 mg daily | 0
ampicillin/sulbactam 9 g daily | 0
vasodilators | 0
diuretics | 0
fraction of inspired oxygen 80% | 0
positive end expiratory pressure 15 cmH2O | 0
diagnosed with ARDS | 120
extracorporeal membrane oxygenation | 120
intravenous methylprednisolone 1 g daily | 120
prednisolone 60 mg daily | 192
respiratory condition improved by day eight | 192
blood in stool | 192
dual antiplatelet therapy | 192
discontinued extracorporeal membrane oxygenation | 240
extubated | 288
prednisolone tapered to 40 mg daily | 408
respiratory condition worsened | 408
re-intubated | 432
intravenous methylprednisolone 1 g daily | 432
prednisolone reduced to 100 mg daily | 504
prednisolone tapered to 80 mg daily | 672
prednisolone tapered to 60 mg daily | 1008
bloody diarrhea started | 192
bloody diarrhea progressively worsened | 192
colonoscopy on day 22 | 528
multiple large ulcers in sigmoid colon and rectum | 528
biopsy of sigmoid colon ulcer | 528
histopathological examination showed infiltration of neutrophils and lymphocytes | 528
CMV-positive cells in mucosa | 528
CMV pp65 antigenemia test positive | 528
diagnosed with CMV enterocolitis | 528
ganciclovir started | 600
peripheral blood C7-HRP test results improved | 600
continued bloody diarrhea | 600
abdominal pain increased | 1080
abdominal computed tomography revealed free air | 1080
gastrointestinal perforation | 1080
died | 1104
autopsy performed | 1104
full-thickness necrotic intestinal wall tissue | 1104
infiltration of necrotic tissue with ameba | 1104
CMV-positive cells in colon | 1104
Entamoeba histolytica trophozoites detected | 1104
fulminant amebic colitis posthumous diagnosis | 1104
CMV enterocolitis posthumous diagnosis | 1104
68 years old|0
male|0
admitted to the hospital|0
chest pain|-72
acute dyspnea|-72
type 2 diabetes mellitus|0
hypertension|0
oral metformin hydrochloride|0
valsartan|0
hemoglobin A1c of 7.7%|0
history of similar diseases in close relatives denied|0
heart sounds normal|0
coarse crackles in both lungs|0
no other abnormalities detected|0
white blood cell count high|0
C-reactive protein levels high|0
myocardial enzymes lactate dehydrogenase elevated|0
aspartate aminotransferase elevated|0
troponin-T positive|0
anti-HIV antibody test negative|0
chest radiography consolidation in right upper lobe|0
bilateral congestion|0
cardiac infarction|0
bacterial pneumonia|0
percutaneous coronary intervention|0
admitted to intensive care unit|0
oxygen saturation 92%|0
respiratory rate 30 breaths/min|0
intubated|0
invasive mechanical ventilation|0
progressive respiratory failure|0
intravenous antibiotics|0
levofloxacin 500 mg daily|0
ampicillin/sulbactam 9 g daily|0
vasodilators|0
diuretics|0
fraction of inspired oxygen 80%|0
positive end expiratory pressure 15 cmH2O|0
diagnosed with ARDS|120
extracorporeal membrane oxygenation|120
intravenous methylprednisolone 1 g daily|120
prednisolone 60 mg daily|192
respiratory condition improved by day eight|192
blood in stool|192
dual antiplatelet therapy|192
discontinued extracorporeal membrane oxygenation|240
extubated|288
prednisolone tapered to 40 mg daily|408
respiratory condition worsened|408
re-intubated|432
intravenous methylprednisolone 1 g daily|432
prednisolone reduced to 100 mg daily|504
prednisolone tapered to 80 mg daily|672
prednisolone tapered to 60 mg daily|1008
bloody diarrhea started|192
bloody diarrhea progressively worsened|192
colonoscopy on day 22|528
multiple large ulcers in sigmoid colon and rectum|528
biopsy of sigmoid colon ulcer|528
histopathological examination showed infiltration of neutrophils and lymphocytes|528
CMV-positive cells in mucosa|528
CMV pp65 antigenemia test positive|528
diagnosed with CMV enterocolitis|528
ganciclovir started|600
peripheral blood C7-HRP test results improved|600
continued bloody diarrhea|600
abdominal pain increased|1080
abdominal computed tomography revealed free air|1080
gastrointestinal perforation|1080
died|1104
autopsy performed|1104
full-thickness necrotic intestinal wall tissue|1104
infiltration of necrotic tissue with ameba|1104
CMV-positive cells in colon|1104
Entamoeba histolytica trophozoites detected|1104
fulminant amebic colitis posthumous diagnosis|1104
CMV enterocolitis posthumous diagnosis|1104
