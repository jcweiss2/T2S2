67 years old | 0
male | 0
admitted because of dyspnea and rapid atrial fibrillation | 0
coronary heart disease | 0
atrial fibrillation | 0
heart failure | 0
diuretics | 0
milrinone | 0
nitrate | 0
radiofrequency catheter ablation | -72
wide area circumferential ablations | -72
pulmonary vein isolation | -72
discharged from the hospital | 72
chest discomfort | 432
fever | 432
confusion | 432
gazing upwards | 432
mild limb seizures | 432
vomiting | 432
temperature of 41°C | 432
WBC 5.2 × 10⁹/L | 432
hsCRP 18.56 mg/L | 432
supraventricular tachycardia | 432
hypothermia therapy | 432
temperature of 37.9°C | 432
blood pressure 99/73 mm Hg | 432
pulse rate 78 beats/min | 432
AF on ECG | 432
NT-proBNP 1550.00 pg/mL | 432
alanine aminotransferase 21 U/L | 432
cardiac troponin I 3.95 μg/L | 432
WBC 10.58 × 10⁹/L | 432
neutrophil 97.2% | 432
hsCRP 26.0 mg/L | 432
fecal occult blood 3+ | 432
cerebral CT no abnormal findings | 432
pulmonary CT no abnormal findings | 432
CECT suspicious thrombus in left atrial appendage | 432
fasting | 432
gastrointestinal decompression | 432
antibiotic | 432
imipenem/cilastatin | 432
linezolid | 432
regained consciousness | 456
repeated epileptic seizures | 456
cerebral MRI lacuna infarctions | 456
emergency EGD small deep ulcer at 30 cm | 456
esophageal stent implanted | 456
WBC counts decreased | 480
hsCRP decreased | 480
epileptic seizures resolved | 480
acid reflux | 552
fluid food intake | 552
temperature increased | 624
WBC counts increased | 624
cardiac CECT esophageal-mediastinum fistula | 624
encapsulated effusion | 624
pneumatosis behind left atrium | 624
posterior wall of LA depression | 624
mediastinal abscess | 624
atrial-esophageal fistula | 624
surgical repair planned | 624
right thoracotomy incision | 624
membranaceous adhesions | 624
funicular adhesions | 624
white lamellar scars under azygos vein | 624
tight adhesion between esophagus and pericardium | 624
separated carefully | 624
6 mm diameter fistula in anterior wall of esophagus | 624
tight adhesion between LA and pericardium | 624
bleeding at posterior wall of LA | 624
rid-muscle flap repair | 624
pleuroclysis with povidone iodine and saline | 624
transferred to ICU | 624
sepsis | 624
infectious shock | 624
fever | 624
chills | 624
metabolic acidosis | 624
hypotension | 624
tachycardia | 624
oliguria | 624
death | 624
