53 years old | 0
male | 0
presented to emergency department | 0
fever | -192
dry cough | -192
myalgia | -192
progressive shortness of breath | -72
vomiting | -24
nonspecific epigastric discomfort | -24
denied chest pain | 0
no history of recent travel | 0
no contact with suspected or confirmed COVID-19 patients | 0
Type-2 diabetes mellitus | 0
hypertension | 0
inferior MI in 2015 | -144480
refused coronary angiography in 2015 | -144480
severe distress | 0
tachypneic (32/min) | 0
tachycardiac (130 bpm) | 0
normotensive | 0
O2 saturation 93% on CPAP with 100% FIO2 | 0
normal body temperature | 0
severely breathless | 24
hypoxic (SpO2 88%) | 24
crackles in both lung fields | 24
normal cardiac examination | 24
1 mm ST elevation at lead V3 | 24
severe left ventricular systolic dysfunction | 24
left ventricular ejection fraction 35% | 24
segmental wall motion abnormalities | 24
bilateral patchy consolidative changes | 24
air space opacities | 24
intubated | 24
mechanical ventilation for ARDS secondary to pneumonia | 24
mechanical ventilation for acute heart failure | 24
treated as acute heart failure | 24
treated as community-acquired pneumonia | 24
treated as possible ACS | 24
intravenous nitrates | 24
diuretics | 24
antibiotics | 24
oral aspirin 300 mg | 24
clopidogrel 600 mg | 24
enoxaparin 60 mg | 24
noradrenaline 0.5 mcg/kg/min | 24
nasopharyngeal swab PCR positive for CoV-2 | 24
leukocytes 12.8 × 103/uL | 24
lymphocytes 0.5 | 24
C-reactive protein 150 mg/L | 24
ferritin 1979 ug/L | 24
troponin-T high sensitive 527 ng/L | 24
N-terminal-proB-type natriuretic peptide 722 pg/mL | 24
lactic acid 7.2 mmol/L | 24
admitted to COVID9-19 intensive care unit | 24
serial ECG biphasic T wave in V2, V3 | 24
inverted T waves in V4–V6 | 24
peak cTn 1806 at 24 hours | 48
good response to medical therapy | 48
less oxygen requirement | 48
severely agitated | 72
hypotension | 72
severe bradycardia | 72
asystole | 72
return of spontaneous circulation | 72
worsening lactic acidosis | 72
pH 6.8 | 72
lactate 19 mmol/L | 72
oxygen saturation 60% on 100% FIO2 | 72
diffuse ST depression | 72
ST elevation in lead aVR | 72
coronary angiography 6 hours after cardiac arrest | 78
tight stenosis of mid-LAD | 78
normal flow in LAD | 78
tight ostial stenosis of obtuse marginal branch | 78
totally occluded mid-right coronary artery | 78
everolimus-eluting stent deployed at LAD | 78
no attempt to stent other lesions | 78
ECG changes improved after PCI | 78
severe sepsis with bilateral pneumonia | 96
mechanical ventilation | 96
noradrenaline till June 20 | 96
weaned from mechanical ventilation | 240
weaned from vasopressors | 240
clarithromycin | 96
piperacillin/tazobactam | 96
ceftriaxone | 96
lopinavir/ritonavir | 96
favipiravir | 96
plasma protein fraction | 96
hydroxychloroquine | 96
acute kidney injury | 240
acute liver injury | 240
complete recovery of renal function | 264
complete recovery of liver function | 264
normalized inflammatory markers | 264
discharged | 576
