40 years old | 0
    male | 0
    admitted as a trauma alert | 0
    gunshot wound to the upper abdomen | 0
    gunshot wound to the chest | 0
    arrived with Glasgow coma score of 15 | 0
    hemodynamically stable | 0
    focused assessment with sonography positive | 0
    taken emergently to the operating room | 0
    emergent exploratory laparotomy | 0
    repair of ballistic gastric serosal tear | 0
    diagnostic pericardial window | 0
    complex hepatotrhaphy | 0
    liver debridement with argon beam coagulation | 0
    liver packing | 0
    repair of the diaphragm | 0
    right chest tube placement | 0
    multiple ballistic perforations injured the diaphragm | 0
    multiple ballistic perforations injured the liver | 0
    multiple ballistic perforations injured the gastric serosa | 0
    identified tissue damage repaired | 0
    bleeding surgically controlled | 0
    estimated blood loss 1,300 mL | 0
    transferred to the intensive care unit | 0
    still intubated | 0
    5 cm H2O positive end expiratory pressure | 0
    sedated | 0
    plans to return to the OR the following day for closure of the abdomen | 0
    transfused one unit of A+ packed red blood cells | 0
    initial hemoglobin on admission 12.9 g/dL | 0
    spiked a fever | 0.5
    developed hematuria | 0.5
    became hypotensive | 0.5
    received a unit of A+ blood by mistake due to clerical error | 0.5
    stabilized with intravenous hydrocortisone 100 mg | 0.5
    intravenous diphenhydramine 50 mg | 0.5
    intramuscular epinephrine 1:1,000, 0.3 mL | 0.5
    labs returned | 0.5
    clinical deterioration became evident | 0.5
    given multiple liter IV fluid boluses without improvement | 0.5
    direct Coombs test positive | 0.5
    haptoglobin < 5.8 mg/dL | 0.5
    lactate dehydrogenase 1,193 U/L | 0.5
    hemolytic reaction | 0.5
    coagulation parameters worsening | 0.5
    hypotension required norepinephrine drip | 0.5
    preoperative creatinine normal at 1.5 mg/dL | 0
    determined to be having an AHTR | 0.5
    employ an urgent RBCET | 4.5
    RBCET started approximately 4.5 hours after mismatched transfusion | 4.5
    RBCET consisted of five units of type O negative blood for a target hemoglobin goal of 9.0 g/dL | 4.5
    over the next 2 days received five units of fresh frozen plasma | 24
    over the next 2 days received two units of PRBC | 24
    over the next 2 days received one unit of platelets | 24
    creatinine peaked at 2.12 mg/dL 17 hours after mismatched transfusion | 17
    direct Coombs returned negative 9 hours after RBCET | 13.5
    norepinephrine discontinued on day 2 | 48
    clinical and lab parameters stabilized over next 4 days | 96
    required no blood products after day 2 | 48
    hospital course prolonged due to surgical interventions to the abdomen | 0
    discharged in stable condition | 144
    no apparent long-term consequences from the transfusion or exchange | 144
    <|eot_id|>
    