46 years old | 0
female | 0
elective sleeve gastrectomy | 0
obesity | -8760
psoriatic arthritis | -8760
surgical hypoparathyroidism | -8760
hypothyroidism | -8760
total thyroidectomy | -8760
multinodular goitre | -8760
oral calcium carbonate | -8760
calcitriol | -8760
planned sleeve gastrectomy | -4
converted to emergency Roux-en-Y gastric bypass surgery | -4
gastric perforations | -4
friable mucosa | -4
abdominal sepsis | -4
transfer to intensive care | 0
critically low calcium level | 0
ionised calcium 0.78 mmol/L | 0
continuous intravenous calcium gluconate infusion | 0
normocalcaemia | 0
maintenance intermittent IV calcium boluses | 0
prolonged ICU admission | 0
abdominal operations | 0
intravenously medication and nutrition | 0
lost 14 kg | 0
Endocrinology advice | 0
manage hypoparathyroidism | 0
manage hypothyroidism | 0
ionised calcium 1.04 mmol/L | 18
TSH 5.83 mU/L | 14
intravenous triiodothyronine | 14
euthyroidism | 14
high dose intravenous calcium | 42
ionised calcium measured daily | 42
serum phosphate level 1.07 mmol/L | 42
intravenous calcitriol | 42
ceased intravenous calcitriol | 47
intramuscular cholecalciferol | 56
low 1,25(OH)vitamin D3 level | 56
normal renal function | 56
eGFR > 90 mL/min/1.73 m2 | 56
still required intravenous calcium gluconate | 84
additional intravenous calcitriol | 84
reduced calcium gluconate requirements | 84
intramuscular thyroxine | 90
intravenous thyroxine | 94
maintenance schedule | 94
controlled hypocalcaemia | 94
controlled hypothyroidism | 94
recovered sufficiently | 672
recommence oral intake | 672
discharged | 672
normocalcaemia on review | 672
normocalcaemia on review | 840
normocalcaemia on review | 1344
weight 71.8 kg | 1344
BMI 29 kg/m2 | 1344