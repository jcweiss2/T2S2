39 years old | 0
    male | 0
    diabetes mellitus | -24
    dyslipidemia | -24
    oral hypoglycemic agents | -24
    epigastric abdominal pain | -24
    nausea | -24
    vomiting | -24
    elevated white cell count | 0
    hyponatremia | 0
    hyperglycemia | 0
    lactic acidosis | 0
    creatinine elevated | 0
    lipase elevated | 0
    triglyceride elevated | 0
    denied binge drinking | 0
    denied abdominal trauma | 0
    denied recent change in medications | 0
    denied recent procedures | 0
    computed tomography diffuse pancreatitis | 0
    abdominal ultrasound hepatic steatosis | 0
    admitted to intensive care unit | 0
    intravenous fluid resuscitation | 0
    electrolyte management | 0
    intravenous insulin drip | 0
    tachypnea | 72
    altered mental status | 72
    worsening acidosis | 72
    intubated | 72
    respiratory failure | 72
    insulin infusion | 72
    triglycerides remained elevated | 72
    abdominal distension | 72
    oliguria | 72
    renal failure | 72
    creatinine elevated | 72
    plasmapheresis initiated | 48
    plasmapheresis triglycerides improved | 72
    hemodialysis initiated | 96
    bladder pressure serial monitoring | 96
    elevated bladder pressures | 120
    peak airway pressures elevated | 120
    cisatracurium | 120
    decompressive laparotomy | 120
    serous ascitic fluid drained | 120
    saponification noted | 120
    postoperative sepsis | 120
    postoperative delirium | 120
    stabilized | 120
    downgraded to medical floor | 120
    renal function improved | 120
    hemodialysis stopped | 120
    discharged | 120
    icosapent ethyl | 0
    omega 3 fatty acids | 0
    fenofibrate added | 120

    