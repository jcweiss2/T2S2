45 years old | 0  
    woman | 0  
    end-stage heart failure | 0  
    cardiac cirrhosis | 0  
    valvular heart disease | -720  
    New York Heart Association class IV | -720  
    mild jaundice | -720  
    mitral valve replacement | -720  
    tricuspid annuloplasty | -720  
    ischemic kidney injury | -672  
    continuous renal replacement therapy (CRRT) | -672  
    cardiac arrest | -624  
    ventricular fibrillation | -624  
    venoarterial extracorporeal membrane oxygenation (ECMO) | -624  
    admission to our institution | 0  
    severe biventricular dysfunction | 0  
    left ventricular ejection fraction < 5% | 0  
    ECMO conversion to central ECMO | 0  
    ECMO flow rate 3.6–4.1 L/min | 0  
    heparinization for ACT 160–180 s | 0  
    CRRT continued | 0  
    norepinephrine infusion (0.03 µg/kg/min) | 0  
    mean arterial pressure 50–60 mmHg | 0  
    progressive hyperbilirubinemia | 0  
    hepatic fissure widening | 0  
    irregular hepatic contours | 0  
    heterogeneous parenchymal enhancement | 0  
    splenomegaly | 0  
    moderate ascites | 0  
    dilated inferior vena cava | 0  
    congestive hepatopathy | 0  
    tracheostomy | 0  
    remifentanil sedation (0.03 µg/kg/min) | 0  
    atrial fibrillation | 0  
    ventricular response 76 bpm | 0  
    cardiomegaly | 0  
    left lung atelectasis | 0  
    left main bronchus compression | 0  
    total bilirubin 47.3 mg/dl | 0  
    direct bilirubin 36.2 mg/dl | 0  
    aspartate transaminase 92 units/L | 0  
    alanine transaminase 51 units/L | 0  
    creatinine 0.91 mg/dl | 0  
    platelet count 34,000 /µl | 0  
    PT INR 1.49 | 0  
    Child-Pugh class C | 0  
    MELD score 26 | 0  
    emergent CHLT scheduled | 0  
    general anesthesia induced | 0  
    midazolam 2 mg | 0  
    etomidate 8 mg | 0  
    atracurium 50 mg | 0  
    desflurane maintenance | 0  
    mechanical ventilation pressure controlled | 0  
    peak airway pressure 20 cmH2O | 0  
    intra@-arterial monitoring | 0  
    central venous pressure monitoring | 0  
    inferior vena cava pressure monitoring | 0  
    pulmonary arterial pressure monitoring | 0  
    Swan-Ganz catheter | 0  
    right femoral artery catheter | 0  
    right femoral vein catheter | 0  
    9-Fr Advanced Venous Access catheter | 0  
    transesophageal echocardiography probe | 0  
    heart transplant planned | 0  
    liver transplant planned | 0  
    histidine-tryptophan-ketoglutarate solution | 0  
    re-sternotomy | 0  
    left femoral vessel cannulation | 0  
    superior vena cava cannulation | 0  
    CPB established | 0  
    heparin 100 mg | 0  
    modified bicaval technique | 0  
    temporary pacemaker inserted | 0  
    heart rate 90 bpm | 0  
    CPB time 148 min | 0  
    transfused 11 units LDRBC | 0  
    transfused 2 units FFP | 0  
    converted to peripheral ECMO | 0  
    protamine sulfate 100 mg | 0  
    ACT 163 s | 0  
    chest left open | 0  
    liver transplantation initiated | 0  
    subcostal incision | 0  
    liver mobilization | 0  
    substantial hemorrhage | 0  
    massive volume resuscitation | 0  
    bleeding control required | 0  
    piggyback technique | 0  
    anhepatic stage | 0  
    transfused LDRBC targeting Hb 10 g/dl | 0  
    transfused FFP for PT INR >3 | 0  
    transfused platelets for count <50,000 /µl | 0  
    potassium >4.5 mEq/L managed | 0  
    insulin 10 IU | 0  
    5% dextrose 200 ml | 0  
    metabolic acidosis corrected | 0  
    half saline 1 L | 0  
    sodium bicarbonate 80 mEq/L | 0  
    calcium chloride 300 mg | 0  
    glucose control post-reperfusion | 0  
    insulin per Portland protocol | 0  
    reperfusion syndrome 3 min | 0  
    epinephrine 100 µg | 0  
    tranexamic acid 500 mg | 0  
    protamine 50 mg | 0  
    ACT 215 s | 0  
    closure of abdominal incision | 0  
    residual bleeding control | 0  
    sternum closure | 0  
    crystalloid 13,600 ml | 0  
    5% albumin 1,250 ml | 0  
    half saline 3,800 ml | 0  
    LDRBC 32 units | 0  
    cell saver blood 5,500 ml | 0  
    FFP 11 units | 0  
    platelets 4 units | 0  
    cryoprecipitate 5 units | 0  
    no urine output | 0  
    red cell mass loss 7,500 ml | 0  
    postoperative creatinine 0.7 mg/dl | 0  
    dobutamine 5 µg/kg/min | 0  
    norepinephrine 0.05 µg/kg/min | 0  
    vasopressin 0.05 units/min | 0  
    epinephrine 0.05 µg/kg/min | 0  
    transferred to ICU on ECMO | 0  
    anesthesia time 13h15min | 0  
    POD 1 | 24  
    ischemic right hand | 24  
    thromboembolectomy right radial artery | 24  
    thromboembolectomy right brachial artery | 24  
    uncertain Allen's test | 24  
    vasopressor contributing to ischemia | 24  
    ECMO removed on POD 4 | 96  
    norepinephrine 0.1 µg/kg/min | 96  
    norepinephrine tapered over 1 month | 720  
    transaminase normalization | 504  
    prothrombin time normalization | 504  
    bilirubin normalization | 504  
    type II respiratory failure | 24  
    mechanical ventilation >1 month | 720  
    oliguric acute kidney injury | 24  
    CRRT continued | 24  
    improved renal function | 504  
    transition to hemodialysis | 1080  
    hemodialysis discontinued | 1080  
    defective wound healing | 504  
    antibiotic treatment | 504  
    surgical revision | 504  
    transudative ascites | 1440  
    right pleural effusion | 1440  
    daily drainage | 1440  
    abdominal CT findings | 1440  
    chronic liver disease signs | 1440  
    mild periportal edema | 1440  
    septic shock due to catheter infection | 1440  
    normal left ventricular function | 1440  
    reduced right ventricular function | 1440  
    pericardial effusion | 1440  
    discharged at 5 months | 3600  
    stable condition | 3600  
    no allograft rejection | 3600  

