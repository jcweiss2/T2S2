18 years old | 0
female | 0
history of autoimmune hepatitis | 0
unprotected sexual intercourse | -14
fever | 0
chills | 0
nausea | 0
dizziness | 0
heavy menorrhasia | 0
jaundice | 0
scleral icterus | 0
abdominal ascites | 0
anasarca | 0
erythematous vaginal vault | 0
lactic acidosis | 0
creatinine | 0
aspartate transaminase | 0
alanine transaminase | 0
total bilirubin | 0
alkaline phosphatase | 0
total protein | 0
albumin | 0
hemoglobin | 0
leukocytes | 0
platelets | 0
prothrombin time | 0
international normalized ratio | 0
beta-human chorionic gonadotropin test | 0
schistocytes | 0
leukocyte count | 0
neutrophilic predominance | 0
cirrhosis | 0
portal hypertension | 0
splenomegaly | 0
generalized edematous wall thickening of the colon and rectum | 0
intubation | 0
intravenous fluids | 0
blood products | 0
vasopressors | 0
vancomycin | 0
piperacillin-tazobactam | 0
doxycycline | 0
clindamycin | 0
intravenous immunoglobulin | 0
non-blanching ecchymoses | -16
flaccid bullae | -16
dusky violaceous ecchymoses | -36
hemorrhagic bullae | -36
lactate dehydrogenase | -36
fibrinogen | -36
D-dimer | -36
urinalysis | -36
salicylate level | -36
acetaminophen level | -36
Chlamydia trachomatis | -36
Neisseria gonorrhea | -36
urine toxicology screen | -36
peritoneal fluid culture | -36
blood culture | -36
pan-susceptible Streptococcus pneumoniae | -36
progressive hypoxia | -48
shock | -48
death | -48
autopsy | -48
cirrhotic liver | -48
diffuse alveolar damage | -48
abdominal compartment | -48
acute-onset excruciating bilateral lower extremity pain | 0
excruiciating pain | 0
edema | 0
ascites | 0
excruiciating pain persisted | 0
fever persisted | 0
chills persisted | 0
nausea persisted | 0
dizziness persisted | 0
heavy menorrhasia persisted | 0
jaundice persisted | 0
scleral icterus persisted | 0
abdominal ascites persisted | 0
anasarca persisted | 0
erythematous vaginal vault persisted | 0
lactic acidosis persisted | 0
creatinine persisted | 0
aspartate transaminase persisted | 0
alanine transaminase persisted | 0
total bilirubin persisted | 0
alkaline phosphatase persisted | 0
total protein persisted | 0
albumin persisted | 0
hemoglobin persisted | 0
leukocytes persisted | 0
platelets persisted | 0
prothrombin time persisted | 0
international normalized ratio persisted | 0
beta-human chorionic gonadotropin test persisted | 0
schistocytes persisted | 0
leukocyte count persisted | 0
neutrophilic predominance persisted | 0
cirrhosis persisted | 0
portal hypertension persisted | 0
splenomegaly persisted | 0
generalized edematous wall thickening of the colon and rectum persisted | 0
intubation persisted | 0
intravenous fluids persisted | 0
blood products persisted | 0
vasopressors persisted | 0
vancomycin persisted | 0
piperacillin-tazobactam persisted | 0
doxycycline persisted | 0
clindamycin persisted | 0
intravenous immunoglobulin persisted | 0
non-blanching ecchymoses persisted | 0
flaccid bullae persisted | 0
dusky violaceous ecchymoses persisted | 0
hemorrhagic bullae persisted | 0
lactate dehydrogenase persisted | 0
fibrinogen persisted | 0
D-dimer persisted | 0
urinalysis persisted | 0
salicylate level persisted | 0
acetaminophen level persisted | 0
Chlamydia trachomatis persisted | 0
Neisseria gonorrhea persisted | 0
urine toxicology screen persisted | 0
peritoneal fluid culture persisted | 0
blood culture persisted | 0
pan-susceptible Streptococcus pneumoniae persisted | 0
progressive hypoxia persisted | 0
shock persisted | 0
death persisted | 0
autopsy persisted | 0
cirrhotic liver persisted | 0
diffuse alveolar damage persisted | 0
abdominal compartment persisted | 0
pneumococcal vaccination | -4
influenza vaccination | -4
COVID-19 vaccination | -4
acute infectious PF | -36
fulminant S. pneumoniae sepsis | -36
PF | -36