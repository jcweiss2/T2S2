32 years old| 0
    man| 0
    classic Pyoderma gangrenosum|  -43800
    cough|  -96
    sputum|  -96
    dyspnea|  -96
    admitted to the Intensive Care Unit| 0
    received methylprednisolone pulses|  -168
    current medication oral prednisolone| 0
    current medication cyclosporine| 0
    current medication surgical wound therapy| 0
    diagnosis of Pyoderma gangrenosum confirmed by biopsy|  -43800
    respiratory rate 30 breaths/min| 0
    temperature 39°C| 0
    heart rate 150 beats/min| 0
    oxygen saturation below 90%| 0
    large and deeply diffuse necrotic skin lesions on upper limbs| 0
    large and deeply diffuse necrotic skin lesions over chest and back| 0
    dermatology examination skin lesions observed| 0
    initial lung examination unremarkable| 0
    initial heart examination unremarkable| 0
    white blood cell count 9.8 × 10^9/l| 0
    neutrophils 79%| 0
    lymphocytes 22%| 0
    monocytes 3%| 0
    eosinophil 1%| 0
    platelets 25 × 10^9/L| 0
    transthoracic echocardiogram no vegetation| 0
    CT scan of lungs multiple 1-2 cm nodules| 0
    CT scan halo sign| 0
    CT scan air-crescent signs| 0
    CT scan small size left pleural effusion| 0
    respiratory failure developed| 48
    intubated| 48
    mechanically ventilated| 48
    bronchoscopy performed| 48
    bronchoalveolar lavage specimen obtained| 48
    diagnosis of probable invasive pulmonary aspergillosis| 48
    direct microscopy examination endobronchial washing| 48
    direct microscopy examination BAL samples acute branching septate hyphae| 48
    culture of samples Aspergillus flavus| 48
    diagnosis of cutaneous fusariosis| 0
    Fusarium proliferatum isolated from skin lesion biopsy| 0
    polymerase chain reaction assays performed with BAL sample| 0
    polymerase chain reaction assays performed with tissue biopsy| 0
    fungal ITS region of rRNA gene amplified| 0
    fungal ITS region of rRNA gene sequenced| 0
    ITS sequences A. flavus submitted to NCBI GenBank| 0
    ITS sequences F. proliferatum submitted to NCBI GenBank| 0
    voriconazole administered| 0
    linezolid administered| 0
    meropenem administered| 0
    ciprofloxacin administered| 0
    dose adjusted based on creatinine clearance| 0
    treatment failed| 0
    expired| 288
