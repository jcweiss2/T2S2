69 years old | 0
male | 0
resides in southern Saudi Arabia | 0
works as a farmer | 0
uncontrolled type II diabetes | -8760
laparoscopic cholecystectomy | -8760
admitted to the emergency department | 0
left lower abdomen pain | -336
intermittent fever | -8760
weight loss | -8760
paraumbilical and left lower quadrant tenderness | 0
distension | 0
no organomegaly | 0
leucocytosis | 0
neutrophilia | 0
eosinophilia | 0
Haemoglobin of 126 g/L | 0
Platelets of 518 * 10^9/L | 0
C-reactive protein 262.48 mg/L | 0
abdominal x-ray showed faecal impaction | 0
nonspecific distribution of bowel gases | 0
no air under diaphragm | 0
no signs of bowel obstruction | 0
CT abdomen and pelvis with contrast showed multifocal segmental wall thickening | 0
fluid collections suggesting concealed perforations | 0
diagnosis of severe diverticulitis | 0
Piperacillin/Tazobactam | 0
maintained nothing by mouth | 0
symptoms worsened | 96
blood-stained stool | 96
CT abdomen and pelvis with contrast repeated | 96
recurrence of multifocal segmental wall thickening | 96
evidence of concealed perforation | 96
interval increase in size of surrounding collections | 96
Infectious diseases team involved | 96
surgical intervention recommended | 96
biopsy for bacterial, TB, fungal cultures, and histopathology | 96
empiric start of liposomal amphotericin B | 96
Amoxicillin/Clavulanic acid | 96
tigecycline | 96
patient condition worsened | 192
persistently febrile | 192
white blood cells increased | 192
absolute eosinophils count increased | 192
haemoglobin dropped | 192
third abdominal CT with contrast | 192
redemonstration of circumferential wall thickening of the colon | 192
interval increase in size of fluid collection | 192
interval increase in abdominopelvic ascites | 192
surrounding inflammatory changes | 192
operation | 216
faecal peritonitis | 216
multiple colon perforation | 216
small bowel adhesion | 216
adhesions between small bowel and transverse colon | 216
adhesolysis | 216
total colectomy | 216
end ileostomy | 216
placement of two drains | 216
transferred to intensive care unit (ICU) | 216
absolute eosinophils count dropped | 216
haemoglobin dropped | 240
inotropic support | 240
transfused several units of packed red blood cells | 240
minimal ventilator settings | 240
minimal respiratory secretions | 240
abdominal and pelvic CT repeated | 240
no collection found | 240
bacterial tissue culture showed heavy growth of Pseudomonas aeruginosa | 240
carbapenem resistant Klebsiella variicola | 240
blood culture from the central line showed Bacteroides fragilis | 240
fungal tissue culture showed Candida glabrata | 240
histopathology showed extensive inflammation | 240
mixed inflammatory cells | 240
sheets of eosinophils | 240
multiple foci of fungal microorganism | 240
hyphae that are irregularly branched | 240
thin walled | 240
occasionally septated | 240
surrounded by thick eosinophilic cuff | 240
Splendore-Hoeppli phenomenon | 240
patient’s condition deteriorated | 264
passed away | 264
refractory septic shock | 264
Basidiobolus ranarum | 0
Gastrointestinal Basidiobolomycosis (GIB) | 0
subcutaneous infection | 0
infection after a scratch or puncture | 0
infection after ingestion of soil | 0
infection after ingestion of animal feces | 0
infection after ingestion of food contaminated with Basidiobolus ranarum | 0
diffuse erythematous or maculopapular eruption | 0
pruritus | 0
DRESS syndrome | 0 
Note: The time stamps are approximate and based on the information provided in the case report. The time stamps are calculated based on the day of admission being day 0.