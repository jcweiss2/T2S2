845-gram male | 0
24 weeks' gestation | 0
born by emergent cesarean section | 0
limp | 0
blue | 0
without cry | 0
Apgar scores were 1 at 1 min | 0
Apgar scores were 6 at 10 min | 10
intubation | 0
admitted to the neonatal intensive care unit (NICU) | 0
passed meconium on the first day of life | 24
normal physical exam | 24
feeding intolerance | 312
lethargy | 312
moderate abdominal distention | 312
sepsis workup initiated | 312
leukocytosis of 41,500/μL | 312
thrombocytopenia | 312
Candida albicans fungemia | 312
intra-abdominal fluid | 312
inferior right hepatic lobe abscess | 312
abdominal X-rays | 312
paracentesis | 312
brown feculent fluid | 312
pediatric surgery consulted | 312
intestinal perforation suspected | 312
grade III necrotizing enterocolitis | 312
exploratory laparotomy | 312
feculent spillage | 312
necrosed colon identified | 312
cecal perforation | 312
necrosis of the ascending and proximal transverse colon | 312
small bowel examined | 312
liver examined | 312
subhepatic abscess opened and evacuated | 312
right hemicolectomy | 312
end ileostomy with mucus fistula created | 312
abdominal distention | 336
increased oxygen requirement | 336
persistent acidosis | 336
additional exploratory laparotomy | 336
intraabdominal abscess evacuated | 336
peritoneal drain placed | 336
Candida albicans and coagulase negative Staphylococci cultured | 336
pseudohyphae on Hematoxylin and Eosin (H&E) staining | 336
pseudohyphae on Grocott's Methenamine Silver (GMS) staining | 336
antifungals administered | 312
antifungals continued for 10 weeks | 744
fungemia resolved | 744
ostomy takedown | 744
discharged home | 744
good status | 744
tolerating enteral feeds | 744
vaginal candidiasis during pregnancy | 0
bacterial vaginosis during pregnancy | 0
clinical chorioamnionitis | 0
tachycardia | 0
intermittent maternal fevers | 0
Candida albicans colonization | -672
vertical transmission of fungal candida | -672 
systemic candidiasis | 312 
intraabdominal fungal abscess | 336 
intestinal candidiasis | 312 
pathologic intestinal candidiasis | 312 
mucosal invasion with Candida Albicans | 312 
fungal sepsis | 312 
successful surgical outcome | 744 
probiotic administration | 0 
colostrum administration | 0 
necrotizing enterocolitis | 312 
Hirschprung's disease | 0 
mechanical bowel obstruction | 0 
idiopathic causes | 0 
intestinal perforation | 312 
peritonitis | 312 
portal venous air | 0 
respiratory complications | 312 
oxygen demand | 312 
microbiological infection | 312 
paracentesis | 312 
surgical intervention | 312 
laparotomy | 312 
peritoneal drainage | 312 
necrotic tissue removal | 312 
sepsis control | 312 
post-surgical complications reduction | 312 
bowel length preservation | 312 
informed consent | 0 
ethical approval | 0 
authorship | 0 
funding | 0 
registration of research studies | 0 
guarantor | 0 
declaration of competing interest | 0