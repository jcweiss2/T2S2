57 years old | 0
male | 0
admitted to hospital | 0
acute abdomen | 0
nausea | 0
vomiting | 0
incarcerated incisional hernia | 0
body mass index 38.3 kg/m2 | 0
elevated white cell count | 0
elevated CRP | 0
elevated interleukins | 0
elevated creatinine | 0
elevated urea | 0
amiodarone | -672
pantoprazole | -672
bisoprolol | -672
eplerenone | -672
sacubitril/valsartan | -672
eliquis | -672
l-thyroxin | -672
dilated cardiomyopathy | -672
atrial fibrillation | -672
left atrial thrombus | -672
implantable cardioverter defibrillator | -672
radioiodine therapy | -672
prior laparoscopic appendectomy | -672
perforated appendicitis | -672
peritonitis | -672
emergency laparotomy | 0
ischaemic segment of ileum | 0
resection of ischaemic ileal segment | 0
end-to-end ileo-ileostomy | 0
sepsis | 0
cardiopulmonary instability | 0
intensive care | 0
discharged home | 264
resected ileum histology | 0
haemorrhagic mucosa | 0
mural necrosis | 0
well-differentiated NET | 0
immunohistochemistry | 0
CK AE 1/3 positive | 0
synaptophysin positive | 0
chromogranin positive | 0
CD56 positive | 0
grade 1 NET | 0
Ki67 < 1% | 0
mitotic activity 1 mitosis/10 HPF | 0
pT2m | 0
pN0 | 0
pL0 | 0
pV0 | 0
tumour-free resection margins | 0
six-week post-surgery | 504
NET-specific workup | 504
computed tomography | 504
no evidence of neuroendocrine disease | 504
Gallium-68 DOTATATE PET/CT | 504
no increased DOTA-D-Phe1-Tyr3-Thr8-octreotide avidity | 504
plasma chromogranin A elevated | 504
5-hydroxyindole acetic acid normal | 504
denies symptoms associated with carcinoid syndrome | 504
repeat laparotomy | 672
palpation of small bowel | 672
resection of 70 cm of ileum | 672
end-to-end ileo-ileostomy | 672
280 cm of unaffected small intestine | 672
histology | 672
well-differentiated NET | 672
chromogranin positive | 672
synaptophysin positive | 672
somatostatin receptor subtype 2A positive | 672
Ki67 < 2% | 672
pT1m | 672
pN1 | 672
pL0 | 672
pV0 | 672
tumour-free resection margins | 672
9 months follow-up | 1944
alive | 1944
no evidence of disease | 1944