70 years old | 0
male | 0
Nigerian | 0
immigrated to the USA | -8760
controlled hypertension | -8760
insulin-dependent diabetes mellitus | -8760
hyperlipidemia | -8760
sickle cell trait | -8760
statin therapy | -8760
discontinued statin therapy | -672
progressive bilateral upper- and lower-extremity weakness | -216
difficulty rising from a sitting position | -216
fatigue | -216
subjective weight loss | -216
decreased appetite | -216
denies skin changes | -216
denies previous trauma | -216
denies sick contacts | -216
denies recent immobilization/hospitalization | -216
denies dysphagia | -216
denies discoloration of urine | -216
3/5 strength in all 4 extremities | 0
no fever | 0
no rash | 0
no tenderness | 0
no swelling | 0
elevated liver enzymes | 0
elevated CPK | 0
eosinophilia | 0
Hgb 10 g/dl | 0
MCV of 95 fl | 0
autoimmune necrotizing myopathy | 0
methotrexate | 0
prednisone | 0
intravenous immunoglobulin | 0
discharged | 216
lethargy | 216
inability to speak | 216
inability to follow commands | 216
dry cough | 216
fever | 216
diarrhea | 216
deterioration in overall condition | 216
febrile patient | 216
tachypnea | 216
tachycardia | 216
crackles | 216
reduced breath sounds | 216
oral thrush | 216
leukopenia | 216
elevated CPK | 216
ABG showed pH 7.57 | 216
lactic acid | 216
bilateral infiltrates | 216
broad-spectrum antibiotics | 216
severely hypoxic | 240
cardiopulmonary arrest | 240
intubated | 240
hypoxic respiratory failure | 240
severe acidosis | 240
return of spontaneous circulation | 240
bilateral worsening of lower lobe infiltrates | 240
acute respiratory distress syndrome | 240
BAL | 240
BAL specimen culture positive for Strongyloides stercoralis | 240
serology testing for Strongyloides negative | 240
HIV testing negative | 240
stool sample negative for Strongyloides | 240
stool sample positive for Strongyloides | 264
Ivermectin | 264
Albendazole | 264
blood cultures positive for Klebsiella pneumoniae | 264
died | 504