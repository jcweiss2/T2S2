29 years old | 0
female | 0
admitted to the hospital | 0
vomiting | -96
general malaise | -96
atypical chest pain | -96
epigastric pain | -96
polyuria | -720
polydipsia | -720
mild eczema | -720
3 pack-year smoking history | -720
normotensive | 0
blood pressure 141/100 mmHg | 0
sinus tachycardia | 0
heart rate 127 b.p.m. | 0
low temperature | 0
temperature 34.6°C | 0
oxygen saturation 98% | 0
respiratory rate 22 breaths/min | 0
severe high anion gap metabolic acidosis | 0
arterial pH 6.87 | 0
hyperglycaemia | 0
plasma glucose 31.6 mmol/L | 0
capillary ketones 4.6 mmol/L | 0
bicarbonate 2.9 mmol/L | 0
PO2 11.7 kPa | 0
PCO2 1.5 kPa | 0
normal CXR | 0
sinus tachycardia on ECG | 0
no evidence of acute coronary syndrome | 0
hypokalaemia | 0
white cell count 33.09 × 10^9/L | 0
neutrophils 28.43 × 10^9/L | 0
CRP 13.9 mg/L | 0
normal plasma sodium | 0
normal serum creatinine | 0
diagnosed with new-onset type 1 DM | 0
diagnosed with severe DKA | 0
treatment for DKA | 0
potassium replacement | 0
fixed rate insulin infusion | 0
volume expansion with crystalloids | 0
empiric treatment with intravenous amoxicillin/clavulanic acid | 0
desaturated to 88% on room air | 12
commenced on supplemental oxygen | 12
ABG on 3 L of oxygen | 12
PaO2 6.4 kPa | 12
PCO2 2.3 kPa | 12
pH 7.24 | 12
bicarbonate 7.5 mmol | 12
type 1 respiratory failure | 24
bilateral infiltrates on CXR | 24
ARDS-like picture | 24
intubated and ventilated | 24
FiO2 100% | 24
peak end expiratory pressure 15 cm H2O | 24
noradrenaline 40 µg/min | 24
vasopressin 2.4 units/h | 24
lung protective ventilation | 24
venous-venous ECMO | 24
Continuous Veno-Venous Hemofiltration (CVVH) | 24
troponin level rose | 48
peri-myocarditis | 48
reduced ejection fraction 45% | 48
discontinued ECMO | 96
extubated | 168
maintained PaO2 16.7 kPa on FiO2 30% | 168
ejection fraction 50-55% | 240
insulin infusion discontinued | 192
commenced on basal/bolus regimen of subcutaneous insulin | 192
discharged to the endocrine ward | 264
discharged home | 384
HbA1c 58 mmol/mol | 384
strongly positive GAD antibodies | 384
normal cardiac function | 384
troponin <14 ng/L | 384
no shortness of breath | 384
clear chest examination | 384
oxygen saturations 99% on room air | 384