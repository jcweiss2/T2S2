72 years old | 0
Hispanic | 0
female | 0
admitted to the hospital | 0
cirrhosis | -672
autoimmune hepatitis | -672
hepatic encephalopathy | -672
ascites | -672
bilious vomiting | -48
diffuse abdominal pain | -48
oliguria | -48
headache | -48
esophagogastroduodenoscopy | -48
gastritis | -48
grade IV esophageal varices | -48
nadolol | 0
spironolactone | 0
furosemide | 0
azathioprine | 0
esomeprazole | 0
lactulose | 0
temperature of 36.06°C | 0
blood pressure of 82/32 mm Hg | 0
regular pulse of 92 beats/min | 0
lethargy | 0
bibasilar rales | 0
tender abdomen | 0
tense ascites | 0
no jaundice | 0
no lower extremity edema | 0
no focal neurological deficits | 0
white blood count of 9,400 cells/mm3 | 0
bandemia | 0
macrocytic anemia | 0
thrombocytopenia | 0
hemoglobin of 9.6 g/dl | 0
hematocrit of 28.5% | 0
platelets of 116,000/μl | 0
MCV of 115.9 fl | 0
INR of 1.98 | 0
prothrombin time of 16 s | 0
new-onset renal failure | 0
creatinine 5 mg/dl | 0
metabolic acidosis | 0
pH 7.39 | 0
HCO3 13.4 | 0
PCO2 22.8 | 0
PO2 77.8 | 0
lactic acid 6.7 mmol/l | 0
serum ammonia 16 μmol/l | 0
sodium 128 meq/l | 0
potassium 5 meq/l | 0
chloride 101 meq/l | 0
bicarbonate 13 meq/l | 0
BUN 70 mg/dl | 0
abdominal CT scan | 0
cirrhotic liver | 0
splenomegaly | 0
ascites | 0
no ruptured viscus | 0
no obstruction | 0
large volume paracentesis | 0
2 l of serosanguinous ascitic fluid | 0
albumin concentration in the fluid <1 mg/dl | 0
serum albumin 2.6 mg/dl | 0
serum-ascites albumin gradient >1.1 | 0
total white and red cell counts in the ascitic fluid 2,889/mm3 and 20,111/mm3 | 0
urine studies suggestive of prerenal cause | 0
renal function did not improve with aggressive volume resuscitation | 0
urine sodium less than 10 meq/l | 0
both kidneys structurally normal on ultrasound | 0
hepatorenal syndrome | 0
midodrine | 0
octreotide | 0
vancomycin | 0
ceftriaxone | 0
ampicillin-sulbactam | 48
gentamicin | 48
deteriorated clinically | 48
transferred to the intensive care unit | 48
respiratory failure | 48
mechanical ventilation | 48
multiple generalized tonic-clonic seizures | 48
lumbar tap not performed | 48
worsening coagulopathy | 48
comfort measures instituted | 48
died | 96
Listeria sepsis | 96
multi-organ failure | 96