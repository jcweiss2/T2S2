10 years old | 0
male | 0
kidney transplantation | -1680
end-stage kidney disease | -1680
chronic interstitial nephritis | -1680
PU valves | -11520
vesico:ureteric reflux | -11520
resection of PU valves | -8640
bilateral ureteric reimplantation | -8640
growth retardation | -11520
underweight | -11520
mother kidney donation | -1680
kidney transplantation on March 8, 2021 | -1680
no induction therapy | -1680
triple immunosuppression | -1680
serum creatinine 0.5 mg/dL | -1680
prophylaxis for pneumocystis | -1680
prophylaxis for cytomegalovirus | -1680
tacrolimus trough level 8 ng/mL | -1680
tacrolimus dose 1.5 mg twice daily | -1680
prednisolone 5 mg daily | -1680
mycophenolate sodium 180 mg twice daily | -1680
regular follow-up | -1680
linear growth 2 cm | -1680
weight gain 4 kg | -1680
high fever | -48
severe cough | -48
vomiting | -48
no loss of smell | -48
no loss of taste | -48
no diarrhea | -48
normal urine output | -48
family members asymptomatic | -48
weight 22.5 kg | 0
temperature 101°F | 0
respiration 26 per min | 0
pulse 120/min | 0
blood pressure 120/80 mm Hg | 0
SpO2 92% | 0
throat normal | 0
chest clear on auscultation | 0
graft kidney non:tender | 0
rapid antigen test positive | 0
nasopharyngeal swab sent for SARS:CoV:2 RT:PCR | 0
HRCT chest CORADS:6 | 0
TSS 18/25 | 0
admitted to hospital | 0
urinalysis normal | 0
Hb 11.3 g/dL | 0
absolute lymphocyte count 820 cells/mm3 | 0
serum creatinine 0.5 mg/dL | 0
serum glutamic:pyruvic transaminase 48 U/L | 0
CRP 9.3 mg/L | 0
ferritin 203 ng/mL | 0
LDH 403 U/L | 0
procalcitonin 0.11 ng/mL | 0
D:dimer 201 ng/mL | 0
ultrasound scan of graft kidney normal | 0
doppler study of graft kidney normal | 0
blood cultures sent | 0
throat swab cultures sent | 0
tacrolimus trough levels analyzed | 0
qt:PCR for CMV analyzed | 0
qt:PCR for BK virus analyzed | 0
hydration given | 0
antipyretics given | 0
piperacillin:tazobactam started | 0
tacrolimus continued 1.5 mg twice daily | 0
prednisolone continued 5 mg daily | 0
mycophenolate stopped | 0
remdesivir loading dose 5 mg/kg | 24
remdesivir 2.5 mg/kg daily for 4 days | 24
afebrile by sixth day | 144
mild cough continued | 144
oxygen saturations normal | 144
urine output normal | 144
creatinine stable 0.5 mg/dL | 144
liver functions normal | 144
PCR for CMV negative | 144
PCR for BK virus negative | 144
blood cultures sterile | 144
throat swab cultures sterile | 144
tacrolimus level 8 ng/mL | 144
discharged | 192
home:quarantine advised | 192
telehealth follow:up continued | 192
asymptomatic on fifteenth day | 360
renal functions normal | 360
lymphocyte count normal | 360
CRP normal | 360
HRCT chest TSS 3/25 | 360
mycophenolate sodium restarted 180 mg daily | 360
telehealth follow:up continued | 360
father tested positive | 360
mother tested negative | 360
elder sibling tested negative | 360
