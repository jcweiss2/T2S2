admitted to the emergency room for abdominal pain | 0
admitted to the emergency room for ketoacidosis decompensation | 0
admitted to the emergency room for uremic syndrome | 0
conscious patient | 0
hemodynamically stable | 0
dyspneic | 0
febrile at 39,6 °C | 0
right lumbar tenderness | 0
oliguric with diuresis at 300 ml/24h | 0
altered renal function with creatinine at 92 mg/l | 0
urea at 3,1 g/l | 0
K+ at 6.9 mmol/l | 0
Na + at 123 mmol/l | 0
blood sugar at 6.5 g/l | 0
alkaline reserves at 8 mEq/l | 0
infectious syndrome with CRP at 418 mg/l | 0
white blood cells at 26000/ml | 0
hemoglobin at 12,3 g/dl | 0
leucocyturia 320,000 | 0
hematuria at 120,000 | 0
emphysematous pyelonephritis | 0
renal abscess ruptured in the intraperitoneal cavity | 0
pneumoperitoneum | 0
admitted to intensive care | 2
dialysis sessions | 2
insulin therapy | 2
antibiotic therapy based on ceftriaxone plus metronidazole | 2
surgical drainage of abscesses | 48
rise of a right double J stent | 48
decrease of the infectious syndrome | 72
apyrexia | 72
chronic renal failure | 120
discharged on day 10 | 240
on oral antibiotics | 240
abdominopelvic CT showed a clear regression of the bubbles of air | 672
double J catheter was removed | 1008
operated for treatment of right inguinal hernia | -7200
type 1 diabetic | 0 
hypertensive on amlodipine | 0 
no shortness of breath | -1 
denies chest pain | -1 
no visible obstacle | 0 
urinary tract infection due to Pseudomonas Aeruginosa | 48 
ECBU culture | 48 
normal diuresis | 120 
creatinine plateau of 20 mg/l | 120 
follow-up | 672 
abdominopelvic CT | 672 
CT scan control | 672 
septic shock | -5.8 
febrile low back pain | -5.8 
bubbly gas pattern | 0 
gas in the collecting system | 0 
gas in the renal parenchyma | 0 
gas or abscess to the perinephric space | 0 
gas or abscess to the pararenal space | 0 
bilateral EPN | 0 
solitary kidney with EPN | 0 
percutaneous drainage failure | 0 
nephrectomy | 0 
broad-spectrum antibiotic therapy | 2 
surgical treatment | 48 
conservative treatment | 2 
medical intensive care | 2 
urgent percutaneous | 48 
surgical or endoscopic drainage | 48 
vital prognosis | 0 
CT scan | 0 
 Declaration of competing interest | 1008 
no conflict of interest | 1008 
specific financial interests | 1008 
relationships and affiliations | 1008 
subject matter | 1008 
materials discussed | 1008 
manuscript | 1008 
single anatomical right kidney | 0 
single kidney | 0 
right kidney | 0 
emphysematous pyelonephritis complicated | 0 
renal abscess | 0 
intraperitoneal cavity | 0 
pneumoperitoneum | 0 
abdominopelvic scan | 0 
right double J stent | 48 
surgical drainage | 48 
abscesses | 48 
antibiotic therapy | 2 
ceftriaxone | 2 
metronidazole | 2 
ECBU culture | 48 
urinary tract infection | 48 
Pseudomonas Aeruginosa | 48 
intensive care | 2 
dialysis sessions | 2 
insulin therapy | 2 
favorable evolution | 72 
infectious syndrome | 72 
apyrexia | 72 
chronic renal failure | 120 
normal diuresis | 120 
creatinine plateau | 120 
oral antibiotics | 240 
abdominopelvic CT | 672 
clear regression | 672 
bubbles of air | 672 
double J catheter | 1008 
removed | 1008 
type 1 diabetic | 0 
hypertensive | 0 
amlodipine | 0 
right inguinal hernia | -7200 
operated | -7200 
treatment | -7200 
septic shock | -5.8 
febrile low back pain | -5.8 
bubbly gas pattern | 0 
gas in the collecting system | 0 
gas in the renal parenchyma | 0 
gas or abscess to the perinephric space | 0 
gas or abscess to the pararenal space | 0 
bilateral EPN | 0 
solitary kidney with EPN | 0 
percutaneous drainage failure | 0 
nephrectomy | 0 
broad-spectrum antibiotic therapy | 2 
surgical treatment | 48 
conservative treatment | 2 
medical intensive care | 2 
urgent percutaneous | 48 
surgical or endoscopic drainage | 48 
vital prognosis | 0 
CT scan | 0 
 Declaration of competing interest | 1008 
no conflict of interest | 1008 
specific financial interests | 1008 
relationships and affiliations | 1008 
subject matter | 1008 
materials discussed | 1008 
manuscript | 1008 
single anatomical right kidney | 0 
single kidney | 0 
right kidney | 0 
emphysematous pyelonephritis complicated | 0 
renal abscess | 0 
intraperitoneal cavity | 0 
pneumoperitoneum | 0 
abdominopelvic scan | 0 
right double J stent | 48 
surgical drainage | 48 
abscesses | 48 
antibiotic therapy | 2 
ceftriaxone | 2 
metronidazole | 2 
ECBU culture | 48 
urinary tract infection | 48 
Pseudomonas Aeruginosa | 48 
intensive care | 2 
dialysis sessions | 2 
insulin therapy | 2 
favorable evolution | 72 
infectious syndrome | 72 
apyrexia | 72 
chronic renal failure | 120 
normal diuresis | 120 
creatinine plateau | 120 
oral antibiotics | 240 
abdominopelvic CT | 672 
clear regression | 672 
bubbles of air | 672 
double J catheter | 1008 
removed | 1008 
type 1 diabetic | 0 
hypertensive | 0 
amlodipine | 0 
right inguinal hernia | -7200 
operated | -7200 
treatment | -7200 
septic shock | -5.8 
febrile low back pain | -5.8 
bubbly gas pattern | 0 
gas in the collecting system | 0 
gas in the renal parenchyma | 0 
gas or abscess to the perinephric space | 0 
gas or abscess to the pararenal space | 0 
bilateral EPN | 0 
solitary kidney with EPN | 0 
percutaneous drainage failure | 0 
nephrectomy | 0 
broad-spectrum antibiotic therapy | 2 
surgical treatment | 48 
conservative treatment | 2 
medical intensive care | 2 
urgent percutaneous | 48 
surgical or endoscopic drainage | 48 
vital prognosis | 0 
CT scan | 0 
 Declaration of competing interest | 1008 
no conflict of interest | 1008 
specific financial interests | 1008 
relationships and affiliations | 1008 
subject matter | 1008 
materials discussed | 1008 
manuscript | 1008 
single anatomical right kidney | 0 
single kidney | 0 
right kidney | 0 
emphysematous pyelonephritis complicated | 0 
renal abscess | 0 
intraperitoneal cavity | 0 
pneumoperitoneum | 0 
abdominopelvic scan | 0 
right double J stent | 48 
surgical drainage | 48 
abscesses | 48 
antibiotic therapy | 2 
ceftriaxone | 2 
metronidazole | 2 
ECBU culture | 48 
urinary tract infection | 48 
Pseudomonas Aeruginosa | 48 
intensive care | 2 
dialysis sessions | 2 
insulin therapy | 2 
favorable evolution | 72 
infectious syndrome | 72 
apyrexia | 72 
chronic renal failure | 120 
normal diuresis | 120 
creatinine plateau | 120 
oral antibiotics | 240 
abdominopelvic CT | 672 
clear regression | 672 
bubbles of air | 672 
double J catheter | 1008 
removed | 1008 
type 1 diabetic | 0 
hypertensive | 0 
amlodipine | 0 
right inguinal hernia | -7200 
operated | -7200 
treatment | -7200 
septic shock | -5.8 
febrile low back pain | -5.8 
bubbly gas pattern | 0 
gas in the collecting system | 0 
gas in the renal parenchyma | 0 
gas or abscess to the perinephric space | 0 
gas or abscess to the pararenal space | 0 
bilateral EPN | 0 
solitary kidney with EPN | 0 
percutaneous drainage failure | 0 
nephrectomy | 0 
broad-spectrum antibiotic therapy | 2 
surgical treatment | 48 
conservative treatment | 2 
medical intensive care | 2 
urgent percutaneous | 48 
surgical or endoscopic drainage | 48 
vital prognosis | 0 
CT scan | 0 
 Declaration of competing interest | 1008 
no conflict of interest | 1008 
specific financial interests | 1008 
relationships and affiliations | 1008 
subject matter | 1008 
materials discussed | 1008 
manuscript | 1008 
single anatomical right kidney | 0 
single kidney | 0 
right kidney | 0 
emphysematous pyelonephritis complicated | 0 
renal abscess | 0 
intraperitoneal cavity | 0 
pneumoperitoneum | 0 
abdominopelvic scan | 0 
right double J stent | 48 
surgical drainage | 48 
abscesses | 48 
antibiotic therapy | 2 
ceftriaxone | 2 
metronidazole | 2 
ECBU culture | 48 
urinary tract infection | 48 
Pseudomonas Aeruginosa | 48 
intensive care | 2 
dialysis sessions | 2 
insulin therapy | 2 
favorable evolution | 72 
infectious syndrome | 72 
apyrexia | 72 
chronic renal failure | 120 
normal diuresis | 120 
creatinine plateau | 120 
oral antibiotics | 240 
abdominopelvic CT | 672 
clear regression | 672 
bubbles of air | 672 
double J catheter | 1008 
removed | 1008 
type 1 diabetic | 0 
hypertensive | 0 
amlodipine | 0 
right inguinal hernia | -7200 
operated | -7200 
treatment | -7200 
septic shock | -5.8 
febrile low back pain | -5.8 
bubbly gas pattern | 0 
gas in the collecting system | 0 
gas in the renal parenchyma | 0 
gas or abscess to the perinephric space | 0 
gas or abscess to the pararenal space | 0 
bilateral EPN | 0 
solitary kidney with EPN | 0 
percutaneous drainage failure | 0 
nephrectomy | 0 
broad-spectrum antibiotic therapy | 2 
surgical treatment | 48 
conservative treatment | 2 
medical intensive care | 2 
urgent percutaneous | 48 
surgical or endoscopic drainage | 48 
vital prognosis | 0 
CT scan | 0 
 Declaration of competing interest | 1008 
no conflict of interest | 1008 
specific financial interests | 1008 
relationships and affiliations | 1008 
subject matter | 1008 
materials discussed | 1008 
manuscript | 1008 
single anatomical right kidney | 0 
single kidney | 0 
right kidney | 0 
emphysematous pyelonephritis complicated | 0 
renal abscess | 0 
intraperitoneal cavity | 0 
pneumoperitoneum | 0 
abdominopelvic scan | 0 
right double J stent | 48 
surgical drainage | 48 
abscesses | 48 
antibiotic therapy | 2 
ceftriaxone | 2 
metronidazole | 2 
ECBU culture | 48 
urinary tract infection | 48 
Pseudomonas Aeruginosa | 48 
intensive care | 2 
dialysis sessions | 2 
insulin therapy | 2 
favorable evolution | 72 
infectious syndrome | 72 
apyrexia | 72 
chronic renal failure | 120 
normal diuresis | 120 
creatinine plateau | 120 
oral antibiotics | 240 
abdominopelvic CT | 672 
clear regression | 672 
bubbles of air | 672 
double J catheter | 1008 
removed | 1008 
type 1 diabetic | 0 
hypertensive | 0 
amlodipine | 0 
right inguinal hernia | -7200 
operated | -7200 
treatment | -7200 
septic shock | -5.8 
febrile low back pain | -5.8 
bubbly gas pattern | 0 
gas in the collecting system | 0 
gas in the renal parenchyma | 0 
gas or abscess to the perinephric space | 0 
gas or abscess to the pararenal space | 0 
bilateral EPN | 0 
solitary kidney with EPN | 0 
percutaneous drainage failure | 0 
nephrectomy | 0 
broad-spectrum antibiotic therapy | 2 
surgical treatment | 48 
conservative treatment | 2 
medical intensive care | 2 
urgent percutaneous | 48 
surgical or endoscopic drainage | 48 
vital prognosis | 0 
CT scan | 0 
 Declaration of competing interest | 1008 
no conflict of interest | 1008 
specific financial interests | 1008 
relationships and affiliations | 1008 
subject matter | 1008 
materials discussed | 1008 
manuscript | 1008 
single anatomical right kidney | 0 
single kidney | 0 
right kidney | 0 
emphysematous pyelonephritis complicated | 0 
renal abscess | 0 
intraperitoneal cavity | 0 
pneumoperitoneum | 0 
abdominopelvic scan | 0 
right double J stent | 48 
surgical drainage | 48 
abscesses | 48 
antibiotic therapy | 2 
ceftriaxone | 2 
metronidazole | 2 
ECBU culture | 48 
urinary tract infection | 48 
Pseudomonas Aeruginosa | 48 
intensive care | 2 
dialysis sessions | 2 
insulin therapy | 2 
favorable evolution | 72 
infectious syndrome | 72 
apyrexia | 72 
chronic renal failure | 120 
normal diuresis | 120 
creatinine plateau | 120 
oral antibiotics | 240 
abdominopelvic CT | 672 
clear regression | 672 
bubbles of air | 672 
double J catheter | 1008 
removed | 1008 
type 1 diabetic | 0 
hypertensive | 0 
amlodipine | 0 
right inguinal hernia | -7200 
operated | -7200 
treatment | -7200 
septic shock | -5.8 
febrile low back pain | -5.8 
bubbly gas pattern | 0 
gas in the collecting system | 0 
gas in the renal parenchyma | 0 
gas or abscess to the perinephric space | 0 
gas or abscess to the pararenal space | 0 
bilateral EPN | 0 
solitary kidney with EPN | 0 
percutaneous drainage failure | 0 
nephrectomy | 0 
broad-spectrum antibiotic therapy | 2 
surgical treatment | 48 
conservative treatment | 2 
medical intensive care | 2 
urgent percutaneous | 48 
surgical or endoscopic drainage | 48 
vital prognosis | 0 
CT scan | 0 
 Declaration of competing interest | 1008 
no conflict of interest | 1008 
specific financial interests | 1008 
relationships and affiliations | 1008 
subject matter | 1008 
materials discussed | 1008 
manuscript | 1008 
single anatomical right kidney | 0 
single kidney | 0 
right kidney | 0 
emphysematous pyelonephritis complicated | 0 
renal abscess | 0 
intraperitoneal cavity | 0 
pneumoperitoneum | 0 
abdominopelvic scan | 0 
right double J stent | 48 
surgical drainage | 48 
abscesses | 48 
antibiotic therapy | 2 
ceftriaxone | 2 
metronidazole | 2 
ECBU culture | 48 
urinary tract infection | 48 
Pseudomonas Aeruginosa | 48 
intensive care | 2 
dialysis sessions | 2 
insulin therapy | 2 
favorable evolution | 72 
infectious syndrome | 72 
apyrexia | 72 
chronic renal failure | 120 
normal diuresis | 120 
creatinine plateau | 120 
oral antibiotics | 240 
abdominopelvic CT | 672 
clear regression | 672 
bubbles of air | 672 
double J catheter | 1008 
removed | 1008 
type 1 diabetic | 0 
hypertensive | 0 
amlodipine | 0 
right inguinal hernia | -7200 
operated | -7200 
treatment | -7200 
septic shock | -5.8 
febrile low back pain | -5.8 
bubbly gas pattern | 0 
gas in the collecting system | 0 
gas in the renal parenchyma | 0 
gas or abscess to the perinephric space | 0 
gas or abscess to the pararenal space | 0 
bilateral EPN | 0 
solitary kidney with EPN | 0 
percutaneous drainage failure | 0 
nephrectomy | 0 
broad-spectrum antibiotic therapy | 2 
surgical treatment | 48 
conservative treatment | 2 
medical intensive care | 2 
urgent percutaneous | 48 
surgical or endoscopic drainage | 48 
vital prognosis | 0 
CT scan | 0 
 Declaration of competing interest | 1008 
no conflict of interest | 1008 
specific financial interests | 1008 
relationships and affiliations | 1008 
subject matter | 1008 
materials discussed | 1008 
manuscript | 1008 
single anatomical right kidney | 0 
single kidney | 0 
right kidney | 0 
emphysematous pyelonephritis complicated | 0 
renal abscess | 0 
intraperitoneal cavity | 0 
pneumoperitoneum | 0 
abdominopelvic scan | 0 
right double J stent | 48 
surgical drainage | 48 
abscesses | 48 
antibiotic therapy | 2 
ceftriaxone | 2 
metronidazole | 2 
ECBU culture | 48 
urinary tract infection | 48 
Pseudomonas Aeruginosa | 48 
intensive care | 2 
dialysis sessions | 2 
insulin therapy | 2 
favorable evolution | 72 
infectious syndrome | 72 
apyrexia | 72 
chronic renal failure | 120 
normal diuresis | 120 
creatinine plateau | 120 
oral antibiotics | 240 
abdominopelvic CT | 672 
clear regression | 672 
bubbles of air | 672 
double J catheter | 1008 
removed | 1008 
type 1 diabetic | 0 
hypertensive | 0 
amlodipine | 0 
right inguinal hernia | -7200 
operated | -7200 
treatment | -7200 
septic shock | -5.8 
febrile low back pain | -5.8 
bubbly gas pattern | 0 
gas in the collecting system | 0 
gas in the renal parenchyma | 0 
gas or abscess to the perinephric space | 0 
gas or abscess to the pararenal space | 0 
bilateral EPN | 0 
solitary kidney with EPN | 0 
percutaneous drainage failure | 0 
nephrectomy | 0 
broad-spectrum antibiotic therapy | 2 
surgical treatment | 48 
conservative treatment | 2 
medical intensive care | 2 
urgent percutaneous | 48 
surgical or endoscopic drainage | 48 
vital prognosis | 0 
CT scan | 0 
 Declaration of competing interest | 1008 
no conflict of interest | 1008 
specific financial interests | 1008 
relationships and affiliations | 1008 
subject matter | 1008 
materials discussed | 1008 
manuscript | 1008 
single anatomical right kidney | 0 
single kidney | 0 
right kidney | 0 
emphysematous pyelonephritis complicated | 0 
renal abscess | 0 
intraperitoneal cavity | 0 
pneumoperitoneum | 0 
abdominopelvic scan | 0 
right double J stent | 48 
surgical drainage | 48 
abscesses | 48 
antibiotic therapy | 2 
ceftriaxone | 2 
metronidazole | 2 
ECBU culture | 48 
urinary tract infection | 48 
Pseudomonas Aeruginosa | 48 
intensive care | 2 
dialysis sessions | 2 
insulin therapy | 2 
favorable evolution | 72 
infectious syndrome | 72 
apyrexia | 72 
chronic renal failure | 120 
normal diuresis | 120 
creatinine plateau | 120 
oral antibiotics | 240 
abdominopelvic CT | 672 
clear regression | 672 
bubbles of air | 672 
double J catheter | 1008 
removed | 1008 
type 1 diabetic | 0 
hypertensive | 0 
amlodipine | 0 
right inguinal hernia | -7200 
operated | -7200 
treatment | -7200 
septic shock | -5.8 
febrile low back pain | -5.8 
bubbly gas pattern | 0 
gas in the collecting system | 0 
gas in the renal parenchyma | 0 
gas or abscess to the perinephric space | 0 
gas or abscess to the pararenal space | 0 
bilateral EPN | 0 
solitary kidney with EPN | 0 
percutaneous drainage failure | 0 
nephrectomy | 0 
broad-spectrum antibiotic therapy | 2 
surgical treatment | 48 
conservative treatment | 2 
medical intensive care | 2 
urgent percutaneous | 48 
surgical or endoscopic drainage | 48 
vital prognosis | 0 
CT scan | 0 
 Declaration of competing interest | 1008 
no conflict of interest | 1008 
specific financial interests | 1008 
relationships and affiliations | 1008 
subject matter | 1008 
materials discussed | 1008 
manuscript | 1008 
single anatomical right kidney | 0 
single kidney | 0 
right kidney | 0 
emphysematous pyelonephritis complicated | 0 
renal abscess | 0 
intraperitoneal cavity | 0 
pneumoperitoneum | 0 
abdominopelvic scan | 0 
right double J stent | 48 
surgical drainage | 48 
abscesses | 48 
antibiotic therapy | 2 
ceftriaxone | 2 
metronidazole | 2 
ECBU culture | 48 
urinary tract infection | 48 
Pseudomonas Aeruginosa | 48 
intensive care | 2 
dialysis sessions | 2 
insulin therapy | 2 
favorable evolution | 72 
infectious syndrome | 72 
apyrexia | 72 
chronic renal failure | 120 
normal diuresis | 120 
creatinine plateau | 120 
oral antibiotics | 240 
abdominopelvic CT | 672 
clear regression | 672 
bubbles of air | 672 
double J catheter | 1008 
removed | 1008 
type 1 diabetic | 0 
hypertensive | 0 
amlodipine | 0 
right inguinal hernia | -7200 
operated | -7200 
treatment | -7200 
septic shock | -5.8 
febrile low back pain | -5.8 
bubbly gas pattern | 0 
gas in the collecting system | 0 
gas in the renal parenchyma | 0 
gas or abscess to the perinephric space | 0 
gas or abscess to the pararenal space | 0 
bilateral EPN | 0 
solitary kidney with EPN | 0 
percutaneous drainage failure | 0 
nephrectomy | 0 
broad-spectrum antibiotic therapy | 2 
surgical treatment | 48 
conservative treatment | 2 
medical intensive care | 2 
urgent percutaneous | 48 
surgical or endoscopic drainage | 48 
vital prognosis | 0 
CT scan | 0 
 Declaration of competing interest | 1008 
no conflict of interest | 1008 
specific financial interests | 1008 
relationships and affiliations | 1008 
subject matter | 1008 
materials discussed | 1008 
manuscript | 1008 
single anatomical right kidney | 0 
single kidney | 0 
right kidney | 0 
emphysematous pyelonephritis complicated | 0 
renal abscess | 0 
intraperitoneal cavity | 0 
pneumoperitoneum | 0 
abdominopelvic scan | 0 
right double J stent | 48 
surgical drainage | 48 
abscesses | 48 
antibiotic therapy | 2 
ceftriaxone | 2 
metronidazole | 2 
ECBU culture | 48 
urinary tract infection | 48 
Pseudomonas Aeruginosa | 48 
intensive care | 2 
dialysis sessions | 2 
insulin therapy | 2 
favorable evolution | 72 
infectious syndrome | 72 
apyrexia | 72 
chronic renal failure | 120 
normal diuresis | 120 
creatinine plateau | 120 
oral antibiotics | 240 
abdominopelvic CT | 672 
clear regression | 672 
bubbles of air | 672 
double J catheter | 1008 
removed | 1008 
type 1 diabetic | 0 
hypertensive | 0 
amlodipine | 0 
right inguinal hernia | -7200 
operated | -7200 
treatment | -7200 
septic shock | -5.8 
febrile low back pain | -5.8 
bubbly gas pattern | 0 
gas in the collecting system | 0 
gas in the renal parenchyma | 0 
gas or abscess to the perinephric space | 0 
gas or abscess to the pararenal space | 0 
bilateral EPN | 0 
solitary kidney with EPN | 0 
percutaneous drainage failure | 0 
nephrectomy | 0 
broad-spectrum antibiotic therapy | 2 
surgical treatment | 48 
conservative treatment | 2 
medical intensive care | 2 
urgent percutaneous | 48 
surgical or endoscopic drainage | 48 
vital prognosis | 0 
CT scan | 0 
 Declaration of competing interest | 1008 
no conflict of interest | 1008 
specific financial interests | 1008 
relationships and affiliations | 1008 
subject matter | 1008 
materials discussed | 1008 
manuscript | 1008 
single anatomical right kidney | 0 
single kidney | 0 
right kidney | 0 
emphysematous pyelonephritis complicated | 0 
renal abscess | 0 
intraperitoneal cavity | 0 
pneumoperitoneum | 0 
abdominopelvic scan | 0 
right double J stent | 48 
surgical drainage | 48 
abscesses | 48 
antibiotic therapy | 2 
ceftriaxone | 2 
metronidazole | 2 
ECBU culture | 48 
urinary tract infection | 48 
Pseudomonas Aeruginosa | 48 
intensive care | 2 
dialysis sessions | 2 
insulin therapy | 2 
favorable evolution | 72 
infectious syndrome | 72 
apyrexia | 72 
chronic renal failure | 120 
normal diuresis | 120 
creatinine plateau | 120 
oral antibiotics | 240 
abdominopelvic CT | 672 
clear regression | 672 
bubbles of air | 672 
double J catheter | 1008 
removed | 1008 
type 1 diabetic | 0 
hypertensive | 0 
amlodipine | 0 
right inguinal hernia | -7200 
operated | -7200 
treatment | -7200 
septic shock | -5.8 
febrile low back pain | -5.8 
bubbly gas pattern | 0 
gas in the collecting system | 0 
gas in the renal parenchyma | 0 
gas or abscess to the perinephric space | 0 
gas or abscess to the pararenal space | 0 
bilateral EPN | 0 
solitary kidney with EPN | 0 
percutaneous drainage failure | 0 
nephrectomy | 0 
broad-spectrum antibiotic therapy | 2 
surgical treatment | 48 
conservative treatment | 2 
medical intensive care | 2 
urgent percutaneous | 48 
surgical or endoscopic drainage | 48 
vital prognosis | 0 
CT scan | 0 
 Declaration of competing interest | 1008 
no conflict of interest | 1008 
specific financial interests | 1008 
relationships and affiliations | 1008 
subject matter | 1008 
materials discussed | 1008 
manuscript | 1008 
single anatomical right kidney | 0 
single kidney | 0 
right kidney | 0 
emphysematous pyelonephritis complicated | 0 
renal abscess | 0 
intraperitoneal cavity | 0 
pneumoperitoneum | 0 
abdominopelvic scan | 0 
right double J stent | 48 
surgical drainage | 48 
abscesses | 48 
antibiotic therapy | 2 
ceftriaxone | 2 
metronidazole | 2 
ECBU culture | 48 
urinary tract infection | 48 
Pseudomonas Aeruginosa | 48 
intensive care | 2 
dialysis sessions | 2 
insulin therapy | 2 
favorable evolution | 72 
infectious syndrome | 72 
apyrexia | 72 
chronic renal failure | 120 
normal diuresis | 120 
creatinine plateau | 120 
oral antibiotics | 240 
abdominopelvic CT | 672 
clear regression | 672 
bubbles of air | 672 
double J catheter | 1008 
removed | 1008 
type 1 diabetic | 0 
hypertensive | 0 
amlodipine | 0 
right inguinal hernia | -7200 
operated | -7200 
treatment | -7200 
septic shock | -5.8 
febrile low back pain | -5.8 
bubbly gas pattern | 0 
gas in the collecting system | 0 
gas in the renal parenchyma | 0 
gas or abscess to the perinephric space | 0 
gas or abscess to the pararenal space | 0 
bilateral EPN | 0 
solitary kidney with EPN | 0 
percutaneous drainage failure | 0 
nephrectomy | 0 
broad-spectrum antibiotic therapy | 2 
surgical treatment | 48 
conservative treatment | 2 
medical intensive care | 2 
urgent percutaneous | 48 
surgical or endoscopic drainage | 48 
vital prognosis | 0 
CT scan | 0 
 Declaration of competing interest | 1008 
no conflict of interest | 1008 
specific financial interests | 1008 
relationships and affiliations | 1008 
subject matter | 1008 
materials discussed | 1008 
manuscript | 1008 
single anatomical right kidney | 0 
single kidney | 0 
right kidney | 0 
emphysematous pyelonephritis complicated | 0 
renal abscess | 0 
intraperitoneal cavity | 0 
pneumoperitoneum | 0 
abdominopelvic scan | 0 
right double J stent | 48 
surgical drainage | 48 
abscesses | 48 
antibiotic therapy | 2 
ceftriaxone | 2 
metronidazole | 2 
ECBU culture | 48 
urinary tract infection | 48 
Pseudomonas Aeruginosa | 48 
intensive care | 2 
dialysis sessions | 2 
insulin therapy | 2 
favorable evolution | 72 
infectious syndrome | 72 
apyrexia | 72 
chronic renal failure | 120 
normal diuresis | 120 
creatinine plateau | 120 
oral antibiotics | 240 
abdominopelvic CT | 672 
clear regression | 672 
bubbles of air | 672