53 years old| 0  
    male| 0  
    unrestrained driver| 0  
    presented to the trauma bay| 0  
    high-speed head-on motor vehicle collision| 0  
    blood pressure 80/20 mm Hg| 0  
    heart rate 126 beats/min| 0  
    tender distended abdomen| 0  
    no signs of seat belt markings| 0  
    computed tomography scan demonstrated active extravasation from the infrarenal aorta| 0  
    surrounding retroperitoneal hematoma| 0  
    no associated abdominal injuries| 0  
    no spinal injuries| 0  
    bilateral rib fractures| 0  
    pulmonary contusions| 0  
    left ulnar fracture| 0  
    right tibia fracture| 0  
    brought emergently to the operating room| 0  
    treated with two proximal aortic cuffs| 0  
    24 × 58-mm cuff placed distally| 0  
    24 × 39-mm cuff placed proximally| 0  
    inferior mesenteric artery intentionally covered| 0  
    tolerated the procedure well| 0  
    extremity fractures treated by orthopedic surgeon| 0  
    follow-up CT scan within 24 hours demonstrated resolution of extravasation| 24  
    resolution of hematoma| 24  
    gram-positive sepsis| 24  
    pneumonia| 24  
    respiratory failure| 24  
    tracheostomy| 24  
    discharged 15 days after initial operation| 360  
    ambulatory condition| 360  
    one year later without clinical sequelae| 8760  
    follow-up CT scan demonstrates normal aorta| 8760  
    stable graft configuration| 8760  
    