77 year old|0
    female |0
    atrial fibrillation |0
    scheduled for emergency laparotomy |0
    emergency laparotomy |0
    closure of hollow viscous perforation |0
    past medical history unremarkable |0
    no medications |0
    general anaesthesia for laparoscopic appendicectomy |-48
    abdominal pain |-24
    fever |-24
    febrile |0
    pulse 110/min |0
    blood pressure 106/72 mmHg |0
    respiratory rate 20/min |0
    no abnormal heart sounds |0
    no abnormal breath sounds |0
    haemoglobin 11.9 g/dl |-6
    total counts 14,000/mm3 |-6
    13% band forms |-6
    serum sodium 140 mEq/l |-6
    serum potassium 3.6 mEq/l |-6
    platelets 220,000/mm3 |-6
    creatinine 1.4 mg% |-6
    bilateral mild pleural effusion |0
    normal cardia |0
    sinus tachycardia |0
    heart rate 106/min |0
    operating room |0
    ECG heart rate 156/min |0
    atrial fibrillation confirmed |0
    invasive blood pressure 106/72 mmHg |0
    SpO2 93% |0
    intravenous metoprolol |0
    no change in heart rate |0
    defibrillator available |0
    blood pressure stable |0
    trachea intubated |0
    rapid sequence induction |0
    midazolam 1 mg |0
    fentanyl 250 mcg |0
    propofol 60 mg |0
    succinylcholine 60 mg |0
    central line inserted |0
    anaesthesia maintained |0
    air |0
    oxygen |0
    sevoflurane |0
    fentanyl |0
    hydromorphone |0
    rocuronium |0
    intravenous amiodarone 150 mg |0
    heart rate reduced to 80–90/min |0
    blood pressure improved 126/86 mmHg |0
    sinus rhythm |0
    uncompensated metabolic acidosis |0
    bicarbonate 16 mEq/l |0
    respiratory alkalosis |0
    PCO2 26 mmHg |0
    serum potassium 3 mEq/l |0
    intravenous potassium 20 mmol/L |0
    repeat serum potassium 3.4 mEq/l |0
    intraoperative period uneventful |0
    transferred to ICU |0
    IV potassium supplementation 20 mmol/l |0
    IV magnesium sulphate 1 g |0
    serum magnesium 1.2 mg/dl |0
    calcium chloride |0
    serum calcium 6 mg/dl |0
    CRP elevated |0
    procalcitonin elevated |0
    thyroid function tests normal |0
    trachea extubated |12
    sinus rhythm |12
    consultation with cardiologist |12
    aspirin 81 mg started |12
    negative transthoracic echocardiogram |12
    regular follow-up advised |12
    discharged home |12
    low-dose aspirin therapy |12
    
    
    