34 years old | 0
male | 0
admitted to the hospital | 0
poor hygiene | 0
alcohol use disorder | -672
cirrhosis | -672
hypertension | -672
hepatitis B | -672
macrocytic anemia | -672
moderate mitral valve regurgitation | -672
previous Clostridium Difficile infection | -672
stage 2 hypertensive chronic kidney disease | -672
previous episodes of acute renal failure | -672
sepsis | 0
extensive edema of the lower body | 0
conscious | 0
verbal-logical contact preserved | 0
wheezing | 0
rhonchi over the lung fields | 0
dullness at the base of the left lung | 0
loud mitral regurgitation murmur | 0
blood pressure 120/80 mmHg | 0
heart rate 100 bpm | 0
body temperature 38.0C | 0
WBC 10.0 × 103/ul | 0
HBG 8.1 g/dl | 0
HCT 25.6 % | 0
PLT 139 × 103/ul | 0
CRP 124 mg/l | 0
Creatinine 1.83 mg/dl | 0
Potassium 4.10 mmol/l | 0
Sodium 130 mmol/l | 0
Albumin 2.5 g/dl | 0
ALT 49 u/l | 0
AST 110 u/l | 0
INR 1.33 | 0
fluid in the pleural cavity | 0
extensive edema of subcutaneous tissue of the lower abdomen and pelvis | 0
no abscess | 0
Mitral Regurgitation with preserved ejection fraction | 0
no other deficits | 0
Ceftazidime | 0
Imipenem/Cilastatin and Vancomycin | 24
blood cultures grew Staphylococcus Epidermidis | 24
wound cultures grew multiple pathogens | 24
skin cultures collected | 24
antibiotic dosage adjusted to Glomerular Filtration Rate (GFR) and dialysis | 24
antibiotic therapy continued | 24
TPN started | 72
Vasopressor support with Norepinephrine | 72
petechiae | 120
bursting blisters oozing with serous content | 120
necrotic changes | 120
pain with movement and palpation | 120
diagnosis of Fournier's Gangrene | 120
transfer to the surgical ward | 120
septic shock | 120
acute renal failure | 120
minimal urine production | 120
CVVHD initiated | 120
first session of CVVHD | 120
four sessions of hemodialysis | 168
first necrosectomy | 168
successful removal of necrotic skin and subcutaneous tissue | 168
FGSI 7 | 168
second necrosectomy | 384
further removal of devitalized tissue | 384
application of sterile dressing with antiseptic solutions | 384
HBOT | 408
thirteen sessions of HBOT | 408
episode of epistaxis from the right nasal sinus | 408
anterior tamponade | 408
completion of HBOT | 504
transfer back to the community hospital | 504
NPWT started | 552
dressing applied on the lower abdomen, right thigh and the anterior surface of the left thigh | 552
general anesthesia | 552
further removal of devitalized tissue | 552
negative pressure dressings fully sealed | 552
discharge of serous-blood content from the wound | 552
negative pressure device set to intermittent mode | 552
NPWT deployed for 16 days | 624
foam changed 4 times | 624
removal of negative pressure dressings | 720
standard sterile dressings impregnated with moisturizing and antimicrobial agents | 720
granulation tissue and wound clearance achieved | 720
qualified for skin transplant | 720
CRP and leukocytes acutely increased | 792
urosepsis | 792
blood and urine cultures positive for Escrichia Coli | 792
antibiotic therapy with Imipenem | 792
vasopressor support | 792
sudden cardiac arrest | 816
death | 816