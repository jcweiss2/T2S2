22 years old | 0
    woman | 0
    type 1 diabetes mellitus | -4320
    poorly controlled type 1 diabetes mellitus | -4320
    presented to the Emergency Department | 0
    fever | -120
    headache | -120
    nausea | -120
    vomiting | -120
    prescribed sumatriptan 50 mg | -216
    home medications: Ademalog insulin | -4320
    home medications: insulin glargine | -4320
    home medications: lisinopril 2.5 mg oral daily | -4320
    purchased 2 cockatiel birds | -4320
    temperature 39.2°C | 0
    pulse 123 beats per minute | 0
    respiratory rate 22 per minute | 0
    blood pressure 131/75 mmHg | 0
    oxygen saturation 100% | 0
    confused | 0
    aphasic | 0
    nuchal rigidity | 0
    right upper-extremity paresis | 0
    negative Kernig’s signs | 0
    negative Brudzinski’s signs | 0
    no papilledema | 0
    white blood cell count 22 K/µL | 0
    hemoglobin 13.8 g/dL | 0
    sodium 129 mEq/L | 0
    potassium 4 mEq/L | 0
    chloride 100 mEq/L |(0)
    bicarbonate 13 mEq/L | 0
    blood urea nitrogen 9 mg/dL | 0
    creatinine 0.89 mg/dL | 0
    creatine phosphokinase 275 U/L | 0
    lactic acid 2.5 mmol/L | 0
    hemoglobin A1c 13.3% | 0
    urine toxicology screen negative | 0
    sinus tachycardia | 0
    computed tomography scan of the head | 0
    started on empiric antibiotics | 0
    vancomycin 1 gram IV twice daily | 0
    ceftriaxone 2 gram IV every 12 hours | 0
    acyclovir 600 milligrams IV every 8 hours | 0
    received 3 liters of isotonic fluids | 0
    lumbar puncture performed | 0
    cloudy cerebrospinal fluid | 0
    cerebrospinal fluid WBC count 2790 cells/µL | 0
    segmented neutrophils 75% | 0
    total protein 163 mg/dL | 0
    glucose 31 mg/dL | 0
    CSF PCR positive for Listeria monocytogenes | 7
    CSF cultures confirmed Listeria | 72
    blood cultures confirmed Listeria | 120
    antimicrobial regimen changed to ampicillin and gentamicin | 7
    admitted to the MICU | 0
    diabetic ketoacidosis | 0
    received 4 liters of isotonic fluids | 0
    initial POCUS hyperdynamic LV function | 24
    repeat echocardiogram showed LV EF 30% | 48
    alertness and aphasia wax and wane | 48
    8-channel EEG no seizure activity | 72
    24-channel EEG no seizure activity | 72
    dark discolored urine | 96
    repeat CPK 27,131 U/L | 96
    CPK peak 299,637 U/L | 144
    aldolase peak 1104 U/L | 144
    non-oliguric | 144
    creatinine at baseline | 144
    rheumatological panel unrevealing | 144
    septic shock | 144
    acute respiratory failure | 144
    new seizure | 144
    intubation | 144
    mechanical ventilation | 144
    vasopressor support | 144
    EEG after seizure treatment | 144
    CPK decline | 144
    received 49 liters of fluids | 240
    vasopressor support for septic shock | 264
    methicillin-resistant Staphylococcus aureus coverage | 264
    Pseudomonas aeruginosa coverage | 264
    mental status improvement | 336
    liberated from mechanical ventilation | 336
    transferred to internal medicine ward | 432
    tachycardic | 456
    short of breath | 456
    CT angiogram showing pulmonary embolism | 456
    transthoracic echocardiogram showing right atrial thrombus | 456
    repeat echocardiogram EF 60% | 480
    interventional radiology-guided thrombectomy | 480
    heparin infusion | 480
    observed in MICU | 528
    transferred to internal medicine ward | 528
    completed 3-week ampicillin course | 504
    normal motor function | 504
    no recurrence of seizures | 504
    discharged on day 23 | 552
    apixaban | 552
    levetiracetam | 552
    no residual neurological deficits | 552
    Listeria meningitis | 0
    Listeria bacteremia | 120
    rhabdomyolysis | 96
    septic cardiomyopathy | 48
    left ventricular dilatation | 48
    right atrial thrombus | 456
    pulmonary embolism | 456
    rehabilitation facility | 552
