23 years old | 0
    female | 0
    ventilated | 0
    ICU admission | 0
    lower uterine segment cesarean section (LUSCS) | -408
    intrauterine death (IUD) | -408
    oligohydramnios | -408
    no fetal cardiac activity | -408
    no fetal movement | -408
    anterior placenta | -408
    oliguric | -408
    drowsy | -408
    jaundice | -408
    high-grade fever | -408
    intubated | -408
    ventilated | -408
    transfused four packed blood cells | -408
    transfused 21 fresh frozen plasmas | -408
    temperature of 38.9°C | 0
    pulse rate of 140/min | 0
    blood pressure of 130/80 mmHg | 0
    SpO2 of 99% | 0
    oxygen-enriched bag ventilation | 0
    icterus | 0
    pallor | 0
    generalized anasarca | 0
    abdominal distention | 0
    scattered rhonchi | 0
    crepitations | 0
    clean abdominal wound | 0
    urinary catheter | 0
    scanty urine | 0
    nasogastric tube | 0
    dark green-colored aspirate | 0
    bleeding per vaginum | 0
    total leukocyte count of 22,000 cu/mm | 0
    polymorphonuclear leukocytosis (84%) | 0
    hemoglobin of 9.3 g/dl | 0
    Prothrombin Time of 17.4 seconds | 0
    PTI Index of 74.7 | 0
    normal renal function tests | 0
    urea of 50 mg/dl | 0
    elevated serum glutamic-oxaloacetic transaminase (220 IU/L) | 0
    elevated serum glutamic pyruvic transaminase (132 IU/L) | 0
    total bilirubin 3.4 mg/dl | 0
    conjugated bilirubin 2.1 mg/dl | 0
    alkaline phosphatase 120 IU/L | 0
    total proteins 4.5 g/L | 0
    albumin 2.0 g/L | 0
    nonreactive viral markers | 0
    24 h urine albumin 2+ positive | 0
    culture and sensitivity of endotracheal secretions | 48
    vasopressor noradrenaline initiated | 48
    inotropic dopamine initiated | 48
    exploratory laparotomy | 72
    intraoperative blood transfusion | 72
    intraoperative blood products | 72
    serosanguineous fluid collection | 72
    persistent hepatic derangement | 72
    hypoproteinemia | 72
    persistent pyrexia (38.9°C–39.4°C) | 72
    polymorphonuclear leukocytosis (25,000–33,000) | 72
    derangement of coagulation | 72
    isolation of P. dispersa | 96
    resistant to standard antimicrobials | 96
    sensitive to tigecycline | 96
    sensitive to colistin | 96
    colistimethate initiated | 96
    persistent fever (38.9°C–39.4°C) | 96
    fibrin degradation products positive | 168
    D-Dimer negative | 168
    blood-stained secretions | 168
    frank blood in secretions | 168
    blood culture negative | 408
    urinary catheter tip culture negative | 408
    pericardial tap culture negative | 408
    ascitic fluid culture negative | 408
    growth of Candida spp. in urine | 408
    vasopressors required | 432
    inotropes required | 432
    ARDS progression | 432
    ventilator support | 432
    renal failure | 432
    multiple dialyses | 432
    red blood cells transfused | 432
    fresh frozen plasma transfused | 432
    total parenteral nutrition | 432
    enteral nutrition | 432
    albumin administered | 432
    cardiac arrest | 432
    cardiopulmonary cerebral resuscitation | 432
    continued intensive care management | 432
    another episode of cardiac arrest | 480
    declared dead | 480

    23 years old | 0  
    female | 0  
    ventilated | 0  
    ICU admission | 0  
    lower uterine segment cesarean section (LUSCS) | -408  
    intrauterine death (IUD) | -408  
    oligohydramnios | -408  
    no fetal cardiac activity | -408  
    no fetal movement | -408  
    anterior placenta | -408  
    oliguric | -408  
    drowsy | -408  
    jaundice | -408  
    high-grade fever | -408  
    intubated | -408  
    ventilated | -408  
    transfused four packed blood cells | -408  
    transfused 21 fresh frozen plasmas | -408  
    temperature of 38.9°C | 0  
    pulse rate of 140/min | 0  
    blood pressure of 130/80 mmHg | 0  
    SpO2 of 99% | 0  
    oxygen-enriched bag ventilation | 0  
    icterus | 0  
    pallor | 0  
    generalized anasarca | 0  
    abdominal distention | 0  
    scattered rhonchi | 0  
    crepitations | 0  
    clean abdominal wound | 0  
    urinary catheter | 0  
    scanty urine | 0  
    nasogastric tube | 0  
    dark green-colored aspirate | 0  
    bleeding per vaginum | 0  
    total leukocyte count of 22,000 cu/mm | 0  
    polymorphonuclear leukocytosis (84%) | 0  
    hemoglobin of 9.3 g/dl | 0  
    Prothrombin Time of 17.4 seconds | 0  
    PTI Index of 74.7 | 0  
    normal renal function tests | 0  
    urea of 50 mg/dl | 0  
    elevated serum glutamic-oxaloacetic transaminase (220 IU/L) | 0  
    elevated serum glutamic pyruvic transaminase (132 IU/L) | 0  
    total bilirubin 3.4 mg/dl | 0  
    conjugated bilirubin 2.1 mg/dl | 0  
    alkaline phosphatase 120 IU/L | 0  
    total proteins 4.5 g/L | 0  
    albumin 2.0 g/L | 0  
    nonreactive viral markers | 0  
    24 h urine albumin 2+ positive | 0  
    culture and sensitivity of endotracheal secretions | 48  
    vasopressor noradrenaline initiated | 48  
    inotropic dopamine initiated | 48  
    exploratory laparotomy | 72  
    intraoperative blood transfusion | 72  
    intraoperative blood products | 72  
    serosanguineous fluid collection | 72  
    persistent hepatic derangement | 72  
    hypoproteinemia | 72  
    persistent pyrexia (38.9°C–39.4°C) | 72  
    polymorphonuclear leukocytosis (25,000–33,000) | 72  
    derangement of coagulation | 72  
    isolation of P. dispersa | 96  
    resistant to standard antimicrobials | 96  
    sensitive to tigecycline | 96  
    sensitive to colistin | 96  
    colistimethate initiated | 96  
    persistent fever (38.9°C–39.4°C) | 96  
    fibrin degradation products positive | 168  
    D-Dimer negative | 168  
    blood-stained secretions | 168  
    frank blood in secretions | 168  
    blood culture negative | 408  
    urinary catheter tip culture negative | 408  
    pericardial tap culture negative | 408  
    ascitic fluid culture negative | 408  
    growth of Candida spp. in urine | 408  
    vasopressors required | 432  
    inotropes required | 432  
    ARDS progression | 432  
    ventilator support | 432  
    renal failure | 432  
    multiple dialyses | 432  
    red blood cells transfused | 432  
    fresh frozen plasma transfused | 432  
    total parenteral nutrition | 432  
    enteral nutrition | 432  
    albumin administered | 432  
    cardiac arrest | 432  
    cardiopulmonary cerebral resuscitation | 432  
    continued intensive care management | 432  
    another episode of cardiac arrest | 480  
    declared dead | 480  
    