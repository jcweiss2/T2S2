42 years old | 0
female | 0
health care provider | 0
admitted to the emergency department | 0
high-grade fever | -48
productive cough | -48
shortness of breath | -48
bony pains | -48
contact with a patient of similar complaints | -48
left nephrectomy | -3600
caesarian section | -3600
abortion | -3600
obese | 0
diabetes mellitus type 2 | 0
Glasgow Coma Scale 15/15 | 0
hemodynamically stable | 0
leukopenia | 0
lymphopenia | 0
bilateral infiltrates on chest x-ray | 0
admitted to the ward | 0
septic screen for MERS-CoV | 0
influenza AB | 0
H1N1 | 0
dengue serology | 0
malaria tests | 0
broad spectrum antibiotics | 0
oseltamivir | 0
admitted to the Intensive Care Unit | 24
extensive bilateral consolidations on chest x-ray | 24
refractory hypoxaemia | 24
elective intubation | 24
mechanical ventilation | 24
Fraction of inspired oxygen 100% | 24
acute respiratory distress syndrome protocol | 24
lung protective strategies | 24
low tidal volume | 24
prone position | 24
tracheal aspirates sent for MERS-CoV | 24
MERS-CoV virus positive | 48
Peginterferon Alpha-2a | 48
ribavirin | 48
intravenous methylprednisolone | 48
Extracorporeal membrane oxygenation treatment contemplated | 72
improvement in respiratory function | 120
weaning trial | 288
sedation cessation | 288
methylprednisolone tapered | 288
Peginterferon Alpha-2a discontinued | 288
ribavirin discontinued | 288
hemodynamically stable | 288
respiratory function improved | 288
radiological features improved | 288
started to wake up | 288
started to move all limbs | 288
polyuric | 312
urine osmolarity 95 | 312
serum osmolarity 341 | 312
urine sodium less than 20 | 312
serum sodium 161 meq/L | 312
chloride 119 meq/L | 312
blood sugar 25 mmol/L | 312
Desmopressin | 312
brain computed tomography | 312
sudden-onset of diabetes insipidus | 312
massive spontaneous intracranial hemorrhage | 312
intra-ventricular extension | 312
tonsillar herniation | 312
unresponsive | 312
Glasgow Coma Scale 3/15 | 312
pupils 3 mm wide with sluggish reaction | 312
CT brain showed right frontal hematoma | 312
subarachnoid hemorrhage | 312
midline shift | 312
subfalcine herniation | 312
normal platelet count | 312
normal coagulation profile | 312
no anti-coagulation treatment | 312
negative blood cultures | 312
neurologists and neurosurgical team review | 312
no surgical intervention | 312
medical supportive measures | 312
lost all brain stem reflexes | 312
pupils became fixed and dilated | 312
follow-up brain CT scan | 312
complete loss of gray and white matter differentiation | 312
large frontal hematoma | 312
complete effacement of extra axial CSF spaces | 312
contrast enhanced CT images | 312
no enhancement of intracranial vessels | 312
computed tomography angiogram | 312
no visualization of Middle cerebral artery | 312
no flow within the posterior circulation | 312
brain death criteria | 312
cardiac arrest | 2664
declared dead | 2664