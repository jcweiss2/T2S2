58 years old | 0
male | 0
admitted to the hospital | 0
hyperpyrexia | -168
dyspnoea | -48
cough | -48
phlegm with blood | -48
history of hypertension | -0
bought a chicken from a local live poultry market | -168
poultry-related exposure | -168
diagnosed with community-acquired pneumonia | -168
antibacterial therapy | -168
condition failed to improve | -168
chest computed tomography scan | -168
multiple ground-glass opacities | -168
consolidation in both lungs | -168
right pleural effusion | -168
transferred to hospital | 0
increased C-reactive protein | 0
procalcitonin | 0
leukopenia | 0
lymphopenia | 0
reduced T lymphocyte subgroups | 0
HIV antibody test negative | 0
arterial blood gas analysis | 0
pH of 7.46 | 0
partial pressure of carbon dioxide | 0
partial pressure of oxygen | 0
severe acute respiratory distress syndrome | 0
endotracheal intubation | 0
mechanical ventilation | 0
antibiotic treatment | 0
moxifloxacin | 0
cefoperazone-sulbactam | 0
corticosteroids | 0
continuous renal replacement therapy | 0
influenza A virus | 0
oseltamivir | 0
veno-venous extracorporeal membrane oxygenation | 96
blood culture yielded Staphylococcus haemolyticus | 96
vancomycin | 96
imipenem/cilastatin | 96
caspofungin | 96
Pseudomonas aeruginosa | 96
CRP and PCT improved | 168
chest X-ray improved | 168
subcutaneous and mediastinal emphysemas | 240
ventilator parameters decreased | 240
emphysemas relieved | 240
BALF retested | 336
influenza A virus still positive | 336
condition deteriorated | 384
chest X-ray worsened | 384
1,3-β-d-glucan test negative | 384
galactomannan test negative | 384
new bacterial co-infections | 384
strong antibacterial drugs | 384
no improvement | 384
BALF and blood cultures positive for C. neoformans | 552
C. neoformans sensitive to flucytosine | 552
fluconazole | 552
voriconazole | 552
amphotericin B | 552
itraconazole | 552
serum cryptococcal capsular polysaccharide antigen test positive | 552
caspofungin ceased | 552
intravenous liposomal amphotericin B | 552
fluconazole | 552
examinations of possible exogenous sources of cryptococcosis negative | 552
C. neoformans infection from initial colonization of respiratory tract | 552
BALF and blood cultures negative for C. neoformans | 672
persistent lung infiltrates | 672
progressive pulmonary fibrosis | 672
ventilator monitoring data showed a constant decrease in tidal volume | 672
BALF and blood cultures positive for multidrug-resistant Stenotrophomonas maltophilia | 960
condition deteriorated | 960
septic shock | 1128
disseminated intravascular coagulation | 1128
multi-organ failure | 1128
died | 1128