78 years old | 0
male | 0
admitted to the hospital | 0
benign prostatic hyperplasia | 0
coronary artery disease | 0
atrial fibrillation | 0
presented to the emergency department | 0
leukocytosis | 0
worsening renal function | 0
hyperkalemia | 0
admitted to the ICU | 0
hemodynamic instability | 0
septic shock secondary to Pseudomonas aeruginosa urinary tract infection | 0
started on cefepime | 0
required vasopressor support | 0
fever of 38.3°C | 168
pustular rash | 168
erythematous base covering upper extremities and trunk | 168
no mucosal involvement | 168
leukocytosis with neutrophilia (8170 neutrophils/µl) | 168
elevated C-reactive protein level (4.15 mg/dL) | 168
chest X-ray obtained | 168
no acute cardiopulmonary abnormality | 168
repeated blood, urine, and pustule cultures for bacteria | 168
negative cultures | 168
persistently hypotensive | 168
repeated CXR | 192
new-onset bilateral interstitial opacities and consolidation | 192
tested for COVID-19 | 192
SARS-CoV-2 RNA nasopharyngeal swab positive | 192
no signs of respiratory distress | 192
no requirement for supplemental oxygen | 192
treated supportively | 192
skin biopsy of the rash | 192
papillary dermal edema | 192
subcorneal/intracorneal pustules | 192
mixed inflammatory infiltrate (lymphocytes, neutrophils, rare eosinophils) | 192
EuroSCAR study group criteria score of 12 (AGEP diagnosis) | 192
cefepime discontinued | 192
treated symptomatically with topical emollients | 192
resolution of exanthem within a few days | 192
post-pustular desquamation | 192
diagnosed with COVID-19 | 192
second reported case of AGEP in COVID-19 patient | 192
COVID-19 infection | 192
vigorous immune response to COVID-19 | 192
concurrent cefepime use | 192
development of AGEP | 192
IL-36 receptor antagonist (IL36RN) gene mutations | 192
lack of lip/oral involvement | 192
cytokine storm | 192
low-grade inflammation in elderly | 192
delayed development of AGEP | 192
cutaneous manifestations of COVID-19 | 192
cephalosporin exposure | 192
genetic predisposition | 192
pro-inflammatory cells and cytokines | 192
resolution after discontinuation of cefepime | 192
