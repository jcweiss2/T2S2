47 years old | 0
male | 0
admitted to the hospital | 0
diabetes mellitus | 0
hypertension | 0
obstructive sleep apnea | 0
BiPAP ventilation | 0
laparoscopic sleeve gastrectomy | 0
complicated hospital course | 0
anastomotic leak | 0
computed tomography-guided aspiration of abdominal collections | 0
closing gastric fistula | 0
closing transverse colon | 0
washing abdomen | 0
repeated peritoneal lavage | 0
peritonitis | 0
sepsis | 0
acute kidney injury | 0
sputum cultures positive for CNSA | 0
no known allergies | 0
vancomycin started | 0
tigecycline started | 0
meropenem started | 0
red-man syndrome | -72
vancomycin infused over 3 hours | 0
peak sample drawn | 144
trough sample drawn | 144
peak level 32.4 mg/L | 144
trough level 24.8 mg/L | 144
dose changed to 1500 mg q24h | 144
predicted peak Cp 19 mg/L | 144
actual peak level 22.7 mg/L | 168
actual trough level 12.5 mg/L | 168
serum creatinine elevated | 0
vancomycin clearance reduced | 0
158 kg | 0
173 cm | 0
MIC 1 mcg/mL | 0
