24 years old | 0
    male | 0
    hyperthyroidism | 0
    noncompliant with methimazole treatment | 0
    presented as a patient to level I trauma facility | 0
    restrained driver in a rollover MVA | 0
    unknown loss of consciousness | 0
    self-extricated from the wreckage | 0
    ambulatory at the scene | 0
    right lower quadrant abdominal pain | 0
    right wrist pain | 0
    consumed ethanol | 0
    heart rate 170 | 0
    blood pressure 156/78 | 0
    temperature not documented | 0
    heart rate 163 | 0
    blood pressure 153/84 | 0
    temperature 37.3°C | 0
    Glascow Coma Score 15 | 0
    anxious | 0
    fine tremor | 0
    hematoma over the left eye | 0
    seat belt sign to the left chest | 0
    right-sided abdominal tenderness to palpation | 0
    left hand abrasions | 0
    right wrist pain without deformity | 0
    no neck abrasions | 0
    no neck contusions | 0
    no goiter present | 0
    focused abdominal sonography for trauma exam negative | 0
    head CT scan negative | 0
    maxillofacial CT scan negative | 0
    chest CT scan negative | 0
    abdomen CT scan negative | 0
    pelvis CT scan negative | 0
    plain radiographs of the extremities negative | 0
    resuscitated with 2 L normal saline | 0
    administered IV lorazepam 2 mg | 0
    administered IV fentanyl 50 mcg | 0
    complete blood count performed | 0
    complete metabolic panel performed | 0
    lactic acid tested | 0
    thyroid studies performed | 0
    ethanol level tested | 0
    rapid urine drug screen performed | 0
    sodium 149 | 0
    potassium 3.4 | 0
    chloride 108 | 0
    carbon dioxide 15 | 0
    anion gap 26 | 0
    BUN 11 | 0
    creatinine 0.51 | 0
    AST 43 | 0
    ALT 58 | 0
    lactic acid 7.6 | 0
    free T4 5.61 | 0
    thyroid stimulating hormone <0.015 | 0
    rapid urine drug screen positive for cannabinoids | 0
    ethanol level 101 | 0
    serum osmolality tested | 0
    ethylene glycol tested | 0
    methanol tested | 0
    serum osmolality 288 | 0
    osmolar gap −6 | 0
    ethylene glycol negative | 0
    methanol negative | 0
    remained hypertensive | 0
    remained tachycardic | 0
    TC suspected | 0
    given methimazole 5 mg | 0
    given propranolol 1 mg injection | 0
    fluid resuscitation continued | 0
    admitted to internal medicine service | 0
    lactic acidosis improved to 0.8 | 168
    sodium 143 | 168
    chloride 109 | 168
    CO2 21 | 168
    anion gap 13 | 168
    AST 24 | 168
    ALT 50 | 168
    blood glucose 102 | 168
    blood glucose 85 | 168
    tachycardia resolved | 24
    hypertension resolved | 24
    continued on methimazole 5 mg 3 times daily | 24
    continued on propranolol 10 mg 3 times daily | 24
    blood cultures negative for growth | 24
    instructed to follow-up with endocrinology | 48
    discharged after 48 hours | 48
    did not follow-up with endocrinology | -4320
    seen again in emergency department 6 months later | -4320
    TC secondary to tonsillitis | -4320
    remained medication noncompliant | -4320
    still yet to follow-up with endocrinology clinic | -4320

    