69 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
Child–Pugh class C cirrhosis | 0 | 0 | Factual
fell on his left side | -1 | -1 | Factual
Glasgow coma score 15/15 | 0 | 0 | Factual
vital signs within normal limits | 0 | 0 | Factual
left hip tenderness | 0 | 0 | Factual
no ecchymosis to the abdomen, flank or thigh | 0 | 0 | Negated
undisplaced fracture of his left acetabulum | 0 | 0 | Factual
liver dysfunction | 0 | 0 | Factual
pH 7.271 | 0 | 0 | Factual
base excess minus 7.3 | 0 | 0 | Factual
PT 18.2 | 0 | 0 | Factual
INR-1.5 | 0 | 0 | Factual
APTT ratio 1.42 | 0 | 0 | Factual
platelets 73 | 0 | 0 | Factual
bilirubin 63 mmol/l | 0 | 0 | Factual
Hb 124 g/l | 0 | 0 | Factual
intravenous cannula inserted | 0 | 0 | Factual
warmed Hartmanns one litre infusion commenced | 0 | 0 | Factual
referred to the Orthopaedic on call team | 1 | 1 | Factual
blood pressure dropped to 75/51 mm Hg | 2 | 2 | Factual
tachycardic | 2 | 2 | Factual
serum lactate 9 mmol/l | 2 | 2 | Factual
FAST examination revealed intraabdominal fluid | 2 | 2 | Factual
treated for sepsis | 2 | 4 | Factual
intensive care, orthopaedic and general registrar attended the patient | 4 | 4 | Factual
pH 7.227 | 4 | 4 | Factual
base excess of −17.9 | 4 | 4 | Factual
serum lactate of 16.3 mmol/l | 4 | 4 | Factual
Hb 75 g/l | 4 | 4 | Factual
arterial blood pressure 90/60 mm Hg | 4 | 4 | Factual
pulse rate 90/min | 4 | 4 | Factual
left lower abdominal quadrant and upper thigh swollen with ecchymosis | 4 | 4 | Factual
diagnosis of haemorrhagic shock | 4 | 4 | Factual
massive transfusion pathway activated | 4 | 4 | Factual
four units of Blood transfused | 4 | 6 | Factual
four units of FFP transfused | 4 | 6 | Factual
two adult therapeutic doses of platelets transfused | 4 | 6 | Factual
10 units of cryoprecipitate transfused | 4 | 6 | Factual
noradrenaline infusion commenced | 6 | 24 | Factual
pelvic binder in place | 6 | 24 | Factual
CT scan performed | 8 | 10 | Factual
CT abdomen confirmed fracture of the left acetabulum | 10 | 10 | Factual
significant haematoma on left pelvic sidewall | 10 | 10 | Factual
8 mm enhancing nodule suggestive of an internal iliac artery pseudoaneurysm | 10 | 10 | Factual
ill-defined blush of contrast within the haematoma | 10 | 10 | Factual
extra-peritoneal haematoma inseparable from the bladder | 10 | 10 | Factual
cirrhotic liver | 10 | 10 | Factual
6.7 cm infra-renal aortic aneurysm | 10 | 10 | Factual
transferred to intensive care unit | 12 | 12 | Factual
CT Angiogram performed | 48 | 50 | Factual
no arterial bleed | 50 | 50 | Factual
prophylactic embolization recommended | 50 | 50 | Factual
gelfoam embolization of anterior and posterior division segmental branches of the left internal iliac artery | 50 | 52 | Factual
10 lb skeletal traction applied | 52 | 120 | Factual
uncontrollable bleeding from his pin site | 120 | 120 | Factual
pin site removed | 120 | 120 | Factual
continuous pressure applied to the wound | 120 | 120 | Factual
died on 30 January 2017 | 1224 | 1224 | Factual
end stage liver failure | 1200 | 1224 | Factual
hepatic encephalopathy | 1200 | 1224 | Factual