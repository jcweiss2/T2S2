83 years old | 0
female | 0
admitted to the emergency department | 0
fever | 0
vomiting | 0
diffuse abdominal pain | 0
right upper quadrant pain | 0
rheumatoid arthritis | -Inf
atrial fibrillation | -Inf
asthma | -Inf
cerebrovascular disease | -Inf
hysterectomy | -Inf
intestinal obstruction | -Inf
no previous history of gallstones | -Inf
regular medication | -Inf
oral steroids | -Inf
methotrexate | -Inf
clopidogrel | -Inf
omeprazole | -Inf
paracetamol | -Inf
hormone replacement therapy | -Inf
nonsteroidal anti-inflammatory drug | -Inf
tenderness in right upper quadrant | 0
guarding in right upper quadrant | 0
temperature 37.6°C | 0
leukocytosis | 0
C-reactive protein elevated | 0
abnormal liver enzymes | 0
ALT elevated | 0
AST elevated | 0
GGT elevated | 0
total blood bilirubin elevated | 0
plain abdominal radiography | 0
circular gas pattern in gallbladder area | 0
computed tomography | 0
gas in gallbladder wall | 0
gas-fluid level within gallbladder | 0
emergency laparoscopic cholecystectomy | 0
extensive inflammation | 0
necrosis of gallbladder | 0
gallbladder distension | 0
gallbladder puncture | 0
extraction of intraluminal pus | 0
dissection in Calot's triangle | 0
exposure of cystic duct | 0
intraoperative cholangiography | 0
excluded biliary obstruction | 0
cholecystectomy | 0
bubbling from gallbladder wall | 0
resection completed | 0
no complications | 0
no conversion to open surgery | 0
laparoscopic abdominal lavage | 0
drainage | 0
postoperative intravenous antibiotic therapy | 0
unremarkable recovery | 0
discharged | 264
pathological analysis | 264
full-thickness infarctive necrosis | 264
abscess | 264
single small calculus | 264
microbiological analysis | 264
Clostridium perfringens | 264
