67 years old | 0
male | 0
cardiogenic cerebral infarction | -672
chills | 0
right chest pain | 0
admitted to the hospital | 0
body temperature 36.4 °C | 0
blood pressure 82/66 mmHg | 0
pulse rate 110/min | 0
oxygen saturation 90% | 0
respiratory rate 30 breaths/min | 0
right coarse crackles | 0
white blood cell count 9500/μl | 0
neutrophils 7695/μl | 0
platelets 165,000/μl | 0
C-reactive protein 2.59 mg/dl | 0
right S2-infiltration | 0
systemic blood pressure rapidly declined to 60 mmHg | 2
oxygen saturation decreased to 70% | 2
transferred to the intensive care unit (ICU) | 2
mechanical ventilation support | 2
oxygenation not fully recovered | 2
bronchoscopy | 2
large amount of bleeding (>1000 ml) from the right upper bronchus | 2
obstructing the right main bronchus | 2
complete opacification of the right hemithorax | 2
veno-venous extracorporeal membrane oxygenation (v-v ECMO) support | 2
P. aeruginosa identified from bronchial secretion and blood | 2
meropenem and ciprofloxacin | 2
management of systemic infection | 2
withdrawal of v-v ECMO | 336
abscess formation progressed in the right lung | 336
P. aeruginosa empyema | 336
purulent sputum and minor bleeding from the right lung | 336
right pneumonectomy and pleural lavage | 720
P. aeruginosa infection resolved | 720
discharged from the ICU | 876
home whirlpool bath | -672
contaminated aerosol | -672
P. aeruginosa isolated from the whirlpool bathtub | -672
genetically identical to the patient's sample | 0
MLST analysis | 0
whole genome sequencing | 0
phylogenetic analysis | 0
exoenzyme S gene (exoS) | 0
drug resistance genes | 0
virulent factor gene | 0
surgical intervention | 720
necrotizing pneumonia | 0
severe purulent pneumonia | 0
genomic analysis | 0
direct exposure to aerosol contaminated with virulent P. aeruginosa | 0