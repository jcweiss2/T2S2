40 years old | 0
male | 0
admitted to the hospital | 0
shock | 0
flu-like illness | -72
nausea | -72
general malaise | -72
lower abdominal pain | -72
severe diarrhea | -72
administered 500 ml of 5% albumin | -72
administered 1,500 ml/day of saline | -72
consciousness deteriorated | -24
right hemiparesis | -24
temperature of 36.0°C | 0
blood pressure of 95/72 mm Hg | 0
pulse of 160 beats/min | 0
respiratory rate of 25 breaths/min | 0
SpO2 was 100% | 0
jugular vein was collapsed | 0
bilateral radial artery pulses were insufficiently palpable | 0
extremities were cold | 0
whole-blood sample was coagulated easily | 0
hyperviscosity | 0
polycythemia | 0
hypoalbuminemia | 0
severe leukocytosis | 0
elevated creatinine | 0
severe metabolic acidosis | 0
influenza virus types A and B were positive | 0
pericardial effusion | 0
collapsed inferior vena cava | 0
occlusion of the division of the left M2 segment of the middle cerebral artery | 0
diffusion-weighted MR imaging revealed high signal intensity in the MCA territory | 0
acute cerebral infarction | 0
external and internal decompression surgery | 20
midline shift of the head on CT | 20
postoperative intracranial pressure was 9 mm Hg | 20
cerebral edema progression | 20
internal decompression | 32
mechanical ventilation | 0
massive fluid resuscitation | 0
swelling, redness, and heat sensation in the lateral surfaces of the legs | 0
pretibial compartment syndrome | 0
bilateral calf fasciotomy | 0
all samples were negative | 0
toxic shock syndrome was considered | 0
sepsis was considered | 0
anaphylaxis was considered | 0
acute adrenal insufficiency was considered | 0
drug reactions were considered | 0
polycythemia vera was considered | 0
severe right hemiparesis | 48
Broca's aphasia | 48
unable to walk without assistance | 48
theophylline was administered | 48
ISCLS attacks were documented | 720
fasciotomy | 720
monoclonal immunoglobulin was found | 720
immunoelectrophoresis | 720
plasmacytosis was not found | 720
bone marrow aspiration | 720
intravenous infusion of immunoglobulins | 720
corticosteroids | 720
immunosuppressive therapy | 720