22 years old| 0
    African American| 0
    female| 0
    systemic lupus erythematosus (SLE)| -105192
    lupus nephritis| -105192
    cyclophosphamide| -105192
    mycophenolate| -105192
    azathioprine| 0
    prednisone| 0
    hypothyroidism| 0
    hypertension| 0
    myasthenia gravis| 0
    admitted to the intensive care unit| 0
    acute hypoxic respiratory failure| 0
    endotracheal intubation| 0
    mechanical ventilation| 0
    febrile (102.3 °F)| 0
    tachycardia (144 beat per minute)| 0
    decreased breath sounds over the left anterior hemi-thorax| 0
    pneumonia| 0
    respiratory muscle weakness| 0
    myasthenia crisis| 0
    sepsis| 0
    plasmapheresis| 0
    steroids| 0
    antimicrobial agents| 0
    pyridostigmine therapy not immediately instituted| 0
    no improvement despite five cycles of plasmapheresis| 0
    pyridostigmine started later| 0
    hypotensive| 192
    oliguria| 192
    acute renal failure| 192
    acute tubular necrosis (ATN)| 192
    abdominal tenderness| 216
    abdominal computed tomography (CT) scan| 216
    free air in the abdominal cavity| 216
    emergent laparotomy| 216
    peritonitis| 216
    gastric cardia perforation| 216
    perforation repaired| 216
    worsening coagulation panel| 0
    liver function tests worsening| 0
    prothrombin time (PT) normal at admission| 0
    PT increased to 18.1 s| 0
    albumin decreased to 2.1 g/dL| 0
    bilirubin normal| 0
    alkaline phosphatase (AKP) normal| 0
    AST normal (19 units/L)| 0
    ALT normal (16 units/L)| 0
    AKP stable| 0
    bilirubin stable| 0
    AST worsened to 352 units/L| 216
    ALT worsened to 369 units/L| 216
    fulminant hepatic failure| 216
    AST peaked to 1,618 units/L| 240
    ALT peaked to 1,018 units/L| 240
    acute respiratory distress syndrome| 360
    fatal cardiac arrest| 360
    herpes hepatitis| 360
    disseminated herpes| 360
    fulminant hepatic failure due to disseminated herpes| 360
    herpes inclusion bodies in liver parenchyma| 360
    liver enlarged and mottled| 360
    zones of coagulative necrosis| 360
    intra-nuclear ground glass inclusions| 360
    minimal inflammatory response| 360
    pneumonia with ARDS| 360
    gastric perforation with peritonitis| 360
    cessation of plasmapheresis| 240
    plasmapheresis cycles| 0
    
    