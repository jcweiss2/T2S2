58 years old|0
    male|0
    presented to the emergency department|0
    found on the floor of his apartment|0
    unable to provide detailed history|0
    several episodes of loose bowel movements|0
    denied change in stool color|0
    denied blood in the diarrhea|0
    no abdominal pain|0
    no nausea|0
    no vomiting|0
    no recent antibiotics use|0
    no fever|0
    no cough|0
    no chest pain|0
    no dyspnea|0
    not hospitalized within the past year|0
    never traveled outside the United States|0
    diagnosed with Crohn's disease|-350400
    multiple bowel resections|-350400
    not on steroids|0
    treated with Vedolizumab|-5760
    infliximab stopped prior to Vedolizumab|-5760
    emaciated patient|0
    blood pressure 78/50|0
    heart rate 98|0
    respiratory rate 22|0
    temperature 99°F|0
    lung exam crackles over the right lung|0
    unremarkable abdominal exam|0
    unremarkable cardiovascular exam|0
    elevated WBCs count 20.9|0
    neutrophils 96.1%|0
    lymphocytes 0.8%|0
    monocytes 2.3%|0
    eosinophils 0%|0
    chest X ray multiple opacities in the right lung field|0
    IgE level 205|0
    HIV negative|0
    admitted to intensive care unit|0
    management of septic shock|0
    management of pneumonia|0
    started on Vancomycin|0
    started on Aztreonam|0
    started on Levofloxacin|0
    started on vasopressors|0
    clinical picture didn't improve|96
    sputum cultures negative|96
    blood cultures negative|96
    CT of the chest|96
    opacification within the entirety of the right lung|96
    air bronchograms|96
    bronchoscopy on 4th day of admission|96
    normal mucosa without lesions|96
    bronchoalveolar lavage obtained|96
    cultures negative for bacteria|96
    cultures negative for tuberculosis|96
    cultures negative for fungi|96
    bronchial washing cytology acute inflammation|96
    bronchial washing cytology filariform larvae|96
    serology positive for Strongyloides antibodies|96
    started on ivermectin|96
    condition improved significantly|96
    discharged|168
    