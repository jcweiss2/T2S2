72 years old | 0
female | 0
admitted to the emergency department | 0
dyspnea | 0
asthma | -672
congestive heart failure | -672
abdominal examination was normal | 0
no abdominal distension | 0
costophrenic sinuses were obscured on the chest radiograph | 0
no free air under the diaphragm | 0
respiratory failure | 0
hypoxemia | 4
hypotension | 4
intubation | 4
accidental esophageal intubation | 4
abdominal distension | 4
nasogastric tube insertion | 4
peritonitis | 4
hemorrhagic fluid from the nasogastric tube | 4
general surgery consultation | 4
excessive abdominal distension | 4
active hemorrhage from the nasogastric tube | 4
intra-abdominal massive free air | 4
emergency laparotomy | 4
perforation focus on the anterior surface of the lesser curvature of the stomach | 4
active arterial bleeding | 4
repair of the perforation focus | 4
Roseo-Graham omental patch | 4
bleeding ceased | 4
no mass or ulcer at the level of the perforation focus | 4
surgical drain positioned | 4
methylene blue test | 72
drain removed | 72
transferred to the ward | 840
discharged | 840