81 years old | 0
man | 0
arrived at IRCCS Policlinico’s Operative Unit of Vascular Surgery | 0
distal wound abscess | -720
right below-the-knee femoropopliteal composite bypass | -720
critical limb ischemia | -720
methicillin-resistant Staphylococcus aureus (MRSA) infection | -720
femoropopliteal bypass | -720
alcoholic liver disease | 0
atrial fibrillation | 0
no anticoagulation therapy | 0
left carotid stenting | 0
significant asymptomatic stenosis | 0
endovascular exclusion of a left iliac aneurysm | 0
no fever | 0
hemoglobin 12 g/dL | 0
International Normalized Ratio (INR) 1.38 | 0
negative blood cultures | 0
very thin and emaciated | 0
body mass index (BMI) 15 | 0
treatable abdomen | 0
no masses palpable | 0
normal heart examination | 0
normal chest examination | 0
palpable femoral pulses bilaterally | 0
absent popliteal pulses bilaterally | 0
absent tibial pulses bilaterally | 0
patent right femoropopliteal bypass | 0
valid flow at Duplex-scan examination | 0
no exposure of the graft through the infected wound | 0
anticoagulation with low-molecular-weight heparin | 0
intravenous antibiotic therapy with Teicoplanin 400 mg daily | 0
acute limb ischemia | 96
bypass thrombosis | 96
significant increase of white blood cells count | 96
fever | 96
surgical exploration of the popliteal artery | 96
no run-off from tibial vessels | 96
graft removed | 96
right thigh amputation | 96
postoperative course uneventful | 96
normalized white blood cells count | 96
fever disappeared | 96
no additional signs of infection | 96
clean stump wound | 96
continued antibiotic therapy with Teicoplanin | 96
discharged on ninth postoperative day (POD) | 216
rehabilitation referral | 216
pulsatile mass in right neck | 648
pulsatile mass in left groin | 648
dysphagia | 648
hemoptysis | 648
duplex ultrasound of neck | 648
duplex ultrasound of left groin | 648
angio-CT scan | 648
hypodense bulk at common carotid artery | 648
hypodense bulk at bifurcation | 648
pseudoaneurysm extending to ICA | 648
dislocating right internal jugular vein | 648
invading nearby parapharyngeal space | 648
small hematoma enveloping left iliac-femoral passage | 648
flow recorded at duplex ultrasound | 648
re-referred to IRCCS Policlinico’s Operative Unit of Vascular Surgery | 648
no fever | 648
Teicoplanin 200 mg twice daily | 648
INR 5.5 | 648
leukocytosis 14700/uL | 648
anemia (hemoglobin 10.4 g/dL) | 648
huge palpable tender pulsatile mass in right neck | 648
smaller pulsatile mass in left groin | 648
trans-thoracic color-Doppler echocardiography | 648
no valvular source of septic embolism | 648
normal heart ejection fraction 68.1% | 648
referred to operating room | 648
general anesthesia | 648
isolated right common femoral artery | 648
selective right internal carotid angiography | 648
voluminous pseudoaneurysm arising from carotid bifurcation | 648
extended toward parapharyngeal space | 648
invisible external carotid artery | 648
visible superior thyroid artery | 648
placement of 0.035-in hydrophilic stiff wire into ICA | 648
exchanged with 10F sheath | 648
deployment of Fluency PTFE-covered nitinol self-expanding stent | 648
angiographic control showing patency of ICA | 648
complete exclusion of lesion | 648
absence of endoleaks | 648
non-pulsatile mass | 648
surgical right laterocervical incision | 648
evacuated hematoma | 648
PTFE graft wrapped around carotid wall | 648
copiously irrigated incision | 648
closed wound in layers | 648
excised left femoral pseudoaneurysm | 648
reconstructed vessel wall with pericardial patch | 648
admitted to intensive care unit | 648
returned to ward | 648
culture samples of laterocervical mass | 648
culture samples of left femoral pseudoaneurysm | 648
MRSA present | 648
postoperative blood samples negative | 648
urine culture with ESBL Escherichia coli | 648
antibiotic therapy with Ceftriaxone 2 g twice daily | 648
continued Teicoplanin | 648
dual therapy for 4 weeks | 648
healed laterocervical wound | 648
healed groin wounds | 648
no signs of infection recurrence | 648
discharged on POD 15 | 360
acetyl salicylic acid 100 mg daily | 360
low-molecular-weight heparin | 360
rehabilitation referral | 360
angio-CT scan showing stent patency | 360
no endoleaks | 360
no flow impairment at duplex ultrasound | 360
7 months follow-up | 5040
poor general condition | 5040
healed laterocervical wound | 5040
healed inguinal wounds | 5040
patent stent | 5040
approved by institutional review board | 5040
informed consent | 5040
atrial fibrillation |8 0
