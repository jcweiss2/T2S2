62 years old| 0
female | 0
admitted to the hospital| 0
type 2 diabetes mellitus| 0
repaglinide| 0
atypical chest pain| 0
no evidence of coronary disease| 0
superficial phlebitis of the left forearm| -48
backaches| -24
fever| -24
readmitted| 0
Glasgow Coma Scale score 15/15| 0
fully alert| 0
no motor deficit| 0
no neck stiffness| 0
major inflammatory syndrome| 0
C-reactive protein level 47.8 mg/dl| 0
normal white blood cell count| 0
renal function mildly impaired| 0
serum creatinine level 2.1 mg/dl| 0
blood urea nitrogen 84 mg/dl| 0
no evidence of pulmonary infection| 0
no evidence of urinary infection| 0
empirical antimicrobial therapy| 0
amoxicillin| 0
clavulanic acid| 0
initial blood cultures grew S. aureus| 0
antimicrobial therapy changed to vancomycin| 0
switched to oxacillin| 0
corticosteroids not prescribed| 0
dysarthria| 48
drowsiness| 48
polypnea| 48
transferred to intensive care unit| 48
became confuse| 48
disorientated| 48
stiff neck| 48
painful neck| 48
normal clinical examination of cranial nerves| 48
normal peripheral reflexes| 48
no motor deficit| 48
lumbar puncture revealed purulent CSF| 48
CSF white blood cell count 31,800/mm3| 48
CSF glucose 54 mg/dl| 48
CSF lactate 13.5 mmol/l| 48
CSF culture negative| 48
contrast-enhanced brain CT| 48
no specific lesion| 48
no sign of ventriculitis| 48
no sign of venous thrombosis| 48
referred to third hospital| 336
Glasgow Coma Scale score 11/15| 336
intubation| 336
mechanical ventilation| 336
major hypoxemia| 336
MRI performed| 336
cervical spinal cord enlarged| 336
T2-weighted images intramedullary hyperintensity| 336
diffuse leptomeningeal enhancement| 336
focal intramedullary gadolinium enhancements| 336
signal abnormalities extended to medulla oblongata| 336
no significant changes in cerebral hemispheres| 336
no evidence of hydrocephalus| 336
no evidence of brain edema| 336
preserved BAEPs| 336
no cortical SSEPs| 336
normal peripheral activities (P9 and N13 complex)| 336
absence of P14 complex| 336
neurological condition worsened within 2 days| 432
spontaneous breathing disappeared| 432
ventilated in pressure control mode| 432
dysautonomic episodes| 432
hypotension| 432
extreme bradycardia| 432
complete quadriparesis| 432
anesthesia| 432
horizontal ophthalmoplegia| 432
conscious| 432
able to respond to simple questions by vertical eye movements| 432
blood cultures positive for methicillin-sensitive S. aureus| 168
endocarditis ruled out| 168
repeated MRI| 456
signal hyperintensity extended to thoracic spinal cord| 456
T1-weighted imaging signal hypointensity of grey matter| 456
day 21| 504
all brain stem reflexes absent| 504
BAEPs absent| 504
persisting wave I upon left ear stimulation| 504
withdrawal of intensive care therapy| 504
died from cardiocirculatory failure| 504
autopsy performed| 504
macroscopic examination confirmed extensive leptomeningitis| 504
microscopic examination confirmed vasculitis| 504
secondary medullar ischemia| 504
no metastatic areas of S. aureus infection| 504
