68 years old | 0
female | 0
admitted to the emergency room | 0
altered level of consciousness | 0
blood pressure 80/60 mm Hg | 0
pulse rate 112 beats/min | 0
respiratory rate 24 breaths/min | 0
body temperature 34.9°C |0
chronic kidney disease (stage 4) | 0
type 2 diabetes mellitus | -157248
insulin treatment | -87600
acute pyelonephritis admission (February 2015) | -33000
acute pyelonephritis admission (December 2016) | -17520
acute pyelonephritis admission (August 2018) | -2352
resided in a nursing hospital | -2352
non-smoker | 0
no previous history of pulmonary disease | 0
elevated white blood cell count | 0
low hemoglobin | 0
normal platelets | 0
elevated blood urea nitrogen | 0
elevated serum creatinine | 0
septic shock | 0
metabolic acidosis | 0
urine microscopy many WBCs | 0
urine dipstick positive for nitrite | 0
transferred to medical intensive care unit | 0
continuous renal replacement therapy | 0
antibiotics adjusted for renal impairment | 0
dyspnea | 408
chest X-ray atelectasis | 408
urine culture Escherichia coli | 408
negative blood culture | 408
chest CT partial atelectasis | 408
prominent wall thickening and enhancement | 408
no evidence of other pulmonary diseases | 408
bronchoscopy inflammation | 480
bronchoscopy necrosis | 480
AFB stain negative | 480
MTB DNA detection negative | 480
MTB culture negative | 480
bronchoscopic biopsy fungal infection | 480
yeast-like fungus | 480
PAS stain positive | 480
Candida albicans growth | 480
intravenous fluconazole | 480
electrolyte imbalance worsened | 480
uremia worsened | 480
dialysis rejected | 480
do-not-resuscitate order | 888
died | 888
