9 years old | 0
    male | 0
    admitted to the pediatric ICU | 0
    septic shock | 0
    respiratory insufficiency | 0
    mechanical ventilation | 0
    cardiac monitoring | 0
    severe neutropenia | -336
    fever of unknown origin | -336
    broad-spectrum antibiotic therapy | -336
    antifungal therapy | -336
    circular erythematous lesions with necrotic center | -216
    extensive necrosis | -216
    septate hyaline hyphae on biopsy | -216
    Grocott staining showing septate hyphae | -216
    culture confirming Aspergillus niger | -216
    whole body CT scan showing no disseminated infection | -216
    amphotericin B therapy | -216
    fluconazole therapy | -216
    voriconazole added to therapy | -216
    no improvement | -216
    death | 2160
    <|eot_id|>
    