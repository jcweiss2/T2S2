46 years old | 0
female | 0
admitted to the hospital | 0
head trauma | -336
headaches | -504
posterior neck pain | -504
nausea | -504
loss of appetite | -504
blurry vision | -504
HIV/AIDS | -672
chronic hepatitis B infection | -672
cocaine abuse | -672
infectious endocarditis | -672
low-grade fever | 0
hypotension | 0
tachycardia | 0
normal respiratory rate | 0
normal oxygen saturation | 0
cachectic patient | 0
acute distress | 0
anemia | 0
leukopenia | 0
moderate hyponatremia | 0
hypochloremia | 0
elevated creatinine level | 0
hypoalbuminemia | 0
pituitary abscess | 0
central hypothyroidism | 0
secondary adrenal insufficiency | 0
low insulin-like growth factor-1 level | 0
low prolactin level | 0
aggressive intravenous fluid resuscitation | 0
broad-spectrum antibiotics | 0
vancomycin | 0
cefepime | 0
metronidazole | 0
fluconazole | 0
oral levothyroxine | 0
intravenous hydrocortisone | 0
diabetes insipidus | 48
oral desmopressin | 48
high urine output | 48
increased thirst | 48
decreased urine osmolality | 48
increased blood osmolality | 48
decreased size of the mass | 240
thickening of the peripheral wall | 240
marked decrease in the pituitary gland volume | 7920
necrosis | 7920
absence of normal tissue enhancement | 7920
residual small effusion | 7920
persistent central hypothyroidism | 7920
persistent secondary adrenal insufficiency | 7920
secondary hypogonadism | 7920
discontinued desmopressin | 168
normal sodium levels | 168
normal serum osmolality | 168
discharged | 432