62 years old | 0
female | 0
Indian | 0
admitted to the hospital | 0
fatigue | -72
bilateral lower extremity pain | -72
weakness | -72
unable to eat | -48
unable to drink | -48
compliant with immunosuppressive regimen | -72
history of end-stage kidney disease | -2160
history of hypertension | -2160
history of diabetes | -2160
solitary kidney | -2160
deceased donor renal transplantation | -2160
rhabdomyolysis | -2160
calcineurin inhibitor−statin interaction | -2160
denies chest pain | 0
denies cough | 0
denies shortness of breath | 0
denies back pain | 0
denies headache | 0
denies visual symptoms | 0
denies speech difficulties | 0
denies nausea | 0
denies vomiting | 0
denies diarrhea | 0
denies fever | 0
denies chills | 0
denies rigors | 0
pain in thighs | -72
no overlying skin changes | -72
no sick contacts | 0
voiding without difficulty | 0
serum calcium 18.0 mg/dl | 0
ionized calcium 2.26 mmol/l | 0
low parathyroid hormone level | 0
creatinine 3.9 mg/dl | 0
oral calcium dosage increased | -2160
hypocalcemia | -2160
hyperphosphatemia | -2160
pretransplantation serum calcium 9 mg/dl | -2160
pretransplantation serum phosphorus 4.3 mg/dl | -2160
pretransplantation alkaline phosphatase 82 U/l | -2160
pretransplantation magnesium 2 mg/dl | -2160
urinalysis positive for 1+ leukocyte esterase | -2160
urinalysis positive for 2+ protein | -2160
urinalysis pH 5 | -2160
posttransplantation nadir serum creatinine 1.1 mg/dl | -2160
posttransplantation serum calcium 9.3 mg/dl | -2160
posttransplantation serum phosphorus 4.7 mg/dl | -2160
posttransplantation magnesium 1.4 mg/dl | -2160
posttransplantation alkaline phosphatase 65 U/l | -2160
urinalysis positive for 1+ leucocyte esterase | -2160
urinalysis negative for protein | -2160
urinalysis pH 7.0 | -2160
history of recurrent renal calculi | -2160
left native nephrectomy | -3600
thyroidectomy | -2880
multinodular goiter | -2880
incidental removal of 2 adenomatous parathyroid glands | -2880
PTH dropped from 300 pg/ml to 9 pg/ml | -2880
commenced oral calcium carbonate supplementation | -2880
commenced oral calcitriol | -2160
serum calcium within normal limits | -72
stopped proton pump inhibitor | -72
losartan dose up titrated | -72
vigorous saline rehydration | 0
improvement in serum calcium | 24
improvement in ionized calcium | 24
improvement in mental status | 24
i.v. bolus doses of furosemide | 24
forced diuresis | 24
calcium levels continued to correct | 48
mental status improved | 48
no additional measures to reduce serum calcium | 48
AKI slow to resolve | 48
tacrolimus trough levels at target | 48
renal ultrasound revealed new renal calculi | 48
mild hydronephrosis | 48
nuclear medicine renogram showed prompt uptake of tracer | 48
delayed excretion consistent with acute tubular necrosis | 48
no definite evidence of significant obstruction | 48
suppressed PTH | 48
25-OH-vitamin D level 10 ng/ml | 48
PTH-related peptide level 0.9 pmol/l | 48
normal serum protein electrophoresis | 48
serum free light chain ratio 1.14 | 48
thyroid-stimulating hormone elevated | 48
levothyroxine dose increased | 48
urinalysis positive for 1+ protein | 48
became hypocalcemic | 72
calcitriol and calcium carbonate supplementation re-introduced | 72
Escherichia coli urosepsis | 96
critical care admission | 96
antibiotics | 96
i.v. fluid resuscitation | 96
mycophenolate mofetil dose reduced | 96
leukopenia | 96
renal allograft function continued to decline | 120
renal biopsy performed | 120
calcium deposition in the tubules | 120
acute tubular necrosis | 120
interstitial inflammation | 120
borderline rejection | 120
no acute vascular or glomerular changes | 120
oral pulse of prednisone | 120
target tacrolimus trough level increased | 120
mycophenolate mofetil dose increased | 120
serum creatinine returned to baseline | 168
nadir serum creatinine 0.8 mg/dl | 168
no further recurrence of hypercalcemia | 168
PTH level remains suppressed | 168