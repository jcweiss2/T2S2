53 years old | 0
male | 0
hypertension | 0
diabetes mellitus | 0
hypothyroidism | 0
dilated cardiomyopathy | 0
admitted to the hospital | 0
prolonged pyrexia | -336
coronary angiography | -336
fever | -168
standard investigations | -168
routine blood cultures | -168
imaging | -168
transferred to our care | -168
febrile | 0
toxic | 0
early diastolic murmur | 0
hemoglobin 8.3 g/dL | 0
white blood cells 9200 cells/mm3 | 0
platelets 2,23,000/mm3 | 0
serum creatinine level 2.2 mg/dL | 0
erythrocyte sedimentation rate 88 mm/h | 0
urine analysis showed 3-5 red blood cells | 0
raised 24-h urine protein of 1527 mg/24 h | 0
mild hepatosplenomegaly | 0
no evidence of focal lesions in the spleen or liver | 0
mildly prominent pulmonary vasculature | 0
cardiomegaly | 0
no significant lung parenchymal pathology | 0
left ventricular ejection fraction (LVEF) of 30% | -168
normal heart valves | -168
global hypokinesia | -168
mild aortic regurgitation | 0
three discrete small mobile vegetations | 0
no evidence of cusp perforation | 0
no ring abscess | 0
LVEF was 20% | 0
choroidal infiltrates | 0
no evidence of embolization to skin | 0
no evidence of embolization to other organ | 0
antinuclear antibodies (anti-ANA) negative | 0
anti– double stranded antibody (anti-dsDNA) negative | 0
anti–nucleophilic cytoplasmic antibodies (anti-ANCA) negative | 0
complement levels (C3 and C4) within normal range | 0
thyroid profile normal | 0
treated for heart failure | 0
ceftriaxone 1 g twice daily intravenously | 0
routine serial bacterial blood cultures did not show any growth | 0
BACTEC Myco/F Lytic medium demonstrated NTM | 0
linezolid and clarithromycin added | 0
species identification using Line probe assay technique revealed M. abscessus | 0
drug sensitivities obtained | 0
sensitive to amikacin | 0
sensitive to clarithromycin | 0
sensitive to linezolid | 0
sensitive to tobramycin | 0
intermediate sensitivity to cefoxitin | 0
resistant to doxycycline | 0
resistant to imipenem | 0
resistant to cefepime | 0
resistant to ceftriaxone | 0
resistant to minocycline | 0
resistant to amox–clavulanic acid | 0
isoniazid added | 0
ethambutol added | 0
cefoxitin added | 0
defervesced for the first time | 168
linezolid withheld for 10 days | 168
linezolid reinstituted in lower doses | 178
creatinine stabilized at 2.6 mg/dL | 504
dyspnea improved | 504
repeat 2D echo showed increase in LVEF to 40% | 504
valvular vegetations present | 504
blood cultures still grew M. abscessus | 504
aortic valve replacement surgery considered | 504
aortic valve replacement surgery withheld | 504
repeat 2D ECHO at 4 weeks post treatment showed no change in vegetation size | 1008
discharged on request | 1008
developed worsening cardiac failure | 1056
died of pulmonary edema | 1056
died of renal dysfunction | 1056