63 years old | 0
female | 0
diagnosed with papillary thyroid carcinoma | -132432
resection | -132432
radiotherapy | -132432
stenosis of the esophagus | -132432
repeated aspiration | -132432
respiratory insufficiency | -132432
pneumonia | -132432
purulent pleurisy | -132432
pleurectomy | -132432
restrictive ventilation pattern | -132432
recurrent nerve palsy | -132432
percutaneous endoscopic gastrostomy | -175200
tracheostoma | -175200
home ventilation | -175200
decreased mobility | -87600
secondary depression | -87600
stopped talking | -87600
mandible fixation | -87600
inability to open mouth | -87600
stented left axis vertebralis | -52560
stenosis of internal axis carotis | -52560
arterial hypertension | -52560
secondary lactase deficiency | -52560
esophageal stenosis dilation | -52560
referred to University of Erlangen | 0
fistula between esophagus and tracheal membrane | 0
examined by multiple chiefs and consultants | 0
deemed too unstable for open surgery | 0
inability to open mouth | 0
recurrent nerve palsy | 0
referral to surgical intensive care unit | 168
suffering from pneumonia | 168
4-multiresistente gramnegative Pseudomonas aeruginosa | 168
veno+venous extracorporeal membrane oxygenation | 168
partial thromboplastin time of 60 seconds | 168
preseptic status | 168
low ventilation forces | 168
thoracic computed tomography | 192
confirmed big fistula of tracheal membrane | 192
decision to try endobronchial stenting | 192
procedure performed | 216
vv-ECMO partly ineffective | 216
rising septical issues | 216
high volume input of physiological saline | 216
retrograde stenting performed | 216
introduced DLET | 216
modified FS stent | 216
created new stoma for tracheal cannula | 216
secured continuous airway replacement | 216
introduced jagwire | 216
flipped FS stent | 216
fixed stent subcutaneously | 216
regular tracheal cannula introduced | 216
spontaneous breathing work increased | 216
vv-ECMO support reduced | 216
lungs re-aerated | 216
patient woke up | 216
communication with family | 216
infections continued | 216
tidal ventilation of 170 mL per breath | 216
reduction of intravenous saline injection | 216
weaning approaches | 216
decision to reduce vv-ECMO support | 468
death due to pulmonary infection | 468
