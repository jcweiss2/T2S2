70 years old | 0
female | 0
admitted to the intensive care unit | 0
altered sensorium | 0
hypotension | 0
fever | -48
diabetes mellitus type 2 | -6720
essential hypertension | -6720
chronic kidney disease | -6720
hemodialysis | -720
volume overload | -720
worsening renal parameters | -720
tender swellings over both inner thighs and buttocks | -720
punch biopsies declined | -720
confused and disoriented to time, place, and person | 0
no obvious focal neurological deficit | 0
pulse rate 110/min | 0
blood pressure 70/50 mm Hg | 0
SPO2 98% in room air | 0
afebrile | 0
bilateral basal crepitations | 0
violaceous nodules with indurations | 0
retiform purpura | 0
tender to palpation | 0
hemoglobin 6.6 g/dl | 0
total leucocyte count 25.0 thou/cumm | 0
neutrophilic leukocytosis | 0
erythrocyte sedimentation rate 119 mm/1st hour | 0
c-reactive protein 247 mg/L | 0
serum albumin 1.01 g/dl | 0
corrected serum calcium 11.08 mg/dl | 0
serum phosphate 4.95 mg/dl | 0
calcium phosphate product 54.8 | 0
PTH 20.0 pg/ml | 0
creatine phosphokinase 57 U/L | 0
subcutaneous edema | 0
no deep vein thrombosis | 0
subcutaneous fat reticulation | 0
edema | 0
soft tissue changes related to lipodermatosclerosis | 0
metabolically inactive subcutaneous fat stranding | 0
panniculitis | 0
no metabolically active disease | 0
ANA profile negative | 0
p ANCA negative | 0
c ANCA negative | 0
APLA IgM negative | 0
IgG kappa monoclonal band | 0
plasma cell <10% | 0
monoclonal gammopathy of uncertain significance (MGUS) | 0
calciphylaxis | 0
IV antibiotics (meropenem and vancomycin) | 0
antifungal agent (micafungin) | 24
intravenous colistin | 48
sterile blood and urine cultures | 48
calcitonin | 48
zoledronic acid | 48
low calcium dialysate | 48
intravenous vitamin K | 48
punch biopsies | 72
vasculopathic lymphoid infiltrate | 72
focal panniculitis | 72
no specific deposits on diffuse immunofluorescence | 72
intravascular lymphoma | 72
refractory septic shock | 96
intravenous hydrocortisone | 96
deterioration of sensorium | 120
expired | 144