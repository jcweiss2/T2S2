18 years old | 0
male | 0
admitted to the hospital | 0
fever | -72
rash | -72
acne |  -672
minocycline |  -672
increased WBC count | 0
eosinophilia| 0
systemic involvement| 0
diffuse erythematous or maculopapular eruption| 0
pruritis | 0
DRESS syndrome | 0
fever persisted | 0
rash persisted | 0
discharged | 24
DALK | 0
granular dystrophy | -672
deep anterior lamellar keratoplasty | 0
recipient stromal flap partially dissected | -8
air injected into the stroma | -8
donor button cut | -8
donor DM peeled off | -8
donor button sutured | -8
age of donor cornea | -672
donor cornea in situ excision | -672
surgery went well | -8
whitish infiltrates along the graft-host junction | 1
severe anterior chamber reaction | 1
postoperative keratitis | 1
graft removed | 1
replaced by another stromal graft | 1
topical vancomycin started | -3
topical ceftazidime started | -3
Gram-negative Bacilli | 1
intraoperative field contaminated | -8
donor cornea contaminated | -672
residual infectious matter in the recipient cornea | -672
postoperative environment contaminated | -8
multidrug resistant Klebsiella | 1
Klebsiella pneumoniae | 1
imipenem started | 1
infiltrates extended toward center of graft | 4
hypopyon persisted | 4
therapeutic penetrating keratoplasty | 4
infiltrates in host DM | 4
graft clear without infiltrates or hypopyon | 5
imipenem continued | 5
gatifloxacin added | 5
prednisolone drops added | 10
unaided vision 6/60 | 42
unaided vision 6/18 with pin hole | 42
graft clear | 42
anterior segment quiet | 42
intraocular pressure normal | 42
eradication of the pathogen | 42