18 years old | 0
male | 0
obesity | 0
psoriatic arthritis | 0
surgical hypoparathyroidism | 0
hypothyroidism | 0
total thyroidectomy | -20
multinodular goitre | -20
elective sleeve gastrectomy | 0
gastric perforations | 0
emergency Roux-en-Y gastric bypass surgery | 0
abdominal sepsis | 4
transfer to intensive care | 4
nil orally | 4
critically low calcium level | 4
asymptomatic | 4
seizure | -4
arrhythmia | -4
intravenous calcium gluconate infusion | 4
normocalcaemia | 4
prolonged ICU admission | 0
more than 20 abdominal operations | 0
lost 14 kg | 0
intravenous medication and nutrition | 0
endocrinology advice | 0
hypoparathyroidism | 0
hypothyroidism | 0
TSH | 0
5.83 mU/L | 14
intravenous triiodothyronine | 14
euthyroidism | 14
high dose intravenous calcium | 14
ionised calcium | 14
serum phosphate level | 14
1.07 mmol/K | 14
intravenous calcitriol | 14
limited stock | 19
high cost | 19
intramuscular cholecalciferol | 14
1,25(OH)vitamin D3 level | 14
31 pmol/L | 14
renal function | 14
eGFR | 14
> 90 mL/min/1.73 m2 | 14
intravenous calcium gluconate | 14
4.4 mmol five times daily | 14
intravenous calcitriol | 14
1 µg alternate daily | 14
intramuscular thyroxine | 18
600 µg | 18
intravenous thyroxine | 22
200 µg alternate daily | 22
maintenance schedule | 22
hypocalcaemia | 22
hypothyroidism | 22
oral intake | 22
recommence | 22
preoperative calcitriol dose | 22
calcium | 22
1200 mg orally twice daily | 22
normocalcaemia | 22
review | 22
6 weeks | 22
12 weeks | 22
4 months | 22
weighed 71.8 kg | 22
BMI of 29 kg/m2 | 22
calcium replacement | 0
enteral absorption | 0
oral treatment | 0
calcium carbonate | 0
calcitriol | 0
parenteral options | 0
IV Calcitriol | 0
1 µg IV every 4 days | 0
IV Calcium gluconate | 0
4.4 mmol IV 5x daily | 0
Teriparatide | 0
20 µg subcut twice daily | 0
NatPara | 0
50–100 µg subcut daily | 0
hypoparathyroidism | 0
surgical | 0
gastrointestinal disorders | 0
malabsorption | 0
escalating oral doses | 0
gastrostomy tube insertion | 0
pancreatic enzyme supplementation | 0
abdominal sepsis | 0
friable mucosa | 0
gastric bypass surgery | 0
pre-existing hypoparathyroidism | 0
elective bariatric surgery | 0
potential difficulties | 0
managing hypocalcaemia | 0
impaired gastrointestinal absorption | 0
complications | 0
approval of subcutaneous recombinant PTH | 0
hypoparathyroidism in Australia | 0