36 years old | 0
male | 0
admitted to the hospital | 0
snakebite over left foot | -72
anti-snake venom | -72
IV fluids | -72
antibiotics | -72
supportive care | -72
decreased urine output | -48
deranged renal functions | -48
AKI | -48
hemodialysis | -48
brought to our hospital | -24
initial evaluation | 0
stabilization in emergency room | 0
admitted to medical intensive care unit | 0
dull drowsy state | 0
arousable | 0
stable hemodynamic | 0
bilateral decreased air entry | 0
swelling at the site of bite | 0
cellulitis | 0
blister formation | 0
hemoglobin (Hb) 7.6 g/dL | 0
total leucocyte count (TLC) 15,000 | 0
platelets ∼50,000 | 0
normal coagulation profile | 0
aPTT 15 seconds | 0
INR ∼1.19 | 0
bedside clotting time 5 minutes | 0
bleeding time 32 seconds | 0
deranged kidney function tests | 0
urea 167 mg/dL | 0
creatinine 6.17 mg/dL | 0
total CPK ∼52,168 | 0
rhabdomyolysis | 0
transaminitis | 0
SGOT/PT ∼1,985/252 | 0
total bilirubin 4.56 | 0
direct bilirubin 0.64 | 0
indirect bilirubin ∼3.92 | 0
sepsis | 0
procalcitonin 4.79 | 0
oxygen support | 0
intravenous antibiotics | 0
antivenom | 0
acute kidney shutdown | 0
anuric status | 0
hemodialysis | 0
heparin free | 0
ultrafiltration | 0
persistent fall in Hb | 0
multiple blood transfusions | 0
hemolysis | 0
fragmented cells | 0
spherocytes | 0
LDH ∼4,128 | 0
worsening of hypoxemia | 168
bilateral infiltrates on chest X-ray | 168
pleural effusion | 168
HFNC oxygen support | 168
FiO2 requirement 0.4 | 168
hemoptysis | 168
CT chest | 168
multifocal peribronchial air space opacification | 168
ground-glass opacification | 168
moderate pleural effusion | 168
lung collapse | 168
diffuse alveolar hemorrhage | 168
steroids | 168
methylprednisolone 80 mg/day | 168
coagulation profile monitored | 168
INR ∼1.17 | 168
thrombocytopenia recovery | 168
HFNC oxygen support continued | 168
bilateral pleural drain | 168
transudative picture | 168
sterile pleural effusion | 168
echocardiography EF ∼55% | 168
ultrasound abdomen bulky hypoechoic kidneys | 168
reduced CMD | 168
ANA negative | 168
C8-ANCA negative | 168
P-ANCA negative | 168
E. coli in sputum culture | 168
meropenem | 168
no improvement | 168
hemoptysis continued | 168
progressive fall in Hb | 168
persistent AKI | 168
plasma exchange therapy | 480
plasma exchange performed | 480
centrifugation technology | 480
jugular venous access | 480
5% Hum albumin | 480
electrolytes monitoring | 480
fluid balance monitoring | 480
proteins monitoring | 480
coagulation monitoring | 480
improved renal parameters | 480
urine output 25-50 mL/hour | 480
third plex | 504
secondary sepsis | 504
leukocytosis | 504
procalcitonin ∼21 | 504
polymyxin B | 504
elective intubation | 504
type I respiratory failure | 504
five sessions of plasma exchange | 504
intermittent hemodialysis | 504
improved oxygen requirement | 504
settling leukocytosis | 504
renal function improved | 504
creatinine 3.5 mg/dL | 504
urine output 2,100 mL/24 hours | 504
pulmonary hemorrhage settled | 504
minimal tracheal bleed | 504
static Hb | 504
bronchoscopy clear airways | 504
HRCT chest multifocal consolidations | 504
continued antibiotics | 504
supportive care | 504
extubation | 504
low-flow oxygen | 504
hemodynamically stable | 504
clearing infiltrates | 504
residual right basal collapse | 504
discharged | 504
creatinine ∼1.2 | 504
good urine output | 504
cleared chest X-ray | 504
healthy on follow-up | 504
fully recovered AKI | 504
creatinine 0.96 | 504
chest X-ray clear | 504
