65 years old | 0
male | 0
admitted to the hospital | 0
muscular pain in the back of the neck | -144
generalized fatigue | -144
weakness | -144
poor oral intake | -144
loose motion | -144
no weight loss | -144
no significant gastrointestinal symptoms | -144
no cardiorespiratory symptoms | -144
dehydration | 0
jaundice | 0
normal heart sounds | 0
no added murmurs | 0
temperature 39.7 C | 0
increased creatine kinase | 0
troponin T high sensitivity | 0
aspartate aminotransferase | 0
alanine aminotransferase | 0
total bilirubin | 0
direct bilirubin | 0
white blood count | 0
normal chest X-ray | 0
normal ECG | 0
hypertension | 0
diabetes mellitus | 0
chronic renal impairment | 0
obesity | 0
metabolic syndrome | 0
obstructive sleep apnea | 0
cervical and lumbar spondylosis | 0
G6PD deficiency | 0
fever with jaundice | 0
infection-related hepatic dysfunction | 0
hemolytic episode | 0
NSAID treatment | -144
Ceftriaxone | 0
no high temperatures | 24
unconscious | 48
unresponsive | 48
no seizure activity | 48
normal vital signs | 48
normal blood glucose | 48
left hemispheric syndrome | 48
severe hemiparesis | 48
gaze deviation | 48
global aphasia | 48
hemianopia | 48
hypoesthesia | 48
NIHSS score 18 | 48
urgent CT of the brain | 48
no acute changes | 48
left middle cerebral artery ischemic stroke | 48
IV r-tPA | 48
onset to needle 30 min | 48
supervision in ICU | 48
follow-up CT of the brain | 72
new ischemic infarct | 72
no hemorrhagic changes | 72
blood culture positive | 72
Gram-positive Streptococcus species | 72
Gentamicin | 72
bedside TTE | 96
departmental TTE | 96
transesophageal echocardiography | 96
large vegetation | 96
mitral regurgitation | 96
Streptococcus agalactiae | 96
combined therapy | 96
Gentamycin | 96
Vancomycin | 96
follow-up TEE | 576
no fresh vegetations | 576
no abscess | 576
no hemorrhage | 576
no mycotic aneurysms | 576
follow-up CT of the brain | 576
newly developed ischemic area | 576
speech difficulties | 576
right hemiparesis | 576
requiring a cane | 576
discharged | 720