37 years old | 0
male | 0
admitted to the hospital | 0
loss of vision in the left eye | 0
COVID-19 infection | -2160
shortness of breath | -2160
difficulty in breathing | -2160
generalized weakness | -2160
fever | -2160
loss of smell | -2160
loss of taste | -2160
tested for real-time reverse transcription-polymerase chain reaction (RT-PCR) for COVID-19 | -2160
positive RT-PCR | -2160
admitted to the hospital | -2160
inflammatory markers erythrocyte sedimentation rate (ESR) | -2160
C-reactive protein (CRP) | -2160
D-dimers | -2160
ferritin | -2160
interleukin-6 | -2160
Electrocardiogram | -2160
Computed tomography (CT) scan of the chest | -2160
ground-glass opacities with reticulations in bilateral lungs | -2160
viral pneumonia | -2160
condition deteriorated | -2148
shifted to the intensive care unit (ICU) | -2148
intubated | -2148
treated with remdesivir | -2148
treated with azithromycin | -2148
treated with tocilizumab | -2148
plasma transfusion | -2148
supportive care | -2148
recovered from pneumonia | -2136
shifted to the ward | -2136
sudden onset of swelling | -2124
foreign body sensation | -2124
drooping of upper eyelid | -2124
diminution of vision of the left eye | -2124
ophthalmological opinion | -2124
no perception of light | -2124
ptosis | -2124
proptosis | -2124
complete ophthalmoplegia | -2124
severe optic disc edema | -2124
cherry red spot | -2124
retinal whitening | -2124
CRAO | -2124
cavernous sinus thrombosis (CST) | -2124
left diffuse pre-septal and retro-orbital edema | -2124
swollen optic nerve sheath | -2124
asymmetric bulging and filling defect of the left cavernous sinus | -2124
thickened and prominent left optic nerve sheath | -2124
ill-defined soft tissue infiltration at orbital apex | -2124
treated with intravenous steroids | -2112
treated with antibiotics | -2112
treated with anticoagulant | -2112
symptomatic care | -2112
biopsy from the nasal mucosa | -2112
no fungal infection | -2112
discharged | -1080
proptosis recovered | -720
ptosis recovered | -720
ophthalmoplegia recovered | -720
presented with complaints of loss of vision in the left eye | 0
unaided visual acuity of 20/20 on Snellen’s chart | 0
normal color vision | 0
exodeviation of 15° on Hirschberg’s test | 0
grade four relative afferent pupillary defect | 0
anterior segment of both eyes was unremarkable | 0
optic disc atrophy | 0
gliosis | 0
macular pucker | 0
intraocular pressure | 0
applanation tonometry | 0
loss of foveal contour | 0
thinning | 0
hyper-reflective internal limiting membrane | 0
vitreomacular traction | 0
fluid pockets in parafoveal area | 0
visual fields examination | 0
visual evoked potential (VEP) | 0
P100 latency and amplitude | 0
diagnosis of CST with subsequent CRAO and optic neuropathy secondary to COVID 19 infection | 0