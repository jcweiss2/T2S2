31 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
non-smoking | 0 | 0 | Factual
Caucasian | 0 | 0 | Factual
no past medical history | 0 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
sudden-onset severe headache | -840 | -840 | Factual
left arm numbness | -840 | -840 | Factual
cranial computed tomography (CT) scan | -840 | -840 | Factual
grade 2 (Hunt and Hess scale) SAH | -840 | -840 | Factual
no prior history of head injury | 0 | 0 | Factual
uncomplicated pregnancy | 0 | 0 | Factual
uncomplicated vaginal delivery | 0 | 0 | Factual
admitted to the neurosurgical ward | -840 | -840 | Factual
digital subtraction angiography (DSA) | -840 | -840 | Factual
ruptured right middle cerebral artery aneurysm | -840 | -840 | Factual
percutaneous endovascular coil embolization | -840 | -840 | Factual
no permanent neurological deficits | -840 | 0 | Factual
fever | -672 | -672 | Factual
chills | -672 | -672 | Factual
constant abdominal pain | -672 | -672 | Factual
purulent uterine discharge | -672 | -672 | Factual
no urinary symptoms | -672 | -672 | Negated
no respiratory symptoms | -672 | -672 | Negated
blood culture | -672 | -672 | Factual
empiric antibacterial therapy | -672 | -672 | Factual
piperacillin/tazobactam | -672 | -672 | Factual
vancomycin | -672 | -672 | Factual
azithromycin | -672 | -672 | Factual
sepsis | -640 | -640 | Factual
septic shock | -640 | -640 | Factual
transferred to the intensive care unit | -640 | -640 | Factual
body temperature 38.3 °C | -640 | -640 | Factual
invasive blood pressure 90/65 mmHg | -640 | -640 | Factual
heart rate 135/min | -640 | -640 | Factual
arterial oxygen saturation 82 % | -640 | -640 | Factual
mild disorientation | -640 | -640 | Factual
slower capillary refill | -640 | -640 | Factual
coarse rales | -640 | -640 | Factual
sequential organ failure assessment (SOFA) score 4 | -640 | -640 | Factual
hemoglobin 6.8 g/dL | -640 | -640 | Factual
d-dimers 4.58 μg/mL | -640 | -640 | Factual
C-reactive protein 322 mg/L | -640 | -640 | Factual
fibrinogen concentration 6.4 mL | -640 | -640 | Factual
blood culture showed E. coli | -640 | -640 | Factual
E. coli sensitive to piperacillin/tazobactam | -640 | -640 | Factual
chest radiography | -640 | -640 | Factual
pulmonary nodules | -640 | -640 | Factual
CT of the thorax | -640 | -640 | Factual
metastatic lung nodules | -640 | -640 | Factual
transvaginal ultrasound | -640 | -640 | Factual
enlarged uterus | -640 | -640 | Factual
complete loss of zonal anatomy | -640 | -640 | Factual
abdominal magnetic resonance imaging (MRI) | -640 | -640 | Factual
enlarged heterogenous myometrial mass | -640 | -640 | Factual
splenic metastatic lesion | -640 | -640 | Factual
serum β-human chorionic gonadotrophin (β-hCG) 232,085 mUI/mL | -640 | -640 | Factual
suction evacuation and curettage | -640 | -640 | Factual
pathology report confirmed choriocarcinoma | -640 | -640 | Factual
International Federation of Gynecology and Obstetrics (FIGO) modified WHO prognostic scoring system | -640 | -640 | Factual
total score of 12 | -640 | -640 | Factual
high risk of developing resistance to single-drug chemotherapy | -640 | -640 | Factual
multiagent chemotherapy regimen | -640 | -640 | Factual
low-dose etoposide | -640 | -640 | Factual
cisplatin | -640 | -640 | Factual
EMA/CO regimen | -608 | -608 | Factual
etoposide | -608 | -608 | Factual
methotrexate | -608 | -608 | Factual
actinomycin D | -608 | -608 | Factual
cyclophosphamide | -608 | -608 | Factual
vincristine | -608 | -608 | Factual
six cycles of EMA/CO | -608 | 0 | Factual
β-hCG levels plateaued | 0 | 0 | Factual
restaging with MRI of the brain | 0 | 0 | Factual
18F-fluorodeoxyglucose (FDG) positron emission tomography (PET)/CT scan | 0 | 0 | Factual
decreased pulmonary nodules | 0 | 0 | Factual
decreased uterine mass | 0 | 0 | Factual
low standardized uptake value (SUV) | 0 | 0 | Factual
revised FIGO score 7 | 0 | 0 | Factual
EP/EMA regimen | 0 | 0 | Factual
normalization of β-hCG | 168 | 168 | Factual
grade 3 neutropenia | -112 | -112 | Factual
granulocyte colony stimulating factor (G-SCF) | -112 | -112 | Factual
dose reduction of etoposide and actinomycin D | -112 | -112 | Factual
grade 2 alopecia | -112 | -112 | Factual
grade 2 nausea | -112 | -112 | Factual
dexamethasone | -112 | -112 | Factual
ondansetron | -112 | -112 | Factual
grade 2 fatigue | 0 | 0 | Factual
male condoms | 0 | 0 | Factual
follow-up | 0 | 504 | Factual
alive 21 months post diagnosis | 504 | 504 | Factual