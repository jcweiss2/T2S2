66 years old | 0
female | 0
smoker | 0
admitted to the hospital | 0
hypotension | 0
referred to the emergency department | 0
colonoscopy | -504
removal of two serrated polyps | -504
from the descending colon | -504
generalized weakness | -336
fatigue | -336
blood pressure of 60/30 mm Hg | -336
sent to the ED | -336
confused | 0
lethargic | 0
fever for the past 5 days | -120
temperature of 98.1 °F | 0
blood pressure of 74/45 mm Hg | 0
heart rate of 99 beats/min | 0
respiratory rate of 18 breaths/min | 0
conjunctivae were pink | 0
no signs of jaundice | 0
lungs were clear to auscultation bilaterally | 0
heart sounds were audible with no murmurs, rubs, or gallops | 0
abdominal examination revealed diffuse abdominal tenderness | 0
bilateral costovertebral angle tenderness | 0
bowel sounds were present in all four quadrants | 0
WBC count of 28,700/mm3 | 0
left shift | 0
normocytic anemia | 0
hemoglobin level of 8.3 g/dL | 0
liver and renal profiles within the normal physiological ranges | 0
2-L intravenous bolus of normal saline | 0
blood pressure raised to 105/60 mm Hg | 0
blood and urine cultures were obtained | 0
started on ceftriaxone | 0
transferred to the medical intensive care unit | 0
contrast-enhanced computed tomography of the abdomen and pelvis | 0
multiple hepatic and perihepatic fluid collections | 0
suspicious of abscesses | 0
extension under the 12th rib and the lower right flank | 0
loculated fluid collection in the right lower quadrant | 0
other smaller fluid collections | 0
interventional radiology and surgery were urgently consulted | 0
four intraabdominal drains were placed | 0
750 cc of pus was drained | 0
pus was sent to the laboratory for culture | 0
ceftriaxone was discontinued | 24
started on IV meropenem, vancomycin, and metronidazole | 24
culture of the pus showed a heavy growth of Streptococcus constellatus | 72
meropenem and vancomycin were discontinued | 72
started on ceftriaxone in addition to metronidazole | 72
marked improvement in the clinical state of the patient | 72
more alert | 72
improved appetite | 72
decreased abdominal tenderness | 72
marked improvement in her WBC count | 168
decrease in the quantity of fluid being drained from the abdomen | 168
less than 10 cc drained per 24-h period | 168
repeat CT scan of the abdomen and pelvis | 168
marked decrease in the intraabdominal abscess | 168
small residual collection, 2 cm in size, located in the segment 4a of the liver | 168
three out of the four drains were removed | 168
drain in the dome of the liver was left in place | 168
last drain was removed | 336
peripherally inserted central catheter was placed | 336
patient was discharged | 336
repeat of CT of abdomen and pelvis 4 weeks later | 672
complete resolution of the abscesses | 672