27 years old | 0
man | 0
admitted to the hospital | 0
pancytopenia | 0
neutrophils: 0.8×109/L | 0
hemoglobin: 9.4 gr/dl | 0
platelets: 4×109/L | 0
muco-cutaneous hemorrhages | 0
severe aplastic anemia | 0
empirical broad spectrum antibiotherapy | 120
piperacillin–tazobactam | 120
amikacin | 120
febrile neutropenia | 120
fever | 120
fever resolved | 120
oral prednisone | 288
admitted to the intensive care unit | 456
septic shock | 456
prednisone stopped | 456
piperacillin-tazobactam restarted | 480
levofloxacin | 480
recovered | 576
admitted to hematology unit | 576
central venous catheter inserted | 600
fever reappeared | 696
fever persisted | 696
poor clinical condition | 696
diarrhea | 696
abdominal pain | 696
dry cough | 696
left thoracic pain | 696
diffuse bowel thickening | 744
normal liver function tests | 744
CVC removed | 744
left blurred vision | 744
cerebral CT scan normal | 744
cerebral magnetic resonance imaging normal | 744
retinal hemorrhage | 744
echocardiogram excluded fungal endocarditis | 744
clinical condition improved | 792
weekly stool examinations negative | 792
daily blood cultures negative | 792
fever persisted | 1008
no documented infection | 1008
negative galactomannan antigenemia | 1008
allogeneic bone marrow transplantation | 1008
cyclosporine started | 1008
fever resolved | 1008
good clinical condition | 1008
voriconazole replaced by posaconazole | 2016
nausea and vomiting | 2016
liposomal amphotericin B discontinued | 2016
left hospital | 2112
posaconazole secondary prophylaxis | 2112
fever resolved | 2112
vision normalized | 2112
no recurrence of infection | 4-month follow-up
no complications of transplantation | 4-month follow-up
