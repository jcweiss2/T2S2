26 years old | 0
    male | 0
    admitted to the hospital | 0
    generalized abdominal pain | -2160
    infrequent watery diarrhea | -2160
    acute hepatitis A | -2160
    increased liver enzymes | -2160
    high HAV IgG Ab | -2160
    abdominal pain not resolved | -2160
    pain radiating to flanks | -2160
    pain aggravating after food ingestion | -2160
    bloody diarrhea episode | -720
    night sweats | -720
    significant weight loss | -720
    epigastric abdominal pain | 0
    infrequent nausea | 0
    vomiting | 0
    watery diarrhea continued | 0
    past history negative | 0
    no smoking | 0
    no addiction | 0
    stable vital signs | 0
    mild epigastric tenderness | 0
    splenomegaly 14 cm span | 0
    abdominal ultrasonography unremarkable | 0
    moderate splenomegaly | 0
    stool exam RBC | 0
    stool exam no WBC | 0
    gastroenterologist consultation | 0
    rheumatologist consultation | 0
    upper gastrointestinal endoscopy chronic gastritis | 0
    histopathology colon biopsy inflammatory bowel disease | 0
    worsened symptoms | 0
    fever | 0
    several episodes bloody diarrhea | 0
    treated with Mesalazine | 0
    treated with Asacol enema | 0
    treated with antibiotics | 0
    peripheral blood smear aggregated platelets | 0
    Doppler ultrasound portal vein increased diameter 16 mm | 0
    Doppler ultrasound splenic vein increased diameter 11 mm | 0
    Doppler ultrasound normal flow | 0
    Doppler ultrasound normal spectral waves | 0
    Doppler ultrasound normal patency superior mesenteric artery | 0
    abdominopelvic computed tomography mesenteric fat stranding | 0
    abdominopelvic computed tomography thick-walled bowels | 0
    abdominopelvic computed tomography portal vein thrombosis | 0
    abdominopelvic computed tomography superior mesenteric vein thromboses | 0
    intolerable abdominal pain | 0
    diarrhea continued | 0
    generalized tenderness | 0
    rebound tenderness | 0
    guarding | 0
    significant thrombocytopenia 22000 | 0
    peripheral blood smear check | 0
    fibrinogen check | 0
    fibrin degradation products check | 0
    thrombocytopenia corrected | 0
    laparotomy | 0
    laparotomy revealed bloody ascites | 0
    laparotomy revealed colon necrosis | 0
    total colectomy | 0
    ileostomy performed | 0
    histopathology colon necrosis | 0
    histopathology intraluminal thrombosis vascular canals | 0
    critically ill | 48
    hypotension | 48
    dyspnea | 48
    abnormal coagulation studies | 48
    no schistocyte | 48
    thrombocytopenia | 48
    elevated fibrinogen | 48
    elevated fibrin degradation products | 48
    treated with fresh frozen plasma | 48
    died | 48
    Factor V Leiden | 48
    antiphospholipid syndrome | 48
    portal system thrombosis | 48
    
    