76 years old | 0
female | 0
metastatic lung adenocarcinoma | -2160
invasive ductal carcinoma of the right breast | -672
lumpectomy | -672
aromatase inhibitor | -672
20 pack-year tobacco use history | -84000
ceased smoking | -84000
recently traveled to the Southwest United States | -168
no known occupational or environmental exposures | 0
no history of chest radiation | 0
lung cancer diagnosed | -2160
hypoxemia on exertion | -2160
computed tomography showed a right upper lobe mass | -2160
lung and liver metastases | -2160
biopsy of the lung and liver | -2160
metastatic adenocarcinoma | -2160
no actionable mutations | -2160
palliative systemic therapy with carboplatin, pemetrexed, and pembrolizumab | -2160
imaging showed stable disease | -1344
fevers | -72
dyspnea on exertion | -72
cough | -72
CT angiogram of the chest | -72
no pulmonary embolism | -72
confluent regions of consolidation in the lungs bilaterally | -72
small left pleural effusion | -72
bilateral cavitary lung lesions | -72
admitted to the intensive care unit | 0
severe hypoxemic respiratory failure | 0
PaO2/FiO2 ratio of 87 | 0
treated with broad-spectrum antibiotics | 0
worsening hypoxemia on day three | 72
endotracheal intubation | 72
mechanical ventilation | 72
positive end-expiratory pressure titrated | 72
lung protective ventilation | 72
bronchoscopy on day three | 72
thin secretions in the left lower lobe | 72
bronchoalveolar lavage studies | 72
slight neutrophilic predominance | 72
negative microbiology studies | 72
transthoracic echocardiogram | 72
mild symmetric left ventricular hypertrophy | 72
normal right ventricular size and systolic function | 72
no significant valvular disease | 72
no signs of increased filling pressures | 72
no atrial septal defect | 72
invasive diagnostic procedures deferred | 72
immune checkpoint inhibitor pneumonitis suspected | 72
intravenous methylprednisolone | 72
significant desaturations despite treatment | 216
intravenous immunoglobulin | 216
rapid and significant clinical and radiographic improvement | 288
successful extubation | 288
repeat chest CT imaging | 288
marked improvement in severe interstitial abnormality | 288
transitioned to prednisone | 336
supplemental oxygen requirement decreased | 336
weaned to an oxymizer device | 336
discharged | 552
oxygen needs decreased | 1008
exercise tolerance improved | 1008
prednisone decreased | 1008
re-staging CT of the torso | 1008
continued improvement of the predominantly left-sided infiltrate | 1008
remaining bilateral subpleural interstitial fibrotic abnormality | 1008
malignant disease burden stable | 1008