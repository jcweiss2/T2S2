44 years old | 0
obese | 0
woman | 0
inhalation injury | 0
second-to-third degree burn injury | 0
32% total body surface area | 0
referred from previous hospital | 0
burn injury on mucous membranes of lips | 0
burn injury on mucous membranes of mouth | 0
burn injury on mucous membranes of eyes full of edema | 0
intubated with endotracheal tube no 6.5 | 0
depth of placement 22 cm from central incisors | 0
fixed with thread on right lip corner | 0
spontaneous symmetrical breathing | 0
respiratory rate 20 per minute | 0
SpO2 100% with T-piece 10 lpm | 0
blood pressure 128/79 mmHg | 0
heart rate 98 per minute | 0
warm extremities | 0
capillary refill time <2 seconds | 0
no spontaneous bleeding | 0
head and neck edema | 0
burn status head neck 5% | 0
burn status anterior trunk 5% | 0
burn status right arm 9% | 0
burn status left arm 6% | 0
burn status left leg 3% | 0
burn status back 4% | 0
nasogastric tube insertion | 0
brownish fluid obtained | 0
high leucocytes 28880 103/µl | 0
blood glucose 242 mg/dL | 0
low albumin 2.5 gr/dL | 0
sputum culture from tracheal secretions revealed Acinetobacter baumanii | 0
treated with tigecycline | 0
grade II-III burn injury 32% total body surface area | 0
stress ulcer | 0
leucocytosis | 0
treated in ICU | 0
early tracheostomy performed | 0
percutaneous dilatational tracheostomy performed | 0
locating trachea with 10cc syringe | 0
syringe showed signs of air bubble | 0
no bleeding occurred | 0
1-cm incision between second and third tracheal ring | 0
ventilator set to PSV/CPAP PS 10 Peep 5 trig 3 FiO2 50% | 0
intubated successfully | 0
treated in ICU from 23rd February to 2nd March 2022 | 0
percutaneous dilatational tracheostomy to facilitate sputum passage | 0
avoiding ETT obstruction | 0
tangential excision | 0
debridement | 0
PDT performed prior to debridement | 0
maintain patient’s airway | 0
provide easier access for debridement | 0
mouth area heavily plastered | 0
using ETT | 0
25% plasbumin transfusion 100 ml for 2 days | 0
PDT done to secure airway | 0
avoid ETT obstruction due to sputum hypersecretion | 0
length of ventilator day 5 days | 0
discharged from ICU after 7 days | 0
moved to normal ward | 0
still cannulated | 0
able to breathe spontaneously | 0
kept PDT after discharge from ICU | 0
better management of secretions | 0
avoid aspiration | 0
discharged after 2 weeks in normal ward | 0
referred back to first hospital | 0
no follow-up for Pseudomonas infection at PDT site | 0
facial burns | 0
singed facial or nasal hair | 0
soot or carbonaceous material on face | 0
soot or carbonaceous material in sputum | 0
airway blockage signs | 0
inhalation injury confirmed | 0
cost constraints preventing further testing | 0
severe swelling of tongue | 0
severe swelling of epiglottis | 0
severe swelling of aryepiglottic folds | 0
restricted breathing | 0
production of edema due to reactive oxygen species | 0
increased permeability to proteins | 0
fluid resuscitation | 0
airway edema developed | 0
upper airway anatomically distorted | 0
upper airway externally compressed | 0
affect airway care | 0
PDT done early to prevent complications | 0
PDT complications | 0
PDT-related death risk | 0
serious bleeding incidents | 0
unrecognized anatomical variations | 0
unanticipated anatomical variations | 0
use of ultrasound not accessible | 0
PDT performed without ultrasound guidance | 0
early PDT within 18 hours after incident | 0
complicating factors obesity | 0
complicating factors short neck | 0
difficulty finding surgical incision site | 0
patient demonstrated good outcome | 0
low mortality risk | 0
treated on ventilator for 5 days | 0
no pulmonary infections | 0
incision site healed well | 0
moved to medical ward after 7 days in ICU | 0
discharged from hospital | 0
securing airway prioritized | 0
conventional ETT not best option | 0
susceptible to clotting | 0
obstruction due to excessive secretions | 0
PDT chosen over traditional tracheostomy | 0
less invasive | 0
lower complication rate | 0
faster recovery time | 0
early PDT to avoid complications | 0
better outcome | 0
