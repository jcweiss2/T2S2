56 years old | 0
female | 0
admitted to the hospital | 0
abdominal pain | -120
long-standing smoker | 0
no previously diagnosed chronic medical conditions | 0
no recent exposure to any sick contacts | 0
upper respiratory tract infection | -336
tachycardic | 0
hypertensive | 0
afebrile | 0
soft but tender abdomen | 0
white blood cell count elevated | 0
CT angiography of the abdomen and pelvis | 0
infrarenal aortic aneurysm | 0
periaortic hematoma | 0
renal arteries and visceral vessels displayed mild atheromatous changes | 0
blood cultures drawn | 0
ciprofloxacin initiated | 0
cefazolin initiated | 0
emergent open repair | 0
edematous retroperitoneum | 0
adherent duodenum | 0
inflammatory changes in the aorta | 0
periaortic fluid sent for Gram stain | 0
Gram stain reported as moderate polymorphs with no organisms seen | 0
in situ aorto-bi-iliac 12 mm × 7 mm Hemashield graft | 0
transferred to the intensive care unit | 0
continued on ciprofloxacin and cefazolin | 0
acute occlusion of the graft | 24
second surgery | 24
extensive thrombectomy of both limbs of the graft | 24
left iliofemoral bypass | 24
increasing pressors to maintain hemodynamics | 24
antibiotics broadened to include meropenem, vancomycin and fluconazole | 24
hemodialysis for renal failure | 24
culture results from the aneurysm sac reported | 96
aneurysm sac infected with Haemophilus influenzae type B | 96
CT scan revealed evidence of free air under the diaphragm | 456
exploratory laparotomy | 456
perforated colon | 456
gross graft contamination with stool and pus | 456
subtotal colectomy | 456
creation of an end-ileostomy | 456
graft heavily irrigated | 456
bilateral axillofemoral grafts placed | 480
explantation of the infected graft | 480
bowel noted to be edematous and friable | 480
inadvertent enterotomies | 480
tracheostomy | 480
prolonged ventilation | 480
new-onset lumbar plexopathy | 480
recovered slowly | 1968
discharged to the floor from ICU | 1968
antibiotics discontinued | 2184
discharged to her home hospital for planned rehabilitation | 2880