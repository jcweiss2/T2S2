72 years old | 0
male | 0
type-2 diabetes | -8760
diabetic micro- and macro-vascular complications | -8760
painful, red, swollen and hyperthermic left lower leg | -72
admitted to hospital | 0
hemodynamically stable | 0
left foot and lower leg badly swollen and tender | 0
interdigital spaces showed macerated skin with fissures | 0
foot pulses not palpable | 0
ankle brachial index (ABI) 0.8 bilaterally | 0
pallanaesthesia | 0
reduced monofilament sensation | 0
ear-temperature 37.6°C | 0
BP 161/86 mmHg | 0
pulse 96/min | 0
high inflammatory markers | 0
CRP 182 mg/L | 0
leukocytes 15.2 g/L | 0
eGFR 80 mL/min/1.73 m2 | 0
HbA1c 90 mmol/mol | 0
x-ray showed normal osseous structures | 0
minimal effusion in the left upper ankle joint | 0
MRI showed unspecific bone marrow oedema | 0
antibiotic therapy changed to Amoxicillin/clavulanic acid | 24
discharged | 168
presented to different hospital | 168
complaining of acute pain in both distal legs | 168
significant bilateral lower extremity oedema | 168
inflammatory signs restricted to the left lower leg | 168
afebrile | 168
hemodynamically stable | 168
mildly elevated CRP | 168
leucocytes within normal limits | 168
cellulitis of the left lower extremity diagnosed | 168
i.v. antibiotics started | 168
painless second-degree ulcer developed | 168
lateral of the right fifth metatarso-phalangeal (MTP) joint | 168
no clinical signs of infection | 168
concomitant cardiac decompensation | 168
treated with diuretics | 168
x-ray and MRI ruled out osteomyelitis | 168
visibly calcified pedal arteries | 168
more comprehensive vascular review ordered | 168
markedly reduced toe pressures | 168
pathologic pulse wave forms | 168
significantly compromised arterial blood flow | 168
confirmed by bilateral angiography | 168
percutaneous transluminal angioplasty | 168
cardiac recompensation | 168
clinical improvement | 168
discharged | 336
referred to diabetic foot clinic | 336
adequate wound management | 336
offloading | 336
lesion lateral to MTP fifth joint on right did not show progress | 336
complaining about severe pain in left foot | 336
moderate swelling and hyperthermia | 336
no obvious pathology detected | 336
progressive deformity of left ankle joint | 504
ulcerous lesion with purulent drainage | 504
large wound cavity | 504
x-ray confirmed destruction and dislocation of upper ankle joint | 504
hospitalized | 504
assigned to complete bed rest | 504
antibiotic therapy with Co-Amoxicillin | 504
blood cultures showed staphylococcus aureus bacteraemia | 504
antibiotic regimen changed to Cefazolin | 504
acute kidney injury | 504
hemodynamic dysfunction | 504
acute toxic nephritis secondary to Co-Amoxicillin | 504
below knee amputation | 504
rejected by patient | 504
agreed to surgery two weeks later | 518
surgery uneventful | 518
multiorgan dysfunction syndrome developed | 524
died on April 11th, 2019 | 524