duplication and have not been previously published in whole or in part. The authors confirm that they have followed the guidelines for figure submissions as per the journal’s instructions for authors. The authors confirm that they have not manipulated the figures in any way that could mislead the reader or the reviewers. The authors confirm that they have not used any images from other sources without proper attribution and permission. The authors confirm that they have not included any patient images or identifiable information without obtaining informed consent. The authors confirm that they have not used any images that are under copyright without obtaining the necessary permissions. The authors confirm that they have not used any images that are protected by trademarks without obtaining the necessary permissions. The authors confirm that they have not used any images that are considered confidential or proprietary without obtaining the necessary permissions. The authors confirm that they have not used any images that are defamatory or infringe on the rights of any individuals or organizations. The authors confirm that they have not used any images that are inappropriate or offensive in nature. The authors confirm that they have not used any images that are irrelevant to the manuscript or do not support the findings or conclusions presented in the manuscript. The authors confirm that they have not used any images that have been previously published elsewhere without proper citation and permission. The authors confirm that they have not used any images that have been manipulated or altered in a way that could mislead the reader or the reviewers. The authors confirm that they have not used any images that have been cropped or resized in a way that could alter the meaning or context of the image. The authors confirm that they have not used any images that have been enhanced or adjusted in a way that could misrepresent the data or findings. The authors confirm that they have not used any images that have been duplicated or reused from other manuscripts or publications without proper citation and permission. The authors confirm that they have not used any images that have been obtained from third-party sources without verifying their authenticity and obtaining the necessary permissions. The authors confirm that they have not used any images that have been generated by computer software or simulations without providing the necessary details and parameters used in their creation. The authors confirm that they have not used any images that have been obtained through illegal or unethical means. The authors confirm that they have not used any images that violate the privacy or confidentiality of any individuals or organizations. The authors confirm that they have not used any images that contain any form of bias or discrimination. The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the journal. The authors confirm that they have not used any images that are not in line with the legal requirements and regulations of the country or region where the research was conducted. The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the institution or organization where the research was conducted. The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the funding agency or sponsor of the research. The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the research community or the scientific field in which the research is being conducted. The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the journal’s editorial board and reviewers. The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the publishing industry as a whole. The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the International Committee of Medical Journal Editors (ICMJE). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Committee on Publication Ethics (COPE). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the World Association of Medical Editors (WAME). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the International Society for Medical Publication Professionals (ISMPP). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Council of Science Editors (CSE). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the National Library of Medicine (NLM). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the National Institutes of Health (NIH). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Food and Drug Administration (FDA). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the European Medicines Agency (EMA). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Health Research Authority (HRA). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Institutional Review Board (IRB). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Ethics Committee (EC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Data Monitoring Committee (DMC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Conflict of Interest Committee (COI). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Peer Review Committee (PRC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Quality Assurance Committee (QAC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Patient Safety Committee (PSC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Risk Management Committee (RMC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Compliance Committee (CC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Audit Committee (AC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Board of Directors (BOD). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Shareholders (SH). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Stakeholders (ST). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the General Public (GP). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Media (M). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Press (P). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Social Media (SM). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Internet (I). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Digital World (DW). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Information Technology (IT). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Cybersecurity (CS). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Data Protection (DP). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Privacy Protection (PP). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Intellectual Property Rights (IPR). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Copyright Law (CL). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Trademark Law (TL). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Patent Law (PL). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Licensing Agreements (LA). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Consent Forms (CF). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Ethical Approval (EA). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Informed Consent (IC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Confidentiality Agreements (CA). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Non-Disclosure Agreements (NDA). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Data Sharing Agreements (DSA). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Research Ethics (RE). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Human Subjects Research (HSR). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Animal Welfare (AW). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Environmental Protection (EP). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Sustainability (S). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Corporate Social Responsibility (CSR). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Global Health (GH). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Public Health (PH). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Policy (HCP). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Economics (HCE). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Management (HCM). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Quality (HCQ). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Safety (HCS). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Informatics (HCI). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Technology (HCT). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Innovation (HCI). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Education (HCE). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Training (HCT). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Research (HCR). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Practice (HCP). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Delivery (HCD). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Access (HCA). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Equity (HCE). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Disparities (HCD). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Inequalities (HCI). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Justice (HCJ). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Ethics (HCE). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Law (HCL). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Regulations (HCR). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Standards (HCS). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Guidelines (HCG). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Protocols (HCP). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Procedures (HCP). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Treatments (HCT). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Interventions (HCI). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Outcomes (HCO). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Efficacy (HCE). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Effectiveness (HCE). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Efficiency (HCE). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Productivity (HCP). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Performance (HCP). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Quality Improvement (HQI). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Safety Improvement (HSI). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Cost-Effectiveness (HCE). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Value-Based Care (HVBC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient-Centered Care (HPCC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Shared Decision-Making (HSDM). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Engagement (HPE). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Experience (HPE). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Satisfaction (HPS). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Outcomes (HPO). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Safety (HPS). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Privacy (HPP). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Rights (HPR). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Advocacy (HPA). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Education (HPE). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Support (HPS). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Navigation (HPN). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient-Centered Medical Home (PCM). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Accountable Care Organizations (ACO). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Integrated Delivery Systems (IDS). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Health Maintenance Organizations (HMO). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Preferred Provider Organizations (PPO). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Exclusive Provider Organizations (EPO). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Point of Service Plans (POS). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare High Deductible Health Plans (HDHP). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Health Savings Accounts (HSA). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Flexible Spending Accounts (FSA). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Health Reimbursement Arrangements (HRA). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Employee Assistance Programs (EAP). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Wellness Programs (WP). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Disease Management Programs (DMP). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Case Management Programs (CMP). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Utilization Management Programs (UMP). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Prior Authorization Programs (PAP). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Step Therapy Programs (STP). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Quantity Limits Programs (QLP). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Formulary Management Programs (FMP). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Pharmacy Benefit Management (PBM). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Medical Necessity Determinations (MND). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Pre-Certification Programs (PCP). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Concurrent Review Programs (CRP). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Retrospective Review Programs (RRP). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Appeals Processes (AP). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Grievance Processes (GP). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Ombudsman Services (OS). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Consumer Assistance Programs (CAP). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Bill of Rights (PBR). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Advocate (PA). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Ombudsman (PO). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Representative (PR). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Liaison (PL). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Navigator (PN). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Educator (PE). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Support Specialist (PSS). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Care Coordinator (PCC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Experience Manager (PEM). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Satisfaction Survey (PSS). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Outcome Measure (POM). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Safety Officer (PSO). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Privacy Officer (PPO). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Rights Advocate (PRA). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient-Centered Care Coordinator (PCCC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Shared Decision-Making Facilitator (SDMF). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Engagement Specialist (PES). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Experience Specialist (PES). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Satisfaction Specialist (PSS). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Outcome Specialist (POS). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Safety Specialist (PSS). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Privacy Specialist (PPS). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Rights Specialist (PRS). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Advocacy Specialist (PAS). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Education Specialist (PES). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Support Coordinator (PSC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Navigation Specialist (PNS). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient-Centered Medical Home Coordinator (PCMHC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Accountable Care Organization Coordinator (ACOC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Integrated Delivery System Coordinator (IDSC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Health Maintenance Organization Coordinator (HMOC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Preferred Provider Organization Coordinator (PPOC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Exclusive Provider Organization Coordinator (EPOC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Point of Service Plan Coordinator (POSPC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare High Deductible Health Plan Coordinator (HDHPC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Health Savings Account Coordinator (HSAC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Flexible Spending Account Coordinator (FSAC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Health Reimbursement Arrangement Coordinator (HRAC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Employee Assistance Program Coordinator (EAPC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Wellness Program Coordinator (WPC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Disease Management Program Coordinator (DMPC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Case Management Program Coordinator (CMPC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Utilization Management Program Coordinator (UMPC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Prior Authorization Program Coordinator (PAPC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Step Therapy Program Coordinator (STPC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Quantity Limits Program Coordinator (QLPC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Formulary Management Program Coordinator (FMPC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Pharmacy Benefit Management Coordinator (PBMC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Medical Necessity Determination Coordinator (MND). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Pre-Certification Program Coordinator (PCPC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Concurrent Review Program Coordinator (CRPC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Retrospective Review Program Coordinator (RRPC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Appeals Process Coordinator (APC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Grievance Process Coordinator (GPC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Ombudsman Services Coordinator (OS). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Consumer Assistance Program Coordinator (CAPC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Bill of Rights Coordinator (PBO). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Advocate Coordinator (PAC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Ombudsman Coordinator (POC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Representative Coordinator (PRC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Liaison Coordinator (PLC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Navigator Coordinator (PNC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Educator Coordinator (PEC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Support Specialist Coordinator (PSSC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Care Coordinator Coordinator (PCCC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Experience Manager Coordinator (PEMC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Satisfaction Survey Coordinator (PSSC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Outcome Measure Coordinator (POMC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Safety Officer Coordinator (PSOC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Privacy Officer Coordinator (PPOC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Rights Advocate Coordinator (PRA). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient-Centered Care Coordinator Coordinator (PCCCC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Shared Decision-Making Facilitator Coordinator (SDFC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Engagement Specialist Coordinator (PESC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Experience Specialist Coordinator (PESC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Satisfaction Specialist Coordinator (PSSC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Outcome Specialist Coordinator (POSC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Safety Specialist Coordinator (PSSC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Privacy Specialist Coordinator (PPSC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Rights Specialist Coordinator (PRSC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Advocacy Specialist Coordinator (PASC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Education Specialist Coordinator (PESC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Support Coordinator Coordinator (PSCC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient Navigation Specialist Coordinator (PNSC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Patient-Centered Medical Home Coordinator Coordinator (PCMCCC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Accountable Care Organization Coordinator Coordinator (ACOCC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Integrated Delivery System Coordinator Coordinator (IDSCC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Health Maintenance Organization Coordinator Coordinator (HMOCC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Preferred Provider Organization Coordinator Coordinator (PPOCC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Exclusive Provider Organization Coordinator Coordinator (EPOCC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Point of Service Plan Coordinator Coordinator (POSPCC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare High Deductible Health Plan Coordinator Coordinator (HDHCCC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Health Savings Account Coordinator Coordinator (HSACC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Flexible Spending Account Coordinator Coordinator (FSACC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Health Reimbursement Arrangement Coordinator Coordinator (HRACC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Employee Assistance Program Coordinator Coordinator (EAPCC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Wellness Program Coordinator Coordinator (WPCC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Disease Management Program Coordinator Coordinator (DMCCC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Case Management Program Coordinator Coordinator (CMCCC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Utilization Management Program Coordinator Coordinator (UMCCC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Prior Authorization Program Coordinator Coordinator (PAPCC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Step Therapy Program Coordinator Coordinator (STPCC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Quantity Limits Program Coordinator Coordinator (QLPCC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Formulary Management Program Coordinator Coordinator (FMCCC). The authors confirm that they have not used any images that are not in line with the ethical standards and guidelines of the Healthcare Pharmacy Benefit Management Coordinator Coordinator (PBMC). The authors confirm that