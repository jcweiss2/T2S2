86 years old | 0
    female | 0
    right hip replacement | -34560
    brought to emergency room | 0
    altered mental status | 0
    not feeling well | -48
    last hospital visit (orthopedic admission) | -34560
    no history of alcohol use | 0
    no history of smoking | 0
    no history of recreational drug use | 0
    denied specific dietary pattern | 0
    no history of numbness | 0
    no history of tingling | 0
    no history of difficulty in walking | 0
    no history of alteration in bowel habit | 0
    no history of alteration in bladder habit | 0
    no history of weight loss | 0
    no history of gastric surgery | 0
    no history of small bowel surgery | 0
    first episode of such symptoms | 0
    not taking any medication | 0
    no significant family history | 0
    intubated in ER | 0
    respiratory distress | 0
    altered mental status | 0
    tachycardia | 0
    tachypnea | 0
    pulse 110 bpm | 0
    blood pressure 148/100 mm Hg | 0
    respiratory rate 32 per minute | 0
    oxygen saturation 80% | 0
    dehydrated | 0
    no evidence of trauma | 0
    rapid shallow respiration | 0
    wheezing | 0
    mild pedal edema | 0
    WBC count 6.5×10³ per µL | 0
    hemoglobin 3.2 gm/dL | 0
    hematocrit 9.6% | 0
    MCV 127 fL | 0
    platelets 59×10³ per µL | 0
    retic count 7.5% | 0
    corrected retic 1.6% | 0
    LDH 7077 IU/L | 0
    haptoglobin 14 mg/dL | 0
    serum electrolytes within normal limits | 0
    arterial blood gas showing severe metabolic acidosis | 0
    high anion gap 29 mmol/L | 0
    BUN 34 mg/dL | 0
    creatinine 1.9 mg/dL | 0
    serum glucose 93 mg/dL | 0
    osmolality 308 mOsm/L | 0
    lactic acid 20.3 mmol/L | 0
    hyperbilirubinemia | 0
    total bilirubin 3.7 mg/dL | 0
    direct bilirubin 1 mg/dL | 0
    aspartate transaminase 51 IU/L | 0
    alanine transaminase 22 IU/L | 0
    alkaline phosphatase 41 IU/L | 0
    BNP 670 pg/mL | 0
    troponin negative | 0
    INR elevated 2.48 | 0
    PT 29 s | 0
    aPTT 24 s | 0
    toxicology screen negative for ethylene glycol | 0
    toxicology screen negative for salicylates | 0
    toxicology screen negative for alcohol | 0
    serum ketones negative | 0
    imaging scans negative | 0
    mild cardiomegaly | 0
    CT head negative | 0
    CT abdomen negative | 0
    CT PE protocol negative | 0
    admitted to ICU | 0
    altered mental status | 0
    multi-organ dysfunction syndrome | 0
    severe metabolic acidosis | 0
    hemolysis | 0
    managed with intravenous antibiotics | 0
    blood transfusion | 0
    received 3 units of blood | 0
    improved significantly after blood transfusion | 0
    lactic acid normalized within 10 hours | 10
    antibiotics discontinued | 10
    acute kidney injury resolved | 0
    mentation improved | 0
    weaned off ventilator | 48
    fecal occult blood tests negative | 0
    ferritin 588 ng/mL | 0
    TIBC 194 µg/dL | 0
    transferrin 155 mg/dL | 0
    iron saturation 91% | 0
    peripheral smear large RBCs | 0
    hypersegmented neutrophils (6-7 lobes) | 0
    schistocytes 1% | 0
    poikilocytes | 0
    anisocytosis | 0
    mixed picture of megaloblastic anemia | 0
    hemolytic anemia | 0
    vitamin B12 38 pg/mL | 0
    methylmalonic acid 753 nmol/L | 0
    homocysteine 99.3 µmol/L | 0
    anti-parietal antibodies 21.7 units | 0
    anti-intrinsic factor antibodies 4.7 AU/mL | 0
    direct Coombs test negative | 0
    indirect Coombs test negative | 0
    fibrinogen 185 mg/dL | 0
    D-dimer 5170 ng/mL | 0
    serology negative for HIV | 0
    serology negative for hepatitis virus | 0
    diagnosed with pernicious anemia | 0
    diagnosed with pseudo-TTP | 0
    intramedullary hemolysis | 0
    started on parenteral vitamin B12 | 0
    hematological parameters improved | 0
    clinical condition improved | 0
    discharged | 0
    blood parameters improved at discharge | 0
    hemoglobin 8.1 gm/dL | 0
    hematocrit 24.3% | 0
    platelets 292,000 per µL | 0
    MCV 98.9 fL | 0
    WBC 5.9 per µL | 0
    BUN 8 mg/dL | 0
    creatinine 0.7 mg/dL | 0
    total bilirubin 0.7 mg/dL | 0
    haptoglobin 144 mg/dL | 0
    LDH 720 IU/L | 0
    INR 1.11 | 0
    PT 12.9 s | 0
    aPTT 28.1 s | 0
    schistocytes 0% | 0
    D-dimer 5170 ng/mL | 0
