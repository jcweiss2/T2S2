53 years old | 0
male | 0
admitted to the hospital | 0
productive cough | -24
fever | -24
chills | -24
30-pack/year history of cigarette smoking | 0
consumed alcohol in moderation | 0
successfully treated for CAP in another hospital | -720
no other problems | 0
acutely ill | 0
blood pressure 82/46 mmHg | 0
respiratory rate 22 breaths per minute | 0
pulse rate 120 beats per minute | 0
body temperature 40℃ | 0
regular heart rhythm | 0
coarse breathing sounds with crackles on the right lower lung field | 0
white blood cell count of 11,500/mm3 | 0
neutrophils 86.1% | 0
lymphocytes 11.5% | 0
monocytes 1.9% | 0
eosinophils 0.2% | 0
hemoglobin 14.4 g/dL | 0
platelet count 188,000/mm3 | 0
C-reactive protein 1.28 mg/dL | 0
arterial blood gas analysis | 0
pH of 7.47 | 0
pCO2 of 22.4 mmHg | 0
pO2 of 52.5 mmHg | 0
HCO3- of 16 mmol/L | 0
O2 saturation of 89% | 0
blood urea nitrogen (BUN)/creatinine (Cr) level of 9/2.05 mg/dL | 0
serum sodium 139 mmol/L | 0
potassium 4.1 mmol/L | 0
chloride 105 mmol/L | 0
urine sodium 19 mmol/L | 0
urine Cr 222.31 mg/dL | 0
fractional excretion of sodium 0.1% | 0
moderate patchy consolidation in the right lower lobe | 0
sepsis caused by CAP | 0
septic shock | 0
central line catheter inserted | 0
fluid resuscitation | 0
oxygen administered via nasal cannula | 0
cultures of blood, sputum, and urine samples | 0
empiric piperacillin/tazobactam with ciprofloxacin injections | 0
admitted into the intensive care unit | 0
APACHE II score 25 | 0
norepinephrine administered | 2
vasopressin administered | 2
respiratory distress worsened | 16
acute respiratory failure | 16
arterial blood gas analysis | 16
pH of 7.085 | 16
pCO2 of 61.4 mmHg | 16
HCO3- of 19 mmol/L | 16
intubated with mechanical ventilation | 16
FiO2 of 1.0 | 16
positive end expiratory pressure at 14 cmH2O | 16
hypoxia persisted | 16
respiratory and metabolic acidosis continued to deteriorate | 16
follow-up arterial blood gas analysis | 24
pH of 7.096 | 24
pCO2 of 63.7 mmHg | 24
pO2 of 77.6 mmHg | 24
HCO3- of 20 mmol/L | 24
O2 saturation of 89% | 24
follow-up chest radiograph | 24
more exacerbated consolidation in the right lung field | 24
patchy opacities in the left lower lobe | 24
antibiotics switched to meropenem with teicoplanin | 24
oliguria ensued | 28
acute kidney injury | 28
BUN/Cr at 26/3.66 mg/dL | 28
continuous renal replacement therapy | 28
septic shock and acute respiratory failure did not improve | 36
cardiac arrest | 36
cardiopulmonary resuscitation | 36
AB identified in both the culture of sputum and two pairs of blood samples | 36
bacterial sensitivity to antibiotics measured | 36
bacterial isolate susceptible to piperacillin/tazobactam | 36
bacterial isolate susceptible to ceftazidime | 36
bacterial isolate susceptible to cefepime | 36
bacterial isolate susceptible to imipenem | 36
bacterial isolate susceptible to meropenem | 36
bacterial isolate susceptible to gentamicin | 36
bacterial isolate susceptible to tobramycin | 36
bacterial isolate tolerant to ampicillin | 36
bacterial isolate tolerant to amoxacillin/clavulanic acid | 36
bacterial isolate tolerant to cafalotin | 36
bacterial isolate tolerant to cefoxitin | 36
bacterial isolate tolerant to trimethoprim/sulfamethoxazole | 36
bacterial isolate moderately tolerant to cefotaxime | 36
bacterial isolate moderately tolerant to levofloxacin | 36
expired | 36