68 years old | 0
lady | 0
para 3 | 0
postmenopausal bleeding | 0
transvaginal ultrasound scan | 0
endometrial thickness 5 mm | 0
outpatient hysteroscopy | -15
procedure uneventful | -15
cavity normal | -15
ostia normal | -15
endometrial biopsy not possible | -15
patient found procedure painful | -15
abdominal pain | 0
nausea | 0
vomiting | 0
fever | 0
sweats | 0
rigors | 0
tachycardic | 0
hypotensive | 0
oxygen saturation 92% | 0
unremarkable examination | 0
high vaginal swab sent | 0
normal bloods | 0
computed tomography scan requested | 0
desaturating | 0
temperature 38.1°C | 0
blood pressure 84/48 mm Hg | 0
arterial blood gases done | 0
lactate 3.6 | 0
admitted to ITU | 0
septic shock | 0
inotropic support | 0
worsening lactate | 0
augmentin started | 0
metronidazole started | 0
gentamicin stat dose | 0
procalcitonin >10.0 μg/L | 0
metronidazole replaced with gentamicin | 0
fever started coming down | 0
lactate levels decreasing | 0
maximum lactate 4.25 | 0
stepped down to HDU | 72
augmentin replaced by benzylpenicillin | 72
clindamycin added | 72
inotropes stopped | 72
transferred to gynecology ward | 72
afebrile | 72
vitals stable | 72
antibiotics switched to oral | 72
discharged | 192
normal CT scan | 0
no perforation | 0
no pelvic collection | 0
HVS growth beta-hemolytic Group A Streptococci | 0
blood cultures growth GAS | 0
septic shock confirmed | 0
TSS | 0
