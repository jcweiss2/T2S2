29 years old | 0
male | 0
asthma | 0
previous gunshot wound | 0
obesity | 0
tobacco use | 0
auto-parts manufacturing unit worker | 0
admitted to the hospital | 0
dyspnea | 0
cough | 0
fatigue | 0
myalgias | 0
febrile | 0
tachycardic | 0
tachypneic | 0
supplemental oxygen | 0
high work of breathing | 0
productive cough | 0
lymphopenia | 0
thrombocytopenia | 0
unremarkable chest radiograph | 0
transferred to ICU | 0
COVID-19 suspicion | 0
SARS-CoV-2 testing | 0
nasopharyngeal swab | 0
M4 viral tube | 0
State Department of Health and Human Services | 0
RT-PCR | 0
Abbott ID NOW | 0
FDA emergency use authorization | 0
higher flow rates on non-rebreather mask | 72
persistent fevers | 96
tachypnea | 96
new consolidative changes | 96
broad-spectrum antibiotics | 96
hydroxychloroquine | 96
mechanical ventilation | 96
chest x-ray | 192
extensive consolidative infiltrates | 192
PaO2/FiO2 ratio of 59 | 192
ARDS | 192
SARS-CoV-2 positive | 192
septic shock | 240
vasopressor support | 240
cytokine labs | 240
interleukin-6 | 240
tocilizumab | 240
DVTs | 240
enoxaparin | 240
fevers | 240
cooling | 240
neuromuscular blockade | 240
deep sedation | 240
ARDS strategies | 240
low tidal volumes | 240
proning | 240
recruitment maneuvers | 240
diuretics | 240
nitric oxide | 240
vitamin C | 240
high plateau pressures | 240
ECMO center | 240
infection control measures | 240
resource allocation | 240
logistical challenges | 240
desaturation | 408
left-sided tension pneumothorax | 408
chest tube | 408
serosanguineous fluid | 408
blood clots | 408
persistent air leaks | 408
family discussion | 408
poor prognosis | 408
goals of care | 408
code status changed to DNR | 408
comfort measures | 408
asystole | 480
death | 480