35 years old | 0
female | 0
gravida 5 | 0
para 2022 | 0
admitted to the hospital | 0
vaginal bleeding | 0
fevers | -120
headache | -120
neck stiffness | -120
altered mental status | -120
dog bite | -72
fetal intrauterine growth restriction | -336
motor vehicular accident | -7200
splenectomy | -7200
diffuse axonal brain injury | -7200
seizure disorder | -7200
cesarean delivery | -7200
tremulous chills | -120
fevers to 102.7°F | -120
off-balance | -120
slurring her words | -120
new-onset significant fatigue | -120
persistent headache | -120
transient spotting | -120
bright red vaginal bleeding | 0
wound on her index finger | -72
well-healing | -72
no erythema | -72
no swelling | -72
no tenderness | -72
category 2 fetal heart tracing | 0
emergent repeat low transverse cesarean section | 0
neonate admitted to the NICU | 0
respiratory failure | 0
intubation | 0
core temperature lability | 0
stable hemodynamic vitals | 0
platelet count 8×10^9/L | 0
transfused with 2 units of platelet | 0
platelet count 55×10^9/L | 0
thrombophilia | 0
baseline platelet count 400×10^9/L | -7200
schistocytes on peripheral smear | 0
normal ADAMST13 level | 0
sepsis | 0
disseminated intravascular coagulation | 0
normal coagulation studies | 0
normal fibrinogen | 0
normal prothrombin time | 0
normal partial prothrombin time | 0
clindamycin | 0
gentamicin | 0
metronidazole | 0
asplenic patient | 0
immunocompromised patient | 0
cell-mediated immune defenses | 0
encapsulated organisms | 0
Capnocytophaga | 0
bacteremia | 0
sepsis | 0
rabies | -72
rabies prophylaxis | -72
meropenem | 0
carbapenem beta-lactam | 0
broad coverage | 0
gram positive organisms | 0
gram negative organisms | 0
x-ray of the finger | 0
unremarkable | 0
no acute signs of osteomyelitis | 0
tick bite | -720
Coxiella burnetii | -720
Q fever | -720
goat placenta | -720
doxycycline | 0
tick-borne rickettsial diseases | 0
meningeal process | 0
neck stiffness | 0
fluctuating mental status | 0
lumbar puncture | 0
high risk for bleeding | 0
encephalopathy | 0
altered mental status | 0
MRI of the brain | 0
no evidence of encephalitis | 0
no acute intracranial processes | 0
chronic change | 0
prior brain injury | -7200
blood cultures | 0
gram negative bacilli | 0
Capnocytophaga species | 0
IV ertapenem | 0
carbapenem beta-lactam antibiotic | 0
10-day course | 0
Capnocytophaga canimorsus | 0
MALDI-TOF mass spectrometry | 0
16S rRNA sequencing | 0
neonate sent to the NICU | 0
briefly intubated | 0
respiratory distress | 0
discharged to the newborn nursery | 144
blood cultures from the neonate | 0
negative | 0
platelet count recovered | 24
278×10^9/L | 24
IV antibiotics | 0
profound thrombocytopenia | 0
platelet consumption | 0
decreased platelet production | 0
C. canimorsus infection | 0
discharged on the sixth hospital day | 144
completed IV ertapenem therapy | 144
outpatient basis | 144
at home | 144