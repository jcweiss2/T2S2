39 years old | 0
female | 0
chronic kidney disease | -7776
maintenance hemodialysis | -7776
severe PAH | -7776
chronic pulmonary thromboembolism | -7776
progressive breathlessness | -168
abdominal distension | -168
Grade III dyspnea | -168
orthopnea | -168
no fever | -168
no cough | -168
blood pressure 92/46 mmHg | -168
pulse rate 96/min | -168
respiratory rate 36/min | -168
recurrent hypotension | -168
non-tolerance to HD | -168
planned peritoneal dialysis | 0
severe hypotension | 0
altered sensorium | 0
shifted to ICU | 0
drowsy | 0
sluggishly responding to verbal commands | 0
distended neck veins | 0
respiratory distress | 0
active accessory muscles of respiration | 0
loud P2 | 0
pan systolic murmur | 0
soft abdomen | 0
mildly distended abdomen | 0
evidence of free fluid | 0
palpable liver | 0
blood pressure 70/40 mmHg | 0
pulse rate 102/min | 0
respiratory rate 30/min | 0
SpO2 99% | 0
Hemoglobin 12.3 g/dl | 0
total leucocyte count 8600/μL | 0
serum sodium 138 mEq/L | 0
serum potassium 6 mEq/L | 0
blood urea nitrogen 63 mg/dl | 0
creatinine 6.0 mg/dl | 0
hypoxia | 0
hypercarbia | 0
mixed acidosis | 0
pH 7.189 | 0
PaCO2 60.3 mmHg | 0
pO2 52.7 mmHg | 0
HCO3 22.5 mmol/L | 0
BE 6.54 mmol/L | 0
serum lactate 1.92 mmol/L | 0
high D-dimer | 0
high fibrin degradation product | 0
dilated right ventricle | 0
moderate tricuspid regurgitation | 0
severe PAH | 0
PASP 93 mmHg | 0
paradoxical septal motion | 0
decreased RV function | 0
reduced LV compliance | 0
no sepsis | 0
no acute myocardial ischemia | 0
infusion nor-adrenaline | 0
infusion dopamine | 0
empiric broad spectrum antibiotics | 0
low molecular weight heparin | 0
sustained low efficiency dialysis | 0
increased vasopressor requirement | 24
infusion vasopressin | 24
elective intubation | 24
ventilation | 24
pre-intubation ABG | 24
post-intubation ABG | 24
pH 7.18 | 24
PaCO2 60 mmHg | 24
PO2 66.6 mmHg | 24
HCO3 21.9 mmol/L | 24
BE 7.1 mmol/L | 24
pH 7.29 | 24
PaCO2 36.7 mmHg | 24
PO2 80.4 mmHg | 24
HCO3 17.3 mmol/L | 24
BE 8.3 mmol/L | 24
echocardiography | 48
PASP 95 mmHg | 48
iNO started | 72
iNO 5 ppm | 72
iNO 10 ppm | 72
improving hemodynamic parameters | 84
vasopressors tapered down | 84
PD restarted | 120
cumulative negative balance 2 L | 120
blood gasses | 120
pH 7.45 | 120
PaCO2 28.4 mmHg | 120
PO2 136.2 mmHg | 120
HCO3 20 mmol/L | 120
BE 5.3 mmol/L | 120
lactates 1.61 mmol/L | 120
follow-up echocardiography | 144
PASP 73 mmHg | 144
PASP 63 mmHg | 168
vasopressors weaned off | 168
NO withdrawn | 168
extubation | 168
non-invasive ventilation | 168
inspiratory positive airway pressure 12 mmHg | 168
expiratory positive airway pressure 4 mmHg | 168
shifted out of ICU | 240
methemoglobin levels < 1% | 240