67 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
mucosal resection for early gastric cancer | -10080 | -10080 | Factual
partial resection for left lung cancer | -10080 | -10080 | Factual
no heart disease | 0 | 0 | Factual
conventional drugs | 0 | 0 | Factual
collected knee-high wild grass from a riverbed | -240 | -240 | Factual
systemic pain | -168 | 0 | Factual
fatigue | -168 | 0 | Factual
fever | -168 | 0 | Factual
chills | -168 | 0 | Factual
watery diarrhea | -168 | 0 | Factual
loss of appetite | -168 | 0 | Factual
mildly disturbed consciousness | -168 | 0 | Factual
decreased white blood cells (WBC) | -24 | 0 | Factual
decreased platelet counts | -24 | 0 | Factual
elevated hepatic enzyme levels | -24 | 0 | Factual
hepatic dysfunction | -24 | 0 | Factual
hospitalized | 0 | 0 | Factual
height of 169.0 cm | 0 | 0 | Factual
body weight of 52.3 kg | 0 | 0 | Factual
Glasgow Coma Scale of 14: E3, V5, M6 | 0 | 0 | Factual
blood pressure of 130/79 mmHg | 0 | 0 | Factual
heart rate (HR) of 96/min | 0 | 0 | Factual
respiratory rate (RR) of 20/min | 0 | 0 | Factual
O2 saturation (SPO2) of 94% | 0 | 0 | Factual
temperature of 38.9°C | 0 | 0 | Factual
crusted skin lesions on the medial surface of the left thigh | 0 | 0 | Factual
freely movable adenopathy of approximately 2 cm in size | 0 | 0 | Factual
aggregated papules in the right inguinal region | 0 | 0 | Factual
no remarkable head-and-neck or chest abnormalities | 0 | 0 | Factual
no remarkable neurological abnormalities | 0 | 0 | Factual
blood count of 1,300 /μL WBC | 0 | 0 | Factual
platelets of 30,000 /μL | 0 | 0 | Factual
neutrophil count of 899 /μL | 0 | 0 | Factual
lymphocyte count of 342 /μL | 0 | 0 | Factual
activated partial thromboplastin time (APTT) of 48.2 seconds | 0 | 0 | Factual
C-reactive protein (CRP) levels of 1.3 mg/dL | 0 | 0 | Factual
aspartate aminotransferase (AST) of 230 U/L | 0 | 0 | Factual
lactate dehydrogenase (LDH) of 760 U/L | 0 | 0 | Factual
creatine kinase (CK) of 746 U/L | 0 | 0 | Factual
sepsis | 24 | 24 | Possible
febrile neutropenia (FN) | 24 | 24 | Possible
hemophagocytosis | 24 | 24 | Possible
antibiotics | 24 | 168 | Factual
elevated ferritin levels of 15,165 ng/mL | 48 | 48 | Factual
screened for potential antibodies specific for cytomegalovirus and Epstein-Barr virus (EBV) | 48 | 48 | Factual
bone marrow biopsy | 48 | 48 | Factual
hemophagocytosis with fewer mature myeloid series cells and more monocytoid and lymphoid cells | 48 | 48 | Factual
immunohistological examination | 48 | 48 | Factual
high number of CD3- and CD4-positive T cells | 48 | 48 | Factual
MUM-1-positive lymphoid cells | 48 | 48 | Factual
CD68, CD163-positive histiomonocytes | 48 | 48 | Factual
no EBV-encoded small RNAs (EBERs)-positive cells | 48 | 48 | Factual
HLH | 48 | 168 | Factual
prednisolone (PSL) at 60 mg/day | 48 | 288 | Factual
chest pain | 72 | 72 | Factual
shivering | 72 | 72 | Factual
fever of 39.2°C | 72 | 72 | Factual
blood pressure at 88/52 mmHg | 72 | 72 | Factual
HR at 89/min | 72 | 72 | Factual
RR at 24/min | 72 | 72 | Factual
SPO2 at 94% | 72 | 72 | Factual
elevated CK levels at 953 U/L | 72 | 72 | Factual
elevated LDH at 1,405 U/L | 72 | 72 | Factual
high-sensitivity troponin I (TnI) at 271 pg/mL | 72 | 72 | Factual
severe left ventricular dysfunction | 72 | 72 | Factual
electrocardiogram (ECG) showed a slight ST elevation in the V1-2 leads | 72 | 72 | Factual
myocarditis | 72 | 168 | Factual
inotropic agents | 72 | 168 | Factual
water balance management | 72 | 168 | Factual
ventilation management | 72 | 168 | Factual
reverse transcription polymerase chain reaction (RT-PCR) analysis | 96 | 96 | Factual
SFTSV RNA copies/mL of 1.77×106 | 96 | 96 | Factual
infected cells stained positively by an anti-SFTSV-nucleoprotein (N) antibody | 96 | 96 | Factual
steroid pulse therapy | 120 | 120 | Possible
circulatory agonist | 168 | 336 | Factual
ventilator management | 168 | 336 | Factual
ECG showed improvement of ST elevation in the V1-2 leads | 336 | 336 | Factual
serum and confirmed negativity for viremia | 408 | 408 | Factual
released from quarantine | 408 | 408 | Factual
coronary angiography (CAG) | 576 | 576 | Factual
endomyocardial biopsy (EMB) | 576 | 576 | Factual
mildly hypertrophic with mild myofibrillar loss and disarrangement | 576 | 576 | Factual
active mononuclear cell infiltration | 576 | 576 | Factual
increases in the number of CD3-positive T cells | 576 | 576 | Factual
CD68-positive macrophages | 576 | 576 | Factual
tenascin-C expression | 576 | 576 | Factual
discharged | 696 | 696 | Factual
follow-up visit | 744 | 744 | Factual
transthoracic echocardiography showed a slight improvement with an EF of 52.5% | 744 | 744 | Factual
no heart failure | 744 | 744 | Factual