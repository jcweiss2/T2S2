56 years old | 0
female | 0
abnormal vaginal discharge | -336
visited gynecologist | -336
vaginal culture | -336
cervical cytology | -336
endometrial cytology | -336
fever | -10
lower abdominal pain | -10
visited emergency room | 0
blood pressure 71/46 mmHg | 0
tenderness from right upper quadrant to lower abdomen | 0
fluid resuscitation therapy | 0
procalcitonin 75.49 ng/mL | 0
abdominal CT examination | 0
full stomach | 0
edema of small intestine | 0
exploratory laparotomy | 3
purulent ascites | 3
bilateral salpingitis | 3
peritoneal lavage and drainage | 3
intubated | 3
noradrenaline administration | 3
meropenem 1.5 g/day | 3
extubated | 48
noradrenaline tapered | 48
noradrenaline terminated | 72
oral intake started | 96
drainage tube removed | 96
GAS detected in vaginal fluid culture | 120
GAS detected in ascitic fluid culture | 120
intravenous injection of antibiotics stopped | 120
oral levofloxacin prescribed | 120
body temperature rose to 38.1 °C | 120
discharged | 240
condition generally good | 2880
infection did not recur | 2880