30 years old | 0
gravida 1 | 0
para 0 | 0
admitted to hospital | 0
preterm labor | 0
21 weeks gestation | 0
prenatal laboratories unremarkable | 0
negative GBS screen | -120
antenatal steroid course | -72
betamethasone | -72
latency antibiotics | -47
ampicillin | -47
azithromycin | -47
magnesium for neuroprotection | -48
male neonate | 0
23 weeks and 4/7 gestational age | 0
vaginal delivery | 0
prolonged rupture of membranes | -58
0.595 kg birth weight | 0
58%ile | 0
intubation | 0
surfactant | 0
respiratory distress | 0
APGAR score 5, 6, 8 | 0
admitted to NICU | 0
high-frequency oscillator | 0
caffeine | 0
umbilical catheters | 0
evaluation for bacterial infection | 0
ampicillin and gentamicin | 0
discontinued antibiotics | 48
nil per os | 0
total parenteral nutrition | 0
conventional mechanical ventilation | 22
failed ventilation | 60
transferred to facility | 72
leukocytosis | 99
bandemia | 99
septic workup | 99
blood culture | 99
empiric treatment | 99
amoxicillin and cefepime | 99
abdominal discoloration | 99
abdominal radiograph | 99
gasless abdomen | 99
blood culture positive | 108.6
M. morganii | 108.6
line removal | 108.6
full sepsis workup | 120
repeat blood cultures | 120
lumbar puncture | 120
nonsterile urine culture | 120
antibiotic coverage broadened | 120
meropenem and ampicillin | 120
CSF analysis | 120
Enterococcus faecalis | 120
nonsterile urine culture positive | 120
Staphylococcus epidermis | 120
M. morganii | 120
E. faecalis | 120
peripheral culture positive | 120
M. morganii | 120
UVC culture negative | 120
clinically worsened | 192
bilious emesis | 192
abdominal discoloration | 192
abdominal radiograph | 192
free intraperitoneal air | 192
spontaneous intestinal perforation | 192
peritoneal drain | 192
intraoperative peritoneal culture | 192
M. morganii | 192
antibiotic coverage changed | 192
vancomycin and fluconazole | 192
M. morganii sensitivities | 216
meropenem changed | 216
ampicillin and cefepime | 216
placental maternal culture | 0
E. coli | 0
Streptococcus viridans | 0
coagulase negative Staphylococcus | 0
Enterococcus | 0
Bacillus fragilis | 0
Prevotella species | 0
clinically improved | 240
enteral feeds | 240
dexamethasone | 240
extubated | 720
weaned to room temperature | 840
patent ductus arteriosus treated | 840
acetaminophen | 840
bilateral germinal matrix hemorrhages | 840
mildly dilated ventricles | 840
normalized | 1008
corrected full-term cranial ultrasound | 1008
small left-sided periventricular cyst | 1008
stage 2 retinopathy of prematurity | 1008
discharged home | 3024
high-risk infant follow-up clinic | 3024
feeding therapy | 3024
infant development services | 3024
physical therapy | 3024
normal cognitive skills | 3024
expressive language | 3024
fine motor skills | 3024
gross motor skills | 3024
sensory processing | 3024
mild delays in receptive language | 3024
social emotional skills | 3024
outpatient magnetic resonance imaging | 3024
no significant structural or signal abnormality | 3024