64 years old | 0
female | 0
admitted to the hepatobiliary surgery department | 0
severe sepsis | -24
liver abscess | -24
conservative treatment | -24
IV antibiotics | -24
transferred to hospital | 0
past medical history not remarkable | 0
well controlled hypertension | 0
stable vital signs | 0
mild pain | 0
discomfort in the right upper quadrant | 0
discomfort in the flank | 0
denied foreign body ingestion | 0
denied recent trauma | 0
abdominal clinical examination did not reveal any abnormalities | 0
normal white blood cells count | 0
C-reactive protein 48 mg/dL | 0
haemoglobin 9.2 g/dL | 0
hematocrit 24 % | 0
aspartate aminotransferase AST 45.4 IU/L | 0
alanine aminotransferase ALT 49.5 IU/L | 0
CT scan showed hypodense area | -24
CT scan showed linear hyperdense feature | -24
abdominal ultrasonography showed elongated hyperechoic structure | 0
scheduled for selective laparotomy | 0
subcostal incision with midline extension | 12
intraoperative finding of scar on the out surface of segment V | 12
loose adhesions between the first part of the duodenum and the inferior surface of the liver | 12
intraoperative ultrasound scan | 12
located and marked the foreign body | 12
5 cm incision in the liver capsule | 12
finger fracture technique of the hepatic parenchyma | 12
foreign body found to be a toothpick | 12
toothpick measured 5.5 cm-long | 12
embedded in tough fibroid tissue | 12
abdomen closed | 24
no drains used | 24
spent two days on the ward | 24
discharged | 48
ingestion of toothpick | -168
migration of toothpick to the liver | -168
toothpick caused liver abscess | -24
liver abscess diagnosed | -24
treatment with IV antibiotics started | -24
treatment with IV antibiotics ended | 0 
Note: The time stamp for the ingestion of the toothpick and its migration to the liver is an approximation, as the exact time is not provided in the case report. The time stamp of -168 hours is an estimate, assuming the toothpick was ingested 7 days prior to the admission.