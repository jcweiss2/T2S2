68 years old | 0
female | 0
poorly controlled DM | 0
altered mental status | -96
unresponsive | -96
blood sugar 498 | -96
tachycardic | 0
heart rate 169 | 0
hypotensive | 0
blood pressure 86/45 | 0
tachypneic | 0
oxygen saturation 92% | 0
WBC 19.4 thous/mm3 | 0
Na 129 Meq/dL | 0
Cl 92 Meq/dL | 0
creatinine 3.63mg/dL | 0
Co2 10 Meq/L | 0
CRP 40.2 mg/dL | 0
ESR 70mm/hr | 0
glucose 719 mg/dL | 0
lactic acid 3.6 mmol/L | 0
abnormally turbid urine | 0
glucose >1000 | 0
WBCs 10–20 | 0
RBCs 5–10 | 0
4+ bacteria | 0
TNTC of yeast | 0
Candida glabrata | 0
IV micafungin | 0
IV cefepime | 0
DKA protocol | 0
hyperosmolar hyperglycemic state | 0
free air in extraperitoneal space | 0
extraperitoneal bladder perforation | 0
foley catheter placement | 0
intubated | 24
extubated | 120
hypoxia | 144
tachypnea | 144
hypertension | 144
ABG showed Pa. O2 in the 40's | 144
reintubated | 144
heparin | 144
fever | 168
tachycardic | 168
tracheostomy | 240
pressure support | 240
transition to comfort care | 528
multiorgan and respiratory failure | 528
cardiac arrest | 528
passed away | 528
type 2 DM | -672
peripheral artery disease | -672
atherosclerosis | -672
coronary artery disease | -672
mesenteric ischemia | -672
gastroparesis | -672
fibromyalgia | -672
stenting procedure | -672
vascular graft | -672