hypertension | 0
diabetes mellitus | 0
intermittent subjective fever | -96
rigors | -96
generalized headache | -96
altered mentation | -96
body malaise | -96
nausea | -96
vomiting | -96
no history of loss of consciousness | -96
no abdominal pain | -96
no change in stool habits/urine color | -96
no recent trauma or falls | -96
febrile | 0
tachypneic | 0
disoriented | 0
good nutritional status | 0
not jaundiced | 0
not cyanosed | 0
pulse rate of 103 beats/min | 0
respiratory rate of 23 breaths/min | 0
blood pressure of 96/60 mmHg | 0
saturating at 98% on room air | 0
normal vesicular breath sounds | 0
normal abdominal examination | 0
IV resuscitation | 0
analgesia | 0
white blood cell count of 8.2 × 103/μL | 0
hemoglobin of 11.5 g/dL | 0
thrombocytopenia of 46,000/mm3 | 0
elevated creatinine 117 μmol/L | 0
BUN 10.5 mmol/L | 0
slightly low sodium of 131 mmol/L | 0
normal serum electrolytes | 0
normal liver | 0
normal coagulation profile | 0
normal chest X-ray | 0
P. falciparum with high parasitemia | 0
admitted to ICU | 0
intravenous artesunate-based regimen | 0
supportive measures | 0
improvement in clinical status | 72
improvement in lab parameters | 72
shifted to general ward | 72
acute abdomen | 120
progressive abdominal pain | 120
nausea | 120
non-bilious vomiting | 120
anxious | 120
afebrile | 120
diaphoretic | 120
tachycardic | 120
tachypneic | 120
hypotensive | 120
saturating well on room air | 120
slightly distended abdomen | 120
tender on superficial palpation | 120
inaudible bowel sounds | 120
low Hb of 7.1 g/dL | 120
hypoechoic nodular cystic area | 120
splenomegaly | 120
hyperdense intrasplenic hematoma | 120
hypodense subcapsular hematoma | 120
splenic laceration | 120
intraperitoneal free fluid | 120
grade 3 splenic injury | 120
blood products mobilized | 120
adequate resuscitation | 120
explorative laparotomy | 120
splenectomy | 120
2.5 L of frank blood evacuated | 120
enlarged spleen | 120
long laceration on the upper pole | 120
uneventful postoperative period | 168
discharged home | 168
fully recovered | 168