62 years old | 0
male | 0
hypertension | 0
hyperlipidaemia | 0
dizziness | -168
fatigue | -168
nausea | -168
vomiting | -168
syncope | 0
out-of-hospital cardiac arrest | 0
ECG showing ST elevations | 0
ventricular fibrillation | 0
cardiac defibrillation | 0
endotracheal intubation | 0
heart rate of 77 b.p.m. | 0
regular rhythm | 0
hypotension | 0
no lower extremity oedema | 0
extremities were cool to touch | 0
mechanical ventilation | 0
aspirin | 0
ticagrelor | 0
heparin | 0
epinephrine infusion | 0
coronary angiogram | 1
no coronary stenosis | 1
right heart catheterization | 6
elevated right-sided filling pressures | 6
right atrial pressure of 22 mmHg | 6
pulmonary artery pressure 61/28 mmHg | 6
pulmonary capillary wedge pressure 15 mmHg | 6
Fick cardiac index 2.6 L/min/m2 | 6
point-of-care echocardiogram | 6
dilated right ventricle | 6
severely reduced right ventricular function | 6
pulmonary angiography | 6
bilateral pulmonary emboli | 6
EkoSonic endovascular thrombolysis catheters | 6
tissue plasminogen activator | 6
upper and lower extremity Doppler ultrasounds | 6
no evidence of venous thrombosis | 6
formal transthoracic echocardiogram | 6
depressed right ventricular function | 6
computed tomography of chest | 96
bilateral peripheral ground-glass opacities | 96
wedge-shaped opacities in the right lung | 96
pulmonary infarctions | 96
broad-spectrum antibiotics | 96
viral respiratory panel | 96
tracheal aspirate culture | 96
methicillin-resistant Staphylococcus aureus | 96
repeat ECG | 96
sinus rhythm | 96
first-degree atrioventricular block | 96
left axis deviation | 96
incomplete right bundle branch block | 96
prolonged QTc interval | 96
anaemia | 96
CT of chest, abdomen, and pelvis | 96
mediastinal haematoma | 96
persistent ground-glass opacities | 96
COVID-19 testing | 96
positive SARS-CoV-2 | 96
transferred to COVID-19-dedicated intensive care unit | 96
enhanced contact precautions | 96
supportive care | 96
extubated | 192
admitted to inpatient rehabilitation facility | 192
discharged home | 672
lifelong apixaban | 672
mild exertional dyspnoea | 720
improvement of right ventricular dilation and systolic function | 720