52 years old | 0
female | 0
primary hypertension | 0
admitted to the emergency department | 0
diffuse myalgias | -72
fever | -72
cough | -72
temperature 35.9°C | 0
pulse oxygen saturation 99% | 0
heart rate 62 per minute | 0
blood pressure 127/89 mmHg | 0
diffuse muscle pain | 0
creatine kinase levels 15000 IU/L | 0
SARS-CoV-2 RNA positive | 0
L452R mutation | 0
mild pulmonary infiltrates | 0
no pulmonary embolism | 0
Glasgow score 12/15 | 48
temperature 40°C | 48
heart rate 130 per minute | 48
hypotension 70/30 mmHg | 48
anuria | 48
diffuse mottling | 48
oxygen therapy | 48
intravenous saline | 48
intravenous bicarbonate | 48
vasopressor support with Norepinephrine | 48
intubated | 48
mechanically ventilated | 48
renal replacement therapy | 48
Hydrocortisone | 48
antibiotics | 48
preventive anticoagulation by Enoxaparine | 48
cardiorespiratory arrest | 72
resuscitation | 72
death | 117 
myoglobin >30 000 | 48
CPK 100 557 | 0
CPK 101 624 | 48
myoglobinuria | 0
dark colored urine | 0
weakness | 0
wbc 10.11 | 0
lymphocytes 1.32 | 0
CRP 37.8 | 0
d-dimer 2.50 | 0
hypersensitive troponin t 962 | 0
hypersensitive troponin t 2028 | 48
creatinine 129 | 0
Egfr 38 | 0
urea 12.8 | 0
K+ 6.4 | 0
K+ 6.7 | 48
AST 2394 | 0
AST 1978 | 48
ALT 561.8 | 0
ALT 517 | 48
COVID-19 viral load 310 | 0
pneumococcal/legionella antigen urines NEGATIVE | 0
pH 7.43 | 0
pH 7.11 | 48
Po2 98 | 0
Po2 67 | 48
pco2 18 | 0
pco2 34 | 48
hco3- 11.9 | 0
hco3- 10.8 | 48
lactate 6.7 | 0
lactate 15.6 | 48