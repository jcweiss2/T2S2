37 years old | 0
Afro-Caribbean | 0
female | 0
admitted to the hospital | 0
lethargy | -504
myalgia | -504
intermittent chest pain | -504
uncomplicated pregnancy | -10080
acute kidney injury | 0
severe hypercalcaemia | 0
proteinuria | 0
treatment with intravenous fluids | 0
treatment with empirical antimicrobials | 0
transferred to the Intensive Care Unit (ICU) | 24
respiratory support | 24
renal replacement therapy | 24
deterioration | 24
vasculitis | 0
autoimmune disease | 0
sepsis | 0
malignancy | 0
leukocytosis | 0
left shift | 0
no abnormal cells | 0
autoimmune screen negative | 0
respiratory virus panel negative | 0
human immunodeficiency virus negative | 0
hepatitis B and C antibodies negative | 0
parathyroid hormone (PTH) level suppressed | 0
recurrent episodes of narrow- and broad-complex tachycardia | 96
poor global systolic function | 96
no pericardial effusion | 96
no obvious valvular abnormality | 96
treatment with DC cardioversion | 96
treatment with antiarrhythmics | 96
sensitivity to amiodarone | 96
sensitivity to lignocaine | 96
sensitivity to adrenaline | 96
fatal brady-tachy arrhythmia | 100
prolonged cardiac arrest | 100
resuscitation unsuccessful | 100
intracellular calcium deposition in cardiac myocytes | 100
widespread calcification in medium- and small-sized arteries | 100
intra-renal arteries with secondary micro-infarcts | 100
infiltration of lymph nodes by large lymphoid blasts | 100
histiocytic haemophagocytosis | 100
lymphoid blasts stained positively for CD3 and CD25 | 100
parathyroid glands histologically normal | 100
antibodies to human T-cell lymphotropic virus (HTLV) type 1 positive | 100
adult HTLV-related adult T-cell leukaemia-lymphoma (ATLL) | 100
hypercalcaemia | 0
cardiac dysrhythmia | 96
arrhythmias | 96
second- or third-degree atrio-ventricular block | 96
intracellular and extracellular calcium deposition | 100
cardiac contraction and myocardial relaxation impacted | 100
malignant cells not seen in peripheral blood film | 0
ATLL diagnosis | 100
HTLV-1 infection | -10080
vertical transmission during lactation | -10080
hypercalcaemia in 70-80% of patients with ATLL | 100
systemic hypercalcaemia and prodigious myocyte calcification | 100
pro-inflammatory processes | 100
refractory cardiovascular instability | 100
rapid demise | 100