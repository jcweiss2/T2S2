85 years old | 0
male | 0
farmer | 0
active lifestyle | 0
admitted to the hospital | 0
transferred from geriatric medicine unit | 0
underwent intensive treatment | 0
sequelae of C. tetani infection | 0
past medical history included atrial fibrillation | -672
past medical history included benign prostatic hypertrophy | -672
injured his leg while working on his farm | -144
admitted to a local hospital | -144
trismus | -144
hypertonia | -144
treated with immunoglobulins | -144
treated with tetanus vaccination | -144
treated with metronidazole | -144
transferred to ICU | -120
tracheostomy | -120
mechanical ventilation | -120
vasoactive support | -120
respiratory failure | -120
seizures | -120
treated with baclofen | -120
treated with midazolam | -120
treated with diazepam | -120
electroencephalography | -120
severely slow cerebral activity | -120
worsening respiratory function | -96
opacity on chest radiography | -96
peripheral leukocytosis | -96
possible ventilator-associated pneumonia | -96
blood cultures | -96
tracheal secretion samples | -96
tracheal secretions tested positive for Klebsiella pneumoniae | -96
tracheal secretions tested positive for methicillin-sensitive Staphylococcus aureus | -96
antibiotic therapy with piperacillin-tazobactam | -96
transferred to geriatric unit | -72
coma | -72
breathed spontaneously on 4 L/min of supplemental oxygen | -72
via a tracheal cannula | -72
antibiotic therapy switched to linezolid | -60
VAP exacerbation | -60
combined treatment with meropenem | -55
septic shock | -55
gradually awoke | -40
feeding tube removed | -40
cholestasis | -30
acute edematous pancreatitis | -30
endoscopic treatment postponed | -30
urinary tract infection | -20
caused by multidrug-resistant organisms | -20
treated with colistin | -20
treated with amoxicillin-clavulanate | -20
clinical condition improved | 0
considered eligible for rehabilitation | 0
placed in MDRO isolation | 0
required tracheal supplemental oxygen | 0
required bladder catheter | 0
developed pressure ulcers | 0
on the right heel | 0
on the left heel | 0
on the sacrum | 0
on the right elbow | 0
sarcopenic | 0
low handgrip strength | 0
low appendicular skeletal mass | 0
underwent rehabilitation | 24
good compliance | 24
Clostridioides difficile infection | 48
treated with oral vancomycin | 48
atrial fibrillation | 72
third-degree atrioventricular block | 72
heart rate 30 beats/min | 72
transferred to cardiac ICU | 72
underwent single-chamber pacemaker implantation | 72
hyperkinetic delirium | 96
Pseudomonas aeruginosa bloodstream infection | 120
treated with ceftazidime-avibactam | 120
treated with amikacin | 120
tested positive for SARS-CoV-2 | 120
treated with remdesivir | 120
placed on droplet isolation | 120
second recurrence of C. difficile | 144
treated with fidaxomicin | 144
bloodstream infection | 168
due to Candida parapsilosis | 168
due to MSSA | 168
due to Candida tropicalis | 168
treated with caspofungin | 168
treated with cefazolin | 168
tracheostomy closure | 240
performed by ENT specialist | 240
performed by pulmonologist | 240
nutritional supplementation | 240
prescribed to manage malnutrition | 240
prescribed to manage sarcopenia | 240
motor reconditioning | 240
respiratory reconditioning | 240
postural transition training | 240
aided transfers | 240
axial stability | 240
balance improvement exercises | 240
breath-movement coordination exercises | 240
thoracic expansion exercises | 240
girdle opening exercises | 240
inhalation-exhalation exercises | 240
wheelchairs recommended | 240
walkers recommended | 240
rehabilitation follow-up evaluations | 240
ENT follow-up evaluations | 240
geriatric follow-up evaluations | 240
discharged | 720