11 years old | 0
    male | 0
    acute abdominal pain | -24
    pushing another boy in a wheelchair | -24
    pain started | -24
    non-colicky pain | -24
    infra-umbilical region pain | -24
    pain worsened after onset | -24
    intermittent projectile vomiting | -24
    no fever | 0
    no chills | 0
    no diarrhoea | 0
    no bloody stool | 0
    septic appearance | 0
    lethargic | 0
    severely dehydrated | 0
    temperature of 37.5°C | 0
    pulse of 157 bpm | 0
    blood pressure of 97/41 mmHg | 0
    moderately distended abdomen | 0
    generalized guarding | 0
    rebound tenderness | 0
    unremarkable digital rectal examination | 0
    blood urea of 10.3 mmol/l | 0
    serum creatinine of 87 umol | 0
    elevated white cell count of 14,700/mm3 | 0
    hemoglobin of 16.8 g/dl | 0
    fluid resuscitation | 0
    catheterized | 0
    nasogastric tube insertion | 0
    oxygen administered per face mask | 0
    laparotomy | 0
    gangrenous loops of small bowel | 0
    large 8x8 cm mesenteric cyst | 0
    ischemic loops of bowel | 0
    ileo-cecal junction | 0
    gangrenous loop of terminal ileum | 0
    resection of gangrenous bowel | 0
    excision of peritoneal sac | 0
    jejunum to ascending colon anastomosis | 0
    abdomen irrigated | 0
    abdomen closed primarily | 0
    haemodynamically unstable | 0
    inotropic support required | 0
    sepsis concern | 0
    anastomotic leak concern | 0
    short bowel syndrome concern | 0
    intensive care unit management | 0
    inotropic support weaned off | 0
    extubated on day 4 | 96
    broad-spectrum antibiotics continued | 0
    no signs of anastomotic leak | 0
    discharged on day 9 | 216
    six months post-operative follow-up | 4320
    no short-bowel syndrome | 4320
    no significant morbidity | 4320
    histology results not available | 0
    peritoneal encapsulation diagnosis | 0
    gangrenous small bowel resection | 0
    vitamin B12 deficiency risk | 4320
    fat malabsorption risk | 4320
    anemia risk | 4320
    diarrhoea resolved | 4320
    