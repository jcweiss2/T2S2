65 years old | 0
female | 0
admitted to the hospital | 0
abdominal pain | -30
pancreatic head lesion | -30
history of stage IIIA lung cancer | -648
smoking history | -648
hypertension | -648
hypothyroidism | -648
dyslipidemia | -648
spiculated suprahilar RUL nodule | -648
lung-RADS 4X | -648
augmented activity in the RUL mass | -648
NSCLC | -648
adenocarcinoma | -648
lymph node sampling | -648
stage IIIA lung adenocarcinoma | -648
program death ligand-1 expression | -648
surgical resection | -648
carboplatin | -567
paclitaxel | -567
radiation therapy | -567
decrease in the RUL mass | -504
adjuvant immunotherapy | -504
durvalumab | -504
pneumonitis | -456
steroid taper | -456
increase in the RUL mass | -396
increase in the RUL mass | -252
respiratory symptom management | -252
radiation oncology clinic | -252
hematology-oncology clinic | -252
thoracic, abdominal, and pelvic CT scan | -168
stable lung nodules | -168
post-radiation changes | -168
radiation fibrosis | -168
epigastric pain | -30
constipation | -30
loss of appetite | -30
weight loss | -30
abdominal and pelvic CT scan | -30
mass in the head of the pancreas | -30
pancreatic ductal dilatation | -30
endoscopic ultra-sound-guided biopsy | 0
tumor cells | 0
nuclear pleomorphism | 0
prominent nucleoli | 0
irregular nuclear contours | 0
coarse chromatin | 0
CK7 | 0
TTF-1 | 0
Napsin-A | 0
CDX-2 | 0
KOC | 0
synaptophysin | 0
Smad-4 | 0
lung adenocarcinoma | 0
metastasized to the pancreas | 0
liver enzymes | 0
AST | 0
ALT | 0
ALP | 0
total bilirubin | 0
direct bilirubin | 0
CA 19.9 | 0
PET/CT scan | 30
fluorodeoxyglucose-avid mass | 30
SUV max | 30
palliative radiation therapy | 90
carboplatin | 90
pemetrexed | 90
generalized weakness | 120
dyspnea | 120
electrolyte derangements | 120
acute anemia | 120
hemoglobin nadir | 120
transfusion | 120
CT scan of the chest | 120
new left lower lobe nodule | 120
staging PET/CT scan | 180
decreased metabolic activity | 180
metabolic activity | 180
fatigue | 180
pulmonology clinic | 210
rapid response | 210
oxygen supplementation | 210
accessory muscles | 210
blood pressure | 210
heart rate | 210
increased dyspnea | 210
cough | 210
generalized weakness | 210
emergency department | 210
hospital admission | 210
right lung consolidation | 210
loculated pleural effusion | 210
acute hypoxic respiratory failure | 210
sepsis | 210
pneumonia | 210
broad-spectrum antibiotics | 210
vancomycin | 210
azithromycin | 210
cefepime | 210
oxygen supplementation | 210
bilevel-positive airway pressure | 210
altered mentation | 216
worsening hypoxemia | 216
vasopressor support | 216
palliative medicine team | 216
inpatient hospice care | 216
death | 216