77 years old | 0
man | 0
admitted to the hospital | 0
progressive lethargy | 0
shortness of breath | 0
septic shock | 0
hypotension | 0
hypoxia | 0
ventilatory support | 0
vasopressor support | 0
tube thoracostomy | 0
large left pleural effusion | 0
copious amounts of purulent fluid | 0
splenectomy | -8760
chemotherapy | -8760
non-Hodgkin's B-cell lymphoma | -8760
tumor recurrence | -5088
radiation therapy | -5088
progressive dysphagia | -5088
initiation of home TPN | -5088
esophagogastroduodenoscopy | -336
bleeding gastric ulcer | -336
cauterized | -336
chest computed tomography | 0
abdominal computed tomography | 0
oral contrast | 0
upper gastrointestinal series | 0
gastropleural fistula | 0
diagnostic laparoscopy | 0
bulky tumor | 0
laparoscopic GPF takedown | 0
partial sleeve gastrectomy | 0
intraoperative EGD | 0
fistulous tract patched with bovine pericardium mesh | 0
closed suction drain | 0
feeding jejunostomy tube | 0
malignant B-cell lymphoma | 0
quick initial recovery | 0
early extubation | 0
transfer out of the intensive care unit | 0
persistent anorexia | 0
pulmonary complications | 0
prolonged hospital course | 0
failing conservative therapy | 0
left thoracotomy | 0
pulmonary decortication | 0
debridement of an empyema | 0
discharged home | 1080
died | 1080
