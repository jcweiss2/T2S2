62 years old | 0
female | 0
admitted to the hospital | 0
type 2 diabetes mellitus | -672
repaglinide | -672
atypical chest pain | 0
coronary angiography | 0
no evidence of coronary disease | 0
superficial phlebitis | 48
venous perfusion | 48
backaches | 72
fever | 72
readmitted | 96
Glasgow Coma Scale score 15/15 | 96
fully alert | 96
no motor deficit | 96
no neck stiffness | 96
major inflammatory syndrome | 96
C-reactive protein level 47.8 mg/dl | 96
normal white blood cell count | 96
mildly impaired renal function | 96
serum creatinine level 2.1 mg/dl | 96
blood urea nitrogen 84 mg/dl | 96
no pulmonary infection | 96
no urinary infection | 96
amoxicillin | 96
clavulanic acid | 96
empirical antimicrobial therapy | 96
blood cultures grew S. aureus | 96
vancomycin | 96
oxacillin | 96
dysarthria | 120
drowsiness | 120
polypnea | 120
transferred to intensive care unit | 120
confuse | 120
disorientated | 120
stiff neck | 120
painful neck | 120
lumbar puncture | 120
purulent cerebrospinal fluid | 120
white blood cell count 31,800/mm3 | 120
neutrophils 85% | 120
lymphocytes 10% | 120
monocytes 5% | 120
CSF glucose 54 mg/dl | 120
lactate 13.5 mmol/l | 120
contrast-enhanced brain CT | 120
no ventriculitis | 120
no venous thrombosis | 120
Glasgow Coma Scale score 11/15 | 336
intubation | 336
mechanical ventilation | 336
major hypoxemia | 336
magnetic resonance imaging | 336
enlarged spinal cord | 336
T2-weighted images showed intramedullary hyperintensity | 336
diffuse leptomeningeal and focal intramedullary gadolinium enhancements | 336
signal abnormalities extended to medulla oblongata | 336
no hydrocephalus | 336
no brain edema | 336
brain stem auditory evoked potentials preserved | 336
no cortical somatosensory evoked potentials | 336
peripheral activities normal | 336
absence of P14 complex | 336
damage caudal to bulbomedullary junction | 336
neurological condition worsened | 360
spontaneous breathing disappeared | 360
ventilated in pressure control mode | 360
dysautonomic episodes | 360
hypotension | 360
extreme bradycardia | 360
complete quadriparesis | 360
anesthesia | 360
horizontal ophthalmoplegia | 360
conscious | 360
able to respond to simple questions | 360
blood cultures still positive for methicillin-sensitive S. aureus | 360
endocarditis ruled out | 360
MRI repeated | 456
signal hyperintensity extended | 456
necrotic damage | 456
all brain stem reflexes absent | 504
BAEPs absent | 504
wave I persisting | 504
ascendant pontine damage | 504
withdrawal of intensive care therapy | 504
cardiocirculatory failure | 504
death | 504
autopsy | 504
extensive leptomeningitis | 504
vasculitis | 504
secondary medullar ischemia | 504