44 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
admitted to the emergency department | 0 | 0 | Factual
left groin and inner thigh redness | -72 | 0 | Factual
pain | -72 | 0 | Factual
swelling | -72 | 0 | Factual
fever | -72 | 0 | Factual
chills | -72 | 0 | Factual
vomiting | -72 | 0 | Factual
treated with intravenous vancomycin | -24 | -24 | Factual
discharged on oral antibiotics | -24 | -24 | Factual
presented to the ED | 0 | 0 | Factual
afebrile | 0 | 0 | Factual
normotensive | 0 | 0 | Factual
tachycardia | 0 | 0 | Factual
mild tachypnea | 0 | 0 | Factual
left inner thigh and groin induration | 0 | 0 | Factual
morbidly obese | 0 | 0 | Factual
lactate 3.5 mmol/L | 0 | 0 | Factual
WBC 18.2 × 103 per mm3 | 0 | 0 | Factual
hemoglobin 12.3 g/dL | 0 | 0 | Factual
sodium 136 mmol/dL | 0 | 0 | Factual
glucose 225 mg/dL | 0 | 0 | Factual
creatinine 1.8 mg/dL | 0 | 0 | Factual
LRINEC score of 6 | 0 | 0 | Factual
bedside ultrasound performed | 0 | 0 | Factual
subcutaneous thickening | 0 | 0 | Factual
air | 0 | 0 | Factual
fascial fluid | 0 | 0 | Factual
started on intravenous vancomycin and piperacillin/tazobactam | 0 | 0 | Factual
surgery consulted | 0 | 0 | Factual
operative debridement | 0 | 0 | Factual
excision of 15 cm × 23 cm of tissue | 0 | 0 | Factual
septic shock | 0 | 0 | Factual
vasopressors | 0 | 0 | Factual
ventilator dependence | 0 | 0 | Factual
repeat washouts with minor debridements | 0 | 72 | Factual
lactate normalization | 72 | 72 | Factual
WBC down-trending | 72 | 72 | Factual
extubated | 120 | 120 | Factual
transferred to a step-down unit | 120 | 120 | Factual
plastic surgery consulted | 120 | 120 | Factual
wound vacuum-assisted closure (V.A.C.) device placed | 216 | 216 | Factual
transferred to the plastic surgery service | 216 | 216 | Factual
discharged home | 672 | 672 | Factual
skin graft | 672 | 672 | Factual