28 years old | 0
African American male | 0
multiple sclerosis | -168
generalized seizure | 0
midazolam | -1
altered mental status | 0
fever | 0
heart rate of 103 beats per minute | 0
blood pressure of 147/74 mmHg | 0
respiratory rate of 16 | 0
oxygen saturation of 97% | 0
lethargic | 0
cardiopulmonary exam normal | 0
abdominal exam normal | 0
no audible murmurs | 0
no bruits | 0
pulses 2+ in upper and lower extremities | 0
no peripheral edema | 0
no notable skin lesions | 0
elevated white blood cell count | 0
elevated creatinine kinase | 0
elevated lactate | 0
chest radiograph normal | 0
CT scan of head showed hypodensities | 0
blood cultures drawn | 0
urine cultures drawn | 0
broad spectrum antibiotics started | 0
vancomycin | 0
piperacillin/tazobactam | 0
levetiracetum | 0
acetaminophen | 0
medical intensive care team consulted | 0
neurology team consulted | 0
admitted to medical telemetry | 0
plan for TTE | 0
plan for vEEG monitoring | 0
aerobic blood cultures grew gram positive cocci | 48
Staphylococcus pettenkoferi | 72
TTE showed no valvular vegetations | 48
TTE showed no regurgitation | 48
vEEG showed nonconvulsive focal seizures | 48
levetiracetum continued | 48
antibiotic regimen de-escalated | 48
vancomycin continued | 48
ceftriaxone started | 48
fevers persisted | 48
blood cultures showed no growth | 48
TEE performed | 96
TEE showed micro-perforations in left coronary leaflet | 96
TEE showed trace to mild aortic regurgitation | 96
structural heart team consulted | 96
no surgical intervention advised | 96
MRI of brain showed white matter lesions | 120
decision to discontinue antibiotics | 120
antiepileptic regimen titrated | 120
lacosamide started | 120
previous hospitalization | -720
septic shock | -720
CoNS bacteremia | -720
broad spectrum antibiotics | -720
TTE negative for valvular vegetations | -720
lumbar puncture showed no infectious etiology | -720
steroids given for multiple sclerosis flare | -720
discharged from previous hospital | -720
discharged from current hospital | 168
plan for primary care follow-up | 168
plan for neurology follow-up | 168