55 years old | 0
    morbidly obese | 0
    male | 0
    diabetes mellitus | 0
    end-stage renal disease | 0
    hemodialysis | 0
    peripheral vascular disease | 0
    left below knee amputation | 0
    right above knee amputation | 0
    right extra anatomical axillobifemoral bypass graft | 0
    right-sided abdominal pain | -48
    vomiting | -48
    fever | -48
    conscious | 0
    alert | 0
    oriented | 0
    pale | 0
    sick | 0
    temperature of 37.8°C | 0
    blood pressure of 150/90 mmHg | 0
    oxygen saturation of 95% | 0
    distended abdomen | 0
    tympanic abdomen | 0
    right upper quadrant tenderness | 0
    right flank tenderness | 0
    total leukocyte count 20 × 10³ | 0
    hemoglobin 10.7 gm% | 0
    acidotic | 0
    pH 7.33 | 0
    laboratory evidence of end-stage renal disease | 0
    chest X-ray demonstrated air under the right hemi-diaphragm | 0
    evaluated by general surgeon | 0
    impression of perforated viscous | 0
    computed tomography scan with contrast | 0
    right perinephric collection | 0
    extension into right sub-phrenic region | 0
    gas in right collecting system | 0
    gas in urinary bladder | 0
    no gas in renal parenchyma | 0
    right atrial thrombus | 0
    started on parenteral antibiotics | 0
    admitted to intensive care unit | 0
    very high risk for surgical intervention | 0
    trial of percutaneous drainage | 0
    failed percutaneous drainage | 0
    dry collection | 0
    very thick collection | 0
    evaluated by anesthetist | 0
    not fit for general anesthesia | 0
    minimal life-saving procedure | 0
    epidural anesthesia | 0
    sedation | 0
    open drainage | 0
    very thick collection | 0
    foul smelly collection | 0
    loculated perinephric collection | 0
    loculated sub-phrenic collection | 0
    cystoscopy | 0
    abnormal bladder mucosa | 0
    multiple cystic lesions | 0
    air bubbles in bladder | 0
    ureteric Double J stent inserted | 0
    drain collecting system | 0
    urethral catheter | 0
    drain bladder | 0
    reasonably well during procedure | 0
    condition deteriorated | 24
    culture showed Klebsiella pneumoniae extended-spectrum β-lactamase | 24
    condition continued to deteriorate | 48
    died | 48
    severe sepsis | 48
    multiple organ failure | 48