33 weeks gestation | 0
preterm male | 0
precipitous vaginal delivery | 0
acute onset of labor | -1
rupture of membranes | -1
respiratory distress | 0
intubated | 0
mechanically ventilated | 0
surfactant administered | 0
Apgar scores 7 at 1 min | 0
Apgar scores 8 at 5 min | 0
birth weight 1870 g | 0
caffeine administered | 1
ampicillin administered | 1
amikacin administered | 1
concern of neonatal sepsis | 1
hypotensive | 2
normal saline boluses | 2
dobutamine drip | 2
cefepime administered | 3
blood cultures negative | 72
antibiotics discontinued | 72
routine cranial ultrasound normal | 72
echocardiogram normal | 72
initial cranial circumference 31 cm | 72
neurological examination normal | 72
abdominal distention | 144
pain on examination | 144
necrotizing enterocolitis suspected | 144
vancomycin administered | 144
meropenem administered | 144
pneumatosis intestinalis not observed | 144
portal venous gas not observed | 144
blood cultures no pathogen | 144
antimicrobial treatment | 144
enteral feedings started | 144
cranial circumference increased | 432
anterior fontanelle bulging | 432
cefipime administered | 432
hypernatremia | 432
enteral sterile water drip | 432
ventricular puncture | 432
cerebrospinal fluid collected | 432
no leukocytes in CSF | 432
glucose decreased in CSF | 432
protein elevated in CSF | 432
cranial ultrasound significant hydrocephalus | 432
no intraventricular hemorrhage | 432
no mass seen | 432
magnetic resonance imaging | 432
hydrocephalus | 432
apparent right frontoparietal cerebral arteriovenous malformation | 432
MR angiography | 432
large saccular aneurysm of right middle cerebral artery | 432
Candida lusitaniae isolated | 480
methicillin-resistant Staphylococcus epidermidis identified | 480
antimicrobial coverage changed | 480
vancomycin administered | 480
amphotericin B administered | 480
neurosurgery consulted | 480
severe apnea | 504
hypotonia | 504
lethargy | 504
resuscitation failed | 504
rupture of aneurysm suspected | 504
death | 504