35 years old | 0
female | 0
gave birth to healthy twins | 0
in vitro fertilization | -280
facial nerve paresis | -672
severe headache | 24
generalized tonic–clonic seizures | 24
loss of consciousness | 24
arterial blood pressure 195/110 mmHg | 24
heart rate 120 beats/min | 24
provisional diagnosis of eclampsia | 24
transferred to the intensive care unit | 24
antihypertensive therapy | 24
intravenous infusion of magnesium sulphate | 24
ebrantil | 24
20% manitol | 24
diazepam | 24
bilateral vision loss | 48
complete blood count normal | 48
liver function tests normal | 48
clotting parameters normal | 48
electrocardiogram normal | 48
proteinuria 2+ | 48
cortical blindness | 48
mild right-sided facial nerve paresis | 48
multislice computed tomography scan | 48
hypodensity of the posterior white matter | 48
MRI | 72
T2- and fluid-attenuated inversion recovery-weighted images hyperintense signals | 72
vasogenic edema | 72
stabilization of the general condition | 72
moved to an obstetrics clinic | 120
oral antihypertensive medication | 120
enalapril maleate | 120
methyldopa | 120
human albumin | 120
follow-up ophthalmological examinations | 120
significant bilateral improvement of the visual function | 120
best-corrected visual acuity 1.0 | 120
visual field image | 120
peripheral relative scotoma | 120
depressed sensitivity of the paracentral left visual field | 120
follow-up MRI | 192
significant regression of the edema | 192
discrete residual changes over the posterior horns of the side ventricles | 192
discharged from the clinic | 216
oral antihypertensive therapy | 216
physical therapy for the paresis of the facial nerve | 216