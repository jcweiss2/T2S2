61 years old | 0
female | 0
rectal prolapse | 0
hypothyroidism | 0
depression | 0
hypertension | 0
dyslipidemia | 0
esophageal reflux | 0
urinary retention | 0
indwelling urinary catheter | 0
chronic back pain | 0
opioids | 0
two previous vaginal childbirths | 0
prolapsed rectum 20 cm in length | 0
viable mucosa | 0
shallow ulceration | 0
reducible | 0
recurred immediately | 0
preoperative colonoscopy | -168
poor bowel preparation | -168
elective perineal proctosigmoidectomy | 0
malaise | 168
lower abdominal pain | 168
decreased level of consciousness | 168
hypotension | 168
leukocytosis | 168
acute kidney injury | 168
urinalysis positive for nitrates | 168
30+ leukocytes/high power field | 168
urosepsis | 168
blocked urinary catheter | 168
ICU admission | 168
resuscitation with intravenous fluids | 168
vasopressors | 168
rectal prolapse on physical examination | 168
herniating sigmoid colon | 192
necrotic sigmoid colon | 192
emergency Hartmann’s procedure | 192
sacral rectopexy | 192
reduction of prolapse and strangulated sigmoid | 192
perforation of the rectum | 192
ischemic necrosis of the resected sigmoid | 192
viable margins | 192
ICU post-operatively | 192
transfer to surgical ward | 216
recovery | 216
functioning colostomy | 216
normalized bladder function | 216
removal of indwelling catheter | 216
transfer to rehabilitation facility | 504
discharge home | 672
follow-up | 1008