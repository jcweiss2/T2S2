71 years old | 0
female | 0
chronic obstructive pulmonary disease | 0
atrial fibrillation | 0
bladder cancer | 0
type 2 insulin-dependent diabetes mellitus | 0
urinary tract infection | -24
sepsis | -24
admitted to the hospital | 0
home dose of 30 units per day of glargine insulin | -24
insulin sliding scale | -24
blood glucose became unresponsive to home dose of insulin | 0
hyperosmolar hyperglycemic state | 0
normal anion gap | 0
normal pH | 0
normal sodium level | 0
increasing glargine dose | 0
glargine dose substantially increased | 12
blood glucose remained uncontrolled | 12
aspart and NPH boluses | 12
aspart and NPH boluses minimally effective | 12
transitioned to regular insulin drip | 24
regular insulin drip initially helpful | 24
regular insulin drip lost efficacy | 48
insulin drip titrated up to maximum dose of 1620 units | 48
total daily insulin | 48
blood glucose remained above 400mg/dL | 48
test for insulin autoantibodies sent | 48
test for insulin autoantibodies negative | 72
producing neutralizing antibodies to insulin | 72
identified detemir as a possible solution | 72
administered one dose of 40 units of detemir | 96
blood glucose dropped 292mg/dL | 120
detemir titrated to optimal dose | 120
insulin drip down-titrated and discontinued | 120
average daily blood glucose maintained at 181mg/dL | 168
transferred to the ward | 168
discharged to a rehabilitation facility | 216
blood sugars maintained between 100 and 200mg/dL | 216
died during a subsequent hospitalization for acute respiratory failure | 1000