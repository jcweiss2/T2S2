62 years old | 0
male | 0
admitted to the hospital | 0
shortness of breath | 0
altered mental status | 0
hypotensive | 0
hypoxic respiratory failure | 0
intubated | 0
pressors | 0
transferred to the intensive care unit | 0
bilateral infiltrates | 0
right pleural effusion | 0
normal sinus rhythm | 0
new low voltage | 0
old left-axis deviation | 0
hyponatremia | 0
acute kidney injury | 0
leukocytosis | 0
lymphopenia | 0
mildly macrocytic anemia | 0
coagulation panel within normal limits | 0
elevated d-dimer | 0
negative serial troponins | 0
pericardial effusion | 0
tamponade physiology | 0
pericardiocentesis | 0
sanguinous fluid drained | 0
right heart catheterization | 0
nasopharyngeal swab for COVID-19 negative | 0
bronchoalveolar lavage sample positive for COVID-19 | 48
hydroxychloroquine | 48
ribavirin | 48
lopinavir-ritonavir combination | 48
steroids | 48
tocilizumab | 48
anakinra | 48
inhaled epoprostenol | 48
pressor and inotropic support decreased | 120
septic shock | 120
weaned off inotropic and pressor support | 240
thoracentesis | 240
transudative nonbloody fluid drained | 240
bacterial and fungal cultures of pleural fluid negative | 240
renal failure | 240
continuous renal replacement therapy | 240
upper gastrointestinal bleeding | 240
conservative management | 240
lower extremity deep vein thrombosis | 240
extubated | 432
discharged | 672
follow-up chest computed tomography | 672
ground-glass opacities | 672
residual right pleural effusion | 672
coronary artery disease | -8760
drug-eluting stent implantation | -8760
hypertension | -8760
hyperlipidemia | -8760
diabetes mellitus | -8760
chronic obstructive pulmonary disease | -8760
alcoholism | -8760
morbid obesity | -8760
COVID-19 pneumonia | 0 
pericardial effusion caused by COVID-19 | 0 
hemorrhagic pericardial effusion | 0 
cardiac tamponade | 0 
pericardiocentesis | 0 
pericardial fluid analysis | 0 
pericardial fluid cytology | 0 
pericardial fluid cultures | 0 
pleural effusion | 0 
pleural fluid analysis | 240 
pleural fluid cultures | 240 
renal failure requiring continuous renal replacement therapy | 240 
upper gastrointestinal bleeding resolved with conservative management | 240 
lower extremity deep vein thrombosis | 240 
extubation | 432 
discharge | 672 
follow-up | 672 
clinic follow-up chest computed tomography | 672 
bilateral ground-glass opacities | 672 
residual right pleural effusion | 672