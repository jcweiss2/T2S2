67 years old | 0
woman | 0
admitted to the hospital | 0
near-obstructing adenocarcinoma of the right colon | 0
laparoscopic-assisted extended right hemicolectomy | 0
discharged | -120
presented to emergency department | -168
diffuse abdominal pain | -168
hematemesis | -168
subjective fevers | -168
CT abdomen | -168
free intraperitoneal fluid | -168
pneumoperitoneum | -168
broad spectrum antibiotics | -168
exploratory laparotomy | -168
succus | -168
anastomotic leak | -168
anastomosis resected | -168
end ileostomy created | -168
stable vital signs | -168
low grade tachycardia | -168
extubated | -168
persistent obtundation | -168
brought to ICU | -168
oxygen saturation above 95% | -168
supplemental oxygen | -168
oropharyngeal airway | -168
nasopharyngeal airway | -168
failed to regain consciousness | -168
apneic | -168
bag valve mask ventilation | -168
naloxone | -168
glycopyrrolate | -168
neostigmine | -168
no clinical improvement | -168
normal blood glucose | -168
arterial blood gas | -168
respiratory acidosis | -168
pH 7.03 | -168
PCO2 107 | -168
PaO2 375 | -168
re-intubated | -168
hypercapnic respiratory failure | -168
sedating medications held | -168
no neurologic improvement | -168
cerebral imaging | -168
CT head | -168
acute cerebellar herniation | -168
diffuse cerebral edema | -168
neurosurgery consulted | -168
external ventricular drain | -168
maximal medical therapy | -168
hypertonic saline | -168
head elevation 30 degrees | -168
normotension | -168
normoglycemia | -168
levetiracetam | -168
seizure prophylaxis | -168
MRI | -168
PRES diagnosis | -168
neurologic function recovery | 0
discharged to rehabilitation | 792
ileostomy reversal | 3600
pre-operative quality of life | 3600
complete resolution of neurological symptoms | 3600
normalization of neuroimaging | 3600
