82 years old | 0
female | 0
admitted to emergency department | 0
hematemesis | 0
high-grade suspicion of upper gastrointestinal bleeding | 0
decreased hemoglobin | 0
elevated infection signs | 0
leukocyte count 27 × 10^9/L | 0
C-reactive protein 15 mg/dL | 0
soft abdomen | 0
diffuse tenderness | 0
no voluntary guarding | 0
septic shock | 0
hemodynamic instability | 0
loss of vigilance | 0
referred to intensive care unit | 0
need for intubation | 0
gastroscopy | 0
no endoscopic evidence for upper gastrointestinal bleeding | 0
spontaneous penetration of the gallbladder | 0
plenty gallstones in the duodenal bulb | 0
computed tomography | 0
chronic cholecystitis | 0
pneumobilia | 0
gallbladder penetration in the duodenal bulb | 0
entry of gallstones in the intestine | 0
reflective intestinal atony | 0
dilated stomach filled with contrast medium | 0
Bouveret syndrome | 0
open cholecystectomy | 24
gallstone salvage from the duodenum | 24
discharged | 120
diabetes | -720
arterial hypertension | -720
no history of biliary symptoms | 0 
gallstone penetration in the duodenal bulb | 0 
biliary enteric fistula not found | 24 
gallstone ileus | 0 
upper gastrointestinal bleeding suspected | 0 
mechanical removal of impacted stones | 24 
endoscopic removal | 24 
surgical removal | 24 
CT scan | 0 
endoscopy | 0 
informed consent obtained | 0 
no conflict of interest | 0 
no financial support | 0