65 years old | 0
female | 0
admitted to the hospital | 0
recurrent fever | -744
nausea | -168
vomiting | -168
highest body temperature 38 ℃ | -744
neutrophil count 6.96×10^9/L ↑ | 0
monocyte count 0.86×10^9/L ↑ | 0
lymphocyte percentage 14.9% ↓ | 0
red blood cell count 3.17×10^12/L ↓ | 0
hemoglobin content 87 g/L ↓ | 0
hematocrit 0.28 L/L ↓ | 0
average red blood cell hemoglobin concentration 312 g/L ↓ | 0
platelet count 363×10^9/L ↑ | 0
platelet distribution width 8.3 fl ↓ | 0
C-reactive protein (CRP) 52.01 mg/L ↑ | 0
diagnosed with secondary infectious thrombocytopenia | 0
diagnosed with gram-negative bacilli septicemia (Klebsiella pneumoniae) | 0
diagnosed with liver abscess | 0
diagnosed with bilateral lung inflammation | 0
diagnosed with type 2 diabetes | 0
diagnosed with hypertension grade 3 (extremely high risk) | 0
given vancomycin | 0
given caspofungin | 0
given dexamethasone | 0
given posaconazole oral suspension | 0
liver abscess puncture and drainage treatment | 24
inflammatory indexes decreased | 48
light perception disappeared in the left eye | 72
eyelid redness and pain | 72
purulent secretion | 72
repeated fever | 72
left-sided headache | 72
diagnosed with endogenous endophthalmitis (left) | 72
diagnosed with orbital cellulitis (left) | 72
diagnosed with rubeosis iridis (left) | 72
diagnosed with exudative retinal detachment (left) | 72
diagnosed with diabetic retinopathy (right) | 72
intravitreal injection with vancomycin and ceftazidime | 96
symptoms relieved | 120
left eyeball enucleation | 240
fever again after the operation | 264
given moxifloxacin | 264
given sulperazon | 264
temperature elevated again | 288
CT examination | 288
inflammation of both lungs | 288
pericardial effusion | 288
bilateral pleural thickening and effusion | 288
atelectasis in right inferior lobe | 288
liver cyst | 288
liver abscess | 288
right renal cyst | 288
myoma of the uterus | 288
history of hypertension | -8760
highest blood pressure 180/100 mmHg | -8760
oral valsartan | -8760
controlled blood pressure at 140/80 mmHg | -8760
no special history of other systematic diseases | 0
no history of surgery | 0
no history of blood transfusion | 0
no history of drug allergy | 0
diagnosed with sepsis | 0
diagnosed with secondary thrombocytopenia | 0
diagnosed with liver abscess | 0
diagnosed with gram-negative bacilli sepsis (Klebsiella pneumoniae) | 0
diagnosed with infection of lumbar vertebrae | 0
diagnosed with mesenteric panniculitis | 0
diagnosed with pelvic effusion | 0
diagnosed with pericardial effusion | 0
diagnosed with suppurative endophthalmitis (left) | 0
diagnosed with orbital cellulitis (left) | 0
diagnosed with retinal detachment (left) | 0
diagnosed with choroidal detachment (left) | 0
diagnosed with type 2 diabetes retinopathy (right) | 0
diagnosed with cortical senile cataract (right, immature stage) | 0
diagnosed with type 2 diabetes | 0
diagnosed with type 2 diabetes nephropathy stage I | 0
diagnosed with type 2 diabetic peripheral neuropathy | 0
diagnosed with hypertension grade 3 (extremely high risk) | 0
diagnosed with hepatic cyst | 0
diagnosed with renal cyst | 0
diagnosed with hypoproteinemia | 0
diagnosed with coronary atherosclerotic heart disease | 0
diagnosed with lacunar cerebral infarction | 0
diagnosed with moderate anemia | 0
diagnosed with risk of malnutrition | 0
convulsion with unconsciousness | 432
transferred to the respiratory intensive care unit | 432
CT examination | 432
lacunar infarction | 432
encephalomalacia | 432
bilateral pleural effusion | 432
lower lobe of the right lung insufficiently inflated | 432
intracranial infection | 432
lumbar puncture | 432
cerebrospinal fluid (CSF) analysis | 432
microbial metagenomic next-generation sequencing (mNGS) | 432
biochemistry analysis | 432
glucose <1.1 mmol/L ↓ | 432
chlorine 108 mmol/L ↓ | 432
CSF protein >3,000 mg/L ↑ | 432
mNGS results | 432
high sequence of Klebsiella pneumoniae | 432
drug-resistant gene SHV-type beta-lactamases (blaSHV) | 432
given 2 g meropenem q8h prolonged for 3 hours | 432
body temperature improved | 456
blood routine improved | 456
CRP improved | 456
CT examination | 720
pulmonary edema and pleural effusion dissipated and absorbed | 720
CSF analyses | 744
chlorine 119 mmol/L ↓ | 744
micro amount of proteins 1,107 mg/L ↑ | 744
microalbumin 816.3 mg/L ↑ | 744
immunoglobulin G 308.5 mg/L ↑ | 744
α2-macroglobulin 18.5 mg/L ↑ | 744
β2-microglobulin 2.67 mg/L ↑ | 744
discharged from the hospital | 744