60 years old | 0
male | 0
presented to an outside hospital | 0
fever | 0
hypotension | 0
altered mental status | 0
low back pain | -24
epigastric pain | -24
chills | -24
vomiting | -24
disoriented | -24
dusky discoloration of face and extremities | -24
splenectomy in 1974 | -336
complicated cholecystectomy in 2014 | -96
no medications | 0
denied recent travel | 0
denied sick contacts | 0
dog bites | -168
scratches from German shepherd | -168
intravenous fluids | 0
packed red blood cells | 0
levofloxacin | 0
CT scan chest, abdomen, pelvis | 0
bilateral lung parenchymal opacities | 0
acute respiratory distress syndrome | 0
intubated for worsening confusion | 0
intubated for hypoxemia | 0
transferred to our hospital | 0
heavily sedated | 0
mechanically ventilated | 0
blood pressure 80/58 mmHg | 0
heart rate 111 bpm | 0
temperature 38.5°C | 0
coarse breath sounds | 0
absent peripheral pulses | 0
cold, dusky extremities | 0
mottling of the skin | 0
violaceous purpura on thighs | 0
superficial linear scratches | 0
erythema on upper extremities | 0
vasopressors administered | 0
blood cultures collected | 0
white blood cell count 18.0 × 10^9/L | 0
platelet count 14 × 10^9/L | 0
INR 1.7 | 0
fibrinogen 178 mg/dL | 0
creatinine 3.8 mg/dL | 0
lactate 5.6 mmol/L | 0
PaO2 60 mmHg | 0
urinalysis 3 erythrocytes | 0
urinalysis 3 leukocytes | 0
negative leukocyte esterase | 0
positive nitrite | 0
2+ protein | 0
1+ bilirubin | 0
>50 bacteria | 0
broad-spectrum antibiotics | 0
vancomycin | 0
cefepime | 0
ampicillin | 0
doxycycline | 0
acyclovir | 0
CT head negative | 0
lumbar puncture performed | 0
11 nucleated cells/µL | 0
531 erythrocytes/µL | 0
glucose 81 mg/dL | 0
protein 100 mg/dL | 0
CSF Gram stain negative | 0
herpes simplex virus PCR negative | 0
ampicillin discontinued | 0
acyclovir discontinued | 0
continuous renal replacement therapy | 0
Wright's stain neutrophils with bacterial rods | 0
Gram-negative rods confirmed | 0
dog bites history | 0
cefepime changed to piperacillin-tazobactam | 0
ciprofloxacin added | 0
admission blood cultures negative | 0
plasma sent for NGS on day 4 | 96
NGS detected C canimorsus | 96
antibiotic regimen narrowed | 96
blood culture grew Gram-negative rods | 120
MALDI-TOF failed | 120
16S sequencing attempted | 120
Clostridium difficile colitis | 264
Candida tropicalis fungemia | 264
recurrent sepsis | 384
progressive gangrene of extremities | 384
transition to comfort care | 912
died | 960
16S sequencing confirmed C canimorsus | 960
