55 years old | 0
male | 0
admitted to the hospital | 0
work-related accident | -1
pulled into a cement mixer | -1
right lower limb completely torn off | -1
conscious and drowsy | -1
patent airway | -1
injury severity score 75 | -1
blood pressure 70 to 85/40 to 50 mmHg | -1
pulse 120 beats per min | -1
bandaging applied with strong mechanical pressure | -1
intravenous rehydration treatment | -1
oxygen inhalation | -1
open wound over the right costal arch | 0
wound traversing toward the right pubic tubercle | 0
wound extending through the perineum | 0
wound ending near the right sacroiliac joint | 0
skin stripped of skin | 0
peritoneum holding in the abdominal contents | 0
cement and foreign matters covering the wound | 0
displaced extremity cold | 0
displaced extremity extensively crushed | 0
displaced extremity pulseless | 0
fluid resuscitation | 0
tetanus prophylaxis | 0
broad-spectrum antibiotics | 0
computed tomography images | 0
loss of right lower limb | 0
loss of right lower abdominal wall | 0
right ilium, right pubis, and right ischium lost | 0
no intra-abdominal injury | 0
bladder intact | 0
rectum intact | 0
CT angiography | 0
transection of right common iliac vessels | 0
therapeutic strategy developed | 0
general anesthesia | 0
systemic exploration of pelvic wound | 0
gross loss of skin from right lower abdomen | 0
severely contaminated peritoneum | 0
bowel peristalsis observed | 0
right side of scrotum avulsed | 0
exposed testis and spermatic cord extravasated | 0
soft tissue surrounding anus and right ilium missing | 0
sacrum exposed | 0
arterial bleeding observed | 0
right external and internal iliac vessels transected | 0
right external and internal iliac vessels thrombosed | 0
main vessels ligated and sutured | 0
wound washed with saline, hydrogen peroxide, and iodophor diluent | 0
wound left open | 0
VSD device applied | 0
rectal tube applied | 0
packed red blood cells transfused | 0
crystalloids transfused | 0
colloids transfused | 0
mechanical ventilation support | 1
blood transfusion | 1
aggressive fluid resuscitation | 1
broad-spectrum antibiotics | 1
antifungal medication | 1
fever persisted | 1
white blood cell count peaked | 5
pneumothorax in right lung | 5
pneumonia in left lung | 5
closed drainage performed | 5
second operation for debridement | 6
granulation tissue observed | 6
devitalized tissue removed | 6
pus samples collected | 6
repetitive irrigation and debridement | 6
VSD therapy continued | 6
Proteus mirabilis and Providencia alcalifaciens isolated | 6
Pseudomonas aeruginosa isolated | 9
antibiotic regimen changed | 9
diverting colostomy performed | 14
body temperature remained high | 14
body temperature dropped | 25
skin defect well defined | 21
skin defect area 28 x 21 cm2 | 21
psychiatric management | 21
nutritional management | 21
chronic pain management | 21
VSD therapy discontinued | 56
skin defect closed by split-skin graft | 56
patient able to walk with crutches | 70
patient performed squatting maneuvers | 70
patient discharged | 72
semi-laparotomy prosthesis applied | 150
wound healed | 365
patient retired due to disability | 365
patient able to take care of himself | 365
phantom pain | 365
no symptoms of depression | 365