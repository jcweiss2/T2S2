90 years old | 0
male | 0
Caucasian | 0
BMI = 22.7 kg/m2 | 0
mild dementia | -8760
hypertension | -8760
atrial fibrillation | -8760
abdominal pain | -72
nausea | -72
vomiting | -72
diarrhea | -72
antihypertensive medications | -8760
no anticoagulants | -8760
no tobacco | -8760
no ethanol | -8760
no drugs | -8760
colonoscopy examination | -8760
normal colonoscopy | -8760
admitted to the VANTHCS Emergency Department | 0
acute distress | 0
diaphoretic | 0
temperature of 96.6° Fahrenheit | 0
heart rate of 117 beats per minute | 0
blood pressure of 126/72 mm/Hg | 0
irregularly irregular rhythm | 0
abdomen soft | 0
abdomen distended | 0
tenderness to palpation | 0
tenderness localized to the left lower quadrant | 0
hematocrit of 49.1% | 0
hemoglobin of 16.1 g/dL | 0
white count of 7.3 K/uL | 0
creatinine of 1.53 mg/dL | 0
potassium of 3.1 mmol/L | 0
albumin of 3.8 g/dL | 0
liver function tests within normal limits | 0
international normalized ratio (INR) within normal limits | 0
CT exam | 0
inflammation in the mesentery of the small bowel | 0
pneumoperitoneum | 0
admitted to the intensive care unit | 0
intravenous fluids | 0
serial abdominal exams | 0
indwelling bladder catheter | 0
broad-spectrum antibiotics | 0
presumptive diagnosis of diverticulitis | 0
initially responded favorably to fluid resuscitation | 2
initially responded favorably to antibiotic treatment | 2
developed tachycardia | 4
abdominal exam changed from localized to diffuse abdominal tenderness | 4
taken to the operating room | 4
exploratory laparotomy | 4
sigmoid redundant | 4
sigmoid demonstrated no abnormalities | 4
sigmoid diverticula | 4
uninflamed | 4
non-perforated diverticula | 4
appendix normal | 4
cecum normal | 4
right colon normal | 4
evisceration of the bowel | 4
jejunum adherent to the left colon | 4
multiple jejunal diverticula | 4
perforation found in one of them | 4
small bowel resection | 4
hand-sewn anastomosis | 4
recovered well from the operation | 168
discharged to a skilled nursing facility | 168
pathological examination | 168
no malignancy | 168
multiple jejunal diverticula | 168
perforated JD | 168
no enterolith | 168