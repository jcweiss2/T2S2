46 years old | 0
woman | 0
diagnosed with severe community acquired pneumonia | 0
respiratory failure | 0
septic shock | 0
acute renal failure | 0
right subclavian vein central venous line placed | 0
volume resuscitation | 0
vasopressors started | 0
intubated | 0
mechanical ventilation | 0
transferred to medical intensive care unit | 0
left peripherally inserted central venous catheter placed | 24
right femoral central venous line placed | 24
routine chest X-ray performed | 42
guidewire lodged partly in heart detected | 42
bedside ultrasonography performed | 42
guidewire traced in inferior vena cava | 42
guidewire up to level of renal veins | 42
taken to interventional radiology suite | 42
right femoral catheter removed | 42
proximal straight end of guidewire found inside tip of central venous catheter | 42
guidewire grasped | 42
guidewire removed | 42
loss of guidewire inside vessel | 0
failure to adhere to good practice | 0
failure to withdraw guidewire until proximal end comes out of catheter port | 0
failure to hold guidewire while advancing catheter beyond skin entry site | 0
