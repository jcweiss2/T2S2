845-gram male | 0
24 weeks' gestation | 0
born to a 23-year-old gravida two African-American mother | 0
emergent cesarean section | 0
infant arrived limp | 0
infant arrived blue | 0
infant arrived without cry | 0
bacterial vaginosis | -4032
vaginal candidiasis | -4032
clinical chorioamnionitis | -4032
Apgar score 1 at 1 minute | 0
Apgar score 6 at 10 minutes | 0
intubation | 0
admitted to NICU | 0
passed meconium | 0
normal physical exam | 0
feeding intolerance | -312
lethargy | -312
moderate abdominal distention | -312
sepsis workup initiated | -312
leukocytosis 41,500/μL | -312
thrombocytopenia | -312
Candida albicans fungemia | -312
abdominal ultrasound showing intra-abdominal fluid | -312
inferior right hepatic lobe abscess | -312
concern for necrotizing enterocolitis | -312
abdominal X-rays | -312
paracentesis | -312
brown feculent fluid | -312
gasless abdomen on X-rays | -312
pediatric surgery consultation | -312
high suspicion of intestinal perforation | -312
grade III necrotizing enterocolitis | -312
emergent exploratory laparotomy | -312
attending surgeon | 0
3rd year surgical resident | 0
feculent spillage | -312
necrosed colon | -312
cecal perforation | -312
necrosis of the ascending colon | -312
necrosis of the proximal transverse colon | -312
small bowel examined | -312
ligament of Treitz to terminal ileum intact | -312
well-perfused small bowel | -312
abdomen washed out | -312
liver examined | -312
no notable abscess | -312
subhepatic abscess opened | -312
evacuated subhepatic abscess | -312
right hemicolectomy | -312
end ileostomy | -312
mucus fistula | -312
postoperative day 5 | 120
abdominal distention | 120
increased oxygen requirement | 120
persistent acidosis | 120
additional exploratory laparotomy | 120
large intraabdominal abscess | 120
right upper quadrant abscess evacuated | 120
peritoneal drain placement | 120
Candida albicans culture | 120
coagulase negative Staphylococci culture | 120
pathologic examination of resected colon | 120
pseudohyphae on H&E | 120
pseudohyphae on GMS staining | 120
mucosal invasion | 120
fungemia resolved | 2160
ostomy takedown | 2160
discharged home | 2160
tolerating enteral feeds | 2160
systemic Candida infection | 0
antifungal medications initiated | -480
medications continued for 10 weeks | 1680
complete clearance of infection | 1680
clinic follow up | 2160
excellent recuperation | 2160
regular bowel movements | 2160
good feeding tolerance | 2160
