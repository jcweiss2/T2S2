20 years old | 0
G1P1001 | 0
presented to an outside hospital | -720
cough | -720
worsening shortness of breath | -720
15-month history of amenorrhea | -10800
vaginal delivery | -10800
two months of morning sickness | -1440
evaluation for pulmonary embolism | -720
infectious etiologies | -720
beta-HCG of approximately 900,000 mIU/mL | -720
adnexal mass | -720
bilateral diffuse pulmonary nodules | -720
intubated due to hypoxemia | -720
empiric antibiotics | -720
septic shock | -720
ventilatory requirements increased | -720
FiO2/PaO2 ratio of 69 | -720
100% FiO2 | -720
hypercarbia to 80 mmHg | -720
increasing positive end-expiratory pressure | -720
lung-protective ventilatory strategies | -720
paralysis | -720
evaluated by multidisciplinary team | -720
transferred for ECMO cannulation | -720
transesophageal echocardiogram | 0
acute right ventricular failure | 0
severe tricuspid regurgitation | 0
dilated right ventricle | 0
moderate to severe systolic dysfunction | 0
intra-atrial septal bowing | 0
underwent cannulation with dual-lumen RVAD | 0
ECMO circuit | 0
dilation and curettage | 0
heparin infusion | 0
weaned from vasopressors | 3
beta-HCG 917,929 mIU/mL | 0
clinical diagnosis of GTN | 0
FIGO stage III | 0
pulmonary lesions | 0
WHO score 14 | 0
induction chemotherapy cisplatin | 24
induction chemotherapy etoposide | 24
beta-HCG fell to 707,706 mIU/mL | 48
AFP less than 0.6 ng/mL | 48
LDH 670 U/L | 48
inhibin B 20 pg/mL | 48
extubated | 48
ECMO circuit complication | 48
acute oxygenator failure | 48
acute tachycardia | 48
hypoxia | 48
hypotension | 48
vasopressor support | 48
ECMO circuit exchanged | 48
reintubation avoided | 48
final pathology from dilation and curettage | 0
no chorionic villi | 0
no fetal parts | 0
no implantation site | 0
no neoplasm | 0
gestational type endometrium with breakdown | 0
complex multi-cystic left adnexa | -720
CT-guided biopsy of pelvic mass | 144
fragments of corpus luteum cyst | 144
thrombocytopenia | variable
nadir platelet 33 10^3/uL | variable
neutropenia | variable
ANC nadir 35 10^3/uL | variable
delayed subsequent doses of induction chemotherapy | variable
beta-HCG continued to fall | variable
MRI brain negative for metastatic lesions | variable
respiratory status improved | variable
decannulated from ECMO | 240
clot on distal tip of cannula | 240
transthoracic echocardiogram | 240
mobile echodensity on tricuspid valve | 240
beta-HCG fell to 60,862 mIU/mL | 240
transferred out of ICU | 288
platelet counts improved | variable
ANC improved | variable
cycle 2 induction chemotherapy | 384
repeat echocardiogram | variable
1.1 cm mobile echodensity on tricuspid valve | variable
therapeutic enoxaparin | variable
discharged home | 432
returned for cycle 1 day 1 EMA-CO | 720
etoposide 100 mg/m2 | 720
methotrexate 300 mg/m2 | 720
dactinomycin 0.5 mg | 720
cyclophosphamide 600 mg/m2 | 720
vincristine 1 mg/m2 | 720
beta-HCG normalized | 720
filgrastim marrow support | 720
3 additional cycles EMA-CO | variable
surveillance | variable
