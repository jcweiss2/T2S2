86 years old | 0
female | 0
Caucasian | 0
admitted to the Emergency Department | 0
acute respiratory distress | 0
discharged from the inpatient unit | -2
complicated urinary tract infection | -48
hypothyroid disorder | 0
mild dementia | 0
traumatic brain injury | 0
substernal chest pain | 0
shortness of breath | 0
blood pressure 105/74 mm Hg | 0
heart rate 132 | 0
respiratory rate 26 | 0
oral temperature 36.7 °C | 0
oxygen saturation 88% | 0
rapid heart rate | 0
bilateral crackles on auscultation of the lungs | 0
sinus tachycardia | 0
ST-segment depressions in the precordial leads V2 to V5 | 0
hypoxemia | 0
mild metabolic acidosis | 0
moderate pulmonary edema | 0
small pleural effusions bilaterally | 0
white blood cell count 26.89 × 10∗3/μL | 0
troponin I 0.38 ng/mL | 0
troponin I 64.50 ng/mL | 2
treatment for flash pulmonary edema | 0
non-invasive ventilation | 0
aspirin | 0
clopidogrel | 0
atorvastatin | 0
antibiotics | 0
furosemide | 0
nitroglycerin | 0
heparin | 0
admitted to the intensive care unit | 2
transthoracic echocardiography | 2
moderate mitral valve regurgitation | 2
mitral valve stenosis | 2
left heart catheterization | 4
large saddle embolism | 4
non-dominant circumflex coronary artery | 4
intensive medical management | 4
respiratory status deteriorated | 8
cardiopulmonary arrest | 12
death | 12
do-not-resuscitate | -24
do-not-intubate | -24