40 years old | 0
female | 0
high fever | -4320
DLBCL diagnosis | -1440
two R-CHOP treatments | -1440
fever persisted | -1440
rituximab | -1440
cyclophosphamide | -1440
doxorubicin | -1440
vincristine | -1440
prednisone | -1440
body temperature 37.8 ℃ | 0
blood pressure 162/104 mmHg | 0
pulse 147 bpm | 0
respiratory rate 28 breaths/min | 0
shortness of breath | 0
moist rales in both lungs | 0
white blood cell count 7.17 × 10^9/L | 0
red blood cell count 2.86 × 10^12/L | 0
haemoglobin 95 g/L | 0
platelet count 403 × 10^9/L | 0
CRP 277.6 mg/L | 0
bone marrow proliferation active | 0
granulocyte red cell proportion inverted | 0
lymphoid malignant tumour cells 22.5% | 0
CD20 (+) | 0
TDT (-) | 0
body temperature 36.5 °C | 24
oxygen saturation 91.3% | 24
white blood cell count 12.32 × 10^9/L | 24
lymphocyte classification 1.0% | 24
monocyte classification 1.0% | 24
neutrophil classification 97.0% | 24
CRP 79.0 mg/L | 24
chest CT multiple consolidation shadows | 0
chest CT plaques in both lungs | 0
pulmonary edema with inflammation | 0
chest CT consolidation disappeared slightly | 24
Pneumocystis in bronchoalveolar lavage fluid | 0
L. pneumophila in bronchoalveolar lavage fluid | 0
P. jirovecii verified | 0
Legionella culture | 96
isothermal chip amplification | 96
L. pneumophila culture positive | 96
imipenem | 0
tigecycline | 0
carprofen | 0
levofloxacin | 24
compound sulfamethoxazole | 24
endotracheal intubation ventilator | 0
septic shock | 720
B-ultrasound pancreas enlarged | 720
drug-induced pancreatitis | 720
death | 720
