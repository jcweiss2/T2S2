87 years old | 0
female | 0
non-insulin dependent diabetes mellitus | 0
chronic hypertension | 0
coronary artery disease | 0
gastro-oesophageal reflux disease | 0
osteoarthritis | 0
right total knee replacement | 0
cervical spine fixation | 0
severe symptomatic aortic stenosis | 0
TAVI | -216
fever | -90
convulsive seizure | -90
CT brain showed acute ischaemic stroke | -90
transferred to ICU | 0
blood cultures grew Corynebacterium | 0
transoesophageal echocardiogram confirmed post-TAVI infective endocarditis | 0
transferred to France | 8
underwent aortic root and valve replacement | 13
discharged from France | 33
admitted to ICU | 33
intubated for respiratory distress | 33
worsening hypoxaemia | 33
bilateral lower lobe opacities | 33
aspiration pneumonia | 33
normochromic normocytic anaemia | 0
normal leucocyte count | 0
thrombocytopenia | 0
elevated inflammatory markers | 0
low albumin value | 0
normal liver and renal function tests | 0
C-reactive protein 104 mg/L | 0
Corynebacterium species in blood cultures | 0
TTE negative for vegetations | 0
TOE showed large mobile vegetation | 1
aortic root pseudoaneurysm | 1
aortic root abscess | 1
CT angiography showed pseudoaneurysm | 2
multidisciplinary team discussion | 0
infective endocarditis diagnosis | 0
meropenem/levofloxacin and vancomycin treatment | 0
partial response in CRP | 6
febrile | 6
transferred to France for surgery | 8
aortic root and valve replacement with homograft | 13
Corynebacterium amycolatum in blood cultures | 13
post-operative course complicated by chylothorax and septic shock | 13
ventilator-associated pneumonia | 13
percutaneous tracheostomy | 13
transferred back to ICU | 33
Glasgow coma scale 6/15 | 33
lumbar puncture normal | 33
MRI head confirmed previous CT head findings | 33
cervical MRI showed degenerative disease | 33
EEG no seizures | 33
nerve conduction/electromyography showed axonal neuropathy | 33
critical illness polyneuropathy and myopathy | 33
Neurology team consultation | 33
intermittent changes in level of consciousness | 33
Rifampin and daptomycin treatment | 33
meropenem and daptomycin treatment | 33
percutaneous endoscopic gastrostomy | 33
optimized nutrition and physiotherapy | 33
improved and weaned off mechanical ventilation | 33
discharged home | 192
follow-up transthoracic echo showed mild aortic regurgitation | 192
preserved EF | 192
inflammatory markers normal | 192
CRP 4.64 mg/L | 192
afebrile and able to follow simple commands | 540