45 years old | 0
male | 0
received YF vaccine | 0
fever | 168
myalgia | 168
headache | 168
vomiting | 168
treated at emergency department | 168
discharged home | 168
antiemetics | 168
analgesics | 168
antibiotics | 168
ciprofloxacin | 168
metronidazole | 168
worsening of symptoms | 216
jaundice | 216
abdominal pain | 216
conjunctival suffusion | 216
altered mental status | 216
respiratory failure | 216
mechanical ventilation | 216
hemodynamic instability | 216
vasopressors | 216
transferred to ICU | 216
leukocytosis | 216
thrombocytopenia | 216
high levels of alanine aminotransferase | 216
high levels of aspartate aminotransferase | 216
high levels of total bilirubin | 216
high levels of creatinine | 216
high levels of creatine phosphokinase | 216
high prothrombin-time international normalized ratio | 216
antibiotic therapy | 216
ceftriaxone | 216
piperacillin-tazobactam | 216
steroids | 216
methylprednisolone | 216
hemoderivatives transfusion | 216
hemodialysis | 216
negative blood cultures | 216
negative serology for dengue fever | 216
negative serology for leptospirosis | 216
abdominal CT | 216
moderate free fluid in the abdominal cavity | 216
improvement in laboratorial parameters | 216
improvement in haemodynamic parameters | 216
no recovery of conscience | 216
suspension of sedative drugs | 216
CNS CT | 336
small frontal lobe bleeding | 336
electroencephalogram analysis | 336
severe diffuse brain dysfunction | 336
death | 480
necropsy | 480
macro and microgoticular steatosis | 480
hepatocytic necrosis | 480
multifocal lymphocyte perivascular encephalitis | 480
angioinvasive hyalohyphomycosis | 480
fungal embolism | 480
thrombosis of large and medium vessels | 480
fungal endomyocarditis | 480
cardiomyocyte necrosis | 480
fungal brain abscesses | 480
necrotizing encephalitis | 480
PCR-based nucleic acid detection | 480
Aspergillus spp. infection | 480
RT-PCR test for YF virus | 480
YF vaccine virus strain | 480
viscerotropic disease | 0
acute multiple organ system dysfunction | 0
YF vaccine associated-VTD | 0
immunocompetent patient | 0
IA | 216
liver failure | 216
immunoparalysis | 216
acute liver failure | 216
ALF | 216
immunodeficiency state | 216
pro-inflammatory cytokines | 216
monocyte and macrophage dysfunction | 216
hepatic macrophages | 216
local injury | 216
systemic inflammation | 216
immunosuppression | 216
innate and adaptative responses | 216
secondary infections | 216
systemic viral infection | 216
Th1 and Th2 imbalance | 216
CD4/CD8 inversion | 216
cytokine inflammatory cascade | 216
transient immunosuppression state | 216
high severity score | 216
concomitant pulmonary infection | 216
corticosteroid use | 216