38 years old | 0
male | 0
agammaglobulinaemia | 0
non-compliant with immunoglobulin administration | 0
dyspnoea | 0
productive cough | 0
fever | 0
tachycardic | 0
tachypnoeic | 0
febrile | 0
body temperature 38.7°C | 0
blood pressure 78/51 mmHg | 0
oxygen saturation 85% | 0
non-rebreather facial mask | 0
aggressive fluid resuscitation | 0
infiltrates in the left lower lobe | 0
mild left pleural effusion | 0
community-acquired pneumonia | 0
septic shock | 0
ceftriaxone | 0
clarithromycin | 0
haematocrit 38.5% | 0
haemoglobin 11.9 g/dL | 0
white cell count 9050 per μL | 0
neutrophils 88.9% | 0
lymphocytes 8.4% | 0
monocytes 2.0% | 0
eosinophils 0.5% | 0
basophils 0.1% | 0
platelet count 92000 per μL | 0
red cell count 5450000 per μL | 0
mean corpuscular volume 70.7 fL | 0
sodium 135 mmol/L | 0
potassium 4.2 mmol/L | 0
chloride 102 mmol/L | 0
carbon dioxide 20 mmol/L | 0
albumin 35 g/dL | 0
calcium 83 mg/L | 0
phosphorus 25 mg/L | 0
magnesium 12 mg/L | 0
alanine aminotransferase 39 UI/L | 0
aspartate aminotransferase 42 UI/L | 0
prothrombin time 15.8 | 0
international normalized ratio 1.48 | 0
thromboplastin time 40 | 0
lactic acid 2.1 mmol/L | 0
procalcitonin 0.33 ng/mL | 0
C-reactive protein 44.3 ng/mL | 0
B-type natriuretic peptide 136 pg/mL | 0
arterial oxygen pressure 65 mmHg | 0
persistent hypoxaemia | 0
worsening respiratory distress | 0
intensive care unit | 2
sedated | 2
intubated | 2
ventilated | 2
increasing left pleural effusion | 2
chest tube inserted | 2
drained fluid compatible with empyema | 2
norepinephrine | 2
haemodynamic stability | 4
urine output improving | 4
CT scan of the thorax | 48
homogeneous density with air bronchogram | 48
Gram stain of sputum revealed Gram-negative bacilli | 48
aerobic blood cultures grew Gram-negative coccobacilli | 48
A. calcoaceticus identified | 48
intravenous immunoglobulins | 24
C-reactive protein peaked | 48
procalcitonin peaked | 48
antibiotic regimen replaced | 48
colistin | 48
cefepime | 48
patient's condition improved | 72
intravenous pressors stopped | 72
weaned off mechanical ventilation | 72
extubated | 96
minimal left pleural effusion | 96
chest tube removed | 96
colistin and cefepime replaced with ciprofloxacin | 96
discharged | 336
ciprofloxacin 500 mg/day | 336
follow-ups | 672