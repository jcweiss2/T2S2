49 years old | 0
    leucodermal | 0
    presented to emergency department | 0
    non-specific malaise | 0
    feeling of postprandial infarction | 0
    colic-like abdominal pain | -1440
    bloodless diarrhoea | -1440
    asthenia | -720
    edema of lower limbs | -720
    edema of face | -720
    polydipsia | -720
    polyuria | -720
    cutaneous trunk hyperpigmentation | -720
    face hyperpigmentation | -720
    non-productive cough | 0
    no recent weight changes | 0
    hypertension | 0
    lisinopril | 0
    furosemide | 0
    tobacco history | 0
    36 pack-year consumption | 0
    slight alcohol habit | 0
    23 g alcohol/day | 0
    dyslipidaemia | 0
    hyperuricaemia | 0
    statin | 0
    colchicine | 0
    lived in Brazil | 0
    lived in Angola | 0
    lived in Guinea | 0
    mild melanoderma | 0
    apyrexia | 0
    conscious | 0
    temporally oriented | 0
    spatially oriented | 0
    weight 96.6 kg | 0
    height 192 cm | 0
    body mass index 26.2 kg/m² | 0
    cardiac auscultation no changes | 0
    pulmonary auscultation bilateral wheezing | 0
    pulmonary auscultation snoring | 0
    blood pressure 196/76 mmHg | 0
    symmetrical soft edema of lower limbs | 0
    no palpable adenopathies | 0
    severe metabolic alkalosis | 0
    hypokalaemia | 0
    moderate hypoxaemia | 0
    elevated serum ACTH | 0
    elevated urinary cortisol | 0
    chest x-ray bilateral pulmonary opacity | 0
    renal ultrasonographic examination normal | 0
    suprarenal ultrasonographic examination normal | 0
    admitted to Endocrinology Department | 0
    diagnostic hypotheses Cushing’s syndrome | 0
    diagnostic hypotheses ectopic ACTH production | 0
    progression of acute respiratory failure | 24
    admitted to ICU | 24
    diagnosis community-acquired pneumonia | 24
    invasive mechanical ventilation | 24
    empirical medication ceftriaxone | 24
    empirical medication azithromycin | 24
    negative Legionella pneumophila urinary antigen | 24
    negative Streptococcus pneumoniae urinary antigen | 24
    negative multiple PCR tests for gastroenteritis | 24
    swollen duodenal folds | 0
    biopsy of duodenal folds | 0
    inflammatory lamina propria infiltrate with eosinophils | 0
    presence of larvae | 0
    presence of eggs | 0
    Strongyloides stercoralis | 0
    ultrasound-guided liver biopsy | 0
    metastasis of small cell neuroendocrine carcinoma | 0
    immunohistochemical profile suggesting pulmonary origin | 0
    treated with ivermectin | 24
    haemodynamic support | 24
    ventilatory support | 24
    etomidate therapy | 24
    metyrapone therapy | 24
    tracheostomy | 528
    transferred to Pulmonology Department | 840
    died | 1080
    laboratory controls 2 months earlier | -1440
    eosinophilia 8.4% | -1440
    laboratory controls 2 years earlier | -17520
    eosinophilia 7.2% | -17520
    eosinophils 0.4% | 0
    lived in endemic areas | 0
    persistent infection over 10 years | 0
    self-infection phenomenon | 0
    reduced immune capacity | 0
    cerebral intraparenchymal haemorrhage | 0
    diffuse metastasis of carcinoma | 0
    primary lesion in pancreas head | 0
    negative parasitological stool tests | 0
    multiorgan infection | 0
    immunocompromised patient | 0
    appropriate clinical context | 0
    appropriate epidemiological context | 0
    