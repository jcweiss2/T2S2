66 years old | 0
female | 0
admitted to the emergency department | 0
general weakness | -168
poor oral intake | -168
diabetes | -87600
hypertension | -87600
metformin | -87600
glimepiride | -87600
hydrochlorothiazide | -87600
losartan | -87600
atorvastatin | -87600
severe osteoarthritis | -87600
multiple steroid injections | -87600
urinary tract infection | -336
Escherichia coli | -336
ceftriaxone | -336
tazobactam | -336
not on antihypertensive medication | -336
height 152 cm | 0
body weight 57 kg | 0
blood pressure 70/50 mmHg | 0
heart rate 70 beats per minute | 0
respiratory rate 20 per minute | 0
body temperature 36.5°C | 0
decreased skin turgor | 0
decreased tongue turgor | 0
unremarkable pulmonary exam | 0
unremarkable cardiac exam | 0
unremarkable abdominal exam | 0
unremarkable neurologic exam | 0
normal serum creatinine | -336
normal calcium | -336
decreased serum magnesium | 0
fractional excretion of sodium 1.0% | 0
pyuria | 0
hypotension | 0
UTI sepsis diagnosis | 0
admitted to intensive care unit | 0
antibiotics | 0
massive hydration | 0
vital signs stabilized | 48
inflammatory signs normalized | 48
blood pressure normalized | 48
elevated serum calcium | 0
elevated creatinine | 0
poor oral intake persisted | 48
general weakness persisted | 48
saline administration | 72
calcitonin administration | 72
serum calcium decreased | 96
serum calcium increased | 168
contrast-enhanced computed tomography | 168
whole body bone scintigraphy | 168
no evidence of malignancy | 168
negative serum protein electrophoresis | 168
negative urine protein electrophoresis | 168
negative anti-neutrophil cytoplasmic antibody titers | 168
negative tumor marker studies | 168
normal thyroid stimulating hormone | 168
normal free thyroxine | 168
osteopenia | 168
suppressed PTH | 168
undetectable PTH-related peptide | 168
low 25-hydroxy vitamin D | 168
multiple steroid injections history | 168
serum cortisol 2.36 μg/dL | 168
serum ACTH 32.51 pg/mL | 168
inadequate cortisol response | 168
secondary adrenal insufficiency diagnosis | 168
hydrocortisone administration | 240
serum calcium normalized | 312
general weakness improved | 312
anorexia improved | 312
magnesium trended normal | 312
serum calcium maintained | 480
osteoporosis risk | 480
corticosteroid replacement | 480
regular bone mineral density monitoring | 480
lost to follow-up | 480
