32 years old | 0
female | 0
pain in the mid-dorsal region | -672
progressive worsening | -672
weakness in the lower limbs | -24
expansive lesion in the eighth thoracic vertebra | -24
local kyphosis | -24
imminent instability | -24
computed tomography scan | -24
magnetic resonance imaging | -24
involvement of the medullary canal | -24
percutaneous CT-guided core-needle biopsy | -24
diagnosis of giant-cell tumor | -24
total en bloc spondylectomy | 0
posterior-only approach | 0
anterior-column reconstruction | 0
titanium mesh | 0
structural allograft | 0
pedicle screw instrumentation | 0
eighth dorsal nerve routes sacrificed | 0
surgery completed | 5
uneventful surgery | 5
no neurologic deficits | 5
pulmonary rehabilitation protocol | 48
progressive dyspnea | 72
impaired gas exchange | 72
bilateral hemothorax | 72
bilateral thoracentesis | 72
recovery from symptoms | 72
worsening of general status | 456
fever | 456
dyspnea | 456
decreased gas exchange | 456
increase in inflammatory markers | 456
moderate fluid collection in both lungs | 456
empyema | 456
septic state | 456
transfer to intensive care unit | 456
surgical debridement | 504
infected tissues removed | 504
allograft and titanium mesh extracted | 504
iliac crest tricortical autograft | 504
anterior support | 504
posterior pedicle instrumentation kept | 504
drains placed | 504
Enterobacter aerogenes identified | 504
pathogen-directed antibiotic therapy | 504
lower respiratory tract infection | 528
Acinetobacter baumannii identified | 528
septated empyema | 544
anterior and posterior approach | 544
complete drainage | 544
subcutaneous abscess | 560
methicillin-resistant Staphylococcus aureus identified | 560
Pseudomonas aeruginosa identified | 560
posterior open drainage | 560
progressive improvement | 672
discharge from hospital | 1872
custom-molded thoracolumbar brace | 1872
physical therapy | 1872
stable and asymptomatic | 6480
no evidence of infection or tumor relapse | 6480
follow-up imaging studies | 6480
no bone graft resorption | 6480
no instrumentation failure | 6480