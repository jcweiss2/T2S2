30 years old | 0
male | 0
admitted to the emergency department | 0
idiopathic bronchiectasis | -8760
fever | -24
productive cough | -24
chest pain | -24
dyspnea | -24
anosmia | -24
contact with COVID-19 patient | -24
nasopharyngeal swabs | 0
bilateral crackles | 0
SpO2 65% | 0
high flow nasal cannula | 0
FiO2 60% | 0
SpO2 82% | 0
peripheral infiltrates | 0
intubated | 2
mechanical ventilation | 2
COVID-19 confirmed | 2
leukocytosis | 2
lymphocytopenia | 2
increased D-dimer | 2
increased C-reactive protein | 2
increased lactate dehydrogenase | 2
increased ferritin | 2
contrast chest CT scans | 2
pulmonary embolism excluded | 2
bilateral ground-glass opacities | 2
bronchiectasis | 2
empiric therapy for COVID-19 | 2
ribavirin | 2
ceftriaxone | 2
azithromycin | 2
prophylactic anticoagulation | 2
ARDS-net | 2
prone position ventilation | 2
supportive ICU care | 2
Bordetella bronchiseptica | 72
doxycycline | 72
vitamin D deficiency | 72
vitamin D3 supplementation | 72
extubated | 360
RT-PCR for COVID-19 negative | 432
microbiology negative | 432
discharged | 480
monitor pet dog | 480
review vitamin D supplementation | 480