78 years old | 0
male | 0
admitted to physician's office | 0
leg edema | -24
ruptured abdominal aortic aneurysm | -8760
smoking | -14400
widowed | 0
retired public school employee | 0
new onset AF | 0
discharged home | 24
warfarin | 24
digoxin | 24
diuretic therapy | 24
shortness of breath | 24
nonproductive cough | -168
malaise | -504
fatigue | -504
weakness | -504
no fever | 24
no chills | 24
no sweats | 24
temperature 36.8oC | 24
pulse 132/minute | 24
blood pressure 105/56 mmHg | 24
respirations 28/minute | 24
jugular venous distension | 24
irregularly irregular pulse | 24
left-sided rhonchi | 24
bibasilar pulmonary crackles | 24
left lower pulmonary infiltrate | 24
left pleural effusion | 24
cardiomegaly | 24
AF | 24
no ischemic changes | 24
dopamine | 24
diltiazem therapy | 24
intravenous furosemide | 24
intravenous heparin | 24
intubated | 24
transferred to referral hospital | 24
unresponsive | 48
cold mottled skin | 48
temperature 36.6oC | 48
heart rate 108/minute | 48
respiratory rate 15/minute | 48
BP 88/47 mmHg | 48
bilateral pulmonary crackles | 48
irregular rhythm | 48
no murmurs | 48
no gallops | 48
mild edema | 48
no pulses palpable | 48
pH 7.26 | 48
pCO2 26 mm Hg | 48
pO2 299 mm Hg | 48
lactate 6.9 mEq/L | 48
glucose 65 mg/dL | 48
creatinine 7.1 mg/dL | 48
dobutamine | 48
gentamicin | 48
ticarcillin/clavulanate | 48
central venous pressure 7 mm Hg | 48
pulmonary artery pressure 32/21 mm Hg | 48
pulmonary artery wedge pressure 19 mm Hg | 48
moderately decreased left ventricular function | 48
unremarkable cardiac valves | 48
hypotensive | 72
multi-organ failure | 72
died | 72
Streptococcus pneumoniae | 72
near-lobar early organizing pneumonia | 72
empyema | 72
severe coronary and systemic atherosclerosis | 72
near-total old occlusion | 72
old myocardial infarctions | 72
mild stenosis | 72
severe atherosclerosis | 72
heart failure | 24
pneumonia | -168
septic shock | 48
cough | -168
leg edema | -24