61 years old|0
    white woman|0
    Ashkenazi Jewish descent|0
    nausea|-192
    vomiting|-192
    fever|-192
    severe pitting edema in both legs|0
    ascites|0
    splenomegaly|0
    palpable axillary lymph nodes|0
    bilateral pleural effusion|0
    retroperitoneal lymph node enlargement|0
    mild anemia|0
    thrombocytopenia|0
    hypoalbuminemia|0
    elevated C-reactive protein|0
    elevated alkaline phosphatase|0
    elevated gamma-glutamyltranspeptidase|0
    negative HIV serology|0
    negative HTLV-1 virus serology|0
    negative HHV-8 PCR|0
    positive anti-citrullinated protein antibody|0
    normal complement levels|0
    no hypergammaglobulinemia|0
    no monoclonal immunoglobulin|0
    elevated interleukin-6|0
    lymphoid hyperplasia|0
    hyalinization of the germinal center|0
    increased scattered plasma cells|0
    increased number of megakaryocytes with dysplastic features|0
    grade 1 fibrosis|0
    negative JAK2V617F mutation|0
    negative CALR exon 9 mutation|0
    diploid karyotype|0
    renal thrombotic microangiopathy|0
    mesangial expansion|0
    duplication of the glomerular capillary basal membrane|0
    increased fluorodeoxyglucose uptake|0
    worsening of anasarca|168
    worsening renal function|168
    multiple organ failure|168
    mechanical ventilation|168
    vasopressor medications|168
    continuous renal replacement therapy|168
    TAFRO syndrome diagnosis|432
    hemoglobin 8.3|432
    white blood cell count 17.11|432
    platelets 21|432
    alkaline phosphatase 205|432
    gamma-glutamyltranspeptidase 210|432
    creatinine 2.14|432
    C-reactive protein 231.2|432
    interleukin-6 722.6|432
    pulse steroids|432
    tocilizumab|432
    rituximab|432
    improvement in respiratory status|600
    improvement in hemodynamic status|600
    weaned from ventilator support|600
    discontinued vasopressor medications|600
    switched to intermittent hemodialysis|936
    discharged from ICU|1104
    discharged from hospital|2160
    complete resolution of anasarca|2160
    complete resolution of organomegaly|2160
    normalization of hemoglobin|2160
    normalization of platelet counts|2160
    decreasing interleukin-6 levels|2160
    outpatient treatment|2160
    tocilizumab every 3 weeks|2160
    tapered steroids|2160
    PET-CT reduction in lymph node size|720
    resolution of pleural effusion|720
    <|eot_id|>
    61 years old|0
    white woman|0
    Ashkenazi Jewish descent|0
    nausea|-192
    vomiting|-192
    fever|-192
    severe pitting edema in both legs|0
    ascites|0
    splenomegaly|0
    palpable axillary lymph nodes|0
    bilateral pleural effusion|0
    retroperitoneal lymph node enlargement|0
    mild anemia|0
    thrombocytopenia|0
    hypoalbuminemia|0
    elevated C-reactive protein|0
    elevated alkaline phosphatase|0
    elevated gamma-glutamyltranspeptidase|0
    negative HIV serology|0
    negative HTLV-1 virus serology|0
    negative HHV-8 PCR|0
    positive anti-citrullinated protein antibody|0
    normal complement levels|0
    no hypergammaglobulinemia|0
    no monoclonal immunoglobulin|0
    elevated interleukin-6|0
    lymphoid hyperplasia|0
    hyalinization of the germinal center|0
    increased scattered plasma cells|0
    increased number of megakaryocytes with dysplastic features|0
    grade 1 fibrosis|0
    negative JAK2V617F mutation|0
    negative CALR exon 9 mutation|0
    diploid karyotype|0
    renal thrombotic microangiopathy|0
    mesangial expansion|0
    duplication of the glomerular capillary basal membrane|0
    increased fluorodeoxyglucose uptake|0
    worsening of anasarca|168
    worsening renal function|168
    multiple organ failure|168
    mechanical ventilation|168
    vasopressor medications|168
    continuous renal replacement therapy|168
    TAFRO syndrome diagnosis|432
    hemoglobin 8.3|432
    white blood cell count 17.11|432
    platelets 21|432
    alkaline phosphatase 205|432
    gamma-glutamyltranspeptidase 210|432
    creatinine 2.14|432
    C-reactive protein 231.2|432
    interleukin-6 722.6|432
    pulse steroids|432
    tocilizumab|432
    rituximab|432
    improvement in respiratory status|600
    improvement in hemodynamic status|600
    weaned from ventilator support|600
    discontinued vasopressor medications|600
    switched to intermittent hemodialysis|936
    discharged from ICU|1104
    discharged from hospital|2160
    complete resolution of anasarca|2160
    complete resolution of organomegaly|2160
    normalization of hemoglobin|2160
    normalization of platelet counts|2160
    decreasing interleukin-6 levels|2160
    outpatient treatment|2160
    tocilizumab every 3 weeks|2160
    tapered steroids|2160
    PET-CT reduction in lymph node size|720
    resolution of pleural effusion|720