57 years old | 0
male | 0
hyperlipidemia | -672
chronic tobacco use | -672
bilateral foot pain | -24
blue discoloration | -24
coolness | -24
fever | -48
fatigue | -48
abdominal discomfort | -48
nonbloody diarrhea | -48
loss of appetite | -48
dog bite | -168
vaccinated for SARS-CoV-2 | 0
asymptomatic for SARS-CoV-2 | 0
admitted to the hospital | 0
afebrile | 0
blood pressure 93/54 mm Hg | 0
heart rate 85 beats/min | 0
respiration 16 breaths/min | 0
saturation 98% on ambient air | 0
regular heart rhythm | 0
no jugular venous distention | 0
clear breath sounds | 0
small left finger lesion | 0
surrounding erythema | 0
discoloration | 0
lower extremities slightly cyanotic | 0
palpable pulses | 0
extremely sensitive to touch | 0
white blood cell count 18.8 × 10^3/µL | 0
neutrophilic bands of 40.8% | 0
hemoglobin 17.1 gm/dL | 0
platelets 72 × 10^3/µL | 0
ESR 28 mm/hr | 0
CRP 42 mg/dL | 0
sodium 130 mmol/L | 0
carbon dioxide 21 mmol/L | 0
blood urea nitrogen 47 mg/dL | 0
creatinine 3.41 mg/dL | 0
aspartate transaminase 502 IU/L | 0
alanine transaminase 257 IU/L | 0
alkaline phosphatase 136 IU/L | 0
NT-Pro-B Natriuretic peptide 5846 pg/mL | 0
troponin 26.2 ng/dL | 0
creatine kinase 1246 IU/L | 0
PT 12.4 seconds | 0
INR 1.08 | 0
PTT 43 seconds | 0
fibrinogen 380 mg/dL | 0
D-dimer greater than 128 mg/dL | 0
SARS-CoV-2 PCR test negative | 0
urinalysis negative for infection | 0
blood culture positive for gram-negative rods | 0
ECG showed ST-segment elevation | 0
chest discomfort | 20
emergent cardiac catheterization | 20
diffuse mild luminal irregularities | 20
no focal stenosis or occlusion | 20
left ventricular end-diastolic pressure elevated | 20
TTE showed LVEF of 30% | 24
diffuse hypokinesis | 24
grade I diastolic dysfunction | 24
supportive on low-dose norepinephrine | 24
computed tomography of chest and abdomen | 24
bilateral peripheral septal thickening of the lungs | 24
no evidence of pulmonary emboli or lymphadenopathy | 24
magnetic resonance imaging of the brain | 24
small acute punctate infarct of the left parietal lobe | 24
bilateral lower extremity arterial Doppler and ankle/brachial indices | 24
no evidence of stenosis or occlusion | 24
IV methylprednisolone | 24
heparin infusion | 24
cefepime | 24
doxycycline | 24
gabapentin | 24
morphine | 24
autoimmune panel negative | 48
stool cultures negative | 48
serology for syphilis, Lyme, diphtheria, viral hepatitis, and parvovirus negative | 48
IgG for mycoplasma pneumoniae positive | 48
Epstein-Barr Virus capsid and nuclear antigen positive | 48
toxoplasma positive | 48
coxsackievirus positive | 48
influenza A and B positive | 48
troponin peaked at 119 ng/mL | 13
ECG showed worsening ST elevation | 13
renal function recovered | 48
platelet count fell to nadir of 28 × 10^3/µL | 48
evaluated for probable diagnosis of HIT, ITP, HUS, and TTP | 48
developed bluish discoloration to the skin of the toes | 48
treated with IVIG and argatroban | 48
platelet count recovery | 120
repeat TTE showed improved LVEF of 45% | 120
repeat ECG showed normalized ST-segments | 120
incomplete right bundle branch block | 120
discharged | 144