69 years old | 0
severe sepsis | 0
pulseless electrical activity cardiac arrest | 0
cardiopulmonary resuscitation | 0
return of spontaneous circulation | 0
hypotension | 0
tachycardia | 0
fluid boluses | 0
metaraminol boluses | 0
tracheal intubation | 0
mechanical ventilation | 0
severe metabolic acidosis | 0
treatment as per surviving sepsis guidelines | 0
central venous catheter insertion | 0
MAP >70 mmHg | 0
fluid resuscitation | 0
norepinephrine infusion | 0
sustained oliguria | 0
systemic acidosis | 0
CVVH initiation | 0
double lumen hemofiltration catheter insertion | 0
chest radiograph showing catheter tips adjacent | 0
CVVH caused precipitous hypotension | 0
PEA arrest | 0
spontaneous circulation restored | 0
epinephrine bolus | 0
CPR | 0
CVVH recommenced | 0.5
fluid boluses | 0.5
epinephrine boluses | 0.5
norepinephrine infusion increase | 0.5
systolic blood pressure >90 mmHg | 0.5
blood pressure fluctuations | 0.5
CVVH stopped | 0.75
norepinephrine requirement reduced | 0.75
hemodynamic stability restored | 0.75
hemofiltration catheter withdrawal | 0.75
repeat chest radiograph | 0.75
CVVH resumed | 0.75
little hemodynamic instability | 0.75
no significant vasopressor increase | 0.75
anaphylaxis | 0
human and technical errors | 0
hypotension attributed to CVVH | 0
hypovolemia | 0
electrolyte disturbances | 0
vasodilatation | 0
tension pneumothorax | 0
thromboembolism | 0
toxins | 0
cardiac tamponade | 0
critical incident reporting | 0
morbidity and mortality meetings | 0
two person checking | 0
labeling of syringes | 0
prefilled syringes | 0
bar codes | 0
guidelines and protocols | 0
alarm settings | 0
