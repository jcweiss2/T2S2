45 years old | 0
male | 0
low backache | -168
weakness of both lower limbs | -168
urinary retention | -48
constipation | -48
full power in the upper limb | 0
Grade 3 power in the lower limbs | 0
thickened ligamentum flavum | 0
cord oedema | 0
distended abdomen | 0
soft abdomen | 0
no clinical evidence of ascites or organomegaly | 0
bowel sounds present | 0
urinary bladder catheterized | 0
normal pre-operative investigations | 0
admitted for laminectomy and decompression of the spine | 0
induction of anaesthesia | 0
invasive blood pressure monitoring | 0
arterial blood gas monitoring | 0
propofol 140 mg | 0
fentanyl citrate 150 μg | 0
rocuronium bromide 50 mg | 0
trachea intubated | 0
mechanical prophylaxis for deep vein thrombosis | 0
warm air blanket | 0
normal post-induction ABG readings | 0
sevoflurane in 50% O2 in air | 0
propofol infusion at 25 μg/kg/min | 0
vecuronium bromide at 2 mg/h | 0
surgery lasted 5 h | 5
intermittent fentanyl | 0
hydration with IV 3.5 L 0.9% saline | 0
hydration with IV 0.5 L colloid | 0
noradrenaline at 2-4 μg/min | 0
blood loss 250 ml | 0
urine output 250 ml | 0
metabolic acidosis | 2
severe canal stenosis | 2
cord oedema | 2
methylprednisolone started | 2
inadequate motor power | 5
inadequate respiratory effort | 5
repeat ABG showed metabolic acidosis | 5
blood sugar 246 mg% | 5
urine ketone negative | 5
insulin infusion started | 5
shifted to intensive care unit | 5
central venous line inserted | 5
central venous pressure 1-2 cm H2O | 5
overnight fluid therapy | 5
resolved acidosis | 24
resolved oliguria | 24
extubated | 24
kidney function test revealed high normal values | 24
normal serum sodium | 24
normal serum potassium | 24
normal thyroid status | 24
upper limb power almost normal | 24
power in both lower limbs 1/5 | 24
methylprednisolone continued | 24
tense abdominal distension | 30
respiratory distress | 30
respiratory alkalosis | 30
reintubated | 30
ventilated | 30
normal chest X-ray | 30
normal echocardiogram | 30
colonic gaseous distension | 30
Ryle's tube inserted | 30
injection neostigmine started | 30
deranged kidney function test | 48
high-grade fever | 48
blood cultures sent | 48
urine cultures sent | 48
tracheal aspirate sent | 48
antibiotics upgraded | 48
sepsis | 48
pancreatitis profile | 48
serum procalcitonin 4.4 ng/ml | 48
hypocalcaemia | 48
hypoalbuminemia | 48
normal serum amylase | 48
normal serum lipase | 48
factitious hypocalcaemia ruled out | 48
hyperphosphatemia | 48
low parathormones | 48
normal magnesium levels | 48
IV albumin started | 48
refractory hypocalcaemia | 48
high doses of IV calcium | 48
oral calcitriol started | 48
renal functions started to resolve | 72
acidosis started to resolve | 72
abdominal symptoms persisted | 72
digital examination ruled out faecal impaction | 72
decompressive sigmoidoscopy performed | 72
total parenteral nutrition started | 72
gastrointestinal symptoms decreased | 96
procalcitonin decreased | 96
total leucocyte count decreased | 96
serum calcium increased | 96
extubated | 216
reintubated | 234
ventilated | 234
severe tachypnoea | 234
decreased consciousness | 234
pulmonary embolism ruled out | 234
MRI spine did not reveal fresh changes | 234
cerebrospinal fluid analysis ruled out meningitis | 234
tracheostomised | 312
steady improvement | 312
weaned off ventilator | 312
fully conscious | 312
good power in all limbs | 312
normal calcium levels | 312
normal albumin levels | 312
no gastrointestinal symptoms | 312
decannulated | 312
discharged | 312