55 years old | 0
male | 0
admitted to the hospital | 0
multiple myeloma | 0
previous stem cell transplant | 0
recurrence of disease | 0
relapsed multiple myeloma | 0
treatment with carfilzomib | -72
intermittent fevers | -48
dyspnea | -72
productive cough | -72
febrile | 0
tachypneic | 0
tachycardic | 0
decreased breath sounds in right lung base | 0
no rales | 0
no wheezing | 0
pancytopenia | 0
white blood cell count 1.2 × 10^9/l | 0
hemoglobin 53 g/l | 0
platelets 4.0 × 10^9/l | 0
treated with cefepime | 0
treated with azithromycin | 0
continued home medications | 0
acyclovir | 0
allopurinol | 0
fluconazole | 0
pantoprazole | 0
new-onset hypoxia | 0
hypotension | 0
altered mental status | 0
transferred to medical intensive care unit | 0
lactic acid 6.1 mMol/l | 0
arterial blood gas pH 7.40 | 0
arterial blood gas PaCO2 3.3 kPa | 0
arterial blood gas PaO2 11.3 kPa | 0
measured O2sat 94% | 0
intubation | 0
treated with topical endobronchial lidocaine | 0
treated with etomidate | 0
treated with succinylcholine | 0
hypoxia worsened | 24
arterial blood gas pH 7.21 | 24
arterial blood gas PaCO2 3.3 kPa | 24
arterial blood gas PaO2 55.1 kPa | 24
measured O2sat 49% | 24
brownish arterial blood | 24
co-oximetry requested | 24
methemoglobin level 53% | 24
treated with methylthioninium chloride | 24
arterial blood gas methemoglobin 12% | 24.5
arterial blood gas methemoglobin 9% | 25
O2sat >90% | 25
bright red arterial blood | 25
septic shock | 0
bacteremia with Rothia mucilaginosa | 0
succumbed to septic shock | 0
