18 years old | 0
male | 0
sports-related injury to the left shoulder | -936
over a dozen surgical revisions | -936
recurrent and prolonged shoulder infections | -936
Pseudomonas aeruginosa | -936
Sphingomonas paucimobilis | -936
Candida colliculosa | -936
Staphylococcus aureus | -936
left shoulder tendon release and revision | -312
CRPS | -312
severe pain | -312
allodynia | -312
edema | -312
muscle spasms | -312
temperature changes | -312
electromyography (EMG) evaluation | -312
brachial plexus injury | -312
asthma | -312
selective IgG3 deficiency | -312
oral medical management | -312
opioids | -312
antidepressants | -312
antispasmodics | -312
left stellate ganglion blockade | -312
significant symptom relief | -312
continuous cervical epidural infusions | -312
left C6–C7 interlaminar epidural catheter | 0
fluoroscopic guidance | 0
preprocedure labs | 0
complete blood count | 0
complete metabolic panel | 0
creatinine phosphokinase | 0
intravenous vancomycin | -1
placement of the catheter | -1
intrathecal and intravascular placement | -1
1% lidocaine with 1:200,000 epinephrine | -1
epidural infusion of 0.25% bupivacaine with hydromorphone 10 mcg per mL and clonidine 1 mcg per mL | -1
methadone 10 mg twice a day | -1
hydromorphone 4 to 8 mg as needed | -1
diazepam 10 mg 4 times a day | -1
baclofen 20 mg 4 times a day | -1
amitriptyline 100 mg once a day | -1
decrease in pain from 9/10 to 7/10 on the VAS | -1
less muscle spasms | -1
continuous infusion increased to 6 mL per hour | -48
demand dose of 2 mL every 15 minutes | -48
improved sleep | -48
further decrease in LUE spasms and edema | -48
VAS of 5/10 | -48
febrile to 38.1°C | -72
progressive headache | -72
neck pain | -72
increase in temperature to 40.0°C | -72
neurological examination remained unchanged | -72
epidural site was nontender to palpation | -72
blood and urine cultures were sent | -72
chest x-ray was negative | -72
laboratory workup was notable for an increase in white count | -72
cefepime was added empirically to vancomycin | -72
abatement of fever | -72
decrease in white count to 5.9×10^3/μL | -72
MRI of the cervical spine | -72
epidural collection from the inferior margin of C3 to T1 | -72
compressing the left C5 and C6 nerve roots | -72
considerable interstitial edema in the left paraspinal muscles | -72
transfer to the neurosciences intensive care unit (NSICU) | -72
hourly neurological examination | -72
intractable nausea and vomiting | -48
left arm weakness | -48
emergent decompression and evacuation | -48
C3 to C7 cervical laminectomies and C4–C5 and C5–C6 left foraminotomies | -48
intraoperative cultures of the cervical abscess were positive for P aeruginosa | -48
intraoperative cultures of the cervical abscess were susceptible to cefepime | -48
urine and blood cultures from hospital day 6 were negative | -48
vancomycin was stopped | -48
cefepime was continued | -48
resolution of arm weakness | -48
uneventful postoperative course | -48
discharged home on postoperative day 3 | -48
intravenous cefepime for a total of 6 weeks | -48