84 years old | 0
female | 0
Caucasian | 0
height 165 cm | 0
weight 45 kg | 0
admitted to the emergency department | 0
generalized abdominal pain | 0
vomiting | 0
diarrhea | 0
altered general status | 0
respiratory distress | 0
tachypneic | 0
accessory muscles used | 0
febrile | 0
tachycardic | 0
desaturation | 0
hypotensive | 0
arterial blood gases taken | 0
primary metabolic acidosis | 0
anion gap 23 | 0
oxygen saturation increased to 95% | 0
hydration with normal saline | 0
systolic blood pressure increased to 120 mmHg | 0
right upper quadrant tenderness | 0
positive Murphy’s sign | 0
blood cultures taken | 0
urine cultures taken | 0
given Amikacin | 0
given Vancomycin | 0
started on intravenous Tazocin | 0
COVID-19 PCR test taken | 0
negative COVID-19 PCR | 0
inflammatory markers elevated | 0
C-reactive protein 50 | 0
lactate dehydrogenase 240 | 0
ferritin 271.6 | 0
fibrinogen 1017.15 | 0
erythrocyte sedimentation rate 86 | 0
lymphopenic | 0
absolute lymphocytic count 357 | 0
elevated amylase | 0
elevated bilirubin | 0
normal aspartate aminotransferase | 0
normal alanine aminotransferase | 0
CT chest-abdomen-pelvis done | 0
extensive patchy consolidations | 0
air bronchograms | 0
ground glass opacities | 0
COVID-19 pneumonia | 0
gallbladder markedly distended | 0
transverse diameter 4.6 cm | 0
enhancing wall with focal defects | 0
partial necrosis | 0
fat stranding | 0
peri-vesicular fluid | 0
pericholecystic abscesses | 0
acute ischemic gangrenous cholecystitis | 0
scheduled for percutaneous drainage | 0
repeat COVID-19 PCR taken | 0
became hypotensive again | 24
refractory to IV fluids | 24
Dopamine started | 24
systolic blood pressure elevated | 24
deteriorated again | 48
hypotensive | 48
desaturated | 48
double oxygen source used | 48
intubated | 48
cardio-pulmonary arrest | 48
resuscitation failed | 48
pronounced dead | 48
repeat PCR for COVID-19 positive | 48
blood cultures negative | 48
urine culture negative | 48