male | 0
neonate | 0
delivered spontaneously | 0
full term | 0
birth weight 4.098kg | 0
head circumference 35 cm | 0
poor feeding | -72
decreased tone | -72
reflexes noted on exam | -72
admitted to neonatal intensive care unit | -72
sepsis workup | -72
cranial ultrasonography | -72
small right-sided choroid plexus cyst | -72
partial agenesis of corpus collosum | -72
spontaneous myoclonic jerks | -72
stimulus-provoked myoclonic jerks | -72
intermittent hiccups | -72
progressively lethargic | -72
unresponsive | -72
central hypotonia | -72
amino acid analysis of CSF and plasma | -96
liver studies | -96
ammonia level | -96
septic workup negative | -96
bedside electroencephalographic monitoring | -96
abnormal electroencephalographic monitoring | -96
diffuse cortical dysfunction | -96
partial seizures | -96
progressive encephalopathy | -96
respiratory insufficiency | -96
mechanical ventilation | -96
MR imaging of brain | -96
1H-MR spectroscopy | -96
elevated glycine peak | -96
glycine concentration 11.8 mmol | -96
choline concentration 2.47 mmol | -96
creatine concentration 7.66 mmol | -96
N-acetylaspartate concentration 5.74 mmol | -96
lactate concentration 2.45 mmol | -96
elevated lactate peak | -96
CSF glycine level 342 μmol/mL | -120
plasma glycine level 1419 μmol/mL | -120
CS- to-plasma glycine concentration ratio 0.24 | -120
urine organic acid analysis negative | -120
treated with dextromethorphan | -120
treated with phenobarbital | -120
treated with sodium benzoate | -120
level of consciousness improved | 120
extubated from mechanical ventilation | 168
follow-up weekly amino acid analysis | 168
decreased plasma glycine concentrations | 168
periodic elevations | 168
DNA testing | 168
homozygous missense mutation | 168
GLDC gene mutation | 168
glycine-restricted diet | 168
feeding problems | 720
poor growth | 720
recurrent vomiting | 720
seizures | 720