83 years old | 0
male | 0
type 2 diabetes | 0
hypertension | 0
atrial fibrillation | 0
myocardial infarction | 0
admitted to ICU | 0
secondary laparotomic surgery | -48
complications from primary low anterior resection | -48
gas and fecal leakage | -48
perforations in colon transversus closed | -48
sacral abscess evacuated | -48
aspirated during intubation | -48
sedation | -48
hemodynamically stable | -48
respiratory stable | -48
baseline sublingual microcirculatory measurement | 0
cardiac arrest | 12
hypoxia | 12
atelectasis of right lung | 12
cardiopulmonary resuscitation | 12
nor-adrenaline administration | 12
adrenaline administration | 12
vasoactive-inotropic score 99 | 12
systemic hemodynamic variables stabilized | 12
rising serum lactate | 12
declining renal function | 12
urine output 17 mL/24 h | 12
sepsis diagnosis | 12
CRRT with CytoSorb hemoadsorber | 12
microcirculatory measurement | 24
microcirculatory measurement | 36
microcirculatory measurement | 48
microcirculatory measurement | 120
hemoadsorber replacement | 24
lactate levels decreased | 24
VIS decreased | 24
TVD increased | 24
microcirculatory flow index normalized | 24
plugged vessels resolved | 36
brisk flow | 36
improved clinical condition | 36
fluid ultrafiltration initiated | 48
aggressive fluid resuscitation | 48
decline in TVD | 48
blood transfusion | 48
ultrafiltration | 48
improved diffusive capacity | 120
regained consciousness | 168
returned to surgery ward | 456
discharged to nursing facility | 1416
normalized renal function | 1416