85 years old| 0
    male | 0
    admitted to the hospital | 0
    fall at home | -24
    worsening lethargy | -168
    productive cough | -168
    decreased oral intake | -168
    transfusion-dependent chronic myelomonocytic leukaemia type 1 | 0
    type II diabetes mellitus | 0
    atrial fibrillation | 0
    permanent pacemaker | 0
    chronic kidney disease stage III | 0
    hypertension | 0
    permanent suprapubic catheter | 0
    neurogenic bladder | 0
    benign prostatic hypertrophy | 0
    restless leg syndrome | 0
    duodenal ulcers | 0
    hypercholesterolaemia | 0
    renal calculi | 0
    pyelonephritis | 0
    infective endocarditis of the aortic valve | 0
    non-ST elevation myocardial infarction | 0
    polymyalgic rheumatoid arthritis | 0
    chronic obstructive pulmonary disease | 0
    low-grade fever | 0
    blood pressure 131/47 mm Hg | 0
    heart rate 70 bpm | 0
    respiratory rate 21 | 0
    oxygen saturation 93% | 0
    crackles at lung bases bilaterally | 0
    massive splenomegaly | -1440
    acute kidney injury | 0
    creatinine 325 μmol/L | 0
    urea 28 mmol/L | 0
    eGFR 14 mL/min/1.73 m² | 0
    serum glucose 14.2 mmol/L | 0
    haemoglobin 80 g/L | 0
    platelets 103×10⁹/L | 0
    white cell count 40.3×10⁹/L | 0
    neutrophils 22.91×10⁹/L | 0
    monocytes 13.43×10⁹/L | 0
    occasional blasts | 0
    metabolic acidosis | 0
    pH 7.31 | 0
    bicarbonate 14 mmol/L | 0
    lactate 1.3 mmol/L | 0
    anion gap 21 mmol/L | 0
    chest X-ray patchy perihilar opacification | 0
    increased interstitial markings | 0
    chest infection | 0
    urinary infection | 0
    ceftriaxone | 0
    doxycycline | 0
    packed red cells transfusion | 0
    tachypnoea | 8
    desaturation 80% | 8
    blood pressure 159/53 mm Hg | 8
    heart rate 70 bpm | 8
    temperature 39.0°C | 8
    fluid overload | 8
    respiratory crackles to mid-zones bilaterally | 8
    poor urine output | 8
    arterial blood gas pH 7.26 | 24
    bicarbonate 10 mmol/L | 24
    lactate 1.1 mmol/L | 24
    anion gap 19 mmol/L | 24
    eGFR 14 mL/min/1.73 m² | 24
    troponin 42 ng/L | 24
    BNP 1544 ng/L | 24
    C-reactive protein 165 mg/L | 24
    WCC 80.4×10⁹/L | 24
    neutrophils 53.22×10⁹/L | 24
    lymphocytes 6.13×10⁹/L | 24
    monocytes 17.61×10⁹/L | 24
    eosinophils 1.15×10⁹/L | 24
    basophils 0.38×10⁹/L | 24
    sepsis | 24
    transfusion-associated circulatory overload | 24
    pulmonary oedema | 24
    haematologic transformation | 24
    piperacillin–tazobactam | 24
    furosemide | 24
    high-flow nasal prong oxygen | 24
    acidosis persisted | 48
    anion gap 21.3 mmol/L | 48
    renal ultrasound multiple small calculi | 48
    no obstruction | 48
    no hydronephrosis | 48
    urine highly positive for leukocytes | 48
    Candida sp culture | 48
    no eosinophils | 48
    no casts | 48
    no monoclonal immunoglobulin | 48
    no Bence-Jones proteins | 48
    PGA considered | 48
    dicloxacillin withheld | 72
    paracetamol withheld | 72
    blood pyroglutamic acid levels requested | 72
    cephalexin recommended | 72
    acceleration phase of leukaemia | 72
    transformation to CMML-2 | 72
    spontaneous tumour lysis syndrome | 72
    urate 1.28 mmol/L | 72
    phosphate 1.83 mmol/L | 72
    creatinine increase ≥1.5 times upper limit | 72
    Candida orthopsilosis blood cultures | 72
    fluconazole | 72
    acidosis resolved | 168
    bicarbonate 26 mmol/L | 168
    anion gap 14.8 | 168
    renal function stabilized | 168
    GFR 16 mL/min/1.73 m² | 168
    creatinine 292 μmol/L | 168
    WCC 20.1×10⁹/L | 168
    neutrophils 11.28×10⁹/L | 168
    monocytes 5.84×10⁹/L | 168
    basophils 0.20×10⁹/L | 168
    PGA confirmed | 168
    blood pyroglutamic acid 62 μmol/L | 168
    discharge to residential aged care facility | 168
    palliative care | 168
