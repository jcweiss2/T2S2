25 years old | 0 | 0 
female | 0 | 0 
autoimmune hepatitis | 0 | 0 
bilateral lower extremity pain | -168 | 0 
edema | -168 | 0 
ascites | -168 | 0 
fever | -168 | 0 
chills | -168 | 0 
nausea | -168 | 0 
dizziness | -168 | 0 
heavy menorrhagia | -168 | 0 
unprotected sexual intercourse | -336 | -336 
acetaminophen | -10080 | 0 
ibuprofen | -10080 | 0 
azathioprine | -10080 | -672 
prednisone | -10080 | -672 
influenza vaccination | -672 | -672 
COVID-19 vaccination | -672 | -672 
admitted to the hospital | 0 | 0 
hemodynamically unstable | 0 | 0 
blood pressure 67/39 mmHg | 0 | 0 
heart rate 129 beats per minute | 0 | 0 
respirations 33 per minute | 0 | 0 
temperature 35.1 degrees Celsius | 0 | 0 
jaundice | 0 | 0 
scleral icterus | 0 | 0 
abdominal ascites with fluid wave | 0 | 0 
anasarca | 0 | 0 
erythematous vaginal vault | 0 | 0 
minimal discharge | 0 | 0 
fine reticular violaceous patches | 0 | 16 
lactic acidosis | 0 | 0 
lactic acid 13.1 mmol/L | 0 | 0 
creatinine 1.49 mg/dL | 0 | 0 
aspartate transaminase 56 units/L | 0 | 0 
alanine transaminase 62 units/L | 0 | 0 
total bilirubin 3.7 mg/dL | 0 | 0 
direct bilirubin 3.19 mg/dL | 0 | 0 
alkaline phosphatase 213 units/L | 0 | 0 
total protein 5.3 g/dL | 0 | 0 
albumin 1.4 g/dL | 0 | 0 
hemoglobin 5.2 g/dL | 0 | 0 
leukocytes 1.3 k/uL | 0 | 0 
platelets 90 k/uL | 0 | 0 
prothrombin time 37.9 s | 0 | 0 
international normalized ratio 3.9 | 0 | 0 
beta-human chorionic gonadotropin test negative | 0 | 0 
schistocytes | 0 | 0 
paracentesis | 0 | 0 
peritoneal fluid analysis | 0 | 0 
leukocyte count 9821 | 0 | 0 
neutrophilic predominance | 0 | 0 
CT angiography | 0 | 0 
cirrhosis | 0 | 0 
portal hypertension | 0 | 0 
splenomegaly | 0 | 0 
edematous wall thickening of the colon and rectum | 0 | 0 
intubation | 0 | 0 
intravenous fluids | 0 | 48 
blood products | 0 | 48 
vasopressors | 0 | 48 
broad-spectrum antibiotic therapy | 0 | 48 
vancomycin | 0 | 48 
piperacillin-tazobactam | 0 | 48 
doxycycline | 0 | 48 
clindamycin | 0 | 48 
intravenous immunoglobulin | 0 | 0 
large violaceous non-blanching ecchymoses | 16 | 16 
flaccid bullae | 16 | 16 
dusky and violaceous skin | 36 | 36 
bullae | 36 | 36 
lactate dehydrogenase 298 units/L | 16 | 16 
fibrinogen 187 mg/dL | 16 | 16 
D-dimer > 20 mcg/mL | 16 | 16 
urinalysis | 16 | 16 
salicylate level negative | 16 | 16 
acetaminophen level negative | 16 | 16 
Chlamydia trachomatis nucleic acid amplification test negative | 16 | 16 
Neisseria gonorrhea nucleic acid amplification test negative | 16 | 16 
urine toxicology screen negative | 16 | 16 
peritoneal fluid culture negative | 16 | 16 
blood culture positive for Streptococcus pneumoniae | 16 | 16 
progressive hypoxia | 16 | 48 
shock | 16 | 48 
death | 48 | 48 
autopsy | 48 | 48 
cirrhotic liver | 48 | 48 
diffuse alveolar damage | 48 | 48 
serous fluid in the abdominal compartment | 48 | 48 
pneumococcal vaccination | -10080 | -10080