53 years old | 0
male | 0
unrestrained driver | -1
high-speed head-on motor vehicle collision | -1
blood pressure 80/20 mm Hg | 0
heart rate 126 beats/min | 0
tender distended abdomen | 0
no signs of seat belt markings | 0
computed tomography scan | 0
active extravasation from the infrarenal aorta | 0
surrounding retroperitoneal hematoma | 0
bilateral rib fractures | 0
pulmonary contusions | 0
left ulnar fracture | 0
right tibia fracture | 0
no associated abdominal or spinal injuries | 0
endovascular stent grafting | 1
two proximal aortic cuffs | 1
24 × 58-mm cuff placed distally | 1
24 × 39-mm cuff placed proximally | 1
inferior mesenteric artery intentionally covered | 1
follow-up CT scan | 24
resolution of the extravasation and hematoma | 24
gram-positive sepsis | 24
pneumonia | 24
respiratory failure | 24
tracheostomy | 24
discharged | 360
ambulatory condition | 360
follow-up CT scan one year later | 8760
normal aorta | 8760
stable graft configuration | 8760