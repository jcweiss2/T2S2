74 years old | 0  
    female | 0  
    admitted for bilateral total knee replacement arthroplasty | 0  
    degenerative osteoarthritis | 0  
    angina | -17520  
    hypertension | -17520  
    isosorbide-5-mininitrate | -17520  
    atenolol | -17520  
    blood tests within normal ranges | 0  
    biochemistry tests within normal ranges | 0  
    simple chest radiograph with cardiomegaly | 0  
    sinus bradycardia | 0  
    first degree atrioventricular block | 0  
    T wave inversion in leads V2-3 | 0  
    ejection fraction 60% | 0  
    CSE anesthesia | 0  
    bupivacaine injection | 0  
    epidural catheter insertion | 0  
    levobupivacaine test dose | 0  
    oxygen administered via face mask | 0  
    stable vital signs during surgery | 0  
    pulse oxygen saturation 100% | 0  
    arterial blood gas analysis within normal ranges | 0  
    operation time 3 hours 5 minutes | 0  
    anesthesia period 4 hours 25 minutes | 0  
    estimated blood loss 1100 ml | 0  
    urine volume 850 ml | 0  
    hydroxyethyl starch administered | 0  
    Hartmann solution administered | 0  
    packed RBCs administered | 0  
    transported to recovery room | 0  
    oxygen supplied via face mask | 0  
    sensation recovered to 11th thoracic segment | 0  
    pain control with levobupivacaine and fentanyl | 0  
    stable vital signs in recovery room | 0  
    arterial blood gas analysis within normal ranges | 0  
    transported to ward | 0  
    oxygen via nasal cannula | 0  
    pulse oxygen saturation 90% | 0  
    oxygen increased to 5 L/min | 0  
    drowsy mental state | 9  
    no response to calling | 9  
    opens eyes to pain | 9  
    blood pressure normal | 9  
    heart rate normal | 9  
    respiratory rate 20/min | 9  
    pulse oxygen saturation 90% | 9  
    oxygen increased to 7 L/min | 9  
    chest radiography performed | 9  
    brain CT performed | 9  
    bilateral pulmonary effusion | 9  
    no abnormal brain CT findings | 9  
    persistent symptoms | 24  
    brain MRI performed | 24  
    3D pulmonary arteriography performed | 24  
    bilateral small high signal intensity lesions | 24  
    reduced ADC | 24  
    fat embolism suggested | 24  
    no pulmonary embolism findings | 24  
    transferred to stroke unit | 24  
    shallow irregular breathing | 24  
    pulse oxygen saturation 84% | 24  
    eyeball deviation left | 24  
    nystagmus | 24  
    unresponsive to strong stimulation | 24  
    stuporous consciousness | 24  
    intubation | 24  
    oxygen saturation 58% | 24  
    blood pressure 70/40 mmHg | 24  
    transferred to ICU | 24  
    mechanical ventilator | 24  
    blood pressure 95/60 | 24  
    fever 38℃ | 24  
    low molecular weight heparin considered | 24  
    hemoglobin 8.3 g/dl | 24  
    platelets 34,000/µl | 24  
    increased coagulation time | 24  
    packed RBCs transfused | 24  
    platelets transfused | 24  
    inotropics administered | 24  
    diuretics administered | 24  
    ischemic colitis | 72  
    petechial rash | 72  
    low molecular weight heparin initiated | 96  
    stuporous consciousness | 96  
    unimproved neurological symptoms | 96  
    electroencephalogram performed | 120  
    moderate to severe diffuse cerebral dysfunction | 120  
    weaned off ventilator | 168  
    endotracheal tube removed | 312  
    improved respiratory symptoms | 312  
    improved neurological symptoms | 312  
    transferred to general ward | 408  
    multiple brain infarctions resolved | 624  
    discharged | 1056  
