52 years old | 0
female | 0
admitted for D10 neurofibroma excision | 0
pre-operative fasting (solid food) | -7
pre-operative fasting (clear water) | -2
uneventful laminectomy and tumor excision | 0
general anesthesia | 0
prone position | 0
surgery duration | 4
intraoperative fentanyl | 0
paracetamol administration | -0.5
reversal of neuromuscular blockade | 0
extubation | 0
shifted to PACU | 0
nausea | 0.5
abdominal pain | 0.5
agitation | 0.5
tachypnea | 0.5
dry mouth, tongue, lips | 0.5
hypotension | 0.5
tachycardia | 0.5
afebrile | 0.5
blood glucose 464 mg/dl | 0.5
ABG analysis (pH 7.12) | 0.5
high anion gap metabolic acidosis | 0.5
bicarbonate 8 mmol/L | 0.5
base deficit 18 | 0.5
AG 22 | 0.5
potassium 4.2 mmol/L | 0.5
sodium 132 mmol/L | 0.5
urinary glucose | 0.5
urinary ketones | 0.5
serum β-hydroxybutyrate 5.8 mmol/L | 0.5
DKA diagnosis | 0.5
fluid resuscitation (0.9% NS) | 0.5
insulin bolus 6 U | 0.5
continuous insulin infusion | 0.5
electrolyte correction | 0.5
serum amylase 210 U/L | 0.5
lipase 155 U/L | 0.5
resolution of ketoacidosis | 0.5
subcutaneous insulin initiation | 0.5
shifted to ward | 72
HbA1c 7.2% | 72
sterile blood cultures | 72
sterile urine cultures | 72
blood glucose normalization | 72
discharged | 168
pre-operative fasting (solid food) | -168
pre-operative fasting (clear water) | -120
afebrile |C:\Users\yuheng\AppData\Local\Temp\1\2\4\5\7\8\9\a\b\c\d\e\f\10\11\12\13\14\15\16\17\18\19\1a\1b\1c\1d\1e\1f\20\21\22\23\24\25\26\27\28\29\2a\2b\2c\2d\2e\2f\30\31\32\33\34\35\36\37\38\39\3a\3b\3c\3d\3e\3f\40\41\42\43\44\45\46\47\48\49\4a\4b\4c\4d\4e\4f\50\51\52\53\54\55\56\57\58\59\5a\5b\5c\5d\5e\5f\60\61\62\63\64\65\66\67\68\69\6a\6b\6c\6d\6e\6f\70\71\72\73\74\75\76\77\78\79\7a\7b\7c\7d\7e\7f\80\81\82\83\84\85\86\87\88\89\8a\8b\8c\8d\8e\8f\90\91\92\93\94\95\96\97\98\99\9a\9b\9c\9d\9e\9f\a0\a1\a2\a3\a4\a5\a6\a7\a8\a9\aa\ab\ac\ad\ae\af\b0\b1\b2\b3\b4\b5\b6\b7\b8\b9\ba\bb\bc\bd\be\bf\c0\c1\c2\c3\c4\c5\c6\c7\c8\c9\ca\cb\cc\cd\ce\cf\d0\d1\d2\d3\d4\d5\d6\d7\d8\d9\da\db\dc\dd\de\df\e0\e1\e2\e3\e4\e5\e6\e7\e8\e9\ea\eb\ec\ed\ee\ef\f0\f1\f2\f3\f4\f5\f6\f7\f8\f9\fa\fb\fc\fd\fe\ff\<|eot_id|>
