58 years old | 0
female | 0
hyperthyroidism | 0
osteoporosis | 0
COPD | 0
classified for lung transplantation | -672
PaO2 61.2 mmHg | -672
PaCO2 44 mmHg | -672
FEV1 0.44 l | -672
FVC 1.38 l | -672
6-MWT 174 metres | -672
RVSP 36 mmHg | -672
PRA 3% | -672
donor identification | -96
transplantation | 0
anterolateral thoracotomy | 0
transverse sternotomy | 0
implantation of left donor lung | 0
anastomosis of pulmonary artery and vein | 0
ventilation resumed | 0
haemostasis obtained | 0
drains inserted | 0
closure of thorax | 0
ICU stay | 0
plasmapheresis | 24
human immunoglobulin | 24
rituximab | 24
primary graft dysfunction | 72
emphysema of recipient's own lung | 72
C1-esterase | 72
lung volume reduction surgery | 72
prolonged air leakage | 72
infusion of FFP | 72
infusion of PRBCs | 72
infusion of albumin | 72
right lung drainage removed | 168
left lung drainage removed | 840
discharged | 1056
PO2 68.9 mmHg | 1056
PCO2 44.0 mmHg | 1056
FEV1 1.12 l | 1056
FVC 1.38 l | 1056
6-MWT 246 metres | 1056
cyclosporine | 1056
mycophenolate mofetil | 1056
prednisone | 1056
first acute organ rejection episode | 1056
methylprednisolone | 1096
tacrolimus | 1096
Moraxella catarrhalis infection | 1096
amoxicillin with clavulanic acid | 1096
transient renal failure | 1096
ion disorders | 1096
hypoproteinaemia | 1096
leukopaenia | 1096
bronchitis | 1344
Corynebacterium pseudodiphtericum | 1344
Escherichia coli urinary tract infection | 1344
second episode of acute graft rejection | 1344
E. coli sepsis | 1560
ceftazidime | 1560
cytomegalovirus disease | 1560
ganciclovir | 1560
pulmonary embolism | 1560
anxiety disorder | 1560
opipramol | 1560
venlafaxine | 1560
leukopenia | 1560
pantoprazole dose reduced | 1560
mycophenolate mofetil dose reduced | 1560
third episode of acute graft rejection | 1824
Pseudomonas aeruginosa infection | 1824
ciprofloxacin | 1824
ceftazidime | 1824
bilateral otitis | 1824
clindamycin | 1824
budesonide inhalation | 1824
hypogammaglobulinaemia | 1824
human immunoglobulins | 1824
bacterial infections | 2544
Acinetobacter baumanii | 2544
Proteus mirabilis | 2544
Candida albicans | 2544
C. glabrata | 2544
Aspargillus species | 2544
cefuroxime | 2544
imipenem | 2544
ampicillin with sulbactam | 2544
amikacin | 2544
amphotericin B | 2544
itraconazole | 2544
colistin | 2544
drug-induced diabetes | 2544
glimepiride | 2544
insulin therapy | 2544
renal failure | 2544
fourth episode of acute lung rejection | 2544
cytomegalovirus disease | 3024
valganciclovir | 3024
leukopaenia | 3024
fifth episode of rejection | 3024
renal failure | 3024
destabilisation of diabetes | 3024
Acinetobacter baumani | 3024
Klebsiella pneumoniae | 3024
Candida albicans | 3024
ceftazidime | 3024
ciprofloxacin | 3024
ampicillin with sulbactam | 3024
colistin | 3024
metronidazole | 3024
tazobactam | 3024
itraconazole | 3024
nystatin | 3024
anti-HLA antibodies | 3024
depression | 3024
mianserin | 3024
posttraumatic haematoma | 3024
VAC-therapy | 3024
death | 4752