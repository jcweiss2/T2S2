history of PAN | -8760
history of paroxysmal atrial fibrillation | -8760
history of hypertension | -8760
history of dyslipidemia | -8760
history of non-insulin dependent diabetes mellitus | -8760
history of admission for septic shock | -720
scrotal pain | 0
fever of 103°F | 0
fatigue | 0
tachycardia to 130 beats per minute | 0
hypotension to 103/40 mm Hg | 0
broad-spectrum antibiotics consisting of vancomycin and Zosyn | 0
admission under medicine service | 0
worsening kidney function | 24
switch in antibiotics to meropenem | 24
continued to spike fevers | 48
no specific source of an infection found | 48
no focus found on CT chest, abdomen, and pelvis | 48
stopping all antibiotics | 48
macular rash | 168
rash progressed to involve axillary area | 240
rash progressed to involve chest, head, neck, and abdomen | 336
decline of mental status | 336
worsening of skin lesions | 336
element of bullae and vesicles | 336
dermatology team involved | 336
biopsy obtained | 336
initiating local steroid cream | 336
rash became pustular | 504
high grade fever of 109°F | 504
transfer to intensive care unit | 504
protocol of cooling | 504
pulse steroids administered | 504
fever subsided | 534
improvement of rash | 534
decreased progression of sloughing | 534
complete resolution of acute kidney injury | 534
taper in steroids | 534
skin biopsy | 0
urine analysis | 0
CT chest/abdomen/pelvis | 0
CBC/BMP/coagulation | 0
differential diagnosis | 0
Generalized acute pustular psoriasis | 0
Acute generalized exanthematous pustulosis | 0
Drug reaction with eosinophilia and systemic manifestation | 0
Steven Johnson syndrome | 0
Leukocytoclastic vasculitis | 0
Subcorneal pustular dermatosis | 0
Cutaneous candidiasis | 0
final diagnosis of AGEP | 504
initiation of immunosuppressive management | 720
discharge from hospital | 720