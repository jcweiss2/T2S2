57 years old | 0
Hispanic | 0
male | 0
admitted to the hospital | 0
coronary artery disease | -6336
myocardial infarction | -6336
ischemic dilated cardiomyopathy | -6336
pocket infection of his cardiac resynchronization therapy defibrillator | 0
erythema | -144
discomfort | -144
edema | -144
serosanguinous drainage | -144
oral amoxicillin treatment | -144
nonbacteremic | 0
afebrile | 0
severely reduced left ventricular systolic function | 0
ejection fraction of 20%–25% | 0
global hypokinesis of the left ventricle | 0
no evidence of vegetations | 0
leads were scarred to the lateral wall of the superior vena cava | 0
transvenous lead extraction | 0
cardiac resynchronization therapy defibrillator pocket capsule was dissected out | 0
device removed | 0
coronary sinus and right atrial leads were extracted | 0
hypotensive | 0
transesophageal echocardiography revealed a large pericardial effusion | 0
emergency midsternotomy | 0
pericardium was opened | 0
significant amount of blood was seen | 0
bleeding was manually controlled | 0
cardiopulmonary bypass was instituted | 0
5-mm tear in the superior cavoatrial junction | 0
perforation in the right atrium | 0
oozing hematoma at the level of the innominate vein | 0
lesions were repaired | 0
right ventricular lead was capped and abandoned | 0
intra-aortic balloon pump was placed | 0
multiple blood transfusions | 0
coagulopathy | 0
transfusions of cryoprecipitate, platelets, fresh frozen plasma, and factor VII | 0
chest was closed | 0
postoperatively transferred to the intensive care unit | 0
severe cardiogenic shock | 0
multiorgan failure | 0
hypotensive | 0
required large doses of vasopressin, epinephrine, and norepinephrine | 0
hypoxic respiratory failure | 0
mechanical ventilation | 0
liver failure | 0
albumin | 0
multiple blood products | 0
broad-spectrum antibiotics | 0
oliguric | 0
continuous venovenous hemodialysis | 24
acute renal failure | 24
bilateral, symmetrical cyanotic changes | 48
vasopressor administration was stopped | 48
upper- and lower-digit ischemia | 216
dry gangrene | 216
dull pain | 216
no ability to move his fingers and toes | 216
bilateral stiffness | 216
2+ pitting edema | 216
nonexistent capillary refill time | 216
palpable 2+ peripheral pulses | 216
Doppler study showed flat waveforms | 216
intra-aortic balloon pump was removed | 168
endotracheal tube was removed | 168
albumin was discontinued | 264
liver enzymes returned to normal limits | 264
kidney function gradually improved | 984
hemodialysis was stopped | 984
mental status improved | 984
necrotic lesions were treated conservatively | 984
povidone-iodine dressings | 984
debridement | 648
negative-pressure wound therapy | 648
purulent, foul-smelling material | 1296
transferred to our facility | 1296
preoperative transesophageal echocardiography | 1296
diminished ejection fraction of 10%–15% | 1296
laser extraction of his retained lead | 1392
60 mL of pus was drained | 1392
antibiotic regimen | 1392
microbial cultures grew Enterobacter cloacae and Staphylococcus epidermidis | 1392
failed screening for subcutaneous implantable cardioverter-defibrillator | 1392
transvenous implantable cardioverter-defibrillator system was implanted | 1568
evaluation of his hands and feet | 1568
no signs of local infection or wet gangrene | 1568
black skin changes and demarcation lines | 1568
frank mummification of his digits and toes | 1568
discharged | 1848
amputation and debridement of his necrotic feet | 2556
amputation of his fingers is scheduled | 2556