44 years old | 0
male | 0
chronic hepatitis B virus carrier | 0
normal liver function | 0
admitted to the hospital | 0
dry cough | -168
shortness of breath | -168
hypodynamia | -168
frequent coughing | -72
yellow-white sputum | -72
high fever | -72
20-year history of smoking | -72000
approximately twenty cigarettes daily | -72000
temperature of 38.7°C | 0
heart rate of 134/min | 0
respiratory rate of 24/min | 0
blood pressure of 124/70 mmHg | 0
fine crackles in the left lung | 0
patchy high-density shadows with blurred margins | 0
pan-lobar pneumonia | 0
slightly elevated leucocyte count | 0
elevated D-dimer | 0
elevated glucose levels | 0
elevated blood urea nitrogen | 0
elevated creatinine | 0
elevated C reactive protein | 0
elevated procalcitonin | 0
elevated alanine aminotransferase | 0
elevated aspartate aminotransferase | 0
elevated lactic dehydrogenase | 0
elevated creatine kinase | 0
elevated serum total bilirubin | 0
decreased serum albumin | 0
decreased serum sodium | 0
normal pH | 0
normal PaO2 | 0
normal blood lactate | 0
decreased PaCO2 | 0
decreased PO2/FiO2 | 0
intubation | 6
ventilator | 6
delirium | 6
transferred to ICU | 6
respiratory status deteriorated | 6
episodes of significant hypoxemia | 12
hemorrhagic fluid gushed out from tracheal tube | 12
wet and dry rales | 12
ARDS | 12
lung-protective ventilation | 12
deep sedation | 12
analgesia | 12
paralysis using neuromuscular blocker | 12
continuous renal replacement therapy | 12
prone-position ventilation | 12
bilateral pulmonary infiltrates increased | 48
leucocyte count increased | 48
PCT levels increased | 48
VV-ECMO | 48
cannulation | 48
ventilatory parameters adjusted | 48
BALF sample obtained | 48
mNGS detection | 48
IL-6 level elevated | 48
IL-8 level elevated | 48
IL-10 level elevated | 48
intravenous antibiotic therapy continued | 48
moxifloxacin | 48
imipenem and cilastatin sodium | 48
C. abortus detected | 48
PCR assay | 48
doxycycline | 72
azithromycin | 72
imipenem and cilastatin sodium | 72
symptoms improved | 96
inflammation indicators improved | 96
neuromuscular blocker discontinued | 96
norepinephrine dosage down-regulated | 96
pulmonary infiltrates improved | 96
lung compliance improved | 96
liver function deteriorated | 96
serum total bilirubin elevated | 96
discharged | 120
passed away | 128