72 years old | 0
male | 0
high-grade fever | -96
referred to a nearby clinic | -96
wife influenza B infection | -168
two daughters influenza B infection | -168
rapid test positive for influenza B antigens | -96
influenza B virus infection diagnosis | -96
oseltamivir administration | -96
persistent fever | -24
dyspnea at rest | -24
admitted to the hospital | 0
temperature 38.7°C | 0
blood pressure 117/80 mmHg | 0
heart rate 76 beats/min | 0
oxygen saturation 88% on room air | 0
fine crackles in lung fields | 0
white blood cell count 7400/mm³ | 0
C-reactive protein 18.1 mg/dL | 0
aspartate transaminase 91 IU/L | 0
L-lactate dehydrogenase 362 IU/L | 0
creatine kinase 793 IU/L |= 0
Krebs von den Lungen-6 1772 U/mL | 0
arterial blood gas analysis hypoxemia | 0
PaO2 72 Torr | 0
nasal oxygen inhalation 5 L/min | 0
chest radiography ground-glass opacity | 0
chest CT diffuse ground-glass opacity | 0
Gram staining negative | 0
Ziehl-Neelsen staining negative | 0
periodic acid-Schiff stain negative | 0
sputum culture negative | 0
blood cultures negative | 0
high-flow nasal oxygen support | 0
peramivir 600 mg/day | 0
piperacillin/tazobactam 13.5 g/day | 0
levofloxacin 500 mg/day | 0
chest CT reticular shadow worsening | 72
PaO2/FiO2 ratio 83 | 72
severe ARDS diagnosis | 72
mechanical ventilation proposed | 72
high PEEP proposed | 72
refusal of intubation | 72
continued high-flow nasal oxygen | 72
polymyxin B-immobilized hemoperfusion | 72
methylprednisolone 60 mg/day | 144
respiratory status no improvement | 144
reticular infiltrates worsening | 144
noninvasive positive pressure ventilation | 144
cyclophosphamide 500 mg biweekly | 144
condition worsening | 3096
death | 3096
autopsy performed | 3096
diffuse alveolar damage | 3096
hyaline membranes | 3096
no specific abnormality in other organs | 3096
