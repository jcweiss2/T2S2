cactus plant injury | -168
left leg swelling | -168
progressive left leg swelling | -48
worsening of erythema | -48
pain | -48
generally unwell | -48
presentation to ED | 0
admitted to ICU | 0
triple vasopressor support initiated | 0
antibiotics initiated | 0
emergency left lower limb fasciotomy | 0
debridement | 0
below knee amputation | 0
post operatively intubated | 1
oliguria | 1
severe acidosis | 1
left internal jugular vascath insertion | 1
CRRT commenced | 1
ventilation sedation | 1
IVIgG therapy initiated | 1
new onset RAF | 2
remained oliguric | 2
echocardiography | 2
amiodarone loading dose | 2
antibiotics unchanged | 2
CRRT continued | 2
Oxiris filter applied | 2
citrate based anticoagulation circuit applied | 2
sepsis induced coagulopathy | 3
bedside surgical debridement | 3
histopathology consistent with NF | 3
wound culture for MCS | 3
tissue culture | 3
vasopressor support weaning | 3
antibiotics unchanged | 3
CRRT continued | 3
oliguria | 4
new onset purpura | 4
weeping skin tears | 4
ongoing RAF | 4
citrate based CRRT continued | 4
double inotropic support | 4
amiodarone infusion | 4
fulminant hepatic failure | 5
encephalopathy | 5
refractory oliguria | 5
dual inotropic support | 5
antibiotics unchanged | 5
CRRT continued | 5
severely deconditioned | 6
ICU acquired weakness | 6
unarousable | 6
no response to noxious stimuli | 6
sedation weaned off | 6
vasopressor weaned off | 6
antibiotic de-escalation | 6
CRRT continued | 6
hyper-ammonium therapy initiated | 6
PRBCs transfusion | 6
jaundice | 7
hypoactive delirium | 7
new onset lateralizing signs | 7
CT brain | 7
ultrasound abdomen | 7
acute calculous cholecystitis | 7
CRRT continued | 7
anuria | 8
hypotensive | 8
febrile | 8
RAF | 8
significant deterioration | 8
commenced on palliative care pathway | 8
deceased | 8
troponin | 8
ammonia | 8
LFT | 8
CRRT continued | 8
renal recovery assessment | 8
vasopressor support recommenced | 8
antibiotic regimen | 8
digoxin | 8
metoprolol | 8