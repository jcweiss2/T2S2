50 years old | 0
male | 0
admitted to the ICU | 0
no past history | 0
emergency decompressive craniectomy | -192
hematoma removal | -192
spontaneous intracerebral and intraventricular hemorrhage | -192
no neurological recovery | -192
follow-up brain CT | -192
rebleeding | -192
second surgery | -192
transferred to hospital for organ donation | -24
brain death | -24
vital signs: blood pressure 75/50 mmHg | 0
vital signs: heart rate 72 bpm | 0
vital signs: pulse oxygen saturation 75% | 0
fluid administration | 0
continuous intravenous infusion of dopamine | 0
mechanical ventilation support | 0
general edema | 0
pink frothy sputum | 0
rales | 0
bilateral infiltration on chest X-ray | 0
concentric left ventricular hypertrophy | 0
preserved contractility | 0
no pulmonary arterial hypertension | 0
first arterial blood gas analysis | 0
pH 7.310 | 0
PaCO2 40.5 mmHg | 0
PaO2 84.9 mmHg | 0
HCO3- 19.9 mEq/L | 0
base excess -5.9 mEq/L | 0
SaO2 94.3% | 0
NPE | 0
hypoxemia | 0
apnea test | 2
SaO2 85.7% | 2
PaO2 66.7 mmHg | 2
alveolar recruitment maneuvers | 2
SpO2 91-93% | 2
SpO2 96.3% | 2
PaO2 93.4 mmHg | 2
frothy sputum removal | 2
dopamine infusion | 2
systolic pressure 90-120 mmHg | 2
diastolic pressure 50-80 mmHg | 2
HR 80-95 bpm | 2
central venous pressure 11-13 mmHg | 2
diabetes insipidus | 2
metabolic acidosis | 2
hyperglycemia | 2
hypernatremia | 2
fluid supplementation | 2
electrolyte correction | 2
sodium bicarbonate administration | 2
insulin infusion | 2
warm air blanket | 2
body temperature 36℃ | 2
total fluids administered 6280 ml | 10.5
total urine output 3840 ml | 10.5
fluid drained from nasogastric tube 1300 ml | 10.5
brain death declaration | 10.5
transfer to OR | 10.5
oxygen 12 L/min | 10.5
manual ventilation | 10.5
vital signs before transfer: BP 120/70 mmHg | 10.5
vital signs before transfer: HR 75 bpm | 10.5
vital signs before transfer: SpO2 99% | 10.5
vital signs in OR: BP 87/55 mmHg | 10.8
vital signs in OR: HR 100 bpm | 10.8
vital signs in OR: SpO2 80% | 10.8
anesthesia machine connection | 10.8
mechanical ventilation | 10.8
SpO2 91% | 10.8
alveolar recruitment maneuvers | 10.8
PEEP 15 cmH2O | 10.8
PIP 30 cmH2O | 10.8
ABGA | 10.8
pH 7.412 | 10.8
PaCO2 33.0 mmHg | 10.8
PaO2 62.3 mmHg | 10.8
HCO3- 20.5 mEq/L | 10.8
BE -3.6 mEq/L | 10.8
SaO2 90.8% | 10.8
dopamine infusion | 10.8
epinephrine infusion | 10.8
NO inhalation | 11
SpO2 99% | 11.3
ABGA | 11.3
pH 7.270 | 11.3
PaCO2 46.3 mmHg | 11.3
PaO2 328.7 mmHg | 11.3
HCO3- 20.8 mEq/L | 11.3
BE -6.0 mEq/L | 11.3
SaO2 99.5% | 11.3
surgery completion | 13.8
kidney retrieval | 13.8
cardiac arrest | 13.8
death declaration | 13.8