56 years old | 0
female | 0
admitted to the hospital | 0
left hydronephrosis | -672
ureteroscopy for left ureter | -48
laparoscopy for lysis of adhesions around left ureter | -48
abdominal discomfort | -48
abdominal distension | -48
oliguria | -48
irritability | -48
body temperature of 39.4°C | -48
pulse rate at 114 beats per minute | -48
blood pressure declined to 86/59 mm Hg | -48
respiratory rate at 28 breaths per minute | -48
oxygen saturation of 89% under oxygen inhalation | -48
white blood cell count of 15.4 × 10^9/L | -48
neutrophils 95% | -48
lymphocytes 5% | -48
platelet count down to 33 × 10^9/L | -48
blood lactate level of 3.6 mmol/L | -48
base excess of -11.4 | -48
serum creatinine increased to 365.7 μmol/L | -48
alanine aminotransferase (ALT) of 224 U/L | -48
aspartate aminotransferase (AST) of 858 U/L | -48
prothrombin time extended to 24.2 seconds | -48
serum level of C-reactive protein of 180.3 mg/L | -48
procalcitonin (PCT) of 49.17 ng/mL | -48
qSOFA score of 3 points | -48
transferred to the ICU | 0
APACHE II score of 32 | 0
SOFA score of 17 | 0
sepsis diagnosis | 0
Primaxin (imipenem/cilastatin) administration | 0
norepinephrine administration | 0
hydrocortisone administration | 0
supplemental fluids administration | 0
continuous renal replacement therapy | 0
respiratory distress | 24
oxygenation index falling down to 184 mm Hg | 24
endotracheal intubation | 24
mechanical ventilation | 24
white blood cell count peaked at 45.3 × 10^9/L | 48
neutrophils 91.5% | 48
lymphocytes 1.8% | 48
C-reactive protein decrease | 48
PCT decrease | 48
ALT decrease | 48
AST decrease | 48
platelet count increase | 48
liver injury aggravation | 120
total bilirubin (TB) rose to 245.5 μmol/L | 120
direct bilirubin (DB) of 196.6 μmol/L | 120
liver function index indicated liver failure | 120
abdominal ultrasound examination | 120
gallbladder wall edema | 120
hepatitis serology negative | 120
autoantibodies for autoimmune liver diseases negative | 120
hepatoprotective drugs administration | 0
supportive therapies | 0
plasma exchange | 120
plasma exchange volume of 1.5 to 3.0 L per day | 120
plasma exchange rate of 1.0 to 1.2 L per hour | 120
mechanical ventilation stopped | 216
endotracheal tube withdrawn | 216
hemodialysis treatment continued | 216
transfer back to the urology department | 288
serum ALT of 23 U/L | 288
AST of 39 U/L | 288
TB of 99.4 μmol/L | 288
DB of 69.8 μmol/L | 288
liver function returned to normal | 295