48 years old | 0
female | 0
Caucasian | 0
admitted to the hospital | 0
burns to the face | 0
inhalation injury | 0
intubated | 0
diffuse carbonaceous sputum | 0
pale friable mucosa | 0
airway protection | 0
sedation | 0
neuromuscular blockade | 0
severe depression | 0
psychotic features | 0
paliperidone palmitate | 0
paliperidone | 0
citalopram | 0
trazodone | 0
risperidone | 0
clonazepam | 0
no known drug allergies | 0
chronic smoker | 0
substance abuser | 0
urine drug screen negative | 0
mild leukocytosis | 0
afebrile | 0
normotensive | 0
adequate urine output | 0
acute respiratory distress syndrome | 0
pressure control ventilation | 0
tracheostomy | 24
febrile | 48
tachycardia | 48
thick yellow secretions | 120
diffuse rhonchi | 120
worsening right-sided patchy infiltrate | 120
culture from broncheo-alvelolar lavage | 144
gram-positive cocci in clusters | 144
vancomycin | 144
cefepime | 144
MRSA | 144
vancomycin MIC = 2 mg/L | 240
ceftaroline fosamil | 240
Teflaro | 240
inhalational thermal injuries | 240
burn patients | 240
PK characterization | 240
serum concentrations | 240
ceftaroline levels | 288
Cmax | 288
Cmin | 288
T ½ | 288
Vd | 288
AUC0–τ | 288
T > MIC | 288
clearance | 288
burn patient | 288
package insert | 288
serum drug assay | 288
PK/PD | 288
antibiotic therapy | 288
infection | 288
mechanical ventilation | 528
decannulated | 552
psychiatric care facility | 1152
discharged | 1152