60 years old | 0  
    man | 0  
    visited the emergency department | 0  
    fever | 0  
    working on farms | -0  
    close contact with swine | -0  
    fever (up to 39.7°C) | 0  
    no defining abnormal findings in physical examinations | 0  
    no specific findings in laboratory data | 0  
    no specific findings in urinalysis | 0  
    no active lung lesion in chest radiograph | 0  
    mild gas accumulation in erect abdominal imaging | 0  
    no definite obstructive lesion in abdominal computed tomography | 0  
    symptoms improved following hydration | 0  
    use of analgesics | 0  
    discharged from the hospital | 0  
    revisited the emergency department | 24  
    persistent fever | 24  
    dizziness | 24  
    vomiting | 24  
    acutely ill | 24  
    drowsy | 24  
    blood pressure of 70/60 mmHg | 24  
    heart rate of 52 beats/min | 24  
    respiratory rate of 20 breaths/min | 24  
    body temperature of 36.0°C | 24  
    lung sounds clear | 24  
    bowel sounds decreased | 24  
    leukopenia | 24  
    white blood cell count 1.470 × 109/L | 24  
    neutrophils 85% | 24  
    lymphocytes 14% | 24  
    monocytes 1% | 24  
    thrombocytopenia | 24  
    platelet count 40 × 109/L | 24  
    higher urea nitrogen | 24  
    higher creatinine | 24  
    urea nitrogen 30.9 mg/dL | 24  
    creatinine 3.04 mg/dL | 24  
    hyperbilirubinemia | 24  
    total bilirubin 3.35 mg/dL | 24  
    metabolic acidosis | 24  
    pH 7.25 | 24  
    pCO2 30.5 mmHg | 24  
    bicarbonate 13.2 mmol/L | 24  
    no active lung lesion in chest radiograph | 24  
    gas accumulation in supine abdominal imaging | 24  
    erect abdominal imaging not performed | 24  
    meropenem administered | 24  
    vancomycin administered | 24  
    blood sample taken for bacterial culture | 24  
    admitted to the intensive care unit | 24  
    blood pressure of 104/48 mmHg | 6  
    heart rate of 130 beats/min | 6  
    respiratory rate of 22 breaths/min | 6  
    continuous infusion of inotropics | 6  
    dopamine 27 μg/min/kg | 6  
    norepinephrine 1.7 μg/min/kg | 6  
    low dose corticosteroid | 6  
    hydrocortisone 100 mg every 8 hours | 6  
    generalized tonic-clonic seizure | 14  
    peripheral oxygen saturation dropped to <90% | 14  
    oxygen therapy | 14  
    endotracheal intubation performed | 14  
    mechanical ventilator applied | 14  
    peripheral oxygen saturation maintained between 95% and 100% | 16  
    total urine output over 16 hours zero | 16  
    substantial hydration | 16  
    use of diuretics | 16  
    continuous renal replacement therapy initiated | 16  
    aerobic blood cultures showed bacterial growth | 12  
    anaerobic blood cultures showed bacterial growth | 12  
    blood cultures revealed gram-positive cocci | 48  
    organisms identified as S. suis | 96  
    vancomycin replaced with ampicillin/sulbactam | 96  
    meropenem replaced with ampicillin/sulbactam | 96  
    vital signs stabilized after 4 days of treatment | 96  
    dopamine administration tapered | 96  
    norepinephrine administration tapered | 96  
    drowsiness did not improve | 96  
    hydrocortisone changed to dexamethasone 5 mg/day | 96  
    ventilator weaning | 168  
    extubation | 168  
    continuous renal replacement therapy stopped | 168  
    mental status improved | 168  
    difficulty in hearing | 168  
    otoscopic examination revealed no abnormal findings | 168  
    tuning fork examination indicated bilateral sensorineural hearing loss | 168  
    spinal tap performed | 168  
    white blood cell count 7/mm3 | 168  
    red blood cell count 16/mm3 | 168  
    opening pressure within normal range 80 mmH2O | 168  
    CSF glucose 143 mg/dL | 168  
    serum glucose 265 mg/dL | 168  
    protein levels higher 125 mg/dL | 168  
    dexamethasone continued 5 mg/day for 3 days | 168  
    dexamethasone continued 2.5 mg/day for 3 days | 168  
    dexamethasone continued 1 mg/day for 3 days | 168  
    back pain | 240  
    back pain did not respond to analgesic drugs | 240  
    bone marrow signal alteration | 240  
    end plate irregularity of the left first and second lumbar spine levels | 240  
    partially unenhanced lesion in the right iliacus muscle | 240  
    partially unenhanced lesion in the left iliopsoas muscle | 240  
    infective spondylitis | 240  
    intramuscular abscess formation | 240  
    no neurologic abnormality noted | 240  
    multiple abscesses located in area not easily accessible percutaneously | 240  
    medical treatment continued with ampicillin/sulbactam | 240  
    transferred to another hospital | 240  
    back pain improved | 240  
    completed 6-week treatment with antibiotics | 240  
    nearly recovered | 240  
    hearing difficulty | 240  
    regularly visiting otolaryngology outpatient department | 240  
    sepsis | 24  
    septic shock | 24  
    multiple abscess formation | 240  
    septic emboli | 240  
    enterocolitis | 24  
    meningitis | 24  
    bacteremia | 24  
    decreased mental focus | 24  
    seizure | 24  
    labyrinthitis | 168  
    infective spondylitis | 240  
    septic arthritis | 240  
    endocarditis | 240  
    pneumonia | 240  
    peritonitis | 240  
    hearing loss | 168  
    septic emboli | 240  
    spondylodiscitis | 240  

    60 years old | 0  
    man | 0  
    visited the emergency department | 0  
    fever | 0  
    working on farms | -0  
    close contact with swine | -0  
    fever (up to 39.7°C) | 0  
    no defining abnormal findings in physical examinations | 0  
    no specific findings in laboratory data | 0  
    no specific findings in urinalysis | 0  
    no active lung lesion in chest radiograph | 0  
    mild gas accumulation in erect abdominal imaging |/tmp/foo.txt