63 years old | 0
female | 0
admitted to the hospital | 0
general body malaise | -48
diarrhea | -48
vomiting | -48
influenza-like symptoms | -48
confusion | 0
splenectomy | -38760
idiopathic thrombocytopenic purpura | -38760
menometrorhagia | -38760
vaccinated with PPV23 | -6720
fever | 0
hypotension | 0
bradycardia | 0
tachypnea | 0
decreased oxygen saturation | 0
cyanosis | 0
severe sepsis | 0
volume therapy | 0
broad-spectrum antimicrobial therapy | 0
hydrocortisone | 0
white blood cell count | 0
neutrophils | 0
hemoglobin | 0
thrombocytes | 0
C-reactive protein | 0
P-lactate | 0
aB-P-O2 | 0
aB-P-CO2 | 0
aB-pH | 0
Streptococcus pneumococcal urinary antigen test | 0
disseminated intravascular coagulation | 24
microthrombi | 24
blood cultures | 48
S. pneumoniae | 48
antimicrobial treatment | 48
penicillin G | 48
suspicion of endocarditis | 72
trans-thoracic echocardiography | 72
modest hypokinesia | 72
ejection fraction | 72
necrosis of fingertips and toes | 72
renal insufficiency | 72
hemodialysis | 72
antibiotic therapy | 72
ceftriaxone | 72
leucocytes | 96
CRP | 96
fever | 96
tracheal secret | 96
culture | 96
negative | 96
transferred from ICU | 216
antibiotics stopped | 216
serological analysis | 216
pneumococcal isolate | 216
serotype 12F | 216
discharged | 528
oral dicloxacillin | 528
necrotic tissue | 528
wound cultures | 528
Staphylococcus aureus | 528
haemolytic streptococci group C/G | 528
amputated | 7776
readmitted | 10320
severe sepsis | 10320
sepsis regimen | 10320
ceftriaxone therapy | 10320
transesophageal echocardiography | 10320
endocarditis | 10320
aortic valve | 10320
blood cultures | 10320
S. pneumoniae | 10320
antimicrobial treatment | 10320
penicillin G | 10320
conservative treatment | 10320
recovered | 11280
serological tests | 10320
pneumococcal capsule polysaccharides | 10320
serotype 12F | 10320
antibodies | 10320
serological analyses | 10320
antibody response | 10320
hyporesponsiveness | 10320
memory B cell pool | 10320
IgG | 10320
PCP | 10320
Luminex | 10320
median fluorescence intensity | 10320
μg/ml | 10320
geometric mean | 10320
SSI’s in-house reference serum | 10320
titer cut-offs | 10320
vaccination coverage | 10320
antipneumococcal-12F-antibodies | -5184
antipneumococcal-12F-antibodies | 4320
antipneumococcal-12F-antibodies | 11280