9 years old | 0
male | 0
previously healthy | 0
periumbilical abdominal pain | -96
watery diarrhea | -96
vomiting | -96
fever | -96
progressive worsening of the pain | -96
discharged home | -24
analgesics | -24
worsening of previous symptoms | 0
antibiotics | 0
transferred | 0
diagnostic procedures | 0
surgical evaluation | 0
dysuria | 0
oliguria |*0
hemodynamically stable | 0
abdominal pain | 0
signs of peritonitis | 0
fasting | 0
ceftriaxone | 0
metronidazole | 0
maintenance fluid | 0
ultrasound examination inconclusive | 0
hypothesis of MIS-C | 0
serology | 0
RT-PCR nasopharynx/oropharynx swab | 0
persistent abdominal pain | 24
several diarrhea episodes | 24
persistent tachycardia | 24
abdominal CT | 24
perforated appendix | 24
pelvic abscess | 24
appendectomy | 24
exploratory laparotomy | 24
abscess formation | 24
drain placement | 24
anatomopathological examination | 24
ulceration | 24
inflammatory infiltrate | 24
neutrophils | 24
mononuclear cells | 24
hemorrhage | 24
wall necrosis | 24
loss of mucosa | 24
SARS-CoV-2 nucleocapsid protein detected | 24
SARS-CoV-2 molecular detection | 24
admitted to PICU | 24
fluid resuscitation | 24
oxygen support | 24
laboratory tests | 24
echocardiogram | 24
hemodynamically stable | 24
clinical improvement | 24
discharged home | 216
COVID-19 infection confirmed | 24
IgG positive | 24
IgM inconclusive | 24
RT-PCR positive | 24
elevated C-reactive protein | 24
elevated fibrinogen | 24
elevated D-dimer | 24
elevated ferritin | 24
leukocytosis | 24
lymphopenia | 24
elevated INR | 24
elevated troponin | 24
elevated creatine kinase | 24
blood culture negative | 24
virus identification in appendix tissue | 24
MIS-C suspected | 24
clinical support | 24
mild MIS-C confirmed | 24
asymptomatic previous infection | 24
appendicitis as part of MIS-C | 24
acute abdomen | 24
SARS-CoV-2 infection confirmed | 24
GI manifestation considered | 24
clinical management | 24
surgical management | 24
