40 years old| 0
male | 0
admitted to tertiary hospital’s intensive care unit (ICU) | 0
acute ischemic stroke | 0
type 1 diabetes mellitus | -87600
kidney transplant | -87600
diabetic kidney disease | -87600
mechanical ventilation (MV) | 0
agitation during percutaneous thrombectomy | 0
rapid deterioration | 24
aspiration pneumonia | 24
septic shock | 24
increasing vasopressors requirements | 24
increasing respiratory support | 24
transthoracic echocardiography | 24
new onset heart systolic murmur | 24
hypertrophic left ventricle | -87600
no other pathological conditions | -87600
dynamic left ventricular outflow tract obstruction (LVOTO) | 24
severe mitral regurgitation (MR) | 24
systolic anterior motion (SAM) of the mitral valve | 24
mean arterial pressure (MAP) of 65 mmHg | 24
norepinephrine 1.8 μg/kg/min | 24
non-fluid responsive | 24
control assisted ventilation | 24
inspired fraction of O2 (FiO2) = 100% | 24
positive end-expiratory pressure (PEEP) of 15 mm Hg | 24
pressure ventilation mode | 24
suboptimal transthoracic window | 24
transesophageal echocardiography (TOE) | 24
hypertrophic septum (17 mm) | 24
hypercontractile status | 24
maximum intraventricular gradient of 165 mm Hg | 24
severe eccentric MR | 24
SAM of anterior and posterior leaflets of the mitral valve | 24
progressive decreasing PEEP from 15 to 5 cm H2O | 24
deterioration in oxygen saturation | 24
pulmonary congestion | 24
volume unresponsiveness | 24
esmolol bolus (500 μg/kg, 4500 μg) | 24
improvement in hemodynamic state | 24
MAP increase from 65 to 85 mm Hg | 24
norepinephrine dose reduction from 1.8 to 0.9 μg/kg/min | 24
oxygen needs maintained | 24
TOE recorded | 24
critical reduction in intraventricular gradient | 24
SAM of the mitral valve reduction | 24
MR improvement | 24
esmolol perfusion started | 24
starting dose of 50 μg/kg/min | 24
TOE-based guidance | 24
norepinephrine reduction to 0.4 μg/kg/min | 24
FiO2 reduction from 100% to 50% | 24
venous oxygen saturation augmentation | 24
lactate levels decrease | 24
hemorrhagic transformation of previous stroke | 288
neurological deterioration | 288
death | 288
