63 years old | 0
female | 0
admitted to the hospital | 0
liver injury | 0
pancytopenia | 0
rheumatoid arthritis | -29184
Steinbrocker radiographic stage IV | -21888
no history of infectious mononucleosis | -29184
no hypersensitivity to mosquito bites | -29184
cervical lymphadenopathy | -3504
axillary lymphadenopathy | -3504
methotrexate | -3504
infliximab | -3504
lymphoproliferative disease | -3504
lymph nodes regressed | -3504
leukocytoclastic vasculitis | -17520
antineutrophil cytoplasmic antibody-negative pauci"immune crescentic glomerulonephritis | -17520
etanercept | -17520
EBV DNA level 940 copies/106 WBC | -17520
anti-EBV VCA IgG positive | -17520
anti-VCA IgM negative | -17520
anti-EBNA antibody negative | -17520
spleen enlargement | -17520
lymphadenopathy | -17520
high-dose corticosteroid treatment | -17520
etanercept discontinued | -17520
clinical findings improved | -17520
abatacept initiated | -10944
exacerbation of rheumatoid arthritis | -10944
prednisolone 4 mg/day | -10944
mild hepatocellular injury | -10944
recurrent fever | -10944
liver injury | -10944
abatacept administered | -10944
persistent liver injury | -10944
pancytopenia developed | -10944
pulse 101 beats/min | 0
blood pressure 103/52 mmHg | 0
body temperature 37°C | 0
respiratory rate 22 breaths/min | 0
oxygen saturation 99% | 0
Eastern Cooperative Oncology Group Performance Status Grade 4 | 0
right upper quadrant tenderness | 0
white blood cell count 2200/μL | 0
hemoglobin 7.6 g/dL | 0
platelet count 61000/μL | 0
aspartate aminotransferase 411 U/L | 0
alanine aminotransferase 425 U/L | 0
alkaline phosphatase 7883 U/L | 0
γ-glutamyl transpeptidase 1223 U/L | 0
total bilirubin 5.0 mg/dL | 0
C-reactive protein 8.97 mg/dL | 0
ferritin 4980 ng/mL | 0
soluble interleukin-2 receptor 4220 U/mL | 0
IgG 456 mg/dL | 0
albumin 2.4 g/dL | 0
prothrombin time INR 1.16 | 0
cytomegalovirus pp65 antigen positive | 0
Aspergillus galactomannan antigen positive | 0
anti-VCA IgG 1:160 | 0
EBV DNA 1200 copies/106 WBC | 0
anti-VCA IgM negative | 0
anti-EBNA antibody negative | 0
antinuclear antibody negative | 0
antimitochondrial M2 antibody negative | 0
anti-hepatitis A virus IgM negative | 0
anti-hepatitis E virus IgA negative | 0
hepatitis B surface antigen negative | 0
anti-hepatitis B surface antibody negative | 0
anti-hepatitis B core antibody negative | 0
hepatitis C virus RNA negative | 0
(1,3)-β-D-glucan negative | 0
no intra- or extrahepatic bile duct dilatation | 0
multifocal low-density liver lesions | 0
splenomegaly | 0
ascites | 0
mediastinal lymphadenopathy | 0
para-aortic lymphadenopathy | 0
hypocellular bone marrow | 0
hemophagocytosis | 0
EBER negative | 0
hemophagocytic lymphohistiocytosis | 0
hepatitis | 0
ferritin elevated | 0
sIL-2R elevated | 0
systemic inflammatory response syndrome | 0
sepsis suspected | 0
meropenem administered | 0
hematopoietic tumors considered | 0
lymphoid tumors considered | 0
supportive therapy | 0
fever | 0
scattered lung nodules | 0
Aspergillus galactomannan positive | 0
CMV pp65 antigen increased | 0
invasive pulmonary aspergillosis suspected | 0
CMV antigenemia suspected | 0
micafungin administered | 0
ganciclovir administered | 0
died | 648
hepatic failure | 648
liver atrophy | 648
bridging fibrosis | 648
zonal necrosis | 648
atypical lymphocyte infiltration | 648
CD3 positive | 648
CD8 positive | 648
TIA1 positive | 648
CD20 negative | 648
CD56 negative | 648
CD79a negative | 648
CD30 negative | 648
EBER positive | 648
CMV negative | 648
histiocytes with hemophagocytosis | 648
spleen infiltration | 648
lymph node infiltration | 648
bone marrow infiltration | 648
Aspergillus hyphae in lung | 648
chronic active EBV T-cell type | 648
systemic form | 648
recurrent fever | 648
persistent fever | 648
hepatitis | 648
splenomegaly | 648
lymphadenopathy | 648
elevated EBV DNA | 648
EBV-infected cytotoxic T-lymphocytes | 648
