57 years old | 0
    male | 0
    admitted to University Hospital | 0
    paraparesis | -2160
    sensory disturbances in both lower extremities | -2160
    fall | -2160
    L3 burst fracture | 0
    spinal canal compression | 0
    posterior lumbar interbody fusion | 0
    paraparesis improved progressively | 0
    no specific symptoms reported | 0
    neuropathic pain | 0
    transferred to rehabilitation hospital | 0
    conservative treatment for neurogenic pain | 0
    gait training | 0
    no specific complication found | 0
    transferred to emergency department | 0
    fever | -168
    general weakness | -168
    leukocytosis | 0
    Klebsiella pneumoniae isolated from blood culture | 0
    Klebsiella pneumoniae isolated from urine culture | 0
    abdominal ultrasonography | 0
    edema in bilateral renal parenchyma | 0
    hyperechogenicity | 0
    renal failure | 0
    acute pyelonephritis | 0
    no local lesion in renal parenchyma | 0
    decreased blood perfusion | 0
    no extension of renal pelvis or renal calyx | 0
    sepsis | 0
    meropenem administered intravenously | 0
    antibiotic treatment for 13 days | 0
    vital signs stable | 0
    laboratory findings returned to normal | 0
    antibiotics stopped on 15th day | 360
    transferred to rehabilitation medicine department | 384
    comprehensive management of CES | 384
    muscular weakness in both lower limbs | 384
    hip flexor 4/4 (right/left) | 384
    knee extensor 3/3 | 384
    ankle dorsiflexor 3/3 | 384
    hallucis extensor 3/3 | 384
    ankle plantar flexor 2/2 | 384
    tingling sensations | 384
    allodynia | 384
    hyperalgesia | 384
    decreased sensations below third lumbar segment | 384
    sitting independently | 384
    standing up independently | 384
    balanced-level walking requiring moderate assistance | 384
    Modified Barthel Index 76 points | 384
    deep tendon reflex decreased in both lower limbs | 384
    no pathological reflex observed | 384
    anal sphincter tone decreased | 384
    bulbocavernosus reflex decreased | 384
    electrodiagnostic study | 384
    normal sensory nerve conduction in both lower limbs | 384
    slow conduction velocity for bilateral peroneal nerves | 384
    slow conduction velocity for bilateral tibial nerves | 384
    decreased amplitude of compound muscle action potential | 384
    H-reflex delayed latency in bilateral tibial nerves | 384
    somatosensory evoked potential stimulating bilateral tibial nerves | 384
    delayed latencies | 384
    bulbocavernosus reflex stimulating pudendal nerves | 384
    delayed latencies | 384
    needle electromyography | 384
    increased insertional activity | 384
    abnormal spontaneous activity in muscles innervated from L2 to S2 | 384
    bilateral lumbosacral polyradiculopathy | 384
    sacral reflex arc lesion | 384
    CES | 384
    indwelling catheter | 384
    self-voiding 100-200 mL | 384
    residual urine volume 200>300 mL | 384
    voiding sense normal | 384
    voiding desire normal | 384
    no incontinence | 384
    no feeling of residual urine | 384
    no hesitancy | 384
    timed intermittent catheterization | 384
    removal of residual urine | 384
    walking independently on even surface | 384
    comprehensive rehabilitative managements | 384
    drug therapy tramadol 150 mg | 384
    drug therapy gabapentin 900 mg | 384
    muscle strengthening exercises | 384
    functional electrical stimulation for bilateral lower limbs | 384
    gait training | 384
    chills | 528
    fever 38.5℃ | 528
    leukocytes 26,110/µL | 528
    hemoglobin 9.3 g/dL | 528
    platelets 168,000/µL | 528
    Creactive protein 34.32 mg/L | 528
    erythrocyte sedimentation rate 120 mm/h | 528
    BUN/creatinine ratio 30.9/1.6 mg/dL | 528
    no other specific finding | 528
    urinalysis specific gravity 1.016 | 528
    urinalysis pH 6.0 | 528
    albumin (2+) | 528
    glucose (3+) | 528
    ketones (-) | 528
    hemoglobin (1+) | 528
    leukocyte (3+) | 528
    nitrate (-) | 528
    red blood cell 1-4/HPF | 528
    white blood cell >5/HPF | 528
    recurrent acute pyelonephritis | 528
    tazobactam administered intravenously | 528
    Klebsiella pneumoniae isolated from blood culture | 528
    Klebsiella pneumoniae isolated from urine culture | 528
    antibiotic changed to meropenem | 528
    sudden left flank pain | 768
    tenderness during voiding | 768
    10×20 cm-sized mass palpated in left abdomen | 768
    blood pressure 100/60 mmHg | 768
    heart rate 115 beats/min | 768
    respiratory rate 20 breaths/min | 768
    axillary temperature 36.5℃ | 768
    leukocytes 28,900/µL | 768
    hemoglobin 7.1 g/dL | 768
    platelets 158,000/µL | 768
    acute hemorrhage suspected | 768
    prothrombin time 13.7 seconds | 768
    international normalized ratio 1.21 | 768
    activated partial thromboplastin time 35.7 seconds | 768
    BUN/creatinine ratio 43.1/3.5 mg/dL | 768
    no other specific finding | 768
    contrast-enhanced abdominal CT | 768
    pyelonephritis with multifocal low-density lesions in left kidney | 768
    perirenal hemorrhage in perinephric space | 768
    active extravasation of contrast media near perinephric space | 768
    hemorrhage in capsular artery outside renal capsule | 768
    retroperitoneal hematoma in left iliac fossa | 768
    systolic blood pressure decreased 90 mmHg | 768
    declined hemoglobin | 768
    emergent transfusion | 768
    angiography performed | 768
    no tumor found | 768
    no vascular malformation found | 768
    coil embolization performed | 768
    suspicion of progressive hemorrhage in left capsular artery | 768
    transferred to intensive care unit | 768
    conservative treatment for acute renal failure | 768
    acute pyelonephritis | 768
    follow-up abdominal CT | 768
    no active bleeding observed | 768
    embolized capsular artery around anterior cortex of left kidney | 768
    acute pyelonephritis at embolized site | 768
    hemorrhage stopped | 768
    nephrectomy not considered | 768
    surgical hematoma removal | 768
    persistent abdominal pains | 768
    voiding cystourethrography | 768
    no vesicoureteral reflux observed | 768
    failed to void after filling 450 mL contrast medium | 768
    urodynamic study | 768
    strong voiding desire when infused with 500 mL saline | 768
    failed to void due to detrusor areflexia | 768
    oral medications alpha blocker | 768
    oral medications choline agonist | 768
    intermittent self-catheterization five times per day | 768
    urinary retention >500 mL | 768
    no additional UTIs | 768
    no other complications | 768
    transferred to rehabilitation hospital | 768
    <|eot_id|>
    