77 years old | 0  
male | 0  
transferred from a rural hospital | 0  
left iliac fossa pain | -72  
diarrhoea | -72  
nausea | -72  
vomiting | -72  
fevers | -72  
advanced prostate cancer | 0  
bony metastasis | 0  
previous chemotherapy | 0  
previous radiotherapy | 0  
type two diabetes mellitus requiring insulin | 0  
regular abiraterone | 0  
regular prednisolone | 0  
regular flutamide | 0  
regular oxycodone | 0  
regular targin | 0  
sinus tachycardia | 0  
elevated temperature | 0  
diffuse tenderness | 0  
left iliac fossa tenderness | 0  
positive bowel sounds | 0  
low haemoglobin | 0  
low white cell count | 0  
normal coagulation | 0  
normal liver function | 0  
normal lipase | 0  
normal lactate | 0  
grossly thickened small bowel | 0  
portal venous gas in liver | 0  
no peritoneal signs | 0  
conservative treatment | 0  
admitted to Intensive Care | 0  
fluid resuscitation | 0  
intravenous tazocin | 0  
granulocyte-colony stimulating factor | 0  
nasogastric decompression | 0  
no source of infection found | 0  
rising C-reactive protein | 0  
clinical condition deterioration | 0  
exploratory laparotomy performed | 0  
moderate bowel oedema | 0  
no bowel necrosis | 0  
no mesenteric necrosis | 0  
division of adhesions of the jejunum | 0  
division of adhesions of the ileum | 0  
chemotherapy/radiotherapy-related severe enterocolitis | 0  
adhesions | 0  
conservatively managed small bowel obstruction | 0  
transferred back to rural hospital | 648  

    