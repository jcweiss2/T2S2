75 years old | 0
male | 0
Japanese | 0
admitted to the hospital | 0
necrotizing pancreatitis | 0
smoked 40 cigarettes per day for 50 years | -36000
old anterior myocardial infarction | -36000
treated with antibiotics | 0
endoscopic catheter drainage of pancreatic necrosis | 0
bradycardia | 192
dyspnea | 192
body temperature of 38.2°C | 192
blood pressure of 74/52 mmHg | 192
pulse rate of 50 beats per minute | 192
oxygen saturation of 91% on 5 L/min oxygen | 192
elevated white blood cell count | 192
elevated C-reactive protein level | 192
elevated presepsin level | 192
sepsis | 192
elevated fibrin degradation products | 192
high prothrombin time-international normalized ratio | 192
low AT activity | 192
coagulation disorder | 192
new-onset ST elevation in inferior leads | 192
complete atrioventricular block | 192
reduced left ventricular ejection fraction of 25% | 192
local hypokinesia in the inferior wall | 192
local dyskinesia in the anterior wall | 192
acute inferior and old anterior myocardial infarction | 192
cardiogenic-septic shock | 192
septic disseminated intravascular coagulation (DIC) | 192
inserted an intra-aortic balloon pump (IABP) | 192
inserted a temporary pacemaker | 192
coronary angiography | 192
sub-occlusion of the proximal right coronary artery (RCA) | 192
dual antiplatelet agents | 192
bolus of 8,000 units of UFH | 192
intravascular ultrasound (IVUS) | 192
hypoechoic plaque with deep ultrasound attenuation | 192
vulnerable plaque at the culprit lesion without visible thrombus | 192
3.0-mm balloon dilatation | 192
thrombolysis in myocardial infarction grade 3 flow | 192
culprit lesion reoccluded | 194
fresh thrombi | 194
activated clotting time (ACT) was insufficient | 194
heparin resistance (HR) | 194
acquired AT deficiency | 194
administered 2,400 units of AT gamma | 194
additional 5,000 units of UFH | 194
ACT increased to 364 seconds | 194
intravascular thrombi decreased | 194
occluded lesion recanalized | 194
implanted a drug-eluting stent | 194
completed PCI without subsequent thrombus formation | 194
plasma AT activity increased to 74% | 196
platelet count did not decrease after PCI | 196
heparin/platelet factor 4 antibody was not detected | 196
IABP and temporary pacemaker removed | 216
died due to sepsis | 1080