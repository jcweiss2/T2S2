34 years old | 0
female | 0
admitted to the hospital | 0
septicemia | 0
superficial inflammation of the left thigh | 0
swelling of the left thigh | -48
chronic pain in the sacro-iliac joint | -336
oral antibiotic therapy | -48
cefuroxime | -48
temperature 39.4°C | -24
increased inflammation parameters | 0
leukocytes 16.000/µL | 0
c-reactive protein 35 mg/dL | 0
spreading inflammation of the soft tissue | 0
i.v. drug abuse | -672
heroin | -672
hepatitis C | -672
computed tomography scan | 0
abscess of the sacro-iliac joint | 0
abscess of the psoas muscle | 0
magnetic resonance imaging | 0
necrotising fasciitis of the left thigh | 0
radical surgical debridement | 0
fasciectomy of the left thigh | 0
abscess of the sacro-iliac joint opened and drained | 0
antibiotic therapy | 0
tobramycin | 0
ceftriaxone | 0
metronidazole | 0
infection with multi-resistant Pseudomonas aeruginosa | 0
infection with Vancomycin-resistant Enterococcus faecalis | 0
planned second revision with surgical debridement | 48
clean wound | 48
no fasciitis progression | 48
infection in the elbow | 48
open surgical debridement | 48
cerebral septic complications | 48
pulmonary septic complications | 48
non-operative treatment | 48
five further sequential operations | 72
continuous vacuum therapy | 72
split skin graft | 168
intermittent hemodiafiltration | 72
septic acute renal failure | 72
Pseudomonas aeruginosa pneumonia | 72
antibiotics | 72
ceftazidime | 72
tracheotomy | 168
spontaneous breathing | 168
erythrocyte concentrates | 168
thrombocyte concentrates | 168
fresh frozen plasma | 168
prothrombin concentrate | 168
critical-illness polyneuropathy | 720
intensive physiotherapy | 720
discharged | 1440
referred to a speciality rehabilitation center | 1440