67 years old | 0
male | 0
admitted to the hospital | 0
left leg swelling | -168
cactus plant injury | -168
Primary Sclerosing Cholangitis | 0
mild Ulcerative Colitis | 0
deranged liver function tests | 0
presentation to ED | 0
left leg swelling from a recent cactus plant prick | 0
Blood Pressure (BP): 71/41mmHg | 0
Mean Arterial Pressure (MAP): 48mmHg | 0
Respiratory Rate: 36 breaths per minute | 0
Heart Rate (HR): 125 beats per minute | 0
sinus tachycardia | 0
Temperature: 39°C | 0
Oxygen Saturation: 86% with 0.21 FiO2 | 0
admitted to the intensive care unit (ICU) | 0
pH 7.15 | 0
PO2 84 | 0
HCO3 15 | 0
Lactate 7.6 | 0
Sodium (Na) 134 | 0
Urea 7.6 | 0
Creatinine (sCr) 173 | 0
eGFR 27 | 0
White Cell Count (WCC) 13.8 | 0
C-reactive protein (CRP) 22 | 0
Hemoglobin (Hb) 114 | 0
Platelet (Plt) 81 | 0
Liver Function Test (LFT)- Total Bilirubin (Bili) 99 | 0
Alanine transaminase (ALT) 61 | 0
Aspartate aminotransferase (AST) 83 | 0
Alkaline Phosphatase (ALP) 96 | 0
Triple vasopressor support initiated | 0
Noradrenaline 20mcg/min | 0
Adrenaline 20mcg/min | 0
Vasopressin 0.04units/min | 0
Antibiotics: Piperacillin-Tazobactam IV 4.5g | 0
Meropenem IV 2g | 0
Lincomycin IV 600mg | 0
Vancomycin IV 2g | 0
Emergency left lower limb fasciotomy | 0
debridement | 0
below knee amputation | 0
necrotizing fasciitis | 0
LRINEC Score of 5 | 0
extensive left foot and below knee tissue necrosis | 0
dishwasher fluid | 0
liquefied fat | 0
unviable skin and muscle | 0
Histopathology | 0
post operatively | 24
transferred to ICU | 24
intubated | 24
possible re-exploration | 24
oliguria | 24
blood gas showed severe acidosis | 24
left internal jugular vascath insertion | 24
continuous renal replacement therapy (CRRT) | 24
pH 7.28 | 24
Lactate 4.7 | 24
Na 130 | 24
sCr 206 | 24
Hb 89 | 24
Plt 105 | 24
WCC 17 | 24
CRP 78 | 24
International normalized ratio (INR) 2.2 | 24
Activated Partial Thromboplastin Time (APTT) 150 | 24
Initial blood cultures (BCs) isolated Group B Streptococcus pneumoniae (GBSPn) | 24
Ventilation sedation: Propofol 170mg/hr | 24
Fentanyl 40mcg/hr | 24
CRRT (Day 1) on heparin circuit | 24
Renal dose - 30ml/kg/hr | 24
Triple vasopressor support continued | 24
Noradrenaline 23mcg/min | 24
Adrenaline 18mcg/min | 24
Vasopressin 0.04units/min | 24
Antibiotics (MLV): Meropenem IV 2g | 24
Lincomycin IV 600mg | 24
Vancomycin IV 2g | 24
Intravenous Immunoglobin G (IVIgG) therapy 100g | 24
taken back to theatre | 48
confirm source control | 48
viability of the left stump | 48
no evidence of necrotic tissue | 48
Rapid Atrial Fibrillation (RAF) | 48
HR 110bpm | 48
oliguric | 48
pH 7.40 | 48
Lactate 3.9 | 48
Na 131 | 48
sCr 116 | 48
WCC 26 | 48
CRP 105 | 48
Procalcitonin (PCT) 21.18 μg/L | 48
Hb 83 | 48
Plt 63 | 48
INR 3.1 | 48
Fibrinogen 2.4 | 48
Echocardiography: Moderate segmental left ventricular dysfunction | 48
Ejection Fraction 40-45% | 48
Dilated atria bilaterally | 48
Raised Right Atrial Pressure | 48
Amiodarone loading dose 300mg | 48
maintenance dose 900mg | 48
Antibiotics remained unchanged (MLV) | 48
CRRT (Day 2) – AN69 anti-inflammatory heparin laden adsorbing filter | 48
Citrate based anticoagulation circuit | 48
Sepsis Induced Coagulopathy (ISTH -SIC criteria) | 72
bedside surgical debridement | 72
pH 7.31 | 72
Lactate 2.4 | 72
Na 135 | 72
sCr 79 | 72
WCC 27 | 72
CRP 127 | 72
Hb 78 | 72
Plt 50 | 72
INR 2.0 | 72
Histopathology consistent with NF | 72
Wound culture for microscopy culture and sensitivity (MCS) had medium growth of GBSPn | 72
Tissue culture (intraoperatively) had medium growth of GBSPn | 72
Vasopressor support - weaning | 72
Noradrenaline 20mcg/min | 72
Adrenaline weaned off | 72
Vasopressin 2.4units/min | 72
Antibiotics remained unchanged (MLV) | 72
CRRT (Day 3) - ongoing | 72
oliguric | 96
pH 7.36 | 96
Lactate 1.5 | 96
Na 130 | 96
sCr 116 | 96
WCC 33 | 96
CRP 103 | 96
PCT 15.37 | 96
Hb 91 | 96
Plt 53 | 96
INR 1.7 | 96
LFT - Bili 131 | 96
AST 127 | 96
ALP 121 | 96
Double inotropic support | 96
Noradrenaline 20mcg/min | 96
Vasopressin 2.4units/min | 96
Antibiotics remained unchanged (MLV) | 96
CRRT (Day 4) | 96
Amiodarone infusion | 96
fulminant hepatic failure/ encephalopathy | 120
Refractory oliguria | 120
pH 7.39 | 120
Lactate 1.2 | 120
Na 134 | 120
sCr 124 | 120
WCC 39.5 | 120
CRP 74 | 120
Hb 116 | 120
Plt 49 | 120
INR 1.5 | 120
LFT- Bili 139 | 120
AST 69 | 120
ALT 97 | 120
ALP 140 | 120
Dual inotropic support | 120
Noradrenaline 20mcg/min | 120
Vasopressin weaned off | 120
Antibiotics remained unchanged (MLV) | 120
CRRT (Day 5) | 120
severely deconditioned | 144
ICU acquired weakness | 144
unarousable | 144
no response to noxious stimuli | 144
Remained intubated and ventilated | 144
Pressure Support Ventilation | 144
Refractory oliguria | 144
PH 7.44 | 144
Lactate 1.1 | 144
WCC 43.5 | 144
CRP 109 | 144
Hb 90 | 144
Plt 57 | 144
INR 1.5 | 144
LFT - Bili 150 | 144
AST 95 | 144
ALP 154 | 144
Sedation weaned off | 144
Off vasopressor | 144
Noradrenaline weaned off | 144
Antibiotic de-escalation | 144
Lincomycin and Vancomycin ceased | 144
Meropenem IV 2g | 144
CRRT (Day 6) | 144
Hyper-Ammonium Therapy initiated | 144
Rifaximin NGT 550mg | 144
Lactulose NGT 20ml | 144
2 units of PRBCs transfusion | 144
jaundice | 168
Hypoactive delirium | 168
RASS -5 | 168
new onset lateralizing signs | 168
CT Brain: No acute intracranial pathology | 168
Ultrasound abdomen: Acute Calculous Cholecystitis | 168
pH 7.44 | 168
Lactate 1.1 | 168
WCC 44.3 | 168
CRP 109 | 168
Hb 129 | 168
Plt 66 | 168
INR 1.3 | 168
LFT - Bili 235 | 168
AST 75 | 168
ALP 175 | 168
Conjugated Bilirubin 142 | 168
Meropenem IV 2g | 168
CRRT (Day 7) | 168
Anuria | 192
Hypotensive BP 71/33 | 192
MAP 51mmHg | 192
Febrile 39°C | 192
RAF HR 160 | 192
Significant deterioration | 192
commenced on palliative care pathway | 192
deceased shortly post treatment withdrawal | 192
Troponin 616 | 192
Ammonia 158 | 192
LFT - Bili 352 | 192
AST 100 | 192
ALP 299 | 192
CRRT (Day 8) | 192
Renal recovery assessment | 192
challenged with combination of Furosemide IV 250mg and Acetazolamide IV 500mg | 192
Recommenced Vasopressor support | 192
Noradrenaline 2.5mcg/min | 192
Antibiotic regimen: Lincomycin IV 600mg | 192
Meropenem IV 2g | 192
Digoxin IV 500mcg | 192
Metoprolol IV 15mg | 192