80 years old | 0
female | 0
admitted to the hospital | 0
Rathke’s cleft cyst | -720
bilateral reduction in visual acuity | -720
bitemporal hemianopsia | -720
mild bifrontal headache | -720
endoscopic surgery | -720
cyst fenestration | -720
partial cyst wall resection | -720
pedicled nasoseptal flap technique | -720
visual disturbances recovery | -720
recurrence of visual disturbance | -336
bifrontal headaches | -336
anisocoric pupils | -336
fixed mydriasis in the left eye | -336
bitemporal hemianopsia | -336
new endoscopic transnasal transsphenoidal surgery | -336
gross total resection | -336
CSF leak | -336
resurface of the skull base with a nasoseptal flap | -336
postoperative sellar MRI | -336
“reservoir sign” | -336
conservative approach with head elevation | -336
neuro check | -336
stable condition | -288
subtle paraparesis | -192
paraplegia | -168
dorsal spine MRI | -168
T3-T4 intramedullary lesion | -168
emergency thoracic laminectomy | -168
SDAVF | -168
intramedullary hematoma | -168
feeder artery on the right T3 dural sleeve | -168
arterial supply interruption | -168
coagulation of the epidural arteries | -168
vessels draining the dural fistula | -168
huge dilated tortuous spinal vein | -168
draining vein-like varix | -168
thrombosed | -168
shunting point coagulated and divided | -168
intramedullary hematoma evacuation | -168
hematomyelia | -168
neurogenic shock | -144
high doses of norepinephrine | -144
intensive care unit | -144
no signs of CSF rhinorrhea | -144
progressive worsening of neurogenic shock | -96
septic shock | -96
pneumonia | -96
higher doses of vasoactive amines | -96
mean arterial pressure | -96
hypoxic encephalopathy | -48
brain death | -48
brain CT | -48
diffuse white matter hypodensity | 0 
discharge | 240