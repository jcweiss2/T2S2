shortness of breath | -96
fever | -96
dry cough | -96
fatigue | -96
reduced breath sounds in the lower segments of the lungs | 0
oxygen saturation 93% | 0
bilateral peripheral ground-glass attenuation and patchy consolidation on chest CT | 0
nasopharyngeal SARS-CoV-2 RT-PCR test positive | 0
increased temperature | 21
saturation with free breathing decreased to 90% | 21
white cell count 7.93 х 109/ L | 21
hemoglobin 159 g/l | 21
platelet count 468 х 109/l | 21
Westergren ESR 41 mm/h | 21
interleukine 6 102 pg/ml | 21
С-reactive protein 142 mg/l | 21
ferritin 939.92 μg/ml | 21
D-dimer 609 ng/ml | 21
procalcitonin 0.11 ng/ml | 21
treatment with dexamethason | 0
treatment with heparin | 0
treatment with tocilizumab | 0
treatment with acetylcysteine | 0
treatment with pantoprazole | 0
treatment with nadroparin calcium | 0
oxygen supplementation | 0
air and pleural effusion in the right pleural cavity | 360
thoracentesis | 360
thoracostomy | 360
evacuation of 1400 ml of yellowish opaque liquid | 360
linezolid therapy | 360
imipenem/cilastatin therapy | 360
oxygen supplementation with flow rate of 8-10 l/min | 360
daily drainage volume 300-1000 ml | 384
pleural effusion with gas bubbles on chest CT | 432
focal area of subpleural infiltration with a central cavity of destruction | 432
air layer along the anterior chest wall | 432
radiological signs of left side hydropneumothorax | 432
pleural fluid analysis | 432
exudative lymphocytic-rich effusion | 432
growth of Acinetobacter baumannii and Pseudomonas aeruginosa | 432
urine culture positive for Klebsiella pneumonia | 432
needle thoracocentesis | 504
new pleural drainage | 504
air and creamy purulent mass aspirated | 504
serofibrinous hemorrhagic fluid drawn | 504
diagnosis of pleural empyema | 504
transfer to Surgical Department | 504
irrigation of right pleural space with antiseptic solutions | 504
lung expansion by continuous vacuum aspiration | 504
encapsulated pleural effusion | 576
ultrasound-guided puncture | 576
new drainage of pleural cavity | 576
antibiotic therapy with colistimethatum natrium and imipenem/cilastatin | 672
discharge from hospital | 1008
oxygen saturation 97% | 1008
chest CT after chest tube removing | 1008
normal lab test scores | 1008
С-reactive protein 11.7 mg/l | 1008
procalcitonin < 0.1 ng/ml | 1008
negative nasopharyngeal SARS-CoV-2 RT-PCR test | 504