64 years old | 0
male | 0
admitted to the hospital | 0
general weakness | -168
myalgia | -168
abdomal pain | -168
thrombosis of the SMV | -168
fever | -168
headache | -168
CT scan | -168
thrombus in SMV | -168
fat stranding | -168
bowel wall edema | -168
metformin | -12000
glimepiride | -12000
linagliptin | -12000
losartan | -12000
rosuvastatin | -12000
dull pressing pain | 0
mild tenderness | 0
hypo-active bowel sound | 0
white blood cell count 16160 /mL | 0
ESR 86 mm/hr | 0
HS-CRP 16 mg/dL | 0
influenza test | 0
influenza B positive | 0
COVID-19 test | 0
COVID-19 negative | 0
peramivir | 0
low molecular weight heparin | 0
total parenteral nutrition | 0
ceftriaxone | 0
fever | 0
abdominal pain | 0
abdominal discomfort | 48
follow-up CT scan | 192
thrombus size decreased | 192
rivaroxaban | 216
soft diet | 216
transferred to general ward | 240
follow-up CT scan | 360
thrombus markedly reduced | 360
discharged | 384
outpatient follow-up | 720
CT scan | 720
SMV thrombosis not seen | 720