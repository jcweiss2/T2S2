59 years old | 0
male | 0
radical cystoprostatectomy | -12
ileal neobladder reconstruction | -12
G2pT2 bladder cancer | -12
urinary incontinence | -9
urodynamics | -9
small capacity neobladder | -9
high pressures | -9
neobladder augmentation cystoplasty | -12
polycystic kidney disease | 0
urinary tract infection | 0
dyspnea at rest | 0
right loin pain | 0
cachectic | 0
dry mucous membranes | 0
tachypnea | 0
tachycardia | 0
hypotension | 0
leucocytosis | 0
mildly raised C-Reactive Protein | 0
mild hypokalaemia | 0
elevated creatinine | 0
elevated urea | 0
uncompensated metabolic acidosis | 0
normal anion gap | 0
microscopic haematuria | 0
sterile pyuria | 0
sinus tachycardia | 0
confused | 48
lethargic | 48
increasing respiratory distress | 48
worsening hyperchloremic metabolic acidosis | 48
unresponsive | 48
Glasgow Coma Score of 8/15 | 48
sodium bicarbonate 8.4% infusion | 48
regained consciousness | 52
improving metabolic acidosis | 52
discharged with oral sodium bicarbonate | 72
neo-bladder excision | 72
ileal conduit formation | 72
no further episodes of metabolic acidosis | 8760