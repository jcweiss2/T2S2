80 years old | 0
    arterial hypertension | -8640
    dyslipidemia | -8640
    type 2 diabetes mellitus | -8640
    ischemic cardiomyopathy | -8640
    preserved ejection fraction | -8640
    chronic hepatitis B virus infection | -8640
    progressive fatigue | -2160
    malaise | -2160
    anorexia | -2160
    cough | -840
    blood-streaked sputum | -840
    progressive peripheral edema | -840
    denied fever | -840
    denied weight loss | -840
    denied arthralgia | -840
    denied skin rash | -840
    multifocal pneumonia | 0
    acute kidney injury | 0
    serum creatinine 5.69 mg/dL | 0
    baseline serum creatinine 0.99 mg/dL | 0
    iron deficiency anemia | 0
    hemoglobin 7.6 g/dL | 0
    admitted to intensive care unit | 0
    intravenous fluid administration | 0
    empiric amoxicillin-clavulanate | 0
    azithromycin | 0
    switched to piperacillin-tazobactam | 24
    elevated erythrocyte sedimentation rate | 0
    negative ANCA | 0
    negative anti-GBM antibodies | 0
    negative antistreptolysin O antibodies | 0
    normal C3 levels | 0
    normal C4 levels | 0
    chronic HBV infection | 0
    negative anti-HCV | 0
    negative HIV | 0
    microscopic hematuria | 0
    subnephrotic proteinuria | 0
    chest CT bilateral nodular infiltrates | 0
    abdomen CT normal kidneys | 0
    hemoptysis | 24
    bronchoscopy | 24
    bronchoalveolar lavage | 24
    bacterial infection excluded | 24
    mycobacterial infection excluded | 24
    fungal infection excluded | 24
    cytologic analysis alveolar macrophages | 24
    polymorphonuclear cells predominance | 24
    no hemosiderin-laden macrophages | 24
    transferred to our hospital | 72
    pale | 72
    afebrile | 72
    blood pressure 130/70 mm Hg | 72
    pulse rate 87 beats/min | 72
    tachypneic | 72
    oxygen saturation 94% | 72
    chest crackles | 72
    peripheral edema | 72
    no skin rash | 72
    hemoglobin 8 g/dL | 72
    white blood cell count 13.2 × 109/L | 72
    C-reactive protein 79.8 mg/L | 72
    ESR 66 mm/h | 72
    serum creatinine 7.3 mg/dL | 72
    blood urea nitrogen 197 mg/dL | 72
    HBV viral load 337,600 IU/mL | 72
    normal platelet count | 72
    normal coagulation tests | 72
    normal bilirubin | 72
    normal aspartate aminotransferase | 72
    normal alanine aminotransferase | 72
    normal albumin | 72
    normal total serum protein | 72
    no monoclonal peak | 72
    urinalysis 25-50 RBC/hpf | 72
    urinary protein 1.46 g/24h | 72
    chest X-ray diffuse infiltrates | 72
    MPO?ANCA 121.1 U/mL | 24
    PR3?ANCA 312.6 U/mL | 24
    anti-GBM antibody 202 U | 24
    rheumatoid factor 26 IU/mL | 24
    normal C3 | 24
    normal C4 | 24
    negative ANA | 24
    negative cryoglobulins | 24
    negative anti-dsDNA | 24
    IV methylprednisolone | 24
    oral prednisolone | 24
    cyclophosphamide | 24
    plasma exchange | 24
    entecavir | 24
    renal biopsy | 144
    cellular crescents | 144
    focal fibrinoid necrosis | 144
    interstitial fibrosis | 144
    inflammatory infiltrate | 144
    linear IgG deposition | 144
    resolution of hypoxemia | 408
    no cough recurrence | 408
    no blood-streaked sputum | 408
    chest CT resolution | 480
    discharged | 816
    entecavir therapy | 816
    undetectable HBV viral load | 2448
    normal liver ultrasound | 2448
    dialysis-dependent | 2448
    no DAH relapse | 17544
    ANCA negative | 17544
    anti-GBM negative | 17544
    