71 years old | 0
female | 0
admitted to the hospital | 0
unconscious state | 0
history of hypertension | -720
history of ischaemic heart disease | -720
history of peripheral vascular disease | -720
stroke | 0
head computed tomographic scan | 0
inotropic support | 24
septic shock | 24
elevated levels of inflammatory markers | 24
erythrocyte sedimentation rate | 24
C-reactive protein | 24
blood obtained | 24
yeast in both aerobic and anaerobic BacT/ALERT culture bottles | 24
caspofungin administered | 24
died | 72
yeast isolate identified as C. parapsilosis | 24
VITEK 2 yeast identification system | 24
referred to the Mycology Reference Laboratory | 24
CHROMagar Candida | 48
turquoise blue colonies | 48
acetate ascospore agar | 48
long ellipsoidal-shaped ascospores | 48
internally transcribed spacer region of ribosomal DNA amplified and sequenced | 48
DNA sequence data comparisons | 48
Lodderomyces elongisporus type strain | 48
Candida parapsilosis strain | 48
antifungal susceptibility determined | 48
Etest | 48
RPMI 1640 medium | 48
MIC values | 48
amphotericin B | 48
fluconazole | 48
voriconazole | 48
posaconazole | 48
itraconazole | 48
flucytosine | 48
caspofungin | 48
micafungin | 48
hospitalized earlier for lower limb ischaemia | -336
discharged 2 weeks before the current episode | -336
no apparent risk factors | 0
history of heart disease | -720
stroke | 0
no antibiotics | 0
no central lines | 0
inoculation of the yeast from the skin | -72
translocation from the gastrointestinal tract | -72
fungaemia | 24
Lodderomyces elongisporus | 24
bloodstream pathogen | 24
virulence attributes | 24
environmental niche | 24
global prevalence | 24
Mexico | 24
Malaysia | 24
China | 24
Australia | 24
Middle East | 24
Japan | 24
Spain | 24
Korea | 24
endocarditis | 24
diverse clinical conditions | 24
caspofungin before cardiac surgery | 24
amphotericin B plus flucytosine | 24
voriconazole | 24
survived | 72
fluconazole | 24
died | 72
micafungin | 24
survived | 72
caspofungin | 24
died | 72
antifungal therapy | 24
echinocandins | 24
caspofungin | 24
micafungin | 24
antifungal susceptibility | 24
C. parapsilosis complex | 24
reduced susceptibility to echinocandins | 24
Infectious Disease Society of America guidelines | 24
therapeutic use of echinocandins | 24
candidaemia | 24
C. parapsilosis | 24
uncommon yeast pathogens | 24
misidentified | 24
VITEK 2 | 24
C. parapsilosis complex | 24
C. orthopsilosis | 24
C. metapsilosis | 24
L. elongisporus | 24
multiplex PCR assay | 24
Mycology Reference Laboratory | 24
culture collection | 24
sputum of a cancer patient | 24
catheter tip of a patient with fungaemia | 24
bloodstream of a cancer patient | 24
matrix-assisted laser desorption/ionization time-of-flight mass spectrometry | 24
rare yeast species | 24
reduced susceptibility | 24
antifungal agents | 24
prolonged survival of seriously ill patients | 24
intensive care units | 24
broad-spectrum antibiotics | 24
life support systems | 24
intravascular catheters | 24
prophylactic and therapeutic use of antifungal agents | 24
selection pressure | 24
increased colonization | 24
invasive infection | 24
delay in accurate identification | 24
lack of experience | 24
diagnostic and therapeutic challenges | 24
higher mortality rates | 24