30 years old | 0
G1P0 | 0
Hispanic female | 0
presented at 15 weeks gestation | 0
primary complaint of 5-day history of acute, progressive right lower and right upper quadrant abdominal pain | -120
abdominal pain associated with dysuria, nausea and vomiting | -120
emesis progressed to complete oral intolerance for the 12 h preceding presentation | -12
emergency department presentation 3 days prior | -72
diagnosed as acute ‘hyperemesis gravidarum’ | -72
obstetrical ultrasound reported ‘single living intrauterine pregnancy with an estimated gestation age of 13 weeks, 6 ± 8 days’ | -72
fetal heart tones (FHTs) measured 160 bpm | -72
orally challenged successfully | -72
discharged home with oral antibiotics and antiemetics | -72
re-presentation | 0
abdominal pain was reported in the right lower, right upper and left lower quadrants | 0
moderate tenderness to palpation was documented in the right lower quadrant | 0
white blood cell count had increased to 16 200 | 0
ultrasound imaging revealed only ‘dilated fluid filled bowel’ | 0
FHTs were reported at 160 bpm | 0
acute gestational appendicitis was diagnosed | 0
general surgery consultation was requested | 0
clinical diagnosis confirmed | 0
laparoscopic abdominal access was achieved | 0
massive bowel distention and purulent ascites | 0
conversion from laparoscopy to open laparotomy | 0
abscess was discovered that had enveloped the ileocecum | 0
perforation of the appendiceal base with extension into the cecum was readily apparent | 0
cecal necrosis | 0
ileocecectomy was performed | 0
abdomen was irrigated | 0
attempted fascial closure was abandoned | 0
abdominal wall tension secondary to pronounced bowel edema | 0
ACS was diagnosed | 0
abdomen was left open | 0
temporary closure was performed | 0
intubated and transferred to the intensive care unit (ICU) | 0
intravenous antibiotics and resuscitation fluids were provided | 0
consultations were obtained with infectious disease | 0
consultations were obtained with the patient's obstetrician | 0
daily FHTs were determined at bedside by the obstetrician | 0
negative pressure therapy was maintained | 0
peritoneal toilet with inspection of the ileocolic anastomosis was performed on post-operative day 4 | 96
complete integrity of the ileocolic anastomosis | 96
no evidence of bowel necrosis was appreciated | 96
significant bowel edema was noted | 96
temporary abdominal closure was achieved | 96
fascial closure was achieved on post-operative day 6 | 144
skin closure was deferred using a Wound VAC | 144
extubated in the ICU | 144
delayed primary closure of the laparotomy incision was performed on post-operative day 12 | 288
progressed to a regular diet without complications | 288
pathology returned a diagnosis of ‘acute ruptured appendicitis with associated abscess formation and acute serositis’ | 288
discharged home on post-operative day 15 | 360
tocolysis was not indicated | 0
tocolysis was deferred throughout her admission | 0
eventual normal spontaneous vaginal delivery was achieved | 7200
mother reports no incisional hernia development at 5 years following surgery | 26280
daughter has obtained all developmental milestones | 26280
daughter has developed only common childhood illnesses | 26280