Here is the extracted table of events and timestamps:

29 years old | 0
male | 0
admitted to the hospital | 0
muscle and joint pain | -144
general weakness | -144
fever | -144
39°C | -144
pronounced liver dysfunction | -144
total bilirubin 5.7 mg/dl | -144
serum glutamic oxaloacetic transaminase 633 U/L | -144
serum glutamic pyruvate transaminase 412 U/L | -144
gamma-glutamyl transferase 161 U/L | -144
lactate dehydrogenase 1668 U/L | -144
C-reactive protein (CRP) 519 mg/l | -144
procalcitonin 1.28 ng/ml | -144
increased leukocyte levels | -144
massive bilateral pneumonia | -144
intubation | -144
mechanical ventilation | -144
FiO2 100% | -144
SpO2 88.7% | -144
norepinephrine 0.6 μg/kg/min | -144
meropenem 1 g every 8 h IV | -144
azithromycin 500 mg once daily IV | -144
oseltamivir 75 mg, every 12 h p.o. | -144
methylprednisolone 80 mg every 12 h IV | -144
stress ulcer prophylaxis | -144
thromboprophylaxis (UFH) | -144
CRRT started | -168
CytoSorb application | -168
norepinephrine requirements lowered | -168
CRP decreased | -168
leukocyte levels normalized | -168
ventilation parameters improved | -168
lung function improved | -168
ICU delirium | -168
antipsychotics | -168
percutaneous tracheostomy | -168
recovery | -168
transferred to general ward | -168
transferred to rehabilitation clinic | -168
influenza A (H1N1) | -168
dual antibiotic therapy | -168
antiviral therapy | -168
corticosteroids | -168
lung-protective ventilation | -168
prone position | -168
CRRT (Fresenius Medical Care, multiFiltrate) | -168
CVVHDF mode | -168
second CytoSorb application | -168
norepinephrine requirements decreased | -168
CRP levels decreased | -168
leukocyte levels normalized | -168
ventilation parameters improved | -168
lung function improved | -168
vasopressors discontinued | -168
vasopressin not available | -168