64 years old| 0
woman| 0
bipolar depression| 0
diabetes| 0
migraine headaches| 0
known seizure disorder| 0
found unresponsive in a non-air-conditioned room| -2
ambient temperature outside in excess of 90°F (33°C)| -2
home medications include amitriptyline 175 mg daily| -672
cyclobenzaprine 10 mg daily| -672
lurasidone 80 mg daily| -672
benztropine 1 mg three times a day| -672
topiramate extended release 100 mg daily| -672
clonazepam 0.5 mg daily| -672
trazodone 100 mg daily| -672
sitagliptin 25 mg daily| -672
erenumab 70 mg injected monthly| -672
Emergency medical service called| -2
febrile on initial evaluation| -2
cool compresses applied| -2
transported to the hospital| -2
hypotensive (blood pressure 84/42)| 0
febrile with a rectal temperature of 42°C| 0
skin warm and dry| 0
mucous membranes dry| 0
remainder of exam normal| 0
neurological examination responsive only to painful stimuli| 0
no focal neurological deficits| 0
no hyperreflexia| 0
no rigidity| 0
leucocytosis (11,400)| 0
creatine phosphokinase normal| 0
EKG normal| 0
admitted to intensive care unit (ICU)| 0
started on vancomycin and cefepime| 0
blood cultures grew Staphylococcus hominis| 24
core body temperature decreased to less than 38°C| 48
mentation returned to baseline| 48
transferred to medical floor| 48
treated for Staph hominis bacteraemia with 7-day course of vancomycin| 48
discontinue use of cyclobenzaprine on discharge| 168
quick recovery| 168
lack of neurological findings (rigidity, tremors)| 168
severe NEHT with associated bacteraemia determined as cause| 168
initially thought to be severely septic| 0
started on broad spectrum antibiotics| 0
concern for drug-drug interactions| 0
serotonin syndrome considered| 0
low suspicion for serotonin syndrome| 0
blood cultures obtained| 0
toxicology consulted| 0
blood cultures positive for S. hominis| 24
toxicology’s assessment stated NEHT precipitated by multiple anticholinergic medications| 24
mentation improved to baseline| 24
revealed feeling overheated and fatigued for past 2 weeks| -336
no medication changes in past 2 weeks| -336
primary care physician advised to continue current medication regimen| 168
discontinued cyclobenzaprine per toxicology’s recommendation| 168
encouraged to discuss weaning medications| 168
educated about risks of polypharmacy| 168
combination of anticholinergic medications increased susceptibility to NEHT| 0
amitriptyline, trazodone, cyclobenzaprine, benztropine inhibited sweating| 0
topiramate caused hypohydrosis| 0
NEHT diagnosed earlier if core temperature remained elevated| 0
high risk for hyperthermia| 0
high dosage medications may increase risk| 0
Anticholinergic Risk Scale score 9| 0
Naranjo Scale score 4 (possible adverse drug reaction)| 0
counselling on risks of NEHT| 168
medicine reconciliation periodically| 168
vulnerability of patients with psychiatric disorders| 0
increase in emergency department visits during heatwaves| 0
thorough history including medication history necessary| 0
communication with physician and pharmacy| 0
electronic health records with pharmacy fill histories| 0
severe NEHT caused by anticholinergic medications| 0
patients with psychiatric disorders and older adults vulnerable| 0
counsel on NEHT risk during summer months| 168
advised to remain hydrated| 168
advised to avoid high temperature environments| 168
importance of medication reconciliation| 168
patient consent for publication obtained| 0
provenance and peer review not commissioned| 0
64 years old|0
woman|0
bipolar depression|0
diabetes|0
migraine headaches|0
known seizure disorder|0
found unresponsive in a non-air-conditioned room|0
ambient temperature outside in excess of 90°F (33°C)|0
home medications include amitriptyline 175 mg daily|0
cyclobenzaprine 10 mg daily|0
lurasidone 80 mg daily|0
benztropine 1 mg three times a day|0
topiramate extended release 100 mg daily|0
clonazepam 0.5 mg daily|0
trazodone 100 mg daily|0
sitagliptin 25 mg daily|0
erenumab 70 mg injected monthly|0
Emergency medical service called|0
febrile on initial evaluation|0
cool compresses applied|0
transported to the hospital|0
hypotensive (blood pressure 84/42)|0
febrile with a rectal temperature of 42°C|0
skin warm and dry|0
mucous membranes dry|0
remainder of exam normal|0
neurological examination responsive only to painful stimuli|0
no focal neurological deficits|0
no hyperreflexia|0
no rigidity|0
leucocytosis (11,400)|0
creatine phosphokinase normal|0
EKG normal|0
admitted to intensive care unit (ICU)|0
started on vancomycin and cefepime|0
blood cultures grew Staphylococcus hominis|24
core body temperature decreased to less than 38°C|48
mentation returned to baseline|48
transferred to medical floor|48
treated for Staph hominis bacteraemia with 7-day course of vancomycin|48
discontinue use of cyclobenzaprine on discharge|168
quick recovery|168
lack of neurological findings (rigidity, tremors)|168
severe NEHT with associated bacteraemia determined as cause|168
initially thought to be severely septic|0
started on broad spectrum antibiotics|0
concern for drug-drug interactions|0
serotonin syndrome considered|0
low suspicion for serotonin syndrome|0
blood cultures obtained|0
toxicology consulted|0
blood cultures positive for S. hominis|24
toxicology’s assessment stated NEHT precipitated by multiple anticholinergic medications|24
mentation improved to baseline|24
revealed feeling overheated and fatigued for past 2 weeks|-336
no medication changes in past 2 weeks|-336
primary care physician advised to continue current medication regimen|168
discontinued cyclobenzaprine per toxicology’s recommendation|168
encouraged to discuss weaning medications|168
educated about risks of polypharmacy|168
combination of anticholinergic medications increased susceptibility to NEHT|0
amitriptyline, trazodone, cyclobenzaprine, benztropine inhibited sweating|0
topiramate caused hypohydrosis|0
NEHT diagnosed earlier if core temperature remained elevated|0
high risk for hyperthermia|0
high dosage medications may increase risk|0
Anticholinergic Risk Scale score 9|0
Naranjo Scale score 4 (possible adverse drug reaction)|0
counselling on risks of NEHT|168
medicine reconciliation periodically|168
vulnerability of patients with psychiatric disorders|0
increase in emergency department visits during heatwaves|0
thorough history including medication history necessary|0
communication with physician and pharmacy|0
electronic health records with pharmacy fill histories|0
severe NEHT caused by anticholinergic medications|0
patients with psychiatric disorders and older adults vulnerable|0
counsel on NEHT risk during summer months|168
advised to remain hydrated|168
advised to avoid high temperature environments|168
importance of medication reconciliation|168
patient consent for publication obtained|0
provenance and peer review not commissioned|0
