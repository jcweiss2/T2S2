30 years old | 0
Caucasian | 0
female | 0
gravida 2 para 1 | 0
presented at 34 2/7 weeks of gestation | 0
emergency room | 0
preterm labor | 0
no significant past medical history | 0
no surgical history | 0
postpartum depression | 0
denied recent international travel | 0
last travel 2 months prior to delivery | -1440
denied illnesses in 3 months prior to delivery | -2160
no sick contacts in last month prior to delivery | -720
no known positive COVID-19 contacts | -720
denied fever | 0
denied respiratory symptoms | 0
denied fatigue | 0
denied myalgia | 0
denied anosmia | 0
denied cough | 0
adequate prenatal care | 0
no maternal concerns | 0
no fetal concerns | 0
prenatal tests unremarkable | 0
group B Streptococcus status unknown | 0
SARS-CoV-2 testing not done | 0
precipitous vaginal delivery | 0
spontaneous rupture of membranes | 0
no respiratory symptoms before delivery | -240
no respiratory symptoms during delivery | 0
no respiratory symptoms after delivery | 240
no chorioamnionitis | 0
placental pathology assessment not done | 0
newborn vigorous at birth | 0
Apgar score 8 at 1 minute | 0
Apgar score 9 at 5 minutes | 0
skin-to-skin care with mother | 0
respiratory distress (grunting) | 0
transfer to radiant warmer | 0
transfer to newborn nursery | 0
noninvasive respiratory support with Vapotherm | 0
capillary blood gas unremarkable | 0
chest X-ray hazy lung fields | 0
no clear infiltrates | 0
no effusions | 0
CBC normal | 0
differential normal | 0
prematurity | 0
continued need for respiratory support | 0
lack of neonatal intensive care services | 0
transfer to level III NICU | 5
worsening hypercarbia | 5
respiratory support escalated to CPAP | 5
noninvasive positive pressure ventilation | 5
FiO2 21% | 5
improvement | 5
lack of prenatal maternal COVID-19 testing | 0
infant tested for SARS-CoV-2 at 24 hours | 24
SARS-CoV-2 positive at DOL 4 | 96
repeat SARS-CoV-2 test DOL 4 | 96
SARS-CoV-2 positive DOL 6 | 144
parents afebrile | 0
parents asymptomatic | 0
allowed bedside visitation | 0
breastfeeding not done | 0
expressed breast milk | 0
COVID-19 positive on DOL 4 | 96
parental visitation restricted | 96
droplet precautions | 96
contact precautions | 96
parents tested with antigen immunoassay | 96
parents SARS-CoV-2 negative | 96
parents tested with RT-PCR DOL 5 | 120
parents SARS-CoV-2 negative | 120
no parental symptoms | 0
respiratory support weaned | 24
empiric antibiotics (ampicillin, gentamicin) | 0
antibiotics discontinued | 48
sepsis evaluation unremarkable | 0
blood culture unremarkable | 0
CBC unremarkable | 0
C-reactive protein unremarkable | 0
feedings via gavage | 0
discharged at 9 days | 216
full oral feeds | 216
indirect hyperbilirubinemia | 0
phototherapy | 0
positive newborn screen for congenital adrenal hyperplasia | 0
congenital adrenal hyperplasia ruled out | 0
transport team notified | 0
no COVID-19 cases in caretakers | 0
NICU transport team tested for antibodies | 0
antibodies negative | 0
neonatal SARS-CoV-2 infection | 24
respiratory distress at birth | 0
asymptomatic mother | 0
mother negative SARS-CoV-2 tests | 96
