28 years old | 0
male | 0
class III obesity | 0
BMI 70.1 kg/m2 | 0
admitted to hospital | 0
weight gain 80 kg | -8760
worsening edema | -168
dyspnea on exertion | -168
supplemental oxygen | 0
arterial blood gas | 0
pH 7.21 | 0
PaCO2 78 mmHg | 0
PaO2 105 mmHg | 0
HCO3− 30.7 mmol/L | 0
provisional diagnosis of acute cardiac failure | 0
obesity hypoventilation syndrome | 0
noninvasive positive-pressure ventilation therapy | 0
furosemide | 0
worsening hypercapnia | 24
impaired consciousness | 24
admitted to ICU | 24
GCS 14 | 24
blood pressure 128/74 mmHg | 24
heart rate 90 bpm | 24
SpO2 90% | 24
expiratory positive airway pressure 6 cmH2O | 24
inspiratory positive airway pressure 18 cmH2O | 24
facial and leg edema | 24
wheezing on expiration | 24
no heart murmur | 24
mildly elevated inflammatory response | 24
elevated BNP level | 24
arterial blood gas analysis | 24
pH 7.236 | 24
PaCO2 94 mmHg | 24
PaO2 78 mmHg | 24
HCO3 39.1 mmol/L | 24
lactate 4.9 mmol/L | 24
respiratory acidosis | 24
chest radiograph | 24
marked cardiomegaly | 24
enhanced pulmonary vasculature | 24
electrocardiogram | 24
heart rate 80 bpm | 24
sinus rhythm | 24
chest computed tomography | 24
no infiltrative shadow | 24
no pleural effusion | 24
no atelectasis | 24
contrast-enhanced CT | 24
no thrombus in pulmonary artery | 24
intubated | 24
ventilator set to assist/control mode | 24
FIO2 0.6 | 24
ventilation frequency 16/min | 24
pressure control 16 cmH2O | 24
positive end-expiratory pressure 10 cmH2O | 24
PAC placed | 48
mean pulmonary artery pressure 49 mmHg | 48
central venous pressure 10 mmHg | 48
pulmonary artery wedge pressure 18 mmHg | 48
cardiac output 7.8 L/min | 48
cardiac index 2.8 L/min/m2 | 48
diagnosis of pulmonary hypertension | 48
transoesophageal echocardiography | 120
no abnormal left ventricular wall motion | 120
no significant valvular disease | 120
no patent foramen ovale | 120
deep sedation management | 120
continuous administration of muscle relaxants | 120
catheter removed | 240
suspicion of catheter infection | 240
mean pulmonary artery pressure 31 mmHg | 240
noradrenaline administration | 240
muscle relaxants discontinued | 240
spontaneous respiration restored | 240
NAd administration discontinued | 360
hemodynamic stability | 360
extubated | 552
discharged from ICU | 672
discharged from hospital | 2040