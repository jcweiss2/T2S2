34 years old | 0
male | 0
admitted to the intensive care unit | 0
septic shock | 0
multiple organ failure | 0
poor oral intake | 0
fever | 0
altered mental status | 0
anorexia | 0
dyspnea | 0
alcohol use disorder | -6720
immigrated from Sudan | -6720
employed at a meat processing plant | -6720
scleral icterus | 0
dry mucosal membranes | 0
tachycardia | 0
bilateral rales | 0
rhonchi | 0
abdomen soft and nontender | 0
abdomen distended | 0
temperature 35.8 degrees Celsius | 0
heart rate 152 beats per minute | 0
sinus rhythm | 0
respiratory rate of 42 breaths per minute | 0
blood pressure 114/75 mmHg | 0
oxygen saturation 97% | 0
heated high flow nasal cannula oxygen therapy | 0
leukopenia | 0
elevated lactic acid | 0
hyperbilirubinemia | 0
elevated liver enzymes | 0
normal ammonia level | 0
urine toxicology screen positive for benzodiazepines | 0
acute respiratory acidosis | 0
anion gap metabolic acidosis | 0
hypoxic respiratory failure | 0
COVID-19 PCR positive | 0
microangiopathic hemolytic anemia ruled out | 0
multifocal pneumonia | 0
right-sided pleural effusion | 0
cardiac enlargement | 0
severe hepatosplenomegaly | 0
steatosis | 0
gallstones | 0
pericholecystic fluid | 0
enlarged kidneys | 0
mesenteric edema | 0
diffuse abdominal lymphadenopathy | 0
omental nodularity | 0
treated with dexamethasone | 0
remdesivir not used | 0
tocilizumab not used | 0
intubation | 24
escalation of antibiotics | 24
worsening renal function | 24
hemodialysis | 24
infectious work-up negative for human immunodeficiency virus | 24
infectious work-up negative for hepatitis B | 24
infectious work-up negative for hepatitis C | 24
infectious work-up negative for syphilis | 24
infectious work-up negative for histoplasma | 24
infectious work-up negative for aspergillus | 24
infectious work-up negative for cryptococcus | 24
infectious work-up negative for candida | 24
infectious work-up negative for pneumocystis jirovecii | 24
infectious work-up negative for herpes simplex virus 1 and 2 | 24
infectious work-up negative for cytomegalovirus | 24
infectious work-up negative for clostridium difficile | 24
infectious work-up negative for malaria | 24
Epstein Barr virus serology consistent with past exposure and immunity | 24
broad gastrointestinal stool polymerase chain reaction negative | 24
sputum cultures with pan-sensitive Klebsiella Pneumoniae | 24
antibiotics de-escalated | 24
hepatitis A IgM serology positive | 24
interferon-gamma release assay positive | 24
concern for latent versus active tuberculosis | 24
acid-fast bacilli cultures positive | 48
diagnosed with active tuberculosis | 48
four-drug TB therapy initiated | 48
four-drug TB therapy discontinued | 50
rifampin, ethambutol, and pyrazinamide restarted | 50
isoniazid held | 50
levofloxacin started | 50
concern for secondary hemophagocytic lymphohistiocytosis | 72
persistent fever | 72
hepatomegaly | 72
erythropenia | 72
leukopenia | 72
elevated ferritin | 72
elevated triglycerides | 72
hypofibrinogenemia | 72
CXCL9 elevated | 72
soluble IL-1 receptor alpha elevated | 72
bone marrow biopsy planned | 72
bone marrow biopsy deferred | 72
H-score calculated | 72
H-score 233 points | 72
empiric methylprednisolone initiated | 72
etoposide not initiated | 72
tracheostomy | 96
percutaneous endoscopic gastrostomy | 96
tracheostomy removed | 168
percutaneous endoscopic gastrostomy removed | 168
hemodialysis line removed | 168
discharged to a long-term care facility | 168
steroid taper | 168
antituberculosis therapy | 168
rifampin | 168
ethambutol | 168
pyrazinamide | 168
levofloxacin | 168