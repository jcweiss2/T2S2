5 years old | 0
male | 0
presented to the pediatric emergency department | 0
fever | -48
neck pain | -48
odynophagia | -48
headache | -48
nasal congestion | -48
lethargy | -48
no cough | -48
no abdominal pain | -48
no vomiting | -48
no diarrhea | -48
no rash | -48
no sick contacts | -48
no recent travel | -48
mild COVID-19 infection 6 weeks prior | -1008
unvaccinated against COVID-19 | 0
tachycardia | 0
fever (103.4 F) | 0
normal blood pressure | 0
normal respiratory rate | 0
normal oxygen saturation | 0
full range of motion of the neck | 0
no respiratory distress | 0
no stridor | 0
shotty posterior cervical lymphadenopathy | 0
elevated CRP | 0
elevated ESR | 0
lymphopenia | 0
normal WBC | 0
mild hyponatremia | 0
negative rapid antigen testing for group A Streptococcus | 0
negative nasopharyngeal PCR for SARS-CoV-2 | 0
negative influenza A and B | 0
negative respiratory syncytial virus | 0
negative blood cultures | 0
X-ray of the neck showing paravertebral soft tissue swelling | 0
CT of the neck suggested retropharyngeal phlegmonous changes or possible early abscess | 0
bilateral reactive lymphadenopathy | 0
admitted | 0
dexamethasone | 0
IV ampicillin–sulbactam | 0
decreased oral intake | 0
maintenance IV fluids | 0
pediatric ENT consultation | 0
antibiotics without drainage | 0
persistent high-grade fevers | 72
tachycardia | 72
tachypnea | 72
worsening tachycardia | 96
worsening tachypnea | 96
borderline hypotension | 96
ongoing fevers | 96
softer voice | 96
facial edema | 96
increased pain with neck motion | 96
new prominent cardiac gallop | 96
1+ soft pulses | 96
mild hepatomegaly | 96
increased CRP | 96
IV Vancomycin | 96
repeat CT neck | 96
CT chest revealed bilateral pleural effusions | 96
subsegmental atelectasis | 96
periportal edema | 96
mediastinal lymphadenopathy | 96
deterioration leading to PICU transfer | 96
epinephrine infusion | 96
high-flow nasal cannula | 96
suspicion for MIS-C | 96
cardiac echocardiogram showing mild biventricular systolic dysfunction | 96
mild four-chamber dilated chambers | 96
positive SARS-CoV-2 serologies | 96
elevated CRP | 96
elevated troponin | 96
elevated BNP | 96
elevated D-dimer | 96
elevated ferritin | 96
elevated fibrinogen | 96
elevated INR | 96
diagnosis of MIS-C | 96
IVIG | 96
methylprednisolone | 96
enoxaparin | 96
clinical improvement | 144
discharge | 192
repeat cardiac echo | 192
normal cardiac function | 192
normal coronary arteries | 192
prednisolone taper | 192
amoxicillin–clavulanate | 192
aspirin 81 mg | 192
