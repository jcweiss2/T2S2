25 years old | 0
male | 0
admitted to the emergency room | 0
motor vehicle crash | -1
Glasgow coma score 8/15 | 0
electively intubated | 0
mechanical ventilation | 0
whole-body computed tomography (CT) | 0
nondisplaced compression fracture at the ninth and 10th thoracic vertebrae | 0
bilateral basal atelectasis/consolidation | 0
bilateral ground-glass opacities | 0
nondisplaced manubrium sternal fracture | 0
small (0.5 cm) contusion over the spleen | 0
acute left subdural hemorrhage | 0
underlying mild brain edema | 0
right midline shift of approximately 1 cm | 0
emergency decompressive craniectomy | 0
extraventricular drain (EVD) insertion | 0
admitted to the surgical intensive care unit (SICU) | 0
mechanical ventilation | 0
fever | 120
leukocytosis | 120
septic workup | 120
cerebral spinal fluid (CSF) analysis | 120
culture | 120
vancomycin | 120
meropenem | 120
antibiotic regimen adjusted | 168
lipid-formulated amphotericin B | 168
vancomycin | 168
EVD removed | 192
deterioration of consciousness | 216
new CT scan of the brain | 216
active hydrocephalus | 216
worsening midline shift | 216
another EVD inserted | 216
full septic workup | 216
debridement at the cephalic surgical site | 432
ceftazidime | 432
tracheostomy placement | 600
febrile | 600
Glasgow coma scale 8/15 | 600
leukocytosis (14.3 k/µL) | 600
septic screening | 600
CSF culture revealed M. hominis | 600
M. hominis | 600
intravenous ciprofloxacin 400 mg every 8 h | 624
clinically improved | 936
transferred to the general ward | 936
third EVD remained in place | 1080
nasogastric feeding | 1080
tracheostomy | 1080
transferred to another health care facility | 1104
M. hominis identified using MALDI-TOF MS | 624
M. hominis susceptible to tetracycline, fluoroquinolone, clindamycin, chloramphenicol, streptomycin, and gentamicin | 624
M. hominis resistant to beta-lactams, sulfonamides, trimethoprim, and rifampin | 624