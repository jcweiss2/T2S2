33 years old | 0
female | 0
admitted to the University Hospital | 0
shortness of breath | 0
feeling ill | -168
general health deterioration | -168
high fever | -168
SARS-CoV-2 positive | -168
elevated body mass index (34) | 0
no preexisting conditions | 0
respiratory function compromised | 0
severe hypoxemia | 0
endotracheal intubation | 0
mechanical ventilation | 0
high ventilation pressure | 0
poor O2 saturation | 0
veno-venous extracorporeal membrane oxygenation (vvECMO) administered | 0
severe acute respiratory distress syndrome (COVID-19-ARDS) | 0
continuous catecholamines | 0
hemodialysis initiated | 96
ECMO removed | 336
weaning achieved | 360
impaired liver function | 0
elevated liver parameters | 0
elevated cholestasis parameters (bilirubin, GGT, AP) | 0
toxic/ischemic liver injury suspected | 0
ketamine sedation | 0
elevated liver enzymes persisted | 336
elevated bilirubin (1.4 mg/dL) | 336
elevated GGT (1299 U/L) | 336
elevated AP (1883 U/L) | 336
elevated AST (162 U/L) | 336
elevated ALT (119 U/L) | 336
Ursofalk® 1000 mg initiated | 336
computed tomography of abdomen (day 10) | 240
no parenchymal damage | 240
no cholestasis | 240
MRCP on day 47 | 1128
mild stenosis of distal CBD | 1128
suspected stricture of prepapillary CBD | 1128
ERCP on day 60 | 1440
rarefication of intrahepatic bile ducts | 1440
MRCP follow-up on day 105 | 2520
multiple diffuse stricture of CBD | 2520
stricture of intrahepatic biliary tree | 2520
T2-signal changes with restricted diffusion | 2520
cholangetic abscess formation | 2520
MRI follow-up on day 129 | 3096
progressive encapsulated intrahepatic fluid accumulation | 3096
restricted diffusion | 3096
rim-contrast enhancement | 3096
progressive intrahepatic abscess | 3096
persistent elevated inflammatory parameters | 0
elevated CRP (peak 217 mg/L) | 0
worsening general condition | 0
renal failure | 0
hemodialysis three times a week | 0
elevated bilirubin (peak 17.29 mg/dL) | 3336
interdisciplinary meeting | 0
orthotopic liver transplantation discussed | 0
kidney transplantation discussed | 0
deterioration in general health | 0
impaired respiratory function | 0
transplantation plan discarded | 0
SSC-CIP suspected | 0
post-COVID-19 cholangiopathy suspected | 0
remdesivir treatment | 0
Convalescent Plasma Transfusion | 0
antibiotics (Noxafil®, Piperacillin/Tazobactam®, Tygacil®, Curam®) | 0
organ failure (respiratory system, kidneys, liver) | 3696
death | 3696
