33 years old | 0
    woman | 0
    previously healthy | 0
    weighing 70 kg | 0
    brought to the emergency department | 0
    cardiac arrest | 0
    undergoing liposuction of her thighs | -45
    liposuction of mid-back | -45
    harvesting 1.5 L of fat | -45
    procedure lasted 45 minutes | -45
    becoming more somnolent | -44
    blood pressure 170/90 mmHg | -44
    suspected hypoglycemia | -44
    administered oral dextrose solution | -44
    started feeling dizzy | -24
    rapid decline of mental status | -24
    tonic-clonic seizure | -24
    complete loss of consciousness | -24
    EMS arrived | -24
    gasping | -24
    cyanotic | -24
    drooling | -24
    cardiopulmonary arrest during transport | -24
    EMS initiated resuscitation | -24
    arrival to ED | 0
    cardiac monitor showed asystole | 0
    intubated | 0
    resuscitation resumed | 0
    return of spontaneous circulation | 22
    asked for procedure details | 0
    power-assisted liposuction technique | 0
    use of five vials of lidocaine 2% | -45
    total lidocaine dose 5000 mg | -45
    prior abdominal liposuction three months earlier | -2160
    normal sinus rhythm | 22
    no QT prolongation | 22
    corrected QT interval 466 ms | 22
    normal QRS interval 100 ms | 22
    no ST- or T-wave abnormalities | 22
    neurological examination revealed no response | 22
    Glasgow Coma Scale 3T | 22
    pupils equal and reactive | 22
    preserved corneal reflexes | 22
    preserved oculocephalic reflexes | 22
    downward Babinski reflex bilaterally | 22
    arterial blood gas pH 7.34 | 22
    CO2 pressure 39.9 mmHg | 22
    O2 pressure 131 mmHg | 22
    bicarbonate 20.8 mmol/L | 22
    white blood cell count 9.8 × 109/L | 22
    hemoglobin 10.4 g/dL | 22
    platelet count 336 × 106/L | 22
    troponin 0.003 ng/mL | 22
    sodium 144 mmol/L | 22
    potassium 3.5 mmol/L | 22
    chloride 99 mmol/L | 22
    bicarbonate 16 mmol/L | 22
    glucose 346 mg/dL | 22
    blood urea nitrogen 13 mg/dL | 22
    creatinine 1.0 mg/dL | 22
    aspartate aminotransferase 225 IU/L | 22
    alanine aminotransferase 238 IU/L | 22
    γ-glutamyl transpeptidase 12 IU/L | 22
    alkaline phosphatase 55 IU/L | 22
    lactate 17.55 mmol/L | 22
    serum lidocaine level 5.30 µg/mL | 22
    CT scan of brain | 22
    CT angiography of chest | 22
    bilateral consolidations | 22
    aspiration pneumonitis | 22
    no intracranial bleeding | 22
    no pulmonary embolism | 22
    no aortic dissection | 22
    started on antibiotic therapy | 22
    generalized myoclonic jerks | 22
    possible anoxic brain injury | 22
    started on valproic acid | 22
    admitted to ICU | 0
    MRI of brain three days later | 72
    severe hypoxic6 ischemic brain injury | 72
    electrocerebral silence on EEG | 72
    increase in brain edema | 1440
    increased pressure | 1440
    electrolytes disturbances | 1440
    multiple nosocomial infections | 1440
    end-organ damage | 1440
    death secondary to septic shock | 1440
    
    
    