40 years old | 0
male | 0
admitted to the hospital | 0
gunshot wound to the upper abdomen | 0
gunshot wound to the chest | 0
Glasgow coma score of 15 | 0
hemodynamically stable | 0
focused assessment with sonography was positive | 0
taken emergently to the operating room | 0
exploratory laparotomy | 0
repair of a ballistic gastric serosal tear | 0
diagnostic pericardial window | 0
complex hepatotrhaphy | 0
liver debridement with argon beam coagulation | 0
liver packing | 0
repair of the diaphragm | 0
right chest tube placement | 0
multiple ballistic perforations | 0
injured diaphragm | 0
injured liver | 0
injured gastric serosa | 0
estimated blood loss for the procedure | 0
1,300 mL blood loss | 0
transferred to the intensive care unit | 0
intubated | 0
5 cm H2O positive end expiratory pressure | 0
sedated | 0
plans to return to the OR the following day | 0
closure of the abdomen | 0
transfused one unit of A+ packed red blood cells | 0
serial labs were ordered | 0
initial hemoglobin on admission | 0
12.9 g/dL hemoglobin | 0
received a unit of mismatched blood | -0.5
clerical error | -0.5
spiked a fever | 0.5
developed hematuria | 0.5
became hypotensive | 0.5
blood bank notified the floor | 0.5
stabilized with intravenous hydrocortisone | 1
stabilized with intravenous diphenhydramine | 1
stabilized with intramuscular eipnephrine | 1
given multiple liter IV fluid boluses | 1
labs revealed direct Coombs test was positive | 2
IgG interpretation | 2
haptoglobin was < 5.8 mg/dL | 2
lactate dehydrogenase was 1,193 U/L | 2
coagulation parameters were worsening | 2
hypotension required a norepinephrine drip | 2
preoperative creatinine had been normal | 0
1.5 m/dL creatinine | 0
determined to have an AHTR | 2
employed an urgent RBCET | 4.5
RBCET started | 4.5
five units of type O negative blood | 4.5
target hemoglobin goal of 9.0 g/dL | 4.5
received five units of fresh frozen plasma | 24
received two units of PRBC | 24
received one unit of platelets | 24
creatinine peaked at 2.12 mg/dL | 17
direct Coombs returned negative | 9
norepinephrine was discontinued | 48
clinical and lab parameters stabilized | 96
discharged in stable condition | 120
no apparent long-term consequences | 120