73 years old | 0
male | 0
prostatic adenocarcinoma | -18240
prostatectomy | -18240
Gleason score of 8 | -18240
protein specific antigen of 17 ng/ml | -18240
adjuvant radiotherapy | -7300
hormone therapy | -7300
acute urine retention | -72
abdominal pain | -72
hematuria | -72
dysuria | -72
transit disorders | -72
anorexia | -72
asthenia | -72
admitted to the hospital | 0
bladder catheterization | 0
thematic urine with clots | 0
venous line with administration | 0
biological check-up | 0
creatinine at 149 | 0
K at 6.9 | 0
electrocardiogramm | 0
blood cells at 14 000/mm3 | 0
C reactive protein at 450 | 0
CT scan | 0
full bladder with multiple dense formations | 0
air bubbles in the bladder | 0
dense heterogeneous non-decreasing formation at the level of the dome | 0
air bubbles within the formation | 0
parietal defect | 0
subperitoneal effusion | 0
hydroaerobic levels in the bladder | 0
pneumoperitoneum | 0
diffuse infiltration of the mesenteric fat | 0
decision to refer to the operating room | 0
intraperitoneal exploration | 12
discreet dilatation of the bowels | 12
minimal effusion | 12
hematoma through the affected peritoneum | 12
breach in the peritoneum | 12
aspiration of the fluid | 12
removal of the hematoma | 12
bladder breach | 12
necrotic edges | 12
inflamed wall | 12
extraction of the intravesical hematoma | 12
cystorraphy | 12
epiploplasty | 12
placement of a Redon drain | 12
peritoneal closure | 12
renal purification session | 24
favorable evolution | 24
urine began to clear | 24
diuresis of 2400 cc | 24
Redon at 30 cc | 24
biological parameters evolution | 24
creatinine at 83 | 24
K at 5.1 | 24
blood cells at 11 700/mm3 | 24
CRP at 324 | 24
extubation | 48
recovery of consciousness | 48
apyretic | 48
diuresis at 2 L | 48
removal of the Redon | 48
disorder of consciousness | 48
respiratory distress | 48
ventricular tachycardia | 48
cardiorespiratory arrest | 48
death | 48
gangrenous cystitis | 0 
DRESS syndrome | -672 
fever | -72 
rash | -72 
acne |  -672 
minocycline |  -672 
increased WBC count | 0 
eosinophilia | 0 
systemic involvement | 0 
diffuse erythematous or maculopapular eruption | 0 
pruritis | 0 
fever persisted | 0 
rash persisted | 0 
discharged | 24