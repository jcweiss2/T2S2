53 years old | 0
female | 0
admitted to the hospital | 0
chest pain | -72
sudden chest pain | -72
constant chest pain | -72
severe chest pain | -72
fever | -72
leukocytosis | -72
viral illness | -72
costochondritis | -72
cyclobenzaprine | -72
nonsteroidal anti-inflammatory | -72
ibuprofen | -72
normal sinus rhythm | -72
no ischemic changes | -72
blood cultures positive for Staphylococcus aureus | -48
low-grade fever | 0
heart rate above 90 beats per minute | 0
respirations over 20 | 0
septic | 0
Infectious Disease service contacted | 0
IV ceftriaxone 2 g daily | 0
IV vancomycin 1,250 mg twice daily | -48
mild murmur | 0
bacteremia | 0
transthoracic echocardiogram | 0
normal ejection fraction | 0
trivial regurgitation of valves | 0
mild regurgitation of mitral valve | 0
transesophageal echocardiogram not performed | 0
urine cultures negative | 0
urinalysis negative | 0
no sputum production | 0
no cough | 0
good dentition | 0
colonoscopy recommended | 0
chest X-ray performed | 0
new right pleural effusion | 0
CT of chest without contrast | 0
possible non-displaced fracture of sternum | 0
osteomyelitis of sternum | 0
magnetic resonance imaging of chest | 0
osteomyelitis involving manubrium and upper part of sternum body | 0
tender to palpation | 0
no overlying erythema | 0
IV antibiotics | 0
improvement of chest pain | 24
IV ceftriaxone 2 g once daily | 0
ibuprofen | 0
oxycodone/acetaminophen | 0
erythrocyte sedimentation rate 38 mm/hr | 0
C-reactive protein 9.9 mg/L | 0
trend of erythrocyte sedimentation rate and C-reactive protein | 24
no recurrence of infection | 336
persistent chest pain | 336
antinuclear antibody 1:320 centromere pattern | 720
HIV test negative | 0
hepatitis panel negative | 0
elevated liver function | 0
aspartate aminotransferase 103 U/L | 0
alanine aminotransferase 180 U/L | 0
alkaline phosphatase 135 U/L | 0
trend of liver function tests | 24
discharge | 336