25 years old | 0
male | 0
admitted to the hospital | 0
fell into an electroplating pool containing 10% HF and 50% nitric acid | -2
exposed to HF and nitric acid | -2
removed clothes and irrigated with running water | -2
calcium gluconate gel was not applied | -2
sent to the hospital emergency room | -2
complained of mild dyspnea | 0
complained of hoarseness | 0
complained of severe pain in the burn area | 0
erythema | 0
edematous | 0
heart rate of 120 beats/min | 0
respiratory rate of 28 breaths/min | 0
axillary temperature at 37.5° | 0
SaO2 at 92% | 0
blood pressure of 124/78 mm Hg | 0
cutaneous injuries on approximately 60% of the TBSA | 0
third degree burns on approximately 13% of the burn area | 0
deep partial thickness burns | 0
conjunctiva congested and edematous | 0
cornea without ulcer | 0
frequent rinsing with normal saline | 0
levofloxacin eye drops | 0
1% calcium gluconate | 0
nasal and oral mucosa pale | 0
profuse secretions | 0
rinsing with 5% calcium gluconate | 0
tracheotomy | 0
bedside mechanic ventilation | 0
burn areas rinsed with 5% sodium bicarbonate | 0
covered with wet sterile gauze containing 10% calcium gluconate | 0
electrocardiography normal | 0
hypocalcemia | 0
hypomagnesemia | 0
hyperkalemia | 0
fluid resuscitation | 0
intravenous administration of 10% calcium gluconate | 0
intravenous administration of 25% magnesium sulfate | 0
invasive hemodynamic monitoring | 0
ventricular fibrillation | 4
defibrillation | 4
dobutamine | 4
glucocorticoid | 4
antibiotic | 4
oxygenation index deteriorated | 24
hypoxemia worsened | 24
ELWI increased | 24
frothy sputum | 24
pulmonary edema | 24
ECMO | 38
venoarterial ECMO | 38
fiberoptic bronchoscopies | 72
aspiration and lavage | 72
burn wound infections | 120
fiberoptic bronchoscopies | 168
congested, edematous mucosa | 168
weaned off of ECMO | 264
catheter removed | 264
vessels repaired | 264
pulmonary infection | 384
burn wound infections | 384
microbiological identification | 384
antibiotic therapy | 384
weaned off of CRRT | 624
skin grafting | 720
fearful of stopping CRRT | 720
discharged | 2160