25 years old | 0
    male | 0
    admitted to the hospital | 0
    exposure to 10% hydrofluoric acid | -2
    exposure to 50% nitric acid | -2
    whole body soaked in acids | -2
    clothes removed by co-workers | -2
    irrigation with running water for 20 minutes | -2
    calcium gluconate gel not applied | -2
    sent to emergency room | -2
    mild dyspnea | 0
    hoarseness | 0
    severe pain in burn area | 0
    erythema | 0
    edematous | 0
    heart rate 120 beats/min | 0
    respiratory rate 28 breaths/min | 0
    axillary temperature 37.5°C | 0
    SaO2 92% | 0
    blood pressure 124/78 mm Hg | 0
    cutaneous injuries on 60% TBSA | 0
    third degree burns on 13% burn area | 0
    deep partial thickness burns on remaining area | 0
    conjunctiva congested | 0
    conjunctiva edematous | 0
    cornea without ulcer | 0
    eyes rinsed with normal saline for 30 minutes | 0
    levofloxacin eye drops | 0
    1% calcium gluconate every 4 hours | 0
    nasal mucosa pale | 0
    oral mucosa pale | 0
    profuse secretions in oral cavity | 0
    rinsing with 5% calcium gluconate | 0
    hypoxemia | 0
    inhalational injury | 0
    tracheotomy | 0
    bedside mechanical ventilation | 0
    burn areas rinsed with 5% sodium bicarbonate | 0
    covered with wet sterile gauze containing 10% calcium gluconate | 0
    electrocardiography normal | 0
    ionic calcium 0.192 mmol/L | 0
    total calcium 0.72 mmol/L | 0
    magnesium 0.4 mmol/L | 0
    potassium 5.49 mmol/L | 0
    sodium 136.8 mmol/L | 0
    liver function normal | 0
    renal function normal | 0
    continuous cardiac monitoring | 0
    fluid resuscitation | 0
    intravenous administration of 10% calcium gluconate | 0
    intravenous administration of 25% magnesium sulfate | 0
    20 mL intravenous bolus of 10% calcium gluconate | 0
    continuous infusion of calcium gluconate at 6 g/h | 0
    continuous intravenous drip of magnesium sulfate at 1.5 g/h | 0
    invasive hemodynamic monitoring with PICCO | 0
    cardiac index 3.02 L/min/m² | 0
    extravascular lung water index 16 mL/kg | 0
    central venous pressure 5 mm Hg | 0
    systemic vascular resistance index 2213 dyn.s/cm⁵.m² | 0
    global end-diastolic index 450 mL/m² | 0
    CRRT applied | 0
    ventricular fibrillation at 4 hours postexposure | 4
    ventricular fibrillation episodes within next 3 hours | 4-7
    defibrillation successful 10 times | 7
    calcium gluconate administered after defibrillation | 7
    invasive arterial blood pressure 86/48 mm Hg | 7
    cardiac index decreased to 2.5 L/min/m² | 7
    dobutamine administration | 7
    glucocorticoid (methylprednisolone 40 mg q8h) | 0
    antibiotic (piperacillin tazobactam 4.5 g q8h) | 0
    oxygenation index deteriorated (PaO2/FiO2 55.2/1.0) | 24
    hypoxemia worsened | 24
    extravascular lung water index increased to 25 mL/kg | 24
    frothy sputum suctioned | 24
    pulmonary edema confirmed by chest x-ray | 24
    ultrafiltration increased | 24
    PEEP increased | 24
    ECMO initiated at 38 hours postexposure | 38
    venoarterial ECMO | 38
    ECMO flow rate 3.0 L/min | 38
    activated clotting time maintained at 160-200 seconds | 38
    arterial oxygen saturation 98% | 38
    hypoxemia corrected | 38
    fiberoptic bronchoscopy on day 3 | 72
    pale mucus in bronchi | 72
    aspiration and lavage performed | 72
    postirrigation fluid yellow | 72
    burn wound infections on day 5 | 120
    fiberoptic bronchoscopy on day 7 | 168
    congested mucosa | 168
    edematous mucosa | 168
    hemodynamic profile stable on day 11 | 264
    oxygenation improved | 264
    ECMO weaned | 264
    catheter removed | 264
    vessels repaired | 264
    deterioration on day 16 | 384
    pulmonary infection | 384
    burn wound infections | 384
    methicillin-resistant Staphylococcus aureus | 384
    Pseudomonas aeruginosa | 384
    antibiotic therapy with imipenem/cilastin | 384
    antibiotic therapy with vancomycin | 384
    CRRT weaned on day 26 | 624
    skin grafting after 1 month | 720
    CRRT cessation after 2 months | 1440
    discharged without complications after 3 months | 2160
    