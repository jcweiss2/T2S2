81 years old | 0
male | 0
admitted to hospital | 0
faeculent vomiting | 0
change in bowel habit | -504
right-sided rib pain | -504
hip pain | -504
unintentional weight loss | -504
atrial fibrillation | 0
warfarin | 0
hypertension | 0
laparoscopic cholecystectomy | -7920
gallstone disease | -7920
bile spillage | -7920
stone debris spillage | -7920
apyrexial | 0
normotensive | 0
normocardiac | 0
abdominal distension | 0
generalized abdominal pain | 0
right flank pain | 0
right upper quadrant peritonitis | 0
absent bowel sounds | 0
empty rectum | 0
high leucocyte count | 0
C-reactive protein | 0
dilated loops of proximal small bowel | 0
faecal loading | 0
no pneumoperitoneum | 0
abdominal CT scan | 0
bowel dilatation | 0
right sub-hepatic multiloculated collection | 0
pneumobilia | 0
emergency laparotomy | 24
no perforation | 24
purulent right upper quadrant collection | 24
pus aspirated | 24
microbiological culture | 24
abdominal lavage | 24
postoperative improvement | 48
sepsis | 48
intensive care admission | 48
broad-spectrum antibiotic therapy | 48
inotropic support | 48
A. israelii isolated | 192
tazobactam and piperacillin | 192
discharged home | 336
intravenous Tazocin | 336
oral penicillin | 336
persistently raised inflammatory markers | 1008
repeat ultrasound scan | 1008
collection of extra-luminal fluid | 1008
ultrasound-guided drainage | 1008
further 3-month course of oral penicillin | 1008
full recovery | 1512