2 years old | 0
boy | 0
admitted to the hospital | 0
high fever | 0
fever not relieved by antipyretic treatment | 0
febrile (BT 39.2°C) | 0
severely ill | 0
extremely irritable | 0
heart rate 170/min | 0
blood pressure 98/51 mmHg | 0
petechial lesions disseminated on torso and limbs | 0
suspicion of meningococcemia | 0
intravenous fluids | 0
ceftriaxone administration | 0
hypotension | 0
massive IV fluids resuscitation | 0
neurological deterioration | 0
inotropic support | 0
intubation | 0
mechanical ventilation | 0
transfer to PICU | 0
Neisseria meningitidis serogroup B isolation from blood culture | 0
cerebrospinal fluid sample normal | 0
continuation of ceftriaxone | 0
gradual improvement of general conditions | 24
CRP decrease from 345 mg/L to 48.4 mg/L | 24
inotropic agents stopped | 120
extubation | 168
continued fever spikes (BT 38.5°C) | 168
suspicion of hospital acquired infection | 168
broader antibiotic therapy with ceftriaxone, gentamicin, teicoplanin | 168
negative blood and urine cultures | 168
negative lumbar puncture | 168
negative chest X-ray | 168
negative brain MRI | 168
transfer to GPU | 312
stable but still febrile (BT 38.5°C) | 312
presence of cutaneous ulcers | 312
hemoglobin 8.1 g/L | 312
RBC 3,050,000/mm3 | 312
MCV 80.6 fl | 312
WBC count 25,830/mm3 | 312
PMN 16,140/mm3 | 312
PLT count 1,090,000/mm3 | 312
CRP 44.80 mg/L | 312
fever persisted (days 136-20) | 312
fever spikes every 6-8 hours | 504
BT >39°C | 504
CRP 89.70 mg/L | 504
ESR 36 mm/h | 504
Ferritin 173 ug/L | 504
neopterine 31.0 nmol/L | 504
TNF 29.8 ng/L | 504
broader antibiotic therapy with meropenem and teicoplanin | 504
negative cultures | 504
erythematous papular rash | 528
hepatomegaly | 528
bilateral cervical lymphadenopathy | 528
suspicion of viral infection | 600
negative serological tests for Adenovirus, EBV, CMV, Parvovirus B19 | 600
neck ultrasound reactive lymph nodes | 600
suspicion of atypical Kawasaki | 600
normal electrocardiogram | 600
echocardiography showed hyperechogenicity of mitral papillary muscles | 600
IVIG administration (2 g/kg) | 624
IVIG repeated | 672
HB 7.4 g/dL | 696
RBC 3,050,000/mm3 | 696
MCV 76.4 fl | 696
WBC count 23,470/mm3 | 696
PMN 11,050/mm3 | 696
PLT count 98,000/mm3 | 696
LDH 1091 U/L | 696
normal renal function | 696
albumin 31 g/L | 696
AST 86 IU/L | 696
ALT 117 IU/L | 696
GGT 300 U/L | 696
sodium 135 mmol/L | 696
triglycerides 361 mg/dL | 696
prolongation of prothrombin time | 696
prolonged activated partial thromboplastin time | 696
fibrinogen 1 g/L | 696
CRP 64.70 mg/L | 696
vitamin K administration | 696
fresh frozen plasma administration | 696
normalization of coagulation pattern | 696
bone marrow aspirate no hemophagocytic lymphohistiocytosis | 696
conjunctival injection | 720
fissured dry lips | 720
facial edema | 720
feet edema | 720
diagnosis of KD | 720
IVMP administration (30 mg/kg) | 768
CRP decrease to 3.36 mg/L | 840
fever reduction | 840
afebrile | 888
discharge | 888
normal ECG at follow-up | 2160
normal echocardiogram at follow-up | 2160
