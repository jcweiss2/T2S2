46 years old | 0
    male | 0
    admitted to ICU | 0
    severe chronic obstructive pulmonary disease (COPD) | 0
    bronchial asthma | 0
    acute proptosis of both eyes | 0
    clinical picture of acute bilateral proptosis with retracted lids | 0
    history of similar episodes in the past | -4320
    diagnosis of globe luxation | 0
    globe reduction by pressing on superior sclera and pinching upper lid | 0
    previous episodes over past 4–5 years | -35040
    episodes initiated after starting wheezing episodes | -35040
    globe luxation episodes occurred with COPD exacerbations | -35040
    bilateral pseudophakia | 0
    normal pupil | 0
    normal fundus | 0
    axial length 23.8 mm | 0
    CT scan of orbit showing no orbital mass | 0
    CT scan showing proptosed eye with stretched optic nerve | 0
    orbit volume normal | 0
    globe volume normal | 0
    repeated episodes of globe luxation every 2 hours | 0
    bilateral temporary tarsorrhaphy | 48
    respiratory paralysis | 72
    septicemia | 72
    expired on third day | 72
    