58 years old | 0
female | 0
admitted to the hospital | 0
upper respiratory tract infection | -168
cough | -168
occasional shortness of breath | -168
low-grade fevers | -168
decadron 40 mg i.m | -168
antibiotics prescription | -168
antibiotics prescription not filled | -168
shortness of breath worsening | -168
cough worsening | -168
acute airway obstruction | 0
acute epiglottitis | 0
emergently intubated | 0
transferred to intensive care unit | 0
hypotensive (BP 90/76 mmHg) | 0
hypoxemic | 0
ventilator support | 0
vasopressors | 0
chest x-ray bilateral peri-hilar consolidation and infiltrates | 0
CT chest diffuse bilateral interstitial and alveolar infiltrates | 0
CT chest bilateral lower lobe air space consolidation | 0
CT neck diffuse swelling of soft tissues | 0
CT neck loss of fat planes throughout pharyngeal region | 0
CT neck marked thickening of retropharyngeal soft tissue | 0
no loculated fluid collections | 0
minimal cervical adenopathy | 0
leukocytosis (15.8×10^9/L) | 0
borderline hematocrit (44%) | 0
normal platelet count (170.5×10^9/L) | 0
normal sodium (139 mEq/L) | 0
normal renal function (BUN 14 mg/dL, creatinine 1.1 mg/dL) | 0
normal ALT (31 IU/L) | 0
normal AST (17 IU/L) | 0
arterial blood gas pH 7.03 | 0
arterial blood gas PaCO2 46 mmHg | 0
arterial blood gas PaO2 46 mmHg | 0
negative blood cultures | 0
intubated in ICU for approximately one week | 168
endoscopic evaluation unremarkable | 0
started on intravenous solumedrol 40 mg q8h | 0
chest x-rays bilateral infiltrates | 168
negative urine cultures | 0
negative sputum cultures | 0
negative influenza serology | 0
negative parainfluenza serology | 0
negative Brucella serology | 0
negative tuberculosis serology | 0
negative Bordetella pertussis serology | 0
negative Mycoplasma serology | 0
negative Legionella serology | 0
negative Chlamydia pneumoniae serology | 0
started on broad-spectrum antibiotics | 0
started on fluconazole 400 mg daily | 0
extubated | 240
transferred to medical floor | 240
recurrent respiratory distress | 240
necessitating reintubation | 240
ICU readmission | 240
bronchoscopy no abnormalities | 240
bronchoalveolar lavage normal | 240
lung biopsy normal | 240
lower GI hemorrhage | 240
upper endoscopy non-contributory | 240
biopsy not done | 240
planned colonoscopy not performed due to hypotension | 240
KUB showed massive pneumoperitoneum | 240
emergent laparotomy | 240
small bowel perforations | 240
cecal perforation | 240
mucosa ulcers | 240
mucosa edema | 240
invasive fungal elements in submucosal and peritoneal tissue | 240
vascular invasion | 240
fungal hyphae morphology consistent with Mucormycosis | 240
vascular thrombosis | 240
hemorrhage | 240
acute inflammation | 240
necrosis | 240
started on liposomal amphotericin B | 240
started on micafungin | 240
discontinuation of fluconazole | 240
additional intestinal resections | 240
final laparotomy 6 days after initial intervention | 288
near complete intestinal infarction | 288
progressive multiorgan failure | 288
ongoing shock | 288
diffuse intestinal ischemia and infarction | 288
DNR status | 288
withdrawal of care | 288
deceased | 288
