79 years old | 0
woman | 0
presented to the emergency department | 0
acute limb ischemia in left leg | -2
hypertension | 0
atrial fibrillation | 0
non-dialysis-dependent chronic renal failure | 0
acute aortic embolic occlusion | -17520
bilateral femoral catheter embolectomy | -17520
warfarin | -17520
irregular medication use | 0
INR 1.1 | 0
arrhythmic pulse | 0
hypertension (160x110mmHg) | 0
normal femoral, popliteal, pedal pulses on right leg | 0
weak femoral pulse on left leg | 0
no distal pulses on left leg | 0
pain | 0
motor deficit | 0
grade IIb limb ischemia | 0
referred for surgery | 0
diminished creatinine clearance (Cockroft-Gault 12mL/min) | 0
general anesthesia | 0
femoral access | 0
dissection of common, superficial, deep femoral arteries | 0
arteriotomy | 0
4-Fr embolectomy catheter used | 0
thrombi retrieved from deep and superficial femoral arteries | 0
catheter progressed >60cm in superficial femoral artery | 0
no pedal or posterior tibial artery catheter palpation | 0
insignificant back bleeding | 0
decision to perform angiography | 0
CO2 angiography | 0
patent popliteal artery | 0
patent fibular artery | 0
occlusion of mid-third anterior tibial artery | 0
new embolectomy performed | 0
catheter progressed to pedal artery | 0
more thrombi retrieved | 0
control angiography | 0
complete resolution of anterior tibial artery occlusion | 0
contrast up to foot | 0
28mL CO2 used | 0
arteriorraphy performed | 0
popliteal and pedal pulses present | 0
resolution of pallor | 0
resolution of hypothermia | 0
no compartment syndrome | 0
ICU admission until postoperative day 11 | 264
no nephrotoxic agents administered | 264
furosemide-stimulated diuresis | 264
urinary tract infection | 432
deteriorating renal function | 432
uremia | 432
dialysis started on postoperative day 18 | 432
pneumonia | 864
septic shock | 864
vasoactive drugs required for 2 days | 864
unrecovered renal function | 864
discharged to hospice care | 864
pedal pulse present | 864
no limb deficit | 864
chronic dialysis required | 864
