65 years old | 0
    man | 0
    fever | 0
    chills | 0
    loss of consciousness | 0
    no response to physical stimulation | 0
    right limb muscle strength grade 0 | 0
    left limb muscle strength grade 2 | 0
    Babinski’s sign positive on right lower limb | 0
    leukocyte count 17.5×10^9/L | 0
    neutrophil count 16.28×10^9/L | 0
    CRP 84.29 mg/L | 0
    blood cultures grew Streptococcus viridans | 0
    no abnormalities in electrocardiogram | 0
    no abnormalities in myocardial infarction markers | 0
    catheter ablation 2 weeks before presentation |  -336
    refractory atrial fibrillation |  -336
    left craniocerebral infarction | 0
    air emboli in right lobe | 0
    air between left atrium and esophagus | 0
    pericardial effusions | 0
    atrial-esophageal fistula | 0
    sepsis | 0
    cerebral infarction | 0
    urgent surgical operation | 0
    esophageal fistula 35 cm from incisor teeth | 0
    fresh blood in esophageal fistula | 0
    standard posterolateral thoracotomy | 0
    dense adhesions between lower esophagus and pericardium | 0
    necrotic tissues above the fistula | 0
    massive bleeding | 0
    1 cm-diameter defect in posterior wall of left atrium | 0
    4-0 Prolene suture | 0
    autologous pericardial tissue | 0
    3-incision esophagectomy | 0
    simultaneous anastomosis | 0
    intensive care unit monitoring | 0
    anti-infection administration | 0
    nutritional support | 0
    anticoagulation | 0
    supportive treatments | 0
    died of sepsis |  576
    died of multiple organ failure |  576

<|eot_id|>
