55 years old | 0
female | 0
admitted to the hospital | 0
fever | -168
dysuria | -168
malaise | -168
urinary incontinence | -168
difficulty ambulating | -168
worsening back pain | -168
poorly-controlled diabetes mellitus type 2 | 0
hypertension | 0
hyperlipidemia | 0
chronic low back pain | 0
temperature 38.3 °C | 0
blood pressure 186/82 mmHg | 0
pulse 114 beats per minute | 0
respiratory rate 20 breaths per minute | 0
oxygen saturation 98% | 0
mildly confused | 0
lethargic | 0
electrocardiography tracing showed poor R-wave progression | 0
left ventricular hypertrophy | 0
chest X-ray did not show any acute process | 0
white blood cell count was 15,600 per cubic millimeter | 0
87% neutrophils | 0
comprehensive metabolic panel and coagulation studies were normal | 0
urine analysis had 3+ bacteria | 0
blood and urine cultures were obtained | 0
sepsis secondary to a urinary tract infection | 0
ceftriaxone | 0
piperacillin –tazobactam | 24
persistent fever | 24
worsening mentation | 24
transferred to the medical intensive care unit | 24
encephalopathy | 24
generalized weakness | 24
diminished strength | 24
diminished tone | 24
diminished sensation in all extremities | 24
patella tendon reflexes were absent bilaterally | 24
rectal tone was normal | 24
nuchal rigidity | 24
moderate tenderness along the entire spine | 24
gram negative bacilli | 24
vancomycin | 24
meropenem | 24
MRI of the spine with contrast | 24
extensive posterior epidural fluid collection | 24
internal air locules | 24
mass effect on the cord | 24
severe thecal sac stenosis | 24
cervical, thoracic, and lumbar decompression | 48
evacuation and aggressive irrigation of the epidural abscess | 48
ESBL-producing Klebsiella pneumoniae | 48
sensitive to fluoroquinolones | 48
sensitive to gentamicin | 48
sensitive to meropenem | 48
fungal and acid fast cultures were negative | 48
recovery was painstakingly slow | 72
intensive physical and occupational therapy | 72
discharged to a skilled nursing facility | 168
meropenem for a total of 12 weeks | 1008
repeat MRI of the entire spine showed complete resolution of epidural abscess | 1008