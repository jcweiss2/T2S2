55 years old | 0
male | 0
presented to the hospital | 0
severe watery diarrhoea | -5760
opening bowels 8-9 times in 24 h | -5760
no other significant symptoms | 0
normal colonoscopy 3 days prior to admission | -72
no past medical history | 0
no surgical history | 0
no regular medications | 0
no significant family history | 0
non-smoker | 0
lethargic | 0
clinically dehydrated | 0
eGFR of 14 mL/min/1.73 m2 | 0
creatinine of 381 μmol/L | 0
serum potassium 2.5 mmol/L | 0
serum calcium 2.88 mmol/L | 0
normal anion gap metabolic acidosis | 0
pH of 7.16 | 0
base excess of -14.2 mmol/L | 0
lactate 0.8 mmol/L | 0
inflammatory markers within normal range | 0
coeliac serology negative | 0
vasculitis screen negative | 0
stool cultures negative | 0
admitted to intensive care unit | 0
central potassium replacement | 0
aggressive rehydration with i.v. fluids | 0
parenteral nutrition commenced | 0
poor absorption from nasogastric feeding | 0
contrast-enhanced CT scan of abdomen obtained | 0
32-mm heterogenous mass in pancreatic body | 0
multiple hypo-attenuating lesions in liver | 0
hepatic lesions suspicious for metastases | 0
metastatic functional pancreatic neuroendocrine tumour suspected | 0
T2 N0 M1 staging | 0
fasting serum gut hormone profile sent | 0
somatostatin 116 pmol/L | 0
gastrin 47 pmol/L | 0
glucagon 66 pmol/L | 0
chromogranin A 223 pmol/L | 0
chromogranin B >4500 pmol/L | 0
VIP 211 pmol/L | 0
PP 6928 pmol/L | 0
repeat profile with concordant results | 0
ultrasound-guided core biopsy of liver lesion | 0
necrotic tissue | 0
viable tumour cells | 0
CK8/18 expression | 0
synaptophysin expression | 0
CD56 expression | 0
chromogranin A expression negative | 0
well-differentiated grade I neuroendocrine tumour | 0
Ki-67 proliferation index 2.9% | 0
p53 WT expression | 0
i.v. somatostatin analogue infusion initiated | 0
octreotide 12.5 µg/h | 0
diarrhoea settled completely | 0
renal function failed to improve | 0
spike high temperatures | 0
inflammatory markers increased | 0
repeat CT obtained | 0
significant intra-intestinal fluid | 0
blood cultures positive for K lebsiella | 0
blood cultures positive for Enterococcus | 0
autonecrosis of pancreatic primary | 0
autonecrosis of liver lesions | 0
treated for bowel bacteria overgrowth sepsis | 0
ultrafiltration commenced | 0
renal function improved significantly | 0
inflammatory markers settled | 0
stepped down to the ward | 0
discharged | 288
converted to long-acting lanreotide injections | 288
eGFR 54 mL/min/1.73 m2 at discharge | 288
in hospital for 1 month | 288
under investigation for MEN-1 syndrome | 0
serum calcium elevated | 0
parathyroid hormone raised | 0
prolactin levels raised | 0
Gallium-68 DOTA-TATE PET CT | 0
MRI of liver | 0
stable disease | 0
good response to SSA | 0
no evidence of disease beyond pancreas and liver | 0
remain on lanreotide injections for 6 months | 0
repeat Ga68 PET/CT | 0
repeat MRI imaging | 0
plan for surgical resection of primary tumour | 0
plan for debulking of liver lesions | 0
VIPoma suspected | 0
PPoma suspected | 0
no shortness of breath | 0
denies chest pain | 0
no rash | 0
no nausea | 0
no vomiting | 0
no back pain | 0
no flushing | 0
no bloating | 0
no mass-effect symptoms | 0
