53 years old | 0
male | 0
admitted to the hospital | 0
subjective fever | -72
chills | -72
diffuse myalgias | -72
productive cough | -72
pneumonia | 0
Levofloxacin prescribed | 0
discharged home | 0
dyspnea | 24
nausea | 24
emesis | 24
syncope | 24
tachycardia (130 beats/min) | 24
normotensive (131/98 mmHg) | 24
tachypneic (22 breaths/minute) | 24
normal oxygen saturations (99% on room air) | 24
temperature of 37.1 degrees Celsius | 24
white blood cell count (WBC) of 22 × 10^9/L | 24
troponin-t (high sensitivity) 31 ng/L | 24
creatine kinase (CK) 7910 U/L | 24
lactate of 9.7 mmol/L | 24
sinus tachycardia | 24
frequent PVCs | 24
sepsis suspected | 24
blood cultures drawn | 24
IV fluids administered | 24
Piperacillin-Tazobactam administered | 24
transferred to tertiary care centre | 24
heart rate 122 beats per minute | 24
blood pressure 111/88 mmHg | 24
respiratory rate 25 breaths per minute | 24
oxygen saturation 99% | 24
temperature of 36.5 degrees Celsius | 24
bilateral pulmonary crackles | 24
normal heart sounds | 24
jugular venous pressure at 4 cm above sternal angle | 24
no pedal edema | 24
mottled skin | 24
cool extremities | 24
capillary refill time approximately six seconds | 24
benign abdominal exam | 24
unremarkable chest radiograph | 24
CT pulmonary angiogram completed | 24
no pulmonary emboli | 24
pulmonary edema | 24
NT-proBNP 8146 pg/ml | 24
consulted to Cardiology | 24
decompensated heart failure suspected | 24
urgent TTE performed | 24
severe global hypokinesis of the left ventricle | 24
ejection fraction of 15–20% | 24
small pericardial effusion | 24
myocarditis suspected | 24
admitted to Cardiac Intensive Care Unit | 24
treated with Colchicine | 24
treated with high-dose Aspirin | 24
troponin peaked at 3871 ng/L | 24
nasopharyngeal swab completed | 24
influenza antigen testing via PCR | 24
empiric Oseltamivir started | 24
positive for Influenza B (post-admission day three) | 72
increasing dyspnea (post-admission day four) | 96
shortness of breath (post-admission day four) | 96
increased oxygen requirements (post-admission day four) | 96
new right-sided airspace opacity on chest x-ray | 96
Vancomycin added | 96
pain to forearms bilaterally | 96
CK elevated at 8321 U/L | 96
right forearm increased sensitivity | 96
right forearm became firm | 96
compartment pressure of 60 mmHg | 96
bedside right forearm fasciotomy | 96
transferred to Medical-Surgical ICU | 96
hypoxemia worsened (post-admission day four) | 96
intubation (post-admission day four) | 96
heart rate 111 beats per minute (ICU admission) | 96
blood pressure 86/57 mmHg (ICU admission) | 96
MAP of 67 mmHg (ICU admission) | 96
oxygen saturation 97% (ICU admission) | 96
pressure support of 8 cmH20 | 96
FiO2 of 45% | 96
PEEP of 10 cmH20 | 96
respiratory rate 19 breaths per minute (ICU admission) | 96
temperature of 37.1 degrees Celsius (ICU admission) | 96
diffuse bilateral crackles | 96
normal heart sounds (ICU admission) | 96
elevated jugular venous pressure at 6 cm above sternal angle | 96
3+ pitting edema to sacrum | 96
mottled skin (ICU admission) | 96
cool extremities (ICU admission) | 96
Norepinephrine started | 96
Furosemide infusion initiated | 96
Norepinephrine discontinued (post-admission day five) | 120
ejection fraction 60–65% (post-admission day five) | 120
intubated (post-admission day seven) | 168
Oseltamivir continued (post-admission day seven) | 168
blood cultures negative (post-admission day seven) | 168
repeat NP PCR test sent (post-admission day seven) | 168
positive for Influenza B (post-admission day ten) | 240
oliguric (post-admission day ten) | 240
creatinine 416 umol/L | 240
renal failure | 240
rhabdomyolysis | 240
continuous renal replacement therapy (post-admission day ten) | 240
recovery of renal function (post-admission day twelve) | 288
extubated (post-admission day twelve) | 288
transferred to home hospital (post-admission day fifteen) | 360
discharged (post-admission day twenty-four) | 576
no influenza immunization | 0
family history of congenital heart disease | 0
