48 years old | 0
    male | 0
    admitted to the hospital | 0
    fever | -72
    cough | -72
    breathlessness | -72
    type 2 diabetes mellitus | -72
    poor glycemic control | -72
    body temperature 39.7°C | 0
    respiratory rate 28 breaths/min | 0
    heart rate 128 bpm | 0
    blood pressure 100/60 mm Hg | 0
    mucopurulent sputum | 0
    decreased breath sounds on the left lung base | 0
    no bilateral crackles | 0
    total leukocyte count 15.9 G/L | 0
    neutrophil predominance | 0
    platelet 78 G/L | 0
    C-reactive protein 324.6 mg/l | 0
    hemoglobin A1c 9.09% | 0
    small pleural effusion | 0
    consolidated lung base | 0
    Ziehl-Neelsen stain from sputum negative for acid-fast bacilli | 0
    sputum culture | 0
    blood culture | 0
    pleural fluid culture | 0
    Gram-negative bacilli in sputum Gram stain | 0
    abundant white blood cells in sputum Gram stain | 0
    blood culture turbidity after 4 days | 96
    subculture on blood agar and Drigalski agar | 96
    smooth white non-hemolytic colonies on blood agar | 96
    non-fermenting colonies on Drigalski agar | 96
    Gram-negative bacilli on Gram stain | 96
    catalase-positive | 96
    oxidase-positive | 96
    API 20NE identification as Aeromonas salmonicida | 96
    treated with cefoperazone-sulbactam | 0
    treated with azithromycin | 0
    treated with gentamicin | 0
    antibiotics changed to piperacillin-tazobactam | 96
    antibiotics changed to fosfomycin | 96
    antibiotics changed to meropenem | 96
    antibiotics changed to ciprofloxacin | 96
    clinical response improved but unstable | 96
    occasional high fever 40°C | 96
    occasional tachypnea | 96
    continued cough with mucopurulent sputum | 96
    16S rRNA gene sequencing matched B. pseudomallei | 96
    second sputum culture same as previous | 96
    immunochromatographic assay positive for melioidosis | 96
    sensitive to amoxicillin/clavulanic acid | 96
    sensitive to ceftazidime | 96
    sensitive to meropenem | 96
    sensitive to sulfamethoxazole/trimethoprim | 96
    sensitive to piperacillin/tazobactam | 96
    transferred to Hue Central hospital | 96

    48 years old | 0
    male | 0
    admitted to the hospital | 0
    fever | -72
    cough | -72
    breathlessness | -72
    type 2 diabetes mellitus | -72
    poor glycemic control | -72
    body temperature 39.7°C | 0
    respiratory rate 28 breaths/min | 0
    heart rate 128 bpm | 0
    blood pressure 100/60 mm Hg | 0
    mucopurulent sputum | 0
    decreased breath sounds on the left lung base | 0
    no bilateral crackles | 0
    total leukocyte count 15.9 G/L | 0
    neutrophil predominance | 0
    platelet 78 G/L | 0
    C-reactive protein 324.6 mg/l | 0
    hemoglobin A1c 9.09% | 0
    small pleural effusion | 0
    consolidated lung base | 0
    Ziehl-Neelsen stain from sputum negative for acid-fast bacilli | 0
    sputum culture | 0
    blood culture | 0
    pleural fluid culture | 0
    Gram-negative bacilli in sputum Gram stain | 0
    abundant white blood cells in sputum Gram stain | 0
    blood culture turbidity after 4 days | 96
    subculture on blood agar and Drigalski agar | 96
    smooth white non-hemolytic colonies on blood agar | 96
    non-fermenting colonies on Drigalski agar | 96
    Gram-negative bacilli on Gram stain | 96
    catalase-positive | 96
    oxidase-positive | 96
    API 20NE identification as Aeromonas salmonicida | 96
    treated with cefoperazone-sulbactam | 0
    treated with azithromycin | 0
    treated with gentamicin | 0
    antibiotics changed to piperacillin-tazobactam | 96
    antibiotics changed to fosfomycin | 96
    antibiotics changed to meropenem | 96
    antibiotics changed to ciprofloxacin | 96
    clinical response improved but unstable | 96
    occasional high fever 40°C | 96
    occasional tachypnea | 96
    continued cough with mucopurulent sputum | 96
    16S rRNA gene sequencing matched B. pseudomallei | 96
    second sputum culture same as previous | 96
    immunochromatographic assay positive for melioidosis | 96
    sensitive to amoxicillin/clavulanic acid | 96
    sensitive to ceftazidime | 96
    sensitive to meropenem | 96
    sensitive to sulfamethoxazole/trimethoprim | 96
    sensitive to piperacillin/tazobactam | 96
    transferred to Hue Central hospital | 96

    48 years old | 0
    male | 0
    admitted to the hospital | 0
    fever | -72
    cough | -72
    breathlessness | -72
    type 2 diabetes mellitus | -72
    poor glycemic control | -72
    body temperature 39.7°C | 0
    respiratory rate 28 breaths/min | 0
    heart rate 128 bpm | 0
    blood pressure 100/60 mm Hg | 0
    mucopurulent sputum | 0
    decreased breath sounds on the left lung base | 0
    no bilateral crackles | 0
    total leukocyte count 15.9 G/L | 0
    neutrophil predominance | 0
    platelet 78 G/L | 0
    C-reactive protein 324.6 mg/l | 0
    hemoglobin A1c 9.09% | 0
    small pleural effusion | 0
    consolidated lung base |B0
    Ziehl-Neelsen stain from sputum negative for acid-fast bacilli | 0
    sputum culture | 0
    blood culture | 0
    pleural fluid culture | 0
    Gram-negative bacilli in sputum Gram stain | 0
    abundant white blood cells in sputum Gram stain | 0
    blood culture turbidity after 4 days | 96
    subculture on blood agar and Drigalski agar | 96
    smooth white non-hemolytic colonies on blood agar | 96
    non-fermenting colonies on Drigalski agar | 96
    Gram-negative bacilli on Gram stain | 96
    catalase-positive | 96
    oxidase-positive | 96
    API 20NE identification as Aeromonas salmonicida | 96
    treated with cefoperazone-sulbactam | 0
    treated with azithromycin | 0
    treated with gentamicin | 0
    antibiotics changed to piperacillin-tazobactam | 96
    antibiotics changed to fosfomycin | 96
    antibiotics changed to meropenem | 96
    antibiotics changed to ciprofloxacin | 96
    clinical response improved but unstable | 96
    occasional high fever 40°C | 96
    occasional tachypnea | 96
    continued cough with mucopurulent sputum | 96
    16S rRNA gene sequencing matched B. pseudomallei | 96
    second sputum culture same as previous | 96
    immunochromatographic assay positive for melioidosis | 96
    sensitive to amoxicillin/clavulanic acid | 96
    sensitive to ceftazidime | 96
    sensitive to meropenem | 96
    sensitive to sulfamethoxazole/trimethoprim | 96
    sensitive to piperacillin/tazobactam | 96
    transferred to Hue Central hospital | 96

    48 years old | 0
    male | 0
    admitted to the hospital | 0
    fever | -72
    cough | -72
    breathlessness | -72
    type 2 diabetes mellitus | -72
    poor glycemic control | -72
    body temperature 39.7°C | 0
    respiratory rate 28 breaths/min | 0
    heart rate 128 bpm | 0
    blood pressure 100/60 mm Hg | 0
    mucopurulent sputum | 0
    decreased breath sounds on the left lung base | 0
    no bilateral crackles | 0
    total leukocyte count 15.9 G/L | 0
    neutrophil predominance | 0
    platelet 78 G/L | 0
    C-reactive protein 324.6 mg/l | 0
    hemoglobin A1c 9.09% | 0
    small pleural effusion | 0
    consolidated lung base | 0
    Ziehl-Neelsen stain from sputum negative for acid-fast bacilli | 0
    sputum culture | 0
    blood culture | 0
    pleural fluid culture | 0
    Gram-negative bacilli in sputum Gram stain | 0
    abundant white blood cells in sputum Gram stain | 0
    blood culture turbidity after 4 days | 96
    subculture on blood agar and Drigalski agar | 96
    smooth white non-hemolytic colonies on blood agar | 96
    non-fermenting colonies on Drigalski agar | 96
    Gram-negative bacilli on Gram stain | 96
    catalase-positive | 96
    oxidase-positive | 96
    API 20NE identification as Aeromonas salmonicida | 96
    treated with cefoperazone-sulbactam | 0
    treated with azithromycin | 0
    treated with gentamicin | 0
    antibiotics changed to piperacillin-tazobactam | 96
    antibiotics changed to fosfomycin | 96
    antibiotics changed to meropenem | 96
    antibiotics changed to ciprofloxacin | 96
    clinical response improved but unstable | 96
    occasional high fever 40°C | 96
    occasional tachypnea | 96
    continued cough with mucopurulent sputum | 96
    16S rRNA gene sequencing matched B. pseudomallei | 96
    second sputum culture same as previous | 96
    immunochromatographic assay positive for melioidosis | 96
    sensitive to amoxicillin/clavulanic acid | 96
    sensitive to ceftazidime | 96
    sensitive to meropenem | 96
    sensitive to sulfamethoxazole/trimethoprim | 96
    sensitive to piperacillin/tazobactam | 96
    transferred to Hue Central hospital | 96