64 years old | 0
female | 0
admitted to the hospital | 0
severe headache | -24
right periorbital swelling | -24
mid-facial swelling | -24
fever (39°C) | -336
headache | -336
light pain in the right ear | -336
purulent secretion from the ear | -336
swelling of the skin behind the right ear | -336
redness of the skin behind the right ear | -336
tinnitus | -336
hearing disorder | -336
right acute mastoiditis | -336
arterial hypertension | -336
angiotensin-converting enzyme inhibitors | -336
marked right facial swelling | 0
marked periorbital swelling | 0
right blepharoptosis | 0
chemosis | 0
proptosis | 0
visual acuity of 7/12 on the right eye | 0
pain on right eye movement | 0
febrile (38.8°C) | 0
conscious | 0
somnolent | 0
elevated white blood cells count | 0
elevated erythrocyte sedimentation rate | 0
elevated C-reactive protein | 0
normal renal function | 0
normal liver function | 0
negative tests for vasculitis | 0
negative HIV test | 0
negative diabetes test | 0
prothrombin G20210A mutation | 0
normal coagulation profile | 0
normal urinalysis | 0
non-opacification of the right cavernous sinus on MRI | 0
intravenous Ceftriaxone | 0
anticoagulation with Enoxaparin | 0
no corticosteroids | 0
blood culture positive for Streptococcus pneumoniae | 48
severe headache persisted | 72
anorexia | 72
high fever | 72
confusion | 72
shortness of breath | 96
reduced oxygen saturation | 96
right lobar pneumonia | 96
non-invasive mechanical ventilation | 96
Amikacin | 96
Piperacillin-Tazobactam | 96
improvement of symptoms | 168
persistence of lacunar image in right cavernous sinus | 168
diminished periorbital swelling | 168
discharged | 336
oral anticoagulant (Acenocoumarol) | 336
full recovery | 336
