25 years old | 0
housewife | 0
given birth to a 3.1-kg baby girl | 0
pregnancy | -168 (assuming pregnancy duration mentioned as 37 weeks, which is approximately 37*7*24=6216 hours before delivery, but since the delivery is at admission, timestamp is 0, so pregnancy start would be -6216 hours. However, the text states "37th week of her first pregnancy", which implies the pregnancy was 37 weeks long, so the start of pregnancy would be -37*7*24= -6216 hours. However, the patient was admitted after delivery, so delivery is at timestamp 0. Therefore, the pregnancy events before delivery would have negative timestamps.)
spontaneous vaginal delivery | 0
episiotomy | 0
severe pain in the region of her buttocks | 0 (post-delivery, so timestamp 0)
shortness of breath | -21 (sudden onset at 03:00h the next day; assuming "next day" after delivery, so 24 hours later, but she arrived at the emergency department the same day. However, the timestamp for admission is 0, so the onset of shortness of breath was 21 hours before admission (03:00 next day, assuming delivery at 00:00, next day 03:00 would be 27 hours after delivery, but since delivery is timestamp 0, and she arrived at the emergency department after the onset, which would be a negative timestamp. However, the timeline is complex; perhaps the onset was 21 hours before admission.)
worsening pain over her right thigh | -21 (same as shortness of breath)
drowsy | 0
tachypneic | 0
oxygen saturation of 56% on room air | 0
high-flow oxygen supply | 0
tachycardia | 0 (pulse 121 bpm)
afebrile | 0 (36°C)
blood pressure unrecordable | 0
resuscitation with 30 mL/kg normal saline | 0
persistently hypotensive | 0 (blood pressure 56/30 mmHg)
noradrenaline infusion | 0
blood pressure steadied | 0
IV heparin 5000 units | 0 (stat dose)
presumptive diagnosis of pulmonary embolism | 0
IV amoxicillin-clavulanate stat dose | 0
septicemic shock | 0
transferred to tertiary hospital | 0
electively intubated | 0
severe metabolic and lactic acidosis | 0
worsening respiratory distress | 0
120 mL/kg crystalloid given | 0
persistently hypotensive post-intubation | 0
fluid resuscitation | 0
adrenaline | 0
vasopressin | 0
dobutamine | 0
grossly swollen right thigh | 0
extensive blistering ecchymotic patches over right thigh | 0
right thigh extending to right buttock | 0
necrotizing fasciitis of the right thigh | 0
acute kidney injury | 0
rhabdomyolysis | 0
coagulopathy | 0
thrombocytopenia | 0
ischemic hepatitis | 0
IV meropenem | 0
IV clindamycin | 0
IV vancomycin | 0
cultures taken from blood and blister fluid | 0
high vaginal swab for culture | 0
transferred to intensive care unit | 0
orthopedic and surgical opinions sought | 0
extensive wound debridement planned | 0
CT pulmonary angiography | 0
small pulmonary embolism | 0
bedside echocardiography | 0
good contractility | 0
intravenous immunoglobulin | 0 (given on the same day)
file.open("data.txt", ios::in | ios::out);
