25 years old | 0
primigravida | 0
male infant | 0
40 + 2 weeks’ gestation | 0
spontaneous onset of labor | 0
fetal distress | 0
ventouse-assisted delivery | 0
birth weight 3940 grams | 0
required immediate resuscitation with mask ventilation | 0
intubated at 8 minutes of age | 0.13
transferred to the neonatal intensive care unit (NICU) | 0.13
synchronized intermittent positive pressure ventilation (SIPPV) | 0.13
gentamicin 4 mg/kg 24-hourly | 0.13
benzyl penicillin 60 mg/kg 12-hourly | 0.13
neutropenia | 18
significant left shift | 18
elevated C-reactive protein (CRP; 60 mg/L) | 18
elevated procalcitonin (68.55 µg/L) | 18
lumbar puncture | 23
normal cell count | 23
negative for a range of pathogens including meningococcus | 23
placental surface eSwab | 23
light pure growth of an organism | 23
Gram-negative diplococci | 23
Neisseria meningitidis | 23
molecular testing | 23
blood cultures taken from the newborn pre–antibiotic treatment | -0.48
negative | -0.48
heel-prick blood in EDTA | 5.5
detected the presence of N. meningitidis genogroup W DNA | 5.5
acute funisitis (vasculitis of umbilical cord vessels) | 0
chorioamnionitis | 0
benzylpenicillin dosage was decreased | 13.5
changed to cefotaxime 50 mg/kg 12-hourly | 13.5
elevated leucocyte count of 21.1×109/L | -2.5
neutrophil count of 18.1×109/L | -2.5
discharged home from the NICU | 192
contact tracing | 192
chemoprophylaxis with ciprofloxacin | 192
vaccination with quadrivalent conjugate meningococcal vaccine | 192