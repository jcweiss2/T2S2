45 years old | 0
male | 0
admitted to the hospital | 0
swelling in the right lower limb | -120
tenderness | -120
leukocytosis | -120
necrotizing fasciitis | -120
septic shock | -120
central line insertion | 0
volume resuscitation | 0
treatment with antibiotics | 0
extensive debridement | 0
intubated | 0
mechanical ventilation | 0
inotropic support | 0
transferred to ICU | 0
bedside ultrasonography | 1
intraluminal hyperechoic shadow | 1
missed guidewire suspected | 1
X-ray ordered | 1
X-ray confirmed guidewire position | 2
ultrasound examination of central venous line | 2
guidewire found in external part | 2
left femoral central catheter inserted | 3
inotropic infusion pump shifted | 3
right internal jugular line clamped | 3
right internal jugular line removed | 3
guidewire removed | 3
repeat bedside ultrasound | 4
guidewire removal confirmed | 4
discharged | unknown