83 years old | 0
female | 0
weight loss | -2160
dyspepsia | -2160
admitted to the emergency department | 0
abdominal pain lasting three days | -72
fever | -48
hypertension | 0
diabetes mellitus | 0
blood pressure 110/70 mmHg | 0
no history of trauma | 0
no history of surgery | 0
no history of alcoholism | 0
no history of smoking | 0
diminished bowel sounds | 0
distended abdomen | 0
diffuse defense | 0
rebound | 0
sensitivity | 0
white blood cell 10.8 103/ml | 0
hemoglobin 8.1 g/dl | 0
urea 38 mg/dL | 0
creatinine 1.6 mg/dL | 0
potassium 5.7 mmol/L | 0
normal blood amylase level | 0
normal electrocardiogram | 0
free air under the right diaphragm | 0
widespread free abdominal fluid | 0
admitted to the intensive care unit | 0
supportive therapy | 0
midline laparotomy | 0
giant perforation 7x7 cm | 0
abdomen full of pus and fibrin | 0
aspiration of purulent material | 0
peritoneal cavity washed with warm saline | 0
decreased blood pressure | 0
inotropic support with dopamine | 0
biopsies from perforation edges | 0
gastric resection not suitable | 0
narrowed perforation with purse-string sutures | 0
omental flap prepared | 0
transfixed perforation with vicryl sutures | 0
narrowed perforation to 4 cm | 0
methylene blue test | 0
placement of three drains | 0
operation time 40 min | 0
intubated | 0
Meropenem 3*1 gr/iv | 0
reduced white blood cell count | 0
improved pre@-renal failure | 0
decreased inotropic agents | 0
smooth abdomen | 0
no distension | 0
no rigidity | 0
methylene blue test on day 5 | 120
methylene blue test on day 6 | 144
no leakage | 120
no leakage | 144
abdominal drains withdrawn | 144
improvement of peritonitis | 0
improved renal functions | 0
pulmonary problems not recovered | 0
conscious | 0
sedation given up | 0
attempted weaning from mechanical ventilator | 0
acquired pneumonia | 0
died of pulmonary failure | 360
moderately differentiated adenocarcinoma | 0
