18 years old | 0
female | 0
admitted to the hospital | 0
rising levels of human chorionic gonadotropin | 0
intermittent vaginal bleeding | 0
vaginal ultrasound scan | 0
intrauterine pregnancy | 0
surgical evacuation of the uterus | 0
abdominal pain | 24
temperature of 39.5°C | 24
suspecting severe endometritis | 24
metronidazole | 24
benzylpenicillin | 24
gentamicin | 24
deteriorated | 48
saturation fell to 90% | 48
respiratory rate rose to around 40 breaths per minute | 48
temperature peaked at 40.7°C | 48
C-reactive protein rose to around 300 mg/L | 48
leukocytes to around 15 × 10^9/L | 48
moved to the intensive care unit | 48
intubated | 48
CT scan | 48
thrombophlebitis of the internal jugular vein | 48
hepatomegaly | 48
diagnosed with Lemierre's syndrome | 48
benzylpenicillin and gentamicin discontinued | 48
tazocin | 48
clindamycin | 48
metronidazole | 48
heparin injections | 48
respiratory support | 72
antibiotics | 72
discharged | 168