64 years old| 0
    male | 0
    admitted to the hospital | 0
    general weakness | -168
    myalgia | -168
    abdominal pain | -168
    fever | 0
    feeling hot | 0
    headache | 0
    no cough | 0
    no sputum | 0
    no diarrhea | 0
    no vomiting | 0
    hypertension | -43800
    diabetes | -43800
    metformin | -43800
    glimepiride | -43800
    linagliptin | -43800
    losartan | -43800
    rosuvastatin | -43800
    dull pressing pain in the right upper quadrant | 0
    mild tenderness in the right upper quadrant | 0
    hypo-active bowel sound | 0
    no other specific findings in physical examinations | 0
    elevated white blood cell count | 0
    elevated ESR | 0
    elevated HS-CRP | 0
    no rebound tenderness | 0
    SMV thrombosis | 0
    influenza B positive | 0
    COVID-19 negative | 0
    peramivir administered | 0
    ICU admission | 0
    LMWH administered | 0
    no oral intake | 0
    total parenteral nutrition administered | 0
    ceftriaxone administered | 0
    fever persisted until day 2 | 72
    abdominal pain persisted until day 3 | 96
    abdominal discomfort persisted until day 6 | 144
    follow-up CT scan on day 8 | 192
    thrombus decreased | 192
    water intake | 204
    rivaroxaban initiated | 204
    soft diet | 240
    moved to general ward | 240
    third follow-up CT scan on day 16 | 384
    thrombus markedly reduced | 384
    discharged | 384
    negative tumor markers | 0
    negative lupus anticoagulant | 0
    negative rheumatoid factor | 0
    normal protein S activity | 0
    normal protein C activity | 0
    no other suspected underlying diseases | 0
    regular outpatient follow-up visits | 384
    improved symptoms | 384
    SMV thrombosis resolved on day 45 | 1080
    