38 years old | 0
female | 0
pregnant | 0
difficulty walking | -432
right inguinal region pain | -432
lower back pain | -432
low-lying placenta | -144
admitted to Department of Obstetrics | 0
body temperature 36.3°C | 0
pulse rate 83 beats/min | 0
blood pressure 116/50 mmHg | 0
respiratory rate 15 breaths/min | 0
SpO2 98% | 0
lower abdominal pain | 0
massive vaginal bleeding | 0
emergency Caesarean section | 0
transferred to ICU | 0
chest X-ray cardiac dilatation | 0
chest X-ray opacity bilateral lower lung fields | 0
hemoglobin 10.1 g/dL before childbirth | 0
hemoglobin 6.1 g/dL after childbirth | 0
contrast-enhanced CT bilateral pleural effusions | 24
contrast-enhanced CT multiple lung nodules | 24
contrast-enhanced CT multiple liver masses | 24
contrast-enhanced CT multiple osteolytic changes | 24
thrombi splenic vein | 24
thrombi inferior vena cava | 24
thrombi left common iliac vein | 24
SpO2 94% with 5 L/min oxygen | 24
non-invasive positive-pressure ventilation | 24
diuretic administration | 24
transferred to Division of General Medicine | 72
conscious | 72
well-oriented | 72
left hip pain | 72
body temperature 37.1°C | 72
pulse rate 93 beats/min | 72
blood pressure 126/82 mmHg | 72
respiratory rate 25 breaths/min | 72
SpO2 96% with 5 L/nasal cannula | 72
conjunctiva anemia | 72
conjunctiva icteric | 72
rubbery hard lymph nodes | 72
respiratory sounds attenuated bilateral lower lung | 72
bilateral breast engorgement | 72
midline Caesarean scar | 72
WBC 11,470/μL | 72
hemoglobin 7.7 g/dL | 72
hypoalbuminemia 2.1 g/dL | 72
lactate dehydrogenase 4,467 units/L | 72
alkaline phosphatase 1,651 units/L | 72
carcinoembryonic antigen 44.0 ng/dL | 72
carbohydrate antigen 19-9 154.7 U/mL | 72
carbohydrate antigen 125 243.6 U/mL | 72
carbohydrate antigen 15-3 55 U/mL | 72
pleural fluid adenocarcinoma | 168
sputum cytology adenocarcinoma | 168
upper gastrointestinal endoscopy unremarkable | 168
colonoscopy unremarkable | 168
breast ultrasonography unremarkable | 168
placenta normal | 168
stopped breastfeeding | 168
SpO2 deterioration | 312
oxygen therapy changed to nasal high-flow | 312
pleural effusion cell block adenocarcinoma | 312
CK7 positive | 312
thyroid transcription factor-1 positive | 312
napsin A positive | 312
EGFR exon 19 deletion | 408
gefitinib initiated | 408
transferred to Division of Respiratory Medicine | 480
pleural effusion reduced | 480
SpO2 improved | 480
discharged | 1080
outpatient treatment | 1080
ambulatory | 1080
