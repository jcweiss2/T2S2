23 years old | -720
pregnant | -720
Caucasian | -720
female | -720
referred for fetal echocardiogram | -720
congenital heart disease | -720
obstetric anatomy scan | -720
maternal medical history unremarkable | -720
family history unremarkable | -720
fetal echocardiogram | -720
DORV | -720
normally related great arteries | -720
remote VSD | -720
moderate to severe hypoplastic mitral valve | -720
hypoplastic left ventricle | -720
APV | -720
to-and-fro flow | -720
dysplastic and rudimentary pulmonary valve tissue | -720
moderate degree of stenosis | -720
peak velocity 3.0 m/s | -720
severely dilated main and branch pulmonary arteries | -720
right ventricular systolic function below normal | -720
no evidence of ductus arteriosus | -720
counseled regarding complex diagnosis | -720
poor prognosis | -720
polyhydramnios | -720
amnioreduction | -720
genetic analysis of amniotic fluid | -720
22q11.2 deletion | -720
DiGeorge syndrome | -720
delivered at 36 weeks gestation | 0
cesarean section | 0
breech position | 0
premature rupture of membranes | 0
severe polyhydramnios | 0
birth weight 2300 grams | 0
cyanotic | 0
apneic | 0
intubation | 0
initial blood gas pH 7.17 | 0
pCO2 69 | 0
pO2 21 | 0
oxygen saturations 70% | 0
hypoxic | 0
100% fractional inspired oxygen | 0
inhaled nitric oxide | 0
prone positioning | 0
dysmorphic features | 0
22q.11 deletion | 0
to-and-fro murmur | 0
cardiac auscultation | 0
postnatal transthoracic echocardiogram | 0
DORV | 0
sub-aortic VSD | 0
side-by-side great arteries | 0
aortic-mitral fibrous discontinuity | 0
severely hypoplastic mitral valve | 0
minimal antegrade flow | 0
hypoplastic left ventricle | 0
non-apex forming | 0
aortic valve leaflets thickened | 0
dysplastic | 0
normal annular measurements | 0
valve annulus 0.9 cm | 0
aortic sinuses 1.22 cm | 0
no evidence of coarctation of aorta | 0
aortic isthmus 0.4 cm | 0
pulmonary valve leaflets dysplastic | 0
rudimentary | 0
mild valvar stenosis | 0
severe/free insufficiency | 0
to-and-fro flow | 0
main pulmonary artery severely dilated | 0
branch pulmonary arteries severely dilated | 0
left pulmonary artery 7.5 mm | 0
right pulmonary artery 8 mm | 0
right ventricle dilated | 0
hypertrophied | 0
severely depressed systolic function | 0
partially restrictive atrial septum | 0
left to right shunting | 0
refractory cardiogenic shock | 0
severe hypoxemia | 0
surgical intervention | 12
atrial septectomy | 12
branch pulmonary artery plication | 12
over sewing of main pulmonary artery | 12
placement of right 3.5 mm modified Blalock-Taussig-Thomas shunt | 12
failed to separate from cardiopulmonary bypass | 12
extracorporeal membrane oxygenator support | 12
hemothorax | 24
acute kidney injury | 24
continuous renal replacement therapy | 24
profoundly immunocompromised | 24
severe lymphopenia | 24
hypogammaglobinemia | 24
DiGeorge syndrome | 24
septic shock | 24
Serratia marcescens septicemia | 24
abdominal compartment syndrome | 24
abdominal decompression | 24
washout | 24
multi-organ failure | 24
profound neurological impairment | 24
comfort care | 24
died | 744