7 years old | 0
male | 0
admitted with generalized convulsive status epilepticus | 0
high fever | -96
diffuse skin rash | -96
right tibia fracture | -336
seizure | 0
maculopapular rash on face, trunk, extremities | 0
nonpurulent conjunctivitis | 0
cracked, fissured lips | 0
cervical lymphadenopathy | 0
fever of 39°C | 0
negative meningeal signs | 0
Glasgow Coma Scale score 7 | 0
elevated ESR (68 mm/1 h) | 0
elevated CRP (29.6 mg/l) | 0
procalcitonin 0.63 ng/ml | 0
leukocytes 6.8x10^9/l | 0
erythrocytes 4.24x10^12/l | 0
hemoglobin 121 g/l | 0
platelets 181x10^9/l | 0
blood urea nitrogen 5.3 mmol/l | 0
serum creatinine 47.1 umol/l | 0
elevated aspartate transaminase (2.9 ukat/l) | 0
elevated alanine transaminase (2.050 ukat/l) | 0
gamma-glutamyl transferase 0.170 ukat/l | 0
lactate dehydrogenase 11.27 lakatl | 0
CSF WBC 1/mm3 | 0
CSF protein 225 mg/dl | 0
CSF glucose 4.84 mmol/l | 0
chloride 118.0 mmol/l | 0
lactate 2.5 mmol/l | 0
negative blood, CSF, urine cultures | 0
negative serological tests for viruses | 0
positive IgG antibodies to cytomegalovirus, adenovirus | 0
normal CT scan of brain | 0
normal chest X-ray | 0
normal ECG | 0
normal transthoracic echocardiogram | 0
normal cardiac markers | 0
cervical lymph nodes 15 mm bilaterally | 0
EEG showing cerebral dysfunction | 0
admitted to Intensive Care Unit | 0
treated with phenobarbital | 0
treated with ceftriaxone | 0
treated with acyclovir | 0
osmotic therapy with mannitol | 0
febrile on 2nd day | 24
impaired consciousness (GCS 6) | 24
respiratory failure | 24
intubation | 24
mechanical ventilation | 24
brain MRI showing cerebral edema | 24
narrowings of middle cerebral artery | 24
diagnosed with Kawasaki disease | 24
cerebral vasculitis | 24
encephalitis | 24
IVIG therapy started | 24
acetylsalicylic acid started | 24
fever resolved | 48
skin rash disappearance | 48
mild consciousness improvement | 48
extubated on 3rd day | 72
acyclovir discontinued | 72
confusion | 72
irritability | 72
delirium | 72
GCS 8-10 | 72
recurrent fever | 72
brain MRI progression on 6th day | 144
steroid pulse therapy started on 9th day | 216
oral prednisolone started | 216
neurological improvement | 216
full motor recovery on 15th day | 360
cognitive improvement | 360
periungual desquamation in 3rd week | 504
normal repeated echocardiogram | 504
discharged after 45 days | 1080
normal cognitive functions at discharge | 1080
corticosteroids tapered and stopped after 3rd month | 2160
follow-up MRI normalization | 1440
parenchymal atrophy | 1440
cerebral circulation normalization | 1440
no antiepileptic drugs used | 1080
negative follow-up MRI after 2 months | 1440
