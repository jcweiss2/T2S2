70 years old | 0
    female | 0
    hereditary hemorrhagic telangiectasia | 0
    severe pulmonary hypertension | 0
    diastolic heart failure | 0
    mild obstructive sleep apnea | 0
    hyperlipidemia | 0
    gastroesophageal reflux | 0
    hypertension | 0
    scheduled for open radical nephrectomy | 0
    left kidney en bloc removal | 0
    5.4-cm mass localized to the lower pole | 0
    concerning for malignancy | 0
    severe exertional dyspnea three years prior | -26208
    left and right heart catheterization | -26208
    angiographically normal-appearing coronary arteries | -26208
    right coronary artery fistula | -26208
    severe precapillary pulmonary hypertension | -26208
    mean pulmonary artery pressure of 45 mmHG | -26208
    pulmonary capillary wedge pressure 8 mmHG | -26208
    pulmonary vascular resistance 7.8 WU | -26208
    cardiac index 3.0 L/min/m2 | -26208
    started on sildenafil | -26208
    WHO class III symptoms improved to class I or II | -26208
    transthoracic echocardiogram | -26208
    RV enlargement | -26208
    decreased RV function | -26208
    moderate-to-severe eccentric TR | -26208
    moderately-to-severely dilated right atrium | -26208
    Doppler-derived estimated systolic pulmonary artery pressure >100 mmHg | -26208
    low normal left ventricular function | -26208
    pulmonary function testing | -26208
    normal volumes | -26208
    spirometry | -26208
    normal forced vital capacity | -26208
    normal forced expiratory volume | -26208
    normal FEV1/FVC ratio | -26208
    severely reduced diffusing capacity (43% of predicted) | -26208
    frequent epistaxis | 0
    episodes of gastrointestinal bleeding | 0
    arterial venous malformations | 0
    previous intervention with nasal endoscopy | 0
    previous intervention with upper-gastrointestinal endoscopy | 0
    mild OSA treated with CPAP | 0
    heart failure with preserved ejection fraction | 0
    anemia | 0
    30-pound weight loss | 0
    synthetic liver dysfunction | 0
    elevated PT INR | 0
    low albumin | 0
    multidisciplinary perioperative consultation | 0
    risks discussed | 0
    benefits discussed | 0
    alternatives discussed | 0
    increased risk due to severe pulmonary hypertension | 0
    patient consented to proceed with surgery | 0
    likelihood for malignant renal cell carcinoma | 0
    ASA physical status IV | 0
    preoperative transthoracic echocardiography | 0
    chest x-ray | 0
    cardiovascular silhouette at the upper limits of normal | 0
    prominent pulmonary arteries | 0
    continued sildenafil | 0
    good response to sildenafil | 0
    exercise tolerance greater than 4 METS | 0
    partial vs. radical nephrectomy discussed | 0
    elected to have entire left kidney removal | 0
    minimal dyspnea with daily activities | 0
    occasional lightheadedness during exertion | 0
    no angina | 0
    denied significant orthopnea | 0
    denied paroxysmal nocturnal dyspnea | 0
    no significant edema | 0
    no hepatosplenomegaly | 0
    frequent epistaxis episodes secondary to HHT | 0
    1:1 mixing study | 0
    elevated PT/INR of 1.3 | 0
    ordered oral vitamin K | 0
    outpatient workup | 0
    no evidence of decompensated liver disease | 0
    low-grade fibrosis on fibroscan | 0
    continued ferrous sulfate | 0
    continued Lasix | 0
    continued omeprazole | 0
    continued albuterol | 0
    admitted on the day of surgery | 0
    temperature 36.6 C | 0
    blood pressure 138/77 mmHG | 0
    respiratory rate 18/min | 0
    pulse oximetry 96% on room air | 0
    pain 0/10 | 0
    reassuring airway exam | 0
    no bleeding episodes other than frequent epistaxis | 0
    denied new or worsening shortness of breath | 0
    denied chest discomfort | 0
    ECG normal sinus rhythm | 0
    rate 95 | 0
    premature ventricular complexes | 0
    inferior and anterolateral T-wave changes | 0
    hemoglobin 11.2 g/dl | 0
    hematocrit 35.4% | 0
    large-bore IV access | 0
    radial arterial line | 0
    induction of general anesthesia | 0
    supine position | 0
    standard ASA monitors | 0
    adequate pre-oxygenation | 0
    administered IV fentanyl | 0
    administered etomidate | 0
    administered lidocaine | 0
    administered rocuronium | 0
    intubated with 7.0-mm endotracheal tube | 0
    Cormack-Lehane grade I view | 0
    no telangiectasias observed during direct laryngoscopy | 0
    confirmed endotracheal tube position | 0
    stable pulse oximetry | 0
    stable heart rate | 0
    stable arterial blood pressure | 0
    Swan-Ganz catheter placed | 0
    right internal jugular venous 9 fr introducer | 0
    initial pulmonary artery pressure 96/46 mmHG | 0
    mean pulmonary artery pressure 65 mmHG | 0
    systemic arterial pressure 125/74 mmHG | 0
    arterial blood gas pH 7.33 | 0
    pCO2 43 mmHG | 0
    pO2 145 mmHG | 0
    HCO3 22.7 mEq/L | 0
    correction of hypercarbia | 0
    correction of mild acidosis | 0
    initiated inhaled nitric oxide 20 ppm | 0
    improvement in pulmonary artery pressures | 0
    nadir pulmonary artery pressure 67/29 mmHG | 0
    mean pulmonary artery pressure 44 mmHG | 0
    systemic arterial pressure 123/67 mmHG | 0
    fluid balance maintained | 0
    adequate urine output | 0
    blood loss less than 100 cc | 0
    transversus abdominal plane block | 0
    ultrasound guidance | 0
    1:1 mixture of 0.25% bupivacaine and 1.3% liposomal bupivacaine | 0
    total 20 cc local infiltration | 0
    general anesthesia maintained with sevoflurane | 0
    surgical time less than 60 min | 0
    right lateral decubitus position | 0
    flank incision | 0
    hemodynamically stable on inhaled nitric oxide | 0
    final arterial blood gas pH 7.38 | 0
    pCO2 38 mmHG | 0
    pO2 182 mmHG | 0
    50% FiO2 | 0
    transferred to surgical intensive care unit | 0
    inhaled nitric oxide weened over 3 h | 0
    pulmonary artery pressures reached baseline | 0
    cardiac output 3–4 L/min | 0
    no evidence of pulmonary arterial crisis | 0
    extubated on postoperative day 0 | 24
    noninvasive positive pressure ventilation | 24
    weened to nasal cannula | 24
    pulse oximetry saturation 93–96% | 24
    numerical rating scale <4 | 24
    multimodal pain regimen | 24
    PO acetaminophen | 24
    IV acetaminophen | 24
    Ultram | 24
    incremental doses of fentanyl | 24
    return of bowel function | 24
    no nasogastric tube | 24
    tolerated oral diet within 24 h | 24
    transferred to step-down unit on postoperative day 1 | 48
    ambulated with assistance | 48
    discharged to home on postoperative day 3 | 72
    renal cell carcinoma | 72
    clear cell type | 72
    high-grade histologic pathology | 72
    classification pT1bG4 | 72
    clear margins | 72
    resumed normal daily activities | 72
    turned 71 years old during hospitalization | 72
    <|eot_id|>
    