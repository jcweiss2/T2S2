2-month-old | 0
male | 0
admitted to the hospital | 0
mild cough | -24
fever (37.8°C) | -24
malaise | -24
close contact with brother with cold | -24
born very preterm (31 weeks + 5 days) | -1344
low birth weight (1700 grams) | -1344
hospitalized for 25 days after birth | -1344
neonatal pneumonia | -1344
coagulation dysfunction | -1344
intracranial hemorrhage (grade I, absorption phase) | -1344
neonatal pathological jaundice | -1344
vaccinated with Bacillus Calmette-Guerin | -1344
mask oxygen inhalation | -24
piperacillin tazobactam | -24
ambroxol | -24
budesonide + ipratropium bromide atomization | -24
clinical symptoms deteriorated rapidly | -24
tachypnea | -24
low oxygen saturation | -24
transferred to PICU | -24
body temperature 37.3°C | 0
heart rate 172 beats per minute | 0
respiratory rate 56 breaths per minute | 0
blood pressure 96/50 mmHg | 0
puffy nose | 0
triple concave signs | 0
mild cyanosis of the lips | 0
Glasgow Coma Score 13 (E4, V3, M6) | 0
oxygen saturation 93% with oxygen mask | 0
pulmonary auscultation rough breath sounds | 0
wheezing in both lungs | 0
umbilical hernia | 0
anterior fontanelle bulge | 0
low response | 0
screaming after stimulation | 0
chest CT scan multiple plaques, streaks, solid shadows, indistinct reticular shadows in both lungs | 0
brain MRI bilateral frontal, parietal, temporal extracranial spaces slightly wider | 0
no obvious abnormality in brain parenchyma | 0
echocardiography no abnormalities | 0
hemoglobin 84 g/L | 0
red blood cell count 3.05 ×10^12/L | 0
white blood cell count 6.5 ×10^9/L | 0
neutrophil count 3.59 ×10^9/L | 0
lymphocyte count 2.16 ×10^9/L | 0
platelet count 280 ×10^9/L | 0
liver function normal | 0
kidney function normal | 0
respiratory failure | 0
severe pneumonia | 0
septic shock | 0
encephalopathy | 0
meropenem | 0
vancomycin | 0
levetiracetam | 0
deterioration after 3 hours in PICU | 3
worsening dyspnea | 3
groans | 3
gray face | 3
cold limbs | 3
speckles all over the body | 3
bilateral crackles | 3
capillary refill time 5 seconds | 3
oxygen saturation 54% | 3
lactate level 7.07 mmol/L | 3
procalcitonin 14.29 ng/mL | 3
invasive ventilator-assisted ventilation | 3
norepinephrine | 3
mannitol | 3
fructose glycerol | 3
immunoglobulin | 3
fresh frozen plasma | 3
viral nucleic acid in BALF negative | 0
respiratory syncytial virus negative | 0
parainfluenza virus 1 negative | 0
parainfluenza virus 2 negative | 0
parainfluenza virus 3 negative | 0
human adenovirus negative | 0
influenza A negative | 0
influenza B negative | 0
human metapneumovirus negative | 0
rhinovirus negative | 0
boca virus negative | 0
novel coronavirus negative | 0
Mycoplasma pneumoniae serology negative | 0
Chlamydia trachomatis serology negative | 0
cytomegalovirus IgM negative | 0
cytomegalovirus IgG negative | 0
sputum bacterial cultures negative | 0
tuberculin test negative | 0
Bordetella pertussis detected in nasopharyngeal specimen | 0
CSF assay normal | 0
CSF cultures negative | 0
blood m-NGS detected Bordetella pertussis | 0
CSF m-NGS detected Bordetella pertussis | 0
levofloxacin initiated | 48
chest x-ray inflammation gradually absorbed | 288
weaned off mechanical ventilation | 312
discharged | 888
