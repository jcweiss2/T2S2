45 years old | 0
    female | 0
    acute emergency presentation | 0
    severe lower abdominal pain | -12
    bright red per rectal bleeding | -12
    rapid deterioration | -12
    worsening pain | -12
    tachycardia | -12
    high-grade fevers | -12
    right-sided colon cancer diagnosis | -8760
    pelvic side wall lymph node metastases | -8760
    surgery with curative intent | -8760
    R0 resection | -8760
    radiotherapy to pelvis | -168
    adjuvant FOLFOX chemotherapy | -168
    schizophrenia | -8760
    Clozapine 300 mg daily | -8760
    severe constipation | 0
    chemotherapy adverse effects | 0
    nausea | 0
    abdominal discomfort | 0
    constipation | 0
    CT abdomen pelvis | 0
    large volume of pneumoperitoneum | 0
    massive sigmoid faecaloma | 0
    stercoral perforation | 0
    ischaemic changes | 0
    emergency laparotomy | 0
    grossly dilated sigmoid colon | 0
    redundant sigmoid colon | 0
    inspissated faecaloma | 0
    perforation mid to distal sigmoid colon | 0
    necrosis of the wall | 0
    Hartmann’s procedure | 0
    extensive washout | 0
    vasopressor support | 0
    septic shock | 0
    granulocyte colony stimulating factor | 0
    febrile neutropaenia | 0
    Clozapine suspended | 0
    G-CSF given | 0
    neutropenia improved | 0
    recovery post-operatively | 0
    discharged to rehabilitation | 240
    histopathology confirmation | 0
    full thickness perforation | 0
    ischaemic necrosis of mucosa | 0
    massive faecaloma | 0
    stercoral perforation diagnosis | 0
    comorbidities | 0
    adjuvant chemotherapy | 0

