42 years old| 0
    male| 0
    admitted to the intensive care unit| 0
    febrile neutropenia| 0
    septic shock from Escherichia coli bacteremia| 0
    severe anemia| 0
    hemoglobin of 5.1 g/dL| 0
    platelet count of 2 k/uL| 0
    blood transfusions| 0
    platelet transfusions| 0
    respiratory failure| 0
    mechanical ventilation| 0
    blood pressure support with four vasopressors| 0
    intravenous methylprednisolone| 0
    meropenem| 0
    hematemesis| 480
    drop in hemoglobin| 480
    pantoprazole drip| 480
    upper endoscopy| 480
    blood clots in the fundus| 480
    blood clots in the upper body| 480
    ulcers in the gastric antrum| 480
    ulcers in the gastric body| 480
    normal esophagus| 480
    normal duodenum| 480
    chronic active gastritis| 480
    foveolar hyperplasia| 480
    repeat endoscopy| 504
    IV erythromycin| 504
    multiple ulcers| 504
    large blood clot in the fundus| 504
    mesenteric angiography| 504
    empiric left gastric artery embolization| 504
    continued hematemesis| 504
    dropping hemoglobin| 504
    exploratory laparotomy| 504
    distended stomach| 504
    blood filled stomach| 504
    multiple deep ulcerations| 504
    total gastrectomy| 504
    esophagojejunostomy| 504
    jejunostomy tube placement| 504
    hemorrhagic ulcers| 504
    deep ulcerations| 504
    broad aseptate fungi| 504
    variable angle branching| 504
    angioinvasion| 504
    Warthin Starry stain negative for Helicobacter pylori| 504
    immunostaining negative for CMV| 504
    hemodynamically stable| 504
    titrated off blood pressure support medications| 504
    extubated| 504
    sputum cultures grew Aspergillus fumigatus| 504
    amphotericin B| 504
    voriconazole| 504
    PCR revealed Mycotypha microspora| 504
    renal failure| 504
    switched to isavuconazole| 504
    discharged| 504
    posaconazole| 504
    micafungin| 504
    germ cell tumor of the mediastinum| -504
    hemorrhagic pituitary prolactinoma| -504
    left middle cerebral artery thrombotic stroke| -504
    Etoposide| -504
    Ifosfamide| -504
    Cisplatin| -504
    last dose a week before emergency room visit| -168
    prolactinoma controlled on Cabergoline| -504
    lethargy| 0
    extreme weakness| 0
    <|eot_id|>
    