73 years old | 0
established renal failure of unknown cause | 0
poor vessels for primary or secondary vascular access | 0
admitted electively | 0
creation of first-stage brachiobasilic arteriovenous fistula | 0
transferred to haemodialysis | -672
peritoneal dialysis | -672
episode of peritonitis | -672
laparotomy | -672
attempts at re-initiating peritoneal dialysis | -672
unsuccessful | -672
dialysing via tunnelled jugular central venous catheter | -672
jugular catheter in situ for 14 months | -672
co-morbidities | 0
previous metallic mitral valve replacement | 0
requiring therapeutic anticoagulation | 0
hypertension | 0
haematuria of unknown cause | 0
native kidneys never biopsied | 0
medically unfit for renal transplantation | 0
developed diarrhoea | -168
rigours post-dialysis | -168
complained of pain around her line | -168
treatment instigated for presumed catheter-associated bacteraemia | -168
remained septic | -168
swinging fevers | -168
one splinter haemorrhage | -168
new murmur noted | -168
possible vegetation on mitral valve on echocardiogram | -168
blood cultures positive for fully sensitive Staphylococcus aureus | -168
multiple screens for MRSA negative | -168
clinical diagnosis of infective endocarditis | -168
appropriate treatment administered | -168
treatment for endocarditis with antibiotics | -168
continued for next 4 weeks | -168
appeared to respond well | -168
represented feeling non-specifically unwell | -168
routine observations normal | -168
blood investigations normal | -168
rapidly deteriorated | -168
lactic acidosis | -168
complained of mild lower abdominal pain | -168
abdomen soft | -168
no evidence of peritonitis | -168
medical condition continued to deteriorate | -168
developed fast, uncontrolled atrial fibrillation | -168
arterial blood gas pH 7.13 | -168
pO2 103 mmHg | -168
pCO2 17.3 mmHg | -168
lactate 13.3 mmol/L | -168
contrast-enhanced CT angiogram patent celiac and superior mesenteric artery axis | -168
patent portal vein | -168
features consistent with chronic pyelonephritis | -168
possible inflammation in gallbladder fossa | -168
inflammatory oedema in Morrison’s pouch | -168
transferred to intensive care unit | -168
resuscitated | -168
intubated | -168
ventilated | -168
remained haemodynamically stable | -168
metabolic acidosis progressively worsened | -168
arterial lactic acid increased to 20 mmol/L | -168
emergency laparotomy performed | -168
sero-purulent fluid in Morrison’s pouch | -168
macro-nodular liver | -168
normal gallbladder | -168
stomach normal | -168
duodenum normal | -168
pancreas normal | -168
small bowel normal | -168
colon normal | -168
extensive inflammatory change around right kidney | -168
nephrectomy performed | -168
transferred back to intensive care unit | -168
haemofiltered for 4 hours | -168
made speedy recovery | -168
arterial lactic acid returned to normal | -168
discharged to ward | 48
pathology chronic pyelonephritis | 48
sclerosis of glomeruli | 48
atrophy of tubules | 48
cystic dilation containing polymorphs | 48
chronic inflammation | 48
fibrosis of parenchyma | 48
no evidence of renal stones | 48
arterioles hypertensive change | 48
final diagnosis chronic pyelonephritis with peri-renal sepsis | 48
liver biopsy congestive hepatomegaly | 48
discussion peri-renal sepsis | 48
chronic renal failure | 48
emergency nephrectomy | 48
overwhelming MRSA urosepsis | 48
stag horn calculus | 48
pyelonephritis accounts for 3–4 hospital admissions per 10,000 females | 48
normal renal function | 48
incidence in chronic pyelonephritis unknown | 48
chronic kidney disease anuric | 48
diagnosis of renal or peri0-renal sepsis difficult | 48
cross-sectional imaging inconclusive | 48
worsening abdominal pain | 48
severe lactic acidosis | 48
no peritonitis | 48
major intra-abdominal vascular event | 48
metastatic sepsis from infective endocarditis | 48
source of sepsis | 48
absence of common conditions causing acute abdomen | 48
obscure renal or peri-renal sepsis considered | 48
surgical management with nephrectomy necessary | 48
