48 years old | 0
woman | 0
presented to the emergency department | 0
left breast enlargement | -8760
black discoloration of breast skin | -8760
fever | -8760
loss of appetite | -8760
weight loss | -8760
diabetes mellitus | -8760
hypertension | -8760
left breast swollen | 0
dark discoloration of skin | 0
multiple small punched-out ulcers | 0
discharging purulent material | 0
nipple retracted | 0
breast tender | 0
breast warm | 0
breast firm on palpation | 0
left axillary lymph node palpable | 0
marked leukocytosis | 0
prolongation of coagulation profile markers | 0
MRSA positive wound culture | 0
MRSA positive blood culture | 0
emergency surgery | 0
simple mastectomy | 0
died | 48
disseminated intravascular coagulation | 48
septicemia secondary to MRSA | 48
no autopsy | 48
PB-ALCL, giant cell-rich pattern diagnosis | 0
CD30 positive | 0
CD45 positive | 0
CD45RO positive | 0
granzyme B positive | 0
TIA-1 positive | 0
vimentin positive | 0
CD4 positive | 0
CD43 positive | 0
EMA positive | 0
BCL-6 positive | 0
BCL-2 positive | 0
loss of CD1a | 0
loss of CD3 | 0
loss of CD5 | 0
loss of CD8 | 0
loss of CD7 | 0
loss of CD2 | 0
CD20 negative | 0
CD19 negative | 0
CD79a negative | 0
PAX-5 negative | 0
ALK-1 negative | 0
CD15 negative | 0
CD68 negative | 0
pancytokeratins negative | 0
S100 protein negative | 0
desmin negative | 0
SMA negative | 0
HMB-45 negative | 0
P63 negative | 0
E-cadherin negative | 0
MIB-1 (Ki-67) labeling index high (95%) | 0
no previous history of lymphoma | 0
no breast implant | 0
no family history of breast cancer | 0
no family history of lymphoma | 0
no radiological studies | 0
no epidermotropism | 0
no involvement of atrophic ducts and lobules | 0
no autolysis study | 48
So creating the table with events and timestamps separated by |.
