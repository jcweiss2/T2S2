60 years old | 0
female | 0
T2b, N1, M0 squamous cell carcinoma of the right lung | -96
pneumonectomy | -96
mediastinal lymphadenectomy | -96
discharged home | -80
progressive dyspnea | -64
denies cough | -64
denies wheezing | -64
denies chest pain | -64
denies fevers | -64
emergency intubation | -64
intubated | -64
sedated | -64
hypotensive | -64
tachycardic | -64
right pneumonectomy wound site healing well | -64
right thorax dull to percussion | -64
absent right-sided breath sounds | -64
cardiac point of maximal impulse shifted toward the left | -64
tracheal deviation towards the left | -64
cardiac auscultation normal | -64
right lower extremity leg swelling | -64
central line placed | -64
central venous pressure 18 cm H2O | -64
elevated leukocytes | -64
mild normocytic anemia | -64
creatinine 1.8 mg/dL | -64
mild hyperkalemia | -64
elevated lactate | -64
undetectable troponin | -64
complete right hemithorax opacification | -64
left-shift of the mediastinum | -64
moderate left pleural effusion | -64
no pulmonary embolus | -64
severe biatrial compression | -64
no tamponade | -64
no restrictive physiology | -64
no pericardial effusion | -64
normal right and left ventricular function | -64
right distal leg deep venous thromboses | -64
urgent bedside decompressive chest tube placement | -64
bilateral effusions | -64
left chest drained | -64
pleural fluid milky white | -64
elevated triglycerides 1729 mg/dL | -64
hemodynamics improved | -56
came off pressors | -56
extubated | -56
diagnosis of tension chylothorax | -56
lymphangiography | -48
no site of thoracic duct leak | -48
left-sided pleural drainage less than 500 cc/day | -40
clinical status improved | -40
surgical exploration not indicated | -40
pigtail catheter placed in right chest | -40
right hemithorax irrigated with antibiotic solution | -40
right-sided chylothorax secondary to lymphatic leakage | -40
left-sided chylothorax secondary to mediastinal transit of chyle | -40
complete parenteral nutrition started | -40
chest tube drainage monitored | -40
chest drain output decreased | -24
transitioned to medium chain triglyceride diet | -24
no increase in chest drain output | -16
right pigtail catheter removed | -4
left chest tube removed | 0
discharged home | 8
right leg deep venous thrombosis treated with intravenous heparin | -64
heparin-induced thrombocytopenia with thrombosis | -24
alternative parenteral anticoagulation | -24
retrievable inferior vena cava filter placed | -24
discharged home on rivaroxaban | 8
tolerating regular diet without evidence of recurrent chylothorax | 384
completed adjuvant chemotherapy | 384