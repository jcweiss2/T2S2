59 years old | 0
male | 0
complaining of sudden chest pain | -1
collapsed in the ambulance | -1
cardiopulmonary resuscitation | -1
ventricular fibrillation | -1
return of spontaneous circulation | -1
admitted to the hospital | 0
blood pressure 105/78 mm Hg | 0
heart rate 120 beats/min | 0
respiratory rate 20 breaths/min | 0
body temperature 35.8°C | 0
diagnosed with ST-segment elevation myocardial infarction | 0
electrocardiogram | 0
cardiac arrest | 0
veno-arterial ECMO | 0
percutaneous coronary intervention | 0
thrombectomy | 0
sedated using remifentanil | 0
sedated using propofol | 0
hemodynamic status improved | 72
oxygenation improved | 72
VA ECMO decannulation | 72
progressive acute kidney injury | 120
continuous renal replacement therapy | 120
veno-venous ECMO | 168
severe acute respiratory distress syndrome | 168
hospital-acquired pneumonia | 168
weaned off VV ECMO | 384
clinical improvement of pneumonia | 384
agitation | 384
ventilator dyssynchrony | 384
vasopressors tapered | 384
alanine aminotransferase increased | 432
aspartate aminotransferase increased | 432
bundle branch block | 480
increased creatinine kinase | 480
increased CK-MB | 480
increased troponin I | 480
hypotension | 480
increased infusion rate of norepinephrine | 480
increased infusion rate of epinephrine | 480
added vasopressin | 480
acute renal failure | 480
metabolic acidosis | 480
propofol infusion discontinued | 480
propofol-related infusion syndrome suspected | 480
initial serum triglyceride level 369 mg/dl | 0
cortisol level normal | 0
thyroid function tests normal | 0
requirement for vasopressors decreased | 504
vasopressin tapered | 504
CK level continued to elevate | 504
L-carnitine administration started | 552
CK level gradually declined | 576
patient stabilized | 576
discharged from ICU | 1224
transferred to a nursing hospital | 2208