69 years old | 0
male | 0
height 170 cm | 0
weight 80 kg | 0
scheduled for repeated arthroscopic lavage of the right knee | 0
septic arthritis | -336
previous arthroscopic lavage | -336
peripheral arterial occlusive disease | -336
hypertension | 0
type 2 diabetes | 0
atrial fibrillation | -336
flecainide | -336
aspirin | -336
preoperative electrocardiogram | 0
normal sinus rhythm | 0
glycopyrrolate | 0
anesthesia induced | 0
propofol | 0
rocuronium | 0
endotracheal tube | 0
electrocardiogram | 0
pulse oxygen saturation | 0
capnogram | 0
esophageal temperature | 0
invasive arterial pressure | 0
sevoflurane | 0
nitrous oxide | 0
arterial blood gas analysis | 10
pH 7.38 | 10
PaCO2 45.1 mmHg | 10
PaO2 85.7 mmHg | 10
HCO3- 26.0 mEq/L | 10
SaO2 95.5% | 10
FiO2 0.5 | 10
end tidal CO2 24 mmHg | 10
tidal volume increased | 10
arterial blood gas analysis | 30
pH 7.31 | 30
PaCO2 47.0 mmHg | 30
PaO2 75.1 mmHg | 30
HCO3- 23.6 mEq/L | 30
SaO2 92.8% | 30
FiO2 0.5 | 30
phenylephrine | 30
blood pressure dropped | 40
heart rate increased | 40
epinephrine | 40
peinephrine | 40
atropine sulfate | 40
vital signs deteriorated | 40
pulsatile activity disappeared | 40
cardiopulmonary resuscitation | 40
surgery completed | 40
nitrous oxide turned off | 40
sevoflurane turned off | 40
epinephrine | 40
atropine sulfate | 40
arterial blood gas analysis | 48
pH 7.37 | 48
PaCO2 27.8 mmHg | 48
PaO2 63.9 mmHg | 48
HCO3- 15.8 mEq/L | 48
SaO2 90.8% | 48
FiO2 1.0 | 48
external cardiac massage stopped | 48
arterial blood gas analysis | 56
pH 6.96 | 56
PaCO2 63.9 mmHg | 56
PaO2 221.4 mmHg | 56
HCO3- 13.9 mEq/L | 56
SaO2 98.5% | 56
FiO2 1.0 | 56
transthoracic echocardiogram | 50
massive pulmonary embolism | 50
thrombus in right atrium | 50
dilated hypokinetic right ventricle | 50
D-shaped left ventricle | 50
alteplase | 77
recombinant tissue-type plasminogen activator | 77
hemodynamic performance stabilized | 77
no sign of bleeding | 77
external cardiac massage stopped | 103
intensive care unit | 103
blood pressure increased | 103
heart rate | 103
mechanical ventilation | 103
heparin | 115
PT INR 1.65 | 115
aPTT 50-70 seconds | 115
consciousness became alert | 127
endotracheal tube extubated | 127
thrombi disappeared | 159
dilated hypokinetic right ventricle returned to normal | 159
heparin infusion stopped | 215
patient recovered | 215
transferred to medical ward | 215