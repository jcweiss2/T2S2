6 years old | 0
male | 0
fatigue | -120
looks pale | -120
shock | 0
altered consciousness (GCS 12) | 0
heart rate of 135 beats per minute | 0
blood pressure 70/40 mmHg | 0
respiratory rate 40 breaths per minute | 0
temperature 36.5oC | 0
prolonged capillary refill time >2 s | 0
oxygen saturation 83% | 0
receiving oxygen 5 L/minutes via simple mask | 0
no enlargement of the spleen | 0
no enlargement of the liver | 0
fluid resuscitation | 0
transfusion | 0
hemodynamic monitoring | 0
inotropic agent administration | 0
orotracheal intubation | 0
fever | -120
abdominal pain | -120
no history of cough | -120
no breathing difficulties | -120
no bleeding | -120
no rashes | -120
no history of traveling | -120
no contact with COVID-19 patients | -120
active child | -48
symptoms abruptly worsened | -24
laboratory tests | 0
hemoglobin 2.9 g/dL | 0
hematocrit 9.3% | 0
leucocyte 18 × 10^3/μL | 0
basophil 0% | 0
eosinophil 0% | 0
neutrophil band 1% | 0
neutrophil segment 55% | 0
lymphocyte 33% | 0
monocyte 4% | 0
erythrocyte 1.13 × 10^12/L | 0
platelets counts 213 × 10^3/μL | 0
albumin 1.96 g/dL | 0
urea 46.2 g/dL | 0
serum creatinine (S-Cre) 1.15 mg/dL | 0
aspartate transaminase (AST) 510 U/L |0
alanine transaminase (ALT) 173 U/L |0
potassium 6 mmol/L |0
sodium 123 mEq/L |0
C-reactive protein (CRP) 0.09 mg/dL |0
procalcitonin 0.78 ng/mL |0
blood gas analysis pH 6.8 |0
pO2 24.2 mmHg |0
pCO2 27.2 mmHg |0
HCO3 4.8 mmol/L |0
TCO2 5.6 mmol/L |0
BE –2.78 mmol/L |0
SO2 17.3% |0
lactate dehydrogenase 10.6 mmol/L |0
peripheral blood smear normochromic erythrocytes |0
anisopoikilocytosis (ovalocyte, pencil cell) |0
microcytic |0
leukocytic hypersegmentation |0
serum iron 157 mcg/dL |0
Total Iron Binding Capacity (TIBC) 207 mcg/dL |0
ferritin 3985 ng/mL |0
rapid test SARS CoV-2 IgM reactive |0
SARS CoV-2 IgG non-reactive |0
PCR SARS CoV-2 negative |0
IgM anti-dengue reactive |0
IgG anti-dengue non-reactive |0
chest x-ray within normal limits |0
diagnosed with refractory septic shock |0
aggressive fluid resuscitation |0
broad-spectrum antibiotic administration |0
hemodynamic instability |0
multiple organ failure |0
passed away |14
