35 years old | 0
man | 0
history of active intravenous (IV) drug use (IVDU) | 0
presented to local emergency department | -336
back pain | -336
intermittent fever | -336
oral levofloxacin | -336
presented to hospital | 0
admitted | 0
severe back pain | 0
progressively worsening shortness of breath | 0
fatigue | 0
several-week history of fever | 0
blood pressure 129/65 mm Hg | 0
heart rate 110 beats/min | 0
temperature 102 °F | 0
respiratory rate 35 breaths/min | 0
transthoracic echocardiography (TTE) revealed vegetations on tricuspid valve | 24
necrotizing bilateral pneumonia | 48
large retropharyngeal abscess | 48
epidural abscess at T8-T9 | 48
spinal cord compression | 48
past medical history of active IVDU of methamphetamine | 0
chronic hepatitis C | 0
type 2 diabetes mellitus | 0
infective endocarditis (IE) suspected | 0
differential diagnoses included tuberculosis | 0
fungal infection | 0
systemic connective tissue diseases | 0
repeated blood cultures grew methicillin-sensitive Staphylococcus aureus (MSSA) | 384
transesophageal echocardiography revealed severe tricuspid regurgitation | 384
large, mobile vegetations attached to tricuspid valve | 384
right ventricular systolic pressure 50 mm Hg | 384
IV vancomycin | 0
IV ceftriaxone | 0
managed in intensive care unit (ICU) | 0
intubated on mechanical ventilator | 96
IV nafcillin | 96
multidisciplinary approach with otolaryngology and neurosurgery | 192
drainage of abscesses | 192
decompressive laminectomy | 192
bacteremia persisted through hospital day 16 | 384
cardiothoracic surgery consulted | 384
endovascular aspiration therapy recommended | 384
catheter-based aspiration therapy pursued | 384
intracardiac echocardiography (ICE) demonstrated large vegetations on tricuspid valve | 384
improvement in tricuspid valve regurgitation observed | 384
transferred to ICU | 384
successfully extubated | 408
discharged home | 624
IV ampicillin and sulbactam | 624
4-month follow-up echocardiography | 2880
mild tricuspid regurgitation | 2880
avoided tricuspid valve replacement surgery | 2880
