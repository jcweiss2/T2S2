69 years old | 0
male | 0
admitted to the hospital | 0
abdominal pain | -168
nausea-vomiting | -168
fever | -24
mental status change | -24
chronic renal disease | 0
primary hypertension | 0
diabetes mellitus | 0
history of coronary bypass surgery | 0
mildly elevated fever | 0
tachycardia | 0
normal blood pressure | 0
Glasgow coma scale score 11 | 0
tenderness in all four quadrants | 0
abdominal distension | 0
obstipation | -72
decreased bowel sounds | 0
empty rectum | 0
leukocytosis | 0
increased levels of serum C-reactive protein | 0
procalcitonin | 0
elevated creatinine | 0
elevated glucose | 0
elevated lactate | 0
abdominal ultrasound | 0
abdominal tomography | 0
duodenal perforation | 0
free air | 0
abscess in the retroperitoneal space | 0
prophylactic broad-spectrum antibiotics | 0
emergency surgery | 0
appendectomy | 0
drained the abscess | 0
inserted multiple drains | 0
no perforation area detected in the upper gastrointestinal tract | 0
cultures of the abscesses negative | 0
followed up in the intensive care unit | 0
septicemia | 0
discharged | 360
painful swelling | 360
fluctuation | 360
purulent discharge from the left side of his scrotum | 360
fistula orifice in the left scrotum | 360
abdominal tomography | 360
abscess cavity extending from the left retroperitoneal area to the left testis | 360
normal leukocyte | 360
increased levels of serum C-reactive protein | 360
procalcitonin | 360
lactate | 360
percutaneous drainage | 360
broad-spectrum antibiotics | 360
abscess culture negative | 360
control tomography | 377
abscess regressed | 377
discharged | 777