34 years old | 0
female | 0
admitted to the hospital | 0
septicemia | 0
superficial inflammation of the left thigh | 0
swelling of the left thigh | -48
chronic pain in the sacro-iliac joint | -336
oral antibiotic therapy (cefuroxime) | -48
temperature of 39.4°C | -24
increased inflammation parameters | 0
leukocytes 16,000/µL | 0
CRP 35 mg/dL | 0
spreading inflammation of the soft tissue (left thigh) | 0
i.v. drug abuse (heroin) | 0
hepatitis C | 0
computed tomography scan of abdomen and left thigh | 0
abscess of the sacro-iliac joint | 0
abscess of the psoas muscle | 0
magnetic resonance imaging (MRI) | 0
necrotizing fasciitis of the left thigh | 0
radical surgical debridement | 0
fasciectomy of the left thigh | 0
abscess of the sacroD iliac joint opened and drained | 0
transferred to intensive care unit | 0
antibiotic therapy (tobramycin, ceftriaxone, metronidazole) | 0
multiDresistant Pseudomonas aeruginosa infection | 0
VancomycinDresistant Enterococcus faecalis infection | 0
planned second revision with surgical debridement | 48
clean wound | 48
infection in the elbow | 0
open surgical debridement of elbow | 0
cerebral septic complications | 0
pulmonary septic complications | 0
five further sequential operations | 0
continuous vacuum therapy | 0
split skin graft | 0
intermittent hemodiafiltration | 0
septic acute renal failure | 0
Pseudomonas aeruginosa pneumonia | 0
antibiotic therapy (ceftazidime) | 0
tracheotomy | 168
returned to spontaneous breathing | 168
erythrocyte concentrates (16 units) | 0
thrombocyte concentrates (3 units) | 0
fresh frozen plasma (6 units) | 0
prothrombin concentrate (3000 units) | 0
transferred to intermediate care unit (IMC) | 1440
criticalDillness polyneuropathy | 1440
discharged | 2160
referred to rehabilitation center | 2160
physiotherapy | 2160
