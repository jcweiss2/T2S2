41 years old | 0
male | 0
admitted to the hospital | 0
abdominal pain | 0
exploratory laparotomy | 0
perforated appendicitis | 0
intraabdominal abscess | 0
hemangioma | 0
intraabdominal sepsis | 0
reoperated | 0
open abdomen | 0
open abdomen lavages | 0
abdominal wall defect | 0
granulation | -720
epithelization of the defect | -720
reconstruction of the abdominal wall | 0
skin incisions | 0
tissue expanders placement | 0
inflation of tissue expanders | 0
expansion of tissue expanders | 0
removal of expanders | 128
prosthetic mesh placement | 128
suction drains placement | 128
suction drains removal | 132
discharged | 96
follow-up | 720
no signs of mesh infection | 720
no extrusion | 720
no recurrent hernia | 720
no ulceration | 720
no enteric fistula | 720