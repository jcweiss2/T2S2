31 years old | 0
G1P0 | 0
primary infertility | -10368
cystic fibrosis | -10368
preconception counseling | -10368
maternal fetal medicine (MFM) | -10368
genetics | -10368
initiating infertility work-up | -10368
reproductive endocrinology and infertility | -10368
height 5 feet 4 inches | 0
weight 128 pounds | 0
body mass index 22 | 0
ovulation predictor kits | -10368
timed intercourse | -10368
hysterosalpingogram | -10368
normal hysterosalpingogram | -10368
semen analysis | -10368
mild teratospermia (6–8%) | -10368
pelvic ultrasound February 23, 2018 | -10368
antral follicle count (AFC) 30+ | -10368
arcuate uterus | -10368
high AFC | -10368
isolated episode anovulation | -10368
low cycle day 21 progesterone level | -10368
polycystic ovarian syndrome work-up | -10368
serum hormone levels within normal limits | -10368
no clinical signs of hyperandrogenism | -10368
ovulation normally | -10368
cardiology clearance | -10368
pulmonary medicine clearance | -10368
ovulation induction protocol started March 22, 2018 | -10368
letrozole 2.5 mg cycle days 3 to 7 | -10368
cycle day 12 ultrasound | -10368
luteinizing hormone (LH) levels | -10368
progesterone levels | -10368
several cycles of ovulation induction | -10368
intrauterine insemination | -10368
failed intrauterine insemination | -10368
combined oral contraceptive pills (COC) July 21, 2018 to August 21, 2018 | -10368
increase in breast size up to six-cup size in 2 to 4 weeks | -10368
IVF egg retrieval preparation September 2018 | -10368
follicle stimulating hormone (FSH, Follistim) | -10368
FSH combined with LH (Menopur) | -10368
gonadotropin-releasing hormone antagonist (Ganirelix) | -10368
no further breast growth during IVF preparation | -10368
breasts back to baseline within 3 to 5 weeks after COC discontinuation | -10368
estradiol use October 2018 | -10368
no noticeable breast changes with estradiol | -10368
progesterone supplementation November 14, 2018 | -10368
dramatic six-cup size increase in breast size over 1 week | -10368
embryo transfer November 18, 2018 | -10368
vaginal progesterone suppositories | -10368
continued breast growth | -10368
prenatal care at 10 weeks gestational age | 0
14-week visit | 0
significant breast pain | 0
breast ultrasound showed no sonographic abnormalities | 0
referred to Endocrinology | 0
15 weeks (February 11, 2019) laboratories | 0
intact parathyroid hormone (PTH) <6.3 | 0
calcium 10.1 | 0
PTH related peptide 1.2 | 0
normal Vitamin D | 0
prolactin 112.5 | 0
thyroid stimulating hormone (TSH) 0.885 | 0
started on bromocriptine 2.5 mg twice daily | 0
increased bromocriptine to 5 mg twice daily | 0
slower rate of breast enlargement | 0
switched to cabergoline 0.5 mg March | 0
accelerated rate of growth | 0
switched back to bromocriptine 10 mg twice daily | 0
16 weeks | 0
met with surgical oncology (breast surgeon) | 0
19 weeks | 0
met with plastic surgery | 0
not a surgical candidate | 0
size, swelling, increased vascularity of the breast | 0
physical therapy recommended | 0
manual lymphatic drainage (MLD) recommended | 0
16-cup total increase in breast size | 0
slowed rate of growth | 0
21 weeks | 0
superficial skin breakdown on the breast | 0
seeing physical therapy | 0
worsening ability to perform activities of daily living | 0
worsening pain | 0
presented to labor and delivery triage at 23 weeks | 0
uncontrolled pain | 0
started on oxycodone | 0
tylenol for pain control | 0
represented at 24 weeks | 0
admitted to antepartum unit | 0
pain control | 0
pain and discomfort progressed | 0
growth of breast tissue | 0
oxycodone up titrated to maximal doses | 0
physical medicine and rehab consultation | 0
methadone initiation | 0
methadone up titrated to 30 mg twice daily | 0
scheduled tylenol | 0
oxycodone | 0
hydromorphone for breakthrough pain | 0
stable pain control | 0
poor mobility related to pain | 0
deep venous thrombosis prophylaxis with daily enoxaparin | 0
better controlled pain | 0
long-term hospitalization complications | 0
skin breakdown | 0
herniation of breast tissue | 0
superficial wounds on breast | 0
ulcerated wounds | 0
herniated breast tissue | 0
hemorrhaged from exposed venous sinuses | 0
seen by surgical oncology (breast surgery) | 0
seen by plastic surgery | 0
avoidance of surgery during pregnancy | 0
concern for vascular compromise | 0
worsening loss of skin integrity | 0
growing wounds | 0
lymphovenous hypertension of the breast | 0
wound care management | 0
green discoloration of wound discharge | 0
colonization with pseudomonas | 0
topical care with hypochlorous acid (Vashe) | 0
wet to dry dressings | 0
no evidence of superimposed infection | 0
no antibiotics required | 0
manual lymphatic drainage (MLD) performed by mother and husband | 0
compression garment | 0
improved symptoms | 0
venous sinus hemorrhages developed around 27 weeks | 0
anticoagulation discontinued | 0
multiple episodes of hemorrhage (100–300cc) | 0
suture ligation by plastic surgery | 0
betamethasone administration for fetal lung maturity | 0
bilateral IV access | 0
crossmatched for four units of packed red blood cells | 0
hemoglobin optimization with intravenous iron infusions | 0
visual hallucinations | 0
psychiatry consulted | 0
anxiety, panic, exhaustion, delirium | 0
started on venlafaxine | 0
switched to citalopram | 0
stabilized briefly | 0
30 weeks | 0
recurrent breast hemorrhage | 0
requested early delivery | 0
shared decision making | 0
neonatology counseling | 0
induction of labor at 31 weeks | 0
rescue dose of betamethasone | 0
magnesium for fetal neuroprotection | 0
induction of labor | 0
recurrent late decelerations | 0
unresponsive to resuscitative measures | 0
primary C-section | 0
neonate appropriate for gestational age | 0
neonatal intensive care unit stay for 6 weeks | 0
respiratory distress syndrome | 0
continuous positive airway pressure | 0
stage II necrotizing enterocolitis | 0
treated with Zosyn for 1 week | 0
postoperative day 5 | 0
breasts felt softer | 0
compression garment fitting looser | 0
recorded breast size | 0
weaned off methadone | 0
well-controlled pain | 0
no pulmonary complications | 0
discharge home | 0
outpatient follow-up with wound care | 0
outpatient follow-up with plastic surgery | 0
outpatient follow-up with breast surgery | 0
outpatient follow-up with MFM | 0
3-week postpartum visit | 0
fully weaned off all narcotics | 0
no withdrawal symptoms | 0
plastic surgery recommended spontaneous regression | 0
interval breast reduction | 0
significant anxiety | 0
body image issues | 0
2 months postpartum | 0
stabilization of breast size | 0
breast reduction planned | 0
free nipple grafts | 0
breast reduction performed 20 weeks postpartum | 0
4,320 g breast tissue removed left | 0
4,762 g breast tissue removed right | 0
estimated blood loss 500cc | 0
discharged on postoperative day 1 | 0
bilateral Jackson-Pratt drains | 0
Conflict of Interest None declared | 0
