36 years old | 0
female | 0
admitted to the hospital | 0
general body ache | -72
malaise | -48
breathing difficulty | -48
diabetes mellitus type II | 0
obstructive sleep apnea | 0
hypertension | 0
hypothyroidism | 0
morbid obesity | 0
tachycardia | 0
tachypnea | 0
leukocytosis | 0
urinary tract infection | 0
pus cell count | 0
antibiotics | 0
meropenem | 0
vasopressors | 0
fluid resuscitation | 0
mechanical ventilation | 0
intubated | 4
anuric | 6
sequential organ failure assessment | 24
MODS score | 24
acute physiology and chronic health evaluation | 24
septic shock | 0
low perfusion state | 0
multi-organ dysfunction | 0
acute respiratory distress syndrome | 0
acute kidney injury | 0
arterial hypotension | 0
hemoadsorption column | 16
CytoSorb | 16
continuous renal replacement therapy | 16
heparin | 16
activated partial thromboplastin time | 16
inotropic support | 16
intravenous hydrocortisone | 16
noradrenalin | 28
vasopressors weaned out | 28
corticosteroids | 28
urine output increased | 72
ventilator parameters improved | 72
SOFA score | 72
MODS score | 72
APACHE II score | 72
laboratory parameters | 72
CytoSorb therapy | 72
discharged | 96