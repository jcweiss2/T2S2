23 years old | 0
female | 0
gravida 2 | 0
para 1 | 0
previous caesarean section | -672
admitted for induction of labour | 0
cervical ripening balloon catheter inserted | 0
cervical ripening balloon catheter removed | 24
artificial rupture of membranes | 24
oxytocin infusion commenced | 24
epidural anaesthesia | 216
indwelling catheter inserted | 216
full dilatation | 360
passive descent of the foetal head | 360
active pushing commenced | 367
cardiotocograph became pathological | 367
instrumental delivery | 367
indwelling catheter balloon deflated | 367
rosé-coloured haematuria noted | 367
vaginal delivery | 367
low cavity vacuum delivery | 367
right mediolateral episiotomy | 367
baby delivered | 367
Apgar scores of 9 and 10 | 367
postpartum haemorrhage | 367
syntocinon infusion | 367
ergometrine administered | 367
episiotomy laceration suture repair | 367
estimated blood loss 600 mL | 367
indwelling catheter reinserted | 367
clear urine noted | 367
epidural catheter removed | 367
normal micturition | 290
indwelling catheter removed | 290
acute right-flank pain | 780
rebound tenderness | 780
febrile | 780
tachycardic | 780
hypotensive | 780
haemoglobin level 86 | 780
white cell count 6 | 780
venous lactate 1.9 | 780
creatinine 58 | 780
CRP 87 | 780
IV crystalloid | 780
ceftriaxone and metronidazole | 780
gentamicin | 780
CT scan | 810
free fluid in the right retroperitoneal space | 810
urinoma | 810
extravasation of contrast | 810
haemoglobin stable at 86 | 840
haematocrit 0.265 | 840
CRP 76 | 840
creatinine 50 | 840
urine microscopy showed organisms | 840
sepsis from a urinary tract source | 840
transferred to intensive care | 840
IV metaraminol | 840
packed red blood cells given | 840
CT IV pyelogram | 960
contrast extravasation at the level of the right mid ureter | 960
ureteric injury | 960
emergency cystoscopy | 1080
posterior bladder wall ecchymosis | 1080
ureteral orifice normal | 1080
guide wire could not be passed | 1080
right rigid ureteroscopy | 1080
grade III incomplete proximal ureteric rupture | 1080
ureteric stent placed | 1080
persistent fevers | 1080
antibiotics upgraded to IV piperacillin/tazobactam | 1080
urine microscopy positive for E. coli | 1080
stepped down to ward-based care | 1200
discharged home | 240
follow-up cystoscopy | 1008
retrograde pyelogram | 1008
stent removed | 1008