61 years old | 0
female | 0
rheumatoid arthritis | -120 months
primary TKA | -120 months
revision TKA | -6 months
oral prednisone | -6 months
tacrolimus | -6 months
etanercept | -6 months
pain in right knee | 0
PJI | 0
intravenous antibiotic treatment | -24
referred to hospital | 0
septic shock | 0
burning sensations in right knee | 0
redness in right knee | 0
local heat in right knee | 0
swelling in right knee | 0
white blood cell count of 8.1×10^9/L | 0
C-reactive protein level of 19.9 mg/L | 0
aspiration of right knee joint | 0
gram-positive streptococci | 0
Streptococcus dysgalactiae | 0
temperature of 38.2°C | 0
heart rate of 128 beats/min | 0
blood pressure of 56/32 mmHg | 0
hemoglobin of 9.5 g/dL | 0
serum glucose of 99 mg/dL | 0
serum creatinine of 2.93 mg/dL | 0
sodium of 139 mEq/L | 0
radiography of right knee | 0
no osteolytic lesions | 0
no periprosthetic loosening | 0
irrigation | 0
debridement | 0
polyethylene liner exchange | 0
antibiotic therapy | 0
mechanical ventilation | 0
meropenem | 0
vancomycin | 0
clindamycin | 0
continuous hemodiafiltration | 0
nor-adrenaline | 0
noradrenaline application stopped | 120
swelling in right knee | 192
burning sensation in right knee | 192
exudate aspiration | 192
white blood cell count of 60×10^4/μL | 192
positive alpha-defensin test | 192
irrigation | 192
debridement | 192
implant removal | 192
antibiotic spacer placement | 192
inflammatory markers normalized | 432
C-reactive protein of 0.05 mg/L | 432
intravenous antibiotic therapy | 432
ampicillin | 432
clindamycin | 432
cefazolin | 504
bucillamine | 720
busiramine | 720
prednisolone | 720
oral cefalexin | 720
re-revision TKA | 1300
no clinical signs of infection | 1300
no pain in right knee | 1560
no swelling in right knee | 1560
no burning sensation in right knee | 1560
right knee motion | 1560