43 years old | 0
    woman | 0
    presented with fever | -240
    presented with dry cough | -240
    mild respiratory distress | -240
    SpO2 88%-89% | -240
    diagnosed with COVID-19 | -72
    polycystic ovarian disease | 0
    blood pressure 140/90 mmHg | 0
    pulse rate 88 beats/min | 0
    respiratory rate 20 breaths/min | 0
    SpO2 92% | 0
    bilateral decrease in air entry | 0
    total leucocyte count 11650 cells/µL | 0
    neutrophils 88% | 0
    lymphocytes 8% | 0
    CRP 16.44 mg/L | 0
    Pct 9.52 ng/mL | 0
    lactate dehydrogenase 282 IU/L | 0
    ferritin 158 ng/mL | 0
    D-dimer 775.84 ng/mL | 0
    interleukin-6 18.55 pg/mL | 0
    slightly elevated liver enzymes | 0
    normal electrolyte | 0
    normal renal function test | 0
    arterial oxygen partial pressure 39.0 mmHg | 0
    chest CT atypical viral infection | 0
    50% lung involvement | 0
    CTSI score 18/25 | 0
    non-rebreather mask 15 L/min oxygen | 0
    oxygen saturation 100% | 0
    echocardiography ejection fraction 60% | 0
    chest physiotherapy | 0
    incentive spirometry | 0
    IV remdesivir | 0
    IV dexamethasone | 0
    oral doxycycline | 0
    low molecular weight heparin | 0
    multivitamins | 0
    antibiotics | 0
    nebulization | 0
    oxygen requirement decreased | 168
    chest CT repeated | 168
    CTSI score 12/25 | 168
    weaned off oxygen | 288
    reports normalized except Pct | 288
    discharged | 456
    persistently elevated Pct | 456
    neck examination unremarkable | 456
    ultrasonography neck thyroid nodule | 456
    FNAC malignant epithelial neoplasm | 456
    left supraclavicular node metastatic carcinoma | 456
    Ctn 406 pg/mL | 456
    CEA not elevated | 456
    PET-CT thyroid nodule | 456
    MTC confirmed | 456
    COVID-19 pneumonia | 0
    total thyroidectomy | 3360
    central lymph node dissection | 3360
    thyroid nodule 3 cm × 2 cm × 1.5 cm | 3360
    MTC with lymphovascular invasion | 3360
    11/14 lymph nodes positive | 3360
    stage III pT2N1M0 | 3360
    postoperatively elevated Ctn 189 pg/mL | 3360
    PET-CT repeated | 3360
    second radical neck dissection | 3360
    6/16 lymph nodes positive | 3360
    Pct 3.54 ng/mL | 3360
    Ctn 14 pg/mL | 3360
    MEN-2 ruled out | 3360
    levothyroxine 150 mcg/d | 4320
    EBRT | 4320
    no recurrence | 4320
    