44 years old | 0
male | 0
nephrolithiasis | 0
HIV | 0
left flank pain | -120
abdominal pain | -120
painful ejaculation | -120
nausea | -120
vomiting | -120
decreased appetite | -120
subjective fever | -120
chills | -120
utilizing a prostate vibrator | -168
admitted to the emergency department | 0
left flank pain radiated into his left lower abdomen | 0
left flank pain radiated into his left testicle | 0
pain was described as achy to sharp | 0
vitals on arrival to the ED | 0
101.2 °F | 0
blood pressure 92/54 mmHg | 0
respiratory rate of 21 breaths/min | 0
weight of 94.5 kg | 0
SpO2 98% on room air | 0
physical exam | 0
in distress secondary to the pain | 0
diaphoretic | 0
appeared ill | 0
oral mucosa was dry | 0
cardiopulmonary exam | 0
sinus tachycardia | 0
no murmur | 0
clear lungs bilaterally | 0
abdominal exam | 0
left costovertebral angle tenderness | 0
left upper and lower abdominal tenderness to palpation | 0
voluntary guarding | 0
genitourinary exam | 0
tenderness to palpation along the left inguinal canal | 0
left epididymitis | 0
no clinical evidence for abscess | 0
no clinical evidence for cellulitis | 0
no clinical evidence for crepitus to the groin | 0
sepsis protocol initiated | 0
two peripheral IVs were placed | 0
urine/blood cultures were taken | 0
laboratory evaluation started | 0
fluid resuscitation initiated | 0
normal saline 30 mL/kg IV bolus | 0
complete blood count | 0
leukocytosis of 18.2 | 0
neutrophil predominance | 0
hemoglobin of 11.6 | 0
platelet level of 220 bil/L | 0
basic metabolic panel | 0
pre-renal azotemia | 0
blood urea nitrogen (BUN) of 27 mg/dL | 0
creatinine of 1.3 mg/dL | 0
blood glucose of 130 | 0
hepatic function panel | 0
unremarkable | 0
lactic acid of 3.2 | 0
lactic acid of 1.5 | 2
urinalysis | 0
2+ blood | 0
+nitrites | 0
3+ leukocyte esterase | 0
>50 WBCs | 0
3+ bacteria | 0
25–50 RBCs | 0
C-reactive protein 7.1 | 0
ceftriaxone | 0
gentamicin | 0
ultrasound of the scrotum with Doppler | 0
prominent epididymis with increased vascularity | 0
small left hydrocele with scattered internal debris | 0
no evidence for compromised arterial flow | 0
no evidence for abscess formation | 0
CT of the abdomen/pelvis without contrast | 0
left-sided peri-ureteral fat stranding | 0
prominent left seminal vesicle | 0
infiltrative fat stranding predominantly centered around the left hemi-pelvis | 0
multiple prominent pelvic lymph nodes up to 8.1 mm | 0
prominent inguinal lymph nodes up to 6.5 mm | 0
prostate is top-normal in size at 5 cm | 0
central venous catheter | 2
inotropic medication | 2
admitted to the intensive care unit | 2
urine and blood cultures grew Escherichia coli | 24
Escherichia coli was pansusceptible | 24
testing for Chlamydia trachomatis and Neisseria gonorrhoeae DNA | 24
negative | 24
off inotropic medication | 72
hemodynamically stable | 72
tolerating a regular diet | 72
discharged | 96
cefuroxime | 96
1-month follow-up | 720
progressing well | 720
denied any complaints | 720