39 years old | 0
    woman | 0
    type 2 diabetes | -168
    deep vein thrombosis | -168
    gastritis | -168
    schizophrenia | -168
    self-harm | -168
    presented to the medical admissions unit | 0
    right sub-mammary abscess | -168
    spreading cellulitis of the breast | -168
    septic | 0
    pyrexia of 39.2 | 0
    blood pressure of 127/65 | 0
    tachycardia of 110 | 0
    widespread cellulitis involving the nipple | 0
    sub-mammary area cellulitis | 0
    cellulitis spreading to the axilla | 0
    white cell count of 23.8 | 0
    neutrophils 19.9 | 0
    CRP of 428 | 0
    simple cellulitis | 0
    commenced on parenteral antibiotics | 0
    fluid resuscitation | 0
    condition worsened | 72
    intravenous benzyl penicillin | 0
    flucloxacillin | 0
    surgical opinion sought | 72
    evidence of synergistic gangrene | 72
    cellulitis spread | 72
    areas of growing necrotic ulceration | 72
    resuscitation commenced | 72
    antibiotic therapy adjusted to imipenem | 72
    antibiotic therapy adjusted to clindamycin | 72
    taken to theatre within a few hours | 72
    partial mastectomy performed | 72
    wound left open and packed | 72
    postoperative stability on intensive care | 72
    returned to theatre for further debridement | 96
    vacuum dressing applied | 96
    signs of sepsis improved | 120
    returned to the ward | 120
    nutritional supplements continued | 120
    adequate hydration continued | 120
    secondary closure performed | 312
    no further breakdown of remaining tissues | 312
    preoperative cultures taken | 72
    gram positive bacteria identified | 72
    gram negative bacteria identified | 72
    Bacteroides spp identified | 72
    histology confirmed microscopic changes | 72
    abscess formation consistent with gangrene | 72
    no evidence of malignancy | 72
    blood markers of infection progressively improved | 168
    no signs of secondary organ failure | 168
    discharged | 528
    intravenous antibiotics administered for 10 days | 240
    changed to oral antibiotics | 240
    co amoxiclav | 240
    metronidazole | 240
    follow-up arranged | 528
    possibility of reconstruction considered | 528
    