26 years old | 0
female | 0
ulcerative colitis | -672
abdominal pain | 0
fever | 0
bloody diarrhoea | 0
generalised weakness | 0
poorly controlled colitis | -672
mesalazine | -672
6-mercaptopurine | -672
prednisolone | -672
analgesia | 0
intravenous fluids | 0
intravenous steroids | 0
discharged | 0
readmitted | 336
sepsis | 336
tachycardia | 336
hypotension | 336
pyrexia | 336
distended abdomen | 336
tender on palpation | 336
tender on percussion | 336
rebound tenderness | 336
peritonitis | 336
colonic distension | 336
emergent caesarean section | 336
total abdominal colectomy | 336
end ileostomy | 336
discharged | 360
ventilator support | 336
weaned off ventilator | 360
completion proctectomy | 672
ileal reservoir | 672
ileoanal anastomosis | 672
diverting ileostomy | 672
loop ileostomy reversed | 2088
bowel movements | 2160
constitutionally well | 2160
surgical wounds | 2160
toxic megacolon | 336
transmural inflammation | 336
bowel wall erosion | 336
fetal delivery | 336
neonatal intensive care | 336
neonatal progressive care | 360
discharged home | 2400
pathologic examination | 336
optimal healing | 2160
reduced fertility | 2160
growth assessments | 2160
satisfactory recovery | 2400
exacerbation during pregnancy | 336
medical therapy | 336
surgical intervention | 336
loop ileostomy reversal | 2088
abdominal radiograph | 336
colonic mucosa | 336
haemorrhage | 336
intramural inflammation | 336
ileostomy scars | 2088
laparotomy | 336
consent for publication | 0
- 26 years old | 0 (since age is at the time of the main admission)
+ Gender: female | 0
