79 years old | 0
male | 0
COPD | 0
stable ischaemic heart disease | 0
bicytopenia | 0
hernia repair | 0
normocytic, normochromic anemia | 0
decreased reticulocyte response | 0
leukopenia | 0
bone marrow aspirate | 0
mild dysplastic changes | 0
plasmacytosis | 0
trephine | 0
increased CD138+ plasma cells | 0
flow cytometry | 0
nonclonal plasma cells | 0
CD45 positive | 0
CD38 bright | 0
CD138 positive | 0
CD56 negative | 0
CD117 negative | 0
no blasts | 0
no clonal lymphoid infiltrate | 0
dyspnoea | -168
fever | -168
anemia | -168
leukopenia | -168
neutropenic sepsis | -168
pneumonia | -168
mild congestive cardiac failure | -168
acute infective exacerbation of COPD | -168
negative blood culture | -168
negative urine culture | -168
negative stool culture | -168
negative sputum culture | -168
negative TB PCR | -168
negative AFB smears | -168
bilateral pleural effusions | -168
focal consolidation | -168
responded to carbapenem antibiotic | -168
transfusion support | -168
no monoclonal paraprotein | -168
faint IgM band | -168
faint lambda band | -168
negative serum M-band | -168
negative skeletal survey | -168
normal serum calcium | -168
polyclonal lymphoplasmacytoid cells | -168
mild splenomegaly | -168
small volume lymphadenopathy | -168
negative HIV serology | -168
deferred bone marrow studies | -168
fever | 0
broad-spectrum antimicrobials | 0
bilateral pleural effusions | 0
bloody pleural fluid | 0
bronchoscopic evaluation | 0
unremarkable connective tissue disease workup | 0
negative BAL malignancy | 0
negative BAL tuberculosis | 0
atypical plasma cells | 0
fungal elements | 0
Candida | 0
Cryptococcus | 0
negative serum cryptococcal antigen | 0
hypotension | 0
ICU admission | 0
inotropic support | 0
GCSF | 0
Amphotericin B | 0
Ambisome | 0
stable pericardial effusion | 0
deferred pericardiocentesis | 0
CN growth in BAL | 0
fluconazole sensitive | 0
IV Fluconazole | 0
deterioration | 0
death | 0
reexamined bone marrow biopsy | 0
GMS-positive yeast | 0
CN PCR confirmation | 0
chronic disseminated CN infection | 0
pleural effusion | 0
pericardial effusion | 0
lymph node involvement | 0
lung involvement | 0
bone marrow involvement | 0
