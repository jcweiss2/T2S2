28 years old | 0
male | 0
admitted to the hospital | 0
fever | -120
diarrhea | -120
icterus | -120
oliguria | -24
breathlessness | -24
edema of the legs | -24
bilateral lower limb motor weakness | -24
pitting edema legs | 0
sinus tachycardia | 0
tachypnoea | 0
normotension | 0
bilateral basal rales | 0
paraparesis | 0
no sensory or bladder abnormalities | 0
proteinuria | 0
hemoglobin level | 0
total leukocyte count | 0
platelet count | 0
severe renal failure | 0
liver function tests | 0
corrected serum calcium | 0
phosphorus | 0
serum creatinekinase | 0
serum lactate dehydrogenase | 0
urine and blood cultures | 0
serum immunoglobulin M antibodies for leptospira | 0
kidneys echogenic and bulky | 0
computed tomography of the brain | 0
electrocardiogram | 0
chest radiograph | 0
arterial blood gas analysis | 0
hemodialysis | 0
hyperkalemia | 0
metabolic acidosis | 0
injection crystalline penicillin | 24
glucose insulin drip | 24
hypernatremia | 24
water deficit | 48
hepatic encephalopathy | 48
carbohydrate diet | 48
lactulose bowel wash | 48
avoidance of protein diet | 48
renal functions improvement | 216
increase in renal output | 216
maintenance of creatinine | 216
parenteral fluid | 216
central venous pressure monitoring | 216
daily output chart | 216
nosocomial infections | 216
physiotherapy | 216
transferred to general ward | 216
discharged | 504
ambulatory state | 504
improved renal function | 504
improved liver function | 504
Grade 5 motor power | 504