55 years old | 0
female | 0
hepatitis C | 0
intra-venous drug use | 0
alcohol abuse | 0
Child-Pugh B liver cirrhosis | 0
abdominal pain | 0
diarrhoea | 0
fevers | 0
confusion | 0
no history of colonic disease | 0
CT of the abdomen | 0
mildly dilated proximal large bowel | 0
no fat stranding or colonic wall thickening | 0
stool PCR positive for campylobacter species | 0
treatment with azithromycin | 0
treatment with ceftriaxone | 0
treatment with metronidazole | 0
intravenous fluids | 0
electrolyte replacement | 0
aspiration pneumonitis | 24
type 2 myocardial infarction | 24
renal failure | 24
metabolic acidosis | 24
intubation | 24
vasopressors | 24
dialysis | 24
transthoracic echocardiography | 24
lumbar puncture | 24
blood cultures | 24
CT scans of the head, chest, abdomen and pelvis | 24
no alternative source of sepsis | 24
antibiotics escalated to piperacillin/tazobactam | 24
bloody diarrhoea | 384
ongoing refractory multi-organ dysfunction | 384
CT abdomen demonstrated colonic wall thickening | 384
no gross dilatation, intramural gas, free gas or obvious bleeding points | 384
upper endoscopy excluded varices and ulcers | 384
transfer to tertiary hospital | 384
emergent laparotomy | 384
viable mildly dilated colon | 384
clear ascites | 384
no evidence of ischaemia, necrosis or perforation | 384
liver was nodular | 384
remainder of the bowel was normal | 384
flexible sigmoidoscopy demonstrated discontinuous areas of non-bleeding ulcerated mucosa | 384
biopsies were taken | 384
case discussed with intensive care and infectious diseases teams | 384
antibiotics changed to daptomycin, ciprofloxacin, fluconazole and metronidazole | 384
worsening haemodynamic instability | 396
increasing amounts of noradrenaline and vasopressin | 396
re-look laparotomy | 396
grossly dilated colon | 396
no perforation or full thickness ischemia | 396
subtotal colectomy | 396
end ileostomy and distal sigmoid mucous fistula | 396
immediate improvement postoperatively | 396
vasopressin ceased | 396
noradrenaline infusion halved | 396
escalating vasopressor requirements | 420
acidosis | 420
liver failure | 420
respiratory failure | 420
death | 432
histology of pathological specimens showed features of infectious colitis and ischemia | 432
macroscopically, multiple discrete areas of mucosal ulceration | 432
microscopically, the ulcerated mucosa showed congestion, neutrophilic infiltration and fibrin thombi | 432
no architectural distortion and cryptitis and crypt abscesses were not prominent features | 432
features typical for inflammatory bowel disease were absent | 432