Here is the table of events and timestamps:

46 years old | 0
male | 0
ulcerative colitis | 0
malaise | -72
fever | -72
loss of appetite | -72
admitted to the hospital | 0
blood pressure 124/46 mmHg | 0
heart rate 122 beats per min | 0
SpO2 98% in room air | 0
respiratory rate 16/min | 0
body temperature 40.2°C | 0
chills | 0
nausea | 0
cardiac arrest | 0
chest compression | 0
tracheal intubation | 0
ventricular fibrillation | 0
defibrillation | 0
adrenaline | 0
diagnosed with Brugada syndrome | 0
coved-type ST elevation in V1 and V2 | 0
improved with acetaminophen | 0
hypercalcemia | 0
high parathyroid hormone levels | 0
abnormal uptake in the anterior mediastinum | 0
ectopic parathyroid adenoma | 0
tumor resection | 24
ECG with J point elevation | -720
ECG with J point elevation | -720
ECG with coved-type ST elevation in V1 and V2 | -720
ECG with J point elevation | -720
ECG with J point elevation | -720
ECG with coved-type ST elevation in V1 and V2 | -720
fever reoccurred | 120
contrast-enhanced CT scan with liver abscess | 120
changed antibiotics to meropenem and vancomycin | 120
puncture drainage | 120
infection controlled | 168
implantation of an implantable cardioverter defibrillator | 168
discharged | 168
family history of sudden death | -720
endocrinologist examination | 0
nonfunctional pituitary adenomas and nonfunctional adrenal tumors | 168
multiple endocrine neoplasia type 1 | 168