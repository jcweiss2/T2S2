45 years old | 0
man | 0
taken to the emergency ward | 0
giant inguinoscrotal hernia | -10080
refused surgery | -10080
inability to walk | 0
gradually loss of strength | 0
progressive increase of hernia | 0
hernia reached the calves | 0
used a small wagon | -720
ulcer | -720
continuously discharging putrid liquid | -720
systemic inflammatory response syndrome | 0
impairment of coagulation | 0
anemia | 0
severe hyponatremia | 0
complete left-sided pleural effusion | 0
intubation | 0
catecholamine therapy | 0
transferred to the intensive care unit | 0
CT scan | 0
complete dislocation of the small bowel | 0
complete dislocation of the large bowel | 0
descending of the duodenum | 0
descending of the pancreas | 0
intrahepatic cholestases | 0
extrahepatic cholestases | 0
congestion of the right kidney | 0
ureter descended into the hernia sac | 0
ureter dilated up to its return into the abdominal cavity | 0
stabilized | 120
surgery attempted | 120
exploration of the abdominal cavity | 120
signs of peritonitis | 120
purulent liquid in the hernia sac | 120
penis identified intra-abdominally | 120
resection of mobile large bowel | 120
resection of distal parts of the ileum | 120
stabilization | 168
resection of the majority of the hernia sac | 168
inability to close the fascia | 168
inflammatory situation | 168
abdominal cavity reconstructed using absorbable mesh grafts | 168
recovered slowly | 168
mobilization complicated | 168
a priori existing lesion of the nervus peroneus | 168
polyneuropathia | 168
discharged from the hospital | 840
following rehabilitation program | 840
regained the ability to walk | 840
regained the ability to care for himself | 840
refused any further plastic reconstruction | 840
