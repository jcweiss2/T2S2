25 years old | 0
male | 0
Afghan | 0
penetrating sharp injury with nail to left heel | -480
lockjaw | -192
muscle spasms | -192
trismus | 0
opisthotonos | 0
generalized attacks | 0
vaccination history negative | 0
human anti-tetanus immunoglobulin | 0
tetanus-diphtheria toxoid | 0
admitted to ICU | 0
midazolam infusion | 0
morphine infusion | 0
feeding via Nasogastric tube | 0
severe spasms | 0
rhabdomyolysis | 0
hydration | 0
bicarbonate infusion | 0
metronidazole | 0
temperature 38°C | 0
tazocine | 72
ciprofloxacin | 72
urine culture positive | 72
Escherichia coli | 72
intubated | 0
pancronium | 0
percutaneous dilatational tracheostomy | 240
discontinued muscle relaxant | 360
baclofen | 360
sciatic nerve block | 432
extubated | 432
pain score decreased | 432
tachycardia | 0
stable blood pressure | 0
routine laboratory data normal | 0
liver function test normal | 0
Creatine Phosphokinase raised | 0
left ICU | 480