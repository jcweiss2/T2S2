45 years old | 0
female | 0
admitted to the hospital | 0
malaise | -72
upper respiratory tract infection | -72
fever | -72
hypotension | 0
tachycardia | -72
heart rate 250 bpm | 0
vagal maneuvers | 0
IV adenosine | 0
ECG | 0
narrow QRS complex tachycardia | 0
crystalloid | 0
IV diltiazem | 0
electrical cardioversion | 0
IV esmolol | 0
digoxin | 0
magnesium sulfate | 0
amiodarone | 0
oxygen requirements | 0
pulmonary edema | 0
IV furosemide | 0
transfer to tertiary hospital | 0
second loading dose of IV amiodarone | 12
electrical cardioversion | 12
IV lidocaine | 12
procainamide | 12
general anesthetic | 12
intubated | 12
cooled to 35.5°C | 12
esmolol infusion | 12
lidocaine infusion | 12
procainamide infusion | 12
heart rate slowed to 130 bpm | 12
AV dissociation | 12
vasopressin infusion | 24
mean arterial pressure 50 mm Hg | 24
taken to cardiac electrophysiology laboratory | 36
antiarrhythmic infusions discontinued | 36
multipolar catheters placed | 36
tachycardia cycle length 504 ms | 36
AV dissociation | 36
His potentials | 36
HV interval 59 ms | 36
scanning diastole with premature ventricular contractions | 36
atrial beats | 36
ventricular overdrive pacing | 36
retrograde His activation | 36
VHHV response | 36
electroanatomic mapping | 36
limited geometry of basal RV septal region | 36
timing points collected | 36
local sharp potentials | 36
catheter pressure terminated tachycardia | 36
cryoablation considered | 36
radiofrequency ablation | 36
initial lesions delivered | 36
ablation at site of earliest activation | 36
tachycardia terminated | 36
slower junctional beats | 36
insurance lesions delivered | 36
temporary atrial pacing wire | 36
sinus node suppression | 36
Streptococcus pneumoniae grown on sputum cultures | 36
IV antibiotics | 36
discharged | 216
no recurrence of tachycardia | 648
previous medical contacts with unstable tachycardia | -1000
prolonged admission to intensive care unit | -1000
supraventricular tachycardia | -1000
resolved with supportive medical treatment | -1000
beta blockade | -1000