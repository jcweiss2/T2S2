13 years old | 0
    girl | 0
    fever | -72
    loss of appetite | -72
    appendectomy | -72
    discharged | -72
    dehydrated | 0
    tachycardia | 0
    tachypnea | 0
    fever | 0
    axillary temperature 38.8 °C | 0
    blood pressure 120/70 mmHg | 0
    normal cardiac examination | 0
    normal pulmonary examination | 0
    diffusely tender abdomen | 0
    painful rebound test | 0
    present intestinal sounds | 0
    normal intestinal sounds | 0
    hyperemic surgical scar | 0
    abdominal ultrasound | 0
    pericolic abscess | 0
    surgically drained abscess | 0
    abdominal secretion culture positive for multisensitive E. coli | 0
    abdominal secretion culture positive for group G β-hemolytic Streptococcus sp | 0
    ceftriaxone prescribed | 0
    metronidazole prescribed | 0
    abdominal pain | 72
    fever relapsed | 72
    antibiotics changed to vancomycin | 72
    antibiotics changed to ceftazidime | 72
    antibiotics changed to amikacin | 72
    intermittent fever | 72
    abdominal CT ruled out surgical complications | 72
    broad-spectrum antibiotic regimen | 72
    fluconazole added | 72
    hypotensive | 288
    tachycardic | 288
    temperature rose to 39.4 °C | 288
    referred to ICU | 288
    vasoactive drugs required | 288
    hemodynamic stabilization | 288
    negative blood cultures | 288
    negative urine cultures | 0
    normal transthoracic echo Doppler Cardiogram | 0
    progressive respiratory failure | 288
    thrombocytopenia | 480
    hyperbilirubinemia | 480
    enlarged prothrombin time | 480
    altered liver enzymes | 480
    exploratory laparotomy | 528
    third surgical procedure | 528
    loose peritoneal adhesions | 528
    no purulent secretion | 528
    no intestinal perforation | 528
    no bowel necrosis | 528
    multiple organ failure | 528
    required hemodialysis | 528
    frequent blood transfusions | 528
    died | 576
    autopsy performed | 576
    Bogota bag closing peritoneotomy | 576
    mild serohemorrhagic effusion | 576
    non-dehiscent surgical sutures | 576
    no signs of peritonitis | 576
    no intra-abdominal purulent collection | 576
    enlarged liver | 576
    winy-colored liver areas | 576
    yellowish liver parenchyma | 576
    ischemic lobular necrosis | 576
    macrovesicular steatosis | 576
    microvesicular steatosis | 576
    enlarged spleen | 576
    reactive spleen parenchyma | 576
    depleted white pulp | 576
    congested red pulp | 576
    ischemic infarction areas in spleen | 576
    histiocytes phagocytizing red blood cells | 576
    lymphocytes present in spleen | 576
    pancreatic steatonecrosis | 576
    pancreatic ischemic necrosis | 576
    adrenal gland cortical ischemic necrosis | 576
    petechiae on lung surfaces | 576
    petechiae on pericardium | 576
    myocardial hemorrhagic suffusions | 576
    recent pericardial hemorrhage | 576
    recent myocardial hemorrhage | 576
    increased lung volume | 576
    shock lung | 576
    alveolar spaces filled with macrophages | 576
    alveolar spaces filled with fibrin | 576
    alveolar spaces filled with red blood cells | 576
    no hemophagocytosis in lungs | 576
    mediastinal lymphadenitis | 576
    intra-abdominal lymphadenitis | 576
    sinusal histiocytosis | 576
    lymphocytic depletion | 576
    histiocytes with erythrocyte phagocytosis | 576
    CD68-positive histiocytes | 576
    S100-negative histiocytes | 576
    hypercellular bone marrow | 576
    granulocytic series elements | 576
    histiocytes with hemophagocytosis | 576
    hypoxic-ischemic encephalopathy | 576
    acute tubular necrosis | 576
    hemophagocytic syndrome | 576
    triggered by acute appendicitis | 576
    hemodynamic shock | 576
    