78 years old | 0
female | 0
admitted to the hospital | 0
complaining of diarrhea | -336
diarrhea | -336
non-bloody diarrhea | -336
abdominal pain | -72
nausea | -72
non-bloody vomiting | -72
no fever | -72
no headache | -72
no cough | -72
no shortness of breath | -72
no jaw claudication | -72
no joint pain | -72
no visual disturbances | -72
immunized against COVID-19 | -672
type 2 diabetes mellitus | -672
hypertension | -672
CKD 3b A2 | -672
depression | -672
hypertriglyceridemia | -672
anemia with CKD | -672
bilateral cataract surgery | -8760
aspirin | -672
atorvastatin | -672
famotidine | -672
glargine insulin | -672
aspart insulin | -672
metformin | -672
metoprolol tartrate | -672
losartan | -672
torsemide | -672
sertraline | -672
no recent medication changes | -72
former smoker | -0
no alcohol or illicit drug use | -0
temperature 36.3°C | 0
blood pressure 165/67 mmHg | 0
heart rate 104 beats per minute | 0
respiratory rate 16 breaths per minute | 0
oxygen saturation normal | 0
leukocytosis | 0
neutrophilia | 0
lymphopenia | 0
hemoglobin 10.6 g/dL | 0
mild thrombocytosis | 0
lactate 6.4 mmol/L | 0
sodium 135 mmol/L | 0
hypochloremia | 0
hyperkalemia | 0
elevated metabolic acidosis | 0
anion gap elevated | 0
glucose 269 mg/dL | 0
blood urea nitrogen 83 mg/dL | 0
creatinine 8.47 mg/dL | 0
normal liver transaminases | 0
normal total bilirubin | 0
creatine kinase 110 U/L | 0
venous blood gas pH <6.80 | 0
pCO2 17 mmHg | 0
beta-hydroxybutyrate 1.8 mmol/L | 0
urinalysis showed glucose 500 mg/dL | 0
urinalysis showed ketones 80 mg/dL | 0
CT scan of abdomen and pelvis | 0
administered i.v. ceftriaxone | 0
administered Flagyl | 0
2 L NaCl 0.9% fluid bolus | 0
300 mEq bicarbonate bolus | 0
bicarbonate drip | 0
repeat lactate showed increase to 9.6 mmol/L | 2
new imaging of abdomen and pelvis | 2
insulin drip initiated | 2
2-L NaCl 0.9% fluid bolus | 2
confusion | 3
lethargy | 3
hypothermia | 3
sudden painless bilateral vision loss | 3
blood pressure stable | 3
heart rate stable | 3
CT head negative | 3
emergent ophthalmology evaluation | 3
preserved extraocular motility | 3
no evidence of retinopathy | 3
no macular edema | 3
no acute glaucoma | 3
no embolic phenomena | 3
MRI of brain revealed no acute abnormalities | 7
repeated blood work showed worsening lactic acid | 7
venous blood gas analysis showed pH 6.87 | 9
pCO2 29 mmHg | 9
worsening lactic acid | 9
CRRT initiated | 9
hypo-tension | 9
norepinephrine infusion initiated | 9
transthoracic echocardiogram | 9
preserved left ventricular ejection fraction | 9
no segmental wall motion abnormalities | 9
no intracardiac mass or thrombus | 9
volatile serum screen revealed high acetone | 9
negative for methanol, ethanol, and isopropanol | 9
metabolic acidosis and vision started to improve | 11
vision and mental status returned to baseline | 11
hypothermia gradually resolved | 11
bicarbonate infusion discontinued | 11
insulin drip transitioned to subcutaneous insulin | 11
weaned off norepinephrine | 16
infectious diseases work-up remained negative | 48
abdominal exam remained benign | 48
no recurrence of diarrhea | 48
empiric antibiotics discontinued | 48
dialysis discontinued | 66
creatinine improved to 2.93 mg/dL | 66
hyperkalemia resolved | 66
discharged home | 72
adjusted insulin regimen | 72
indefinite discontinuation of metformin | 72