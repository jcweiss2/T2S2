32 years old | 0
male | 0
admitted to the hospital | 0
beating | -1
multiple blunt trauma | -1
Glasgow Coma Scale score was 10 | 0
heart rate was 95 | 0
blood pressure was 120/80 mmHg | 0
loss of consciousness | -1
no nausea | 0
no vomiting | 0
pain on bilateral upper quadrants | 0
no abdominal tenderness | 0
no rebound tenderness | 0
no abdominal rigidity | 0
no hematuria | 0
leukocytosis | 0
hemoglobin level was 14.8 g/dl | 0
AST was 496 U/l | 0
ALT was 940 U/l | 0
direct bilirubin was 0.44 mg/dl | 0
total bilirubin was 0.82 mg/dl | 0
CT scan | 0
right parietal bone depression fracture | 0
free perihepatic fluid | 0
free perisplenic fluid | 0
splenic laceration | 0
abdominal CT scan | 4
increased perihepatic fluid | 4
heterogeneous appearance at falciform ligament | 4
focal enlargement and mural thickening at the second and third part of the duodenum | 4
neurosurgical operation | 4
postoperative follow-up | 24
decreased pain on abdomen | 24
leukocyte count decreased to 15,800×10^6 /ml | 24
AST had become 2265 U/l | 24
ALT had become 2224 U/l | 24
Hgb was 9.5 g/dl | 24
tachycardia | 48
tenderness on four quadrants of abdomen | 48
total bilirubin was 24.63 mg/dl | 48
direct bilirubin was 10.8 mg/dl | 48
urea was 48 mg/dl | 48
creatinine was 0.93 mg/dl | 48
amylase was 214 U/l | 48
exploratory laparotomy | 48
bile in abdomen | 48
common hepatic duct fully transected | 48
cholecystectomy | 48
drain placed to common hepatic duct | 48
multiple drains placed inside the abdomen | 48
operation ended | 48
abdominal drains removed | 120
discharged | 240
biliary drain changed for percutaneous biliary drainage | 720
second operation | 840
Roux-en-Y hepaticojejunostomy | 840
discharged | 850
full recovery | 850