19 years old | 0
male | 0
admitted to the hospital | 0
intermittent fever | -240
shortness of breath | -240
New York Heart Association class III | -240
blood culture positive for methicillin-susceptible Staphylococcus aureus | -240
administered broad-spectrum antibiotics | -240
transesophageal echocardiogram | -240
Sievers type I bicuspid aortic valve | -240
moderate aortic insufficiency | -240
vegetation attached on the ventricular side of the aortic leaflet | -240
vegetation attached to the A2 segment of mitral valve | -240
mitral regurgitation | -240
aortomitral pseudoaneurysm | -240
magnetic resonance imaging of the brain | -240
septic emboli | -240
subarachnoid hemorrhage | -240
aneurysm in the right pre-central sulcus | -240
no neurologic manifestations | -240
multidisciplinary team discussion | -12
planned for urgent cardiac surgery | -12
consented for bioprosthetic valve | -12
cardiac exposure via sternotomy | 0
aorta and both cavae cannulated | 0
cardiopulmonary bypass initiated | 0
cardioplegic arrest achieved | 0
aortic valve excised | 0
aortomitral aneurysm debrided | 0
MV approached via left atriotomy | 0
anterior mitral leaflet vegetations excised | 0
perforation repaired using a bovine pericardial patch | 0
left ventricular cavity and aortomitral area irrigated with antibiotic solution | 0
porcine aortic root prosthesis sized | 0
prosthesis turned inside-out | 0
prosthesis placed inside the left ventricular outflow tract | 0
prosthesis depth secured with sutures | 0
prosthetic rim sutured to aortic annulus | 0
annulus at the noncoronary cusp reconstructed with bovine pericardial strip | 0
prosthesis everted back to normal orientation | 0
coronary ostia reimplanted | 0
distal graft to ascending aorta anastomosis completed | 0
intraoperative TEE demonstrated normal functioning aortic root prosthesis | 0
mild central leak in the MV | 0
successful repair of aortomitral defect | 0
separated from cardiopulmonary bypass | 0
no rhythm abnormalities | 0
uneventful postoperative stay in the intensive care unit | 12
microbiology result of the excised tissue negative | 12
received 6 weeks of intravenous flucloxacillin | 12
discharged | 432
no neurologic deficits at the time of discharge | 432
completely well at 6 weeks follow-up | 1008