76 years old | 0
female | 0
diabetic | 0
altered mental status | 0
found down in a pool of blood and urine | 0
gross hematuria | 0
Foley catheter placement | 0
afebrile | 0
blood urea nitrogen of 110 mg/dL | 0
serum creatinine of 3.4 mg/dL | 0
thrombocytopenia | 0
leukocytosis with left shift | 0
blood culture produced gram-negative rods | 24
Escherichia coli | 24
non-contrast Computed Tomography (CT) | 0
status post bilateral nephrectomy | 0
retroperitoneal extraluminal air | 0
air within the lumen of the bladder | 0
bladder wall thickening | 0
severe sepsis | 0
hyperosmolar hyperglycemic non-ketotic syndrome | 0
acute kidney injury | 0
fluid resuscitation | 0
glucose control | 0
administration of antibiotics | 0
pressor support | 0
stabilized overnight | 24
anuric | 24
multisystem organ dysfunction | 24
multiple inotropic agents | 24
review of CT imaging by the Urology team | 24
diagnosis of bilateral emphysematous pyelonephritis | 24
emergent bilateral nephrectomy considered | 24
conservative approach chosen | 24
cystoscopy with bilateral retrograde pyelogram | 48
placement of ureteral stents | 48
gross purulent discharge | 48
interventional radiology consulted | 72
bilateral percutaneous renal abscess drains placed | 72
no significant output or improvement | 96
expired | 120