28 years old | 0
    male | 0
    presented to the emergency department | 0
    fever | -120
    diarrhea | -120
    icterus | -24
    oliguria | -24
    breathlessness | -24
    edema of the legs | -24
    bilateral lower limb motor weakness | -24
    no sensory involvement | -24
    no bladder involvement | -24
    pitting edema legs | 0
    icterus | 0
    sinus tachycardia | 0
    pulse 120/min | 0
    tachypnea | 0
    respiratory rate 32/min | 0
    normotension | 0
    blood pressure 120/80 mm Hg | 0
    bilateral basal rales | 0
    paraparesis | 0
    Grade 1/5 motor power | 0
    no sensory abnormalities | 0
    no bladder abnormalities | 0
    no meningeal signs | 0
    deep tendon reflexes normal | 0
    sensory system plantar response normal | 0
    transferred to ICU | 0
    proteinuria | 0
    red blood cells in urine | 0
    pus cells in urine | 0
    hemoglobin 12.5 g/dL | 0
    total leukocyte count 6800 cells/cubic mm | 0
    platelet count 75000/cubic mm | 0
    severe renal failure | 0
    blood urea 198 mg/dL | 0
    serum creatinine 4.8 mg/dL | 0
    sodium 152 meq/L | 0
    potassium 6.9 meq/L | 0
    total bilirubin 8.8 mg/dL | 0
    direct bilirubin 4.7 mg/dL | 0
    aspartate aminotransferase 201 U/L | 0
    alanine aminotransferase 167 U/L | 0
    alkaline phosphatase 57 U/L | 0
    serum total protein 5.6 g/dL | 0
    albumin 2.6 g/dL | 0
    corrected serum calcium 8.8 mg/dL | 0
    phosphorus 4.5 mg/dL | 0
    serum creatine kinase 670 U/L | 0
    serum lactate dehydrogenase 142 U/L | 0
    urine culture sterile | 0
    blood culture sterile | 0
    serum IgM antibodies for leptospira positive | 0
    titer IgM antibodies for leptospira 60 U/ml | 0
    kidneys echogenic | 0
    kidneys bulky on ultrasonography | 0
    computed tomography of the brain normal | 0
    electrocardiogram sinus tachycardia | 0
    tall tented T waves suggestive of hyperkalemia | 0
    chest radiograph bilateral diffuse infiltrates | 0
    arterial blood gas analysis metabolic acidosis | 0
    pH 6.9 | 0
    SpO2 96% | 0
    PaO2 82 mmHg | 0
    PaCO2 35 mm Hg | 0
    HCO3 8 mEq/L | 0
    admitted to ICU | 0
    hemodialysis for acute renal failure | 0
    hemodialysis to control hyperkalemia | 0
    hemodynamic stability | 0
    MRI of spinal cord normal | 0
    nerve conduction velocity bilateral lumbosacral polyradiculopathy | 0
    no evidence of myopathy on EMG | 0
    CSF study no cells | 0
    CSF normal sugar | 0
    CSF normal proteins | 0
    CSF no organism on staining | 0
    persistence of paraparesis after correcting hyperkalemia | 0
    leptospirosis manifesting with Weil's syndrome | 0
    leptospirosis manifesting with paraparesis | 0
    antibiotic treatment with crystalline penicillin | 0
    nine cycles of hemodialysis | 0
    hyperkalemia corrected | 24
    hypernatremia corrected | 48
    prevention of hepatic encephalopathy | 0
    carbohydrate diet | 0
    lactulose bowel wash | 0
    avoidance of protein diet | 0
    renal functions started improving | 216
    increased renal output | 216
    maintenance of creatinine without dialysis | 216
    parenteral fluid based on CVP monitoring | 0
    daily output chart | 0
    precautions against nosocomial infections | 0
    physiotherapy | 0
    transferred to general ward | 216
    discharged | 504
    improved renal function | 504
    improved liver function | 504
    Grade 5 motor power in both lower limbs | 504
    