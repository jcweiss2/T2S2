fatigue | -72
anosmia | -72
dyspnea | -72
SpO2 levels 55% | -72
nasal cannula oxygen therapy | -72
SpO2 levels improved to 75% | -72
chest radiography | -48
bilateral lung infiltrates | -48
RT-PCR swab tested positive for SARS-CoV-2 infection | -48
admitted in a COVID-19 infirmary unit | 0
non-invasive ventilation support | 0
intubation | 12
invasive mechanical ventilation | 12
ventral decubitus positioning | 12
Escherichia coli detected on sputum culture | 48
methicillin-sensitive Staphylococcus aureus detected on sputum culture | 48
superinfection | 48
amoxicillin prescribed | 48
blood culture revealed methicillin-resistant Staphylococcus aureus | 48
methicillin-resistant Staphylococcus aureus dismissed | 48
steady clinical improvement | 96
extubation | 120
discharged | 168
retrosternal thoracalgia | 168
thoracalgia irradiating to the left upper limb | 168
abduction limited due to pain | 168
external rotation limited due to pain | 168
soft tissue swelling of the shoulder and arm | 168
fever | 168
increased levels of C-reactive protein | 168
hemoculture negative | 168
urine culture negative | 168
chest radiograph performed | 168
thoracic CT performed | 168
typical changes compatible with sequelae of Covid-19 pneumonia | 168
admitted for further investigation and treatment planning | 168
gentamicin prescribed | 168
gentamicin administered | 168
thoracic CT with intravenous contrast administration | 216
scapulohumeral synovitis | 216
intra-muscular collections | 216
glenohumeral joint fluid | 216
bilateral shoulder magnetic resonance imaging (MRI) with intravenous contrast administration | 240
infraspinatus fossa collections | 240
subscapular fossa collections | 240
capsular thickening | 240
increased signal intensity post-gadolinium administration | 240
septic arthritis | 240
rotator cuff collections | 240
myonecrosis | 240
aspiration of the infraspinatus fossa collection | 264
seropurulent fluid | 264
drainage catheter | 264
drainage catheter removed | 264
evaluation of the aspirate | 264
negative results for Mycobacterium tuberculosis | 264
negative results for anaerobic and aerobic bacteria | 264
improvement of left shoulder range of motion | 288
physical rehabilitation exercises | 288
transferred to another hospital | 288
indication to continue physical therapy and rehabilitation exercises | 288