60 years old | 0
    woman | 0
    small median abdominal incisional hernia | -43680
    laparotomic appendectomy | -43800
    acute appendicitis | -43800
    peritoneal abscess | -43800
    abdominal wall bulging in right quadrants | 0
    xipho-pubic scar | 0
    umbilicus | 0
    14 mm diameter tumefaction | 0
    ultrasound scan confirmed diagnosis | 0
    abdominoplasty | 0
    incisional hernia repair | 0
    open keel technique | 0
    xipho-pubic scar excised | 0
    dissection of umbilicus | 0
    supra-umbilical hernia sac | 0
    linear median incision along sub"umbilical linea alba | 0
    preperitoneal plane assessment | 0
    limited viscerolysis | 0
    abdominal wall defect corrected | 0
    rectus abdominis muscle plasty | 0
    Vicryl 1.0 stitches | 0
    umbilicus reconstruction using Santanelli technique | 0
    two Redon type surgical drains placed | 0
    weak peristalsis | 48
    resumption of intestinal flow | 48
    afebrile | 0
    good general conditions | 0
    deambulation started | 48
    bowels open for gas | 72
    bowels open for faeces | 72
    postoperative course uneventful | 0
    normal bowel function | 0
    drains removed | 96
    discharged | 96
    first follow-up | 96
    clean healing wound | 96
    deterged and dressed wound | 96
    four follow-up visits | 120
    stitches removed | 552
    fever episode | 696
    epigastric bulg | 696
    median epigastric bulg | 696
    xipho/umbilical region ballottement | 696
    erythema of overlying skin | 696
    pain during abdominal wall palpation | 696
    60 cc pus drained | 696
    cavity cleaned | 696
    subcutaneous abscess in epigastric region | 696
    purulent material collected | 696
    microbiological testing | 696
    Streptococcus anginosus positive | 696
    antibiotic therapy with Levoxacin 500 mg | 696
    persistent pain | 744
    xipho/umbilical bulge draining purulent exudate | 744
    dyspnoea after rinsing | 744
    chest X-ray showing sub-diaphragmatic free gas | 744
    abdominal CT scan confirming free endoperitoneal gas | 744
    intestinal perforation | 744
    exploratory laparotomy | 744
    plastic peritonitis | 744
    extended right and transverse colectomy | 744
    perforation located | 744
    abscessing mass located | 744
    ileal loops damaged | 744
    right monolateral salpingo-ovariectomy | 744
    temporary ileostomy | 744
    histological examination | 744
    resected small intestines | 744
    resected right colon | 744
    resected right ovary | 744
    resected right Fallopian tube | 744
    haemorrhagic serositis of distal ileum and caecum | 744
    ischaemic necrosis | 744
    ulceration in right colon | 744
    transferred to ICU | 744
    Metronidazole administered | 744
    Levofloxacin administered | 744
    Imipenem administered | 744
    Tigecicline administered | 744
    Fluconazole administered | 744
    ileostomy reversal surgery | 2016
    discharged after reversal | 2016
    
    60 years old | 0
    woman | 0
    small median abdominal incisional hernia | -43680
    laparotomic appendectomy | -43800
    acute appendicitis | -43800
    peritoneal abscess | -43800
    abdominal wall bulging in right quadrants | 0
    xipho-pubic scar | 0
    umbilicus | 0
    14 mm diameter tumefaction | 0
    ultrasound scan confirmed diagnosis | 0
    abdominoplasty | 0
    incisional hernia repair | 0
    open keel technique | 0
    xipho-pubic scar excised | 0
    dissection of umbilicus | 0
    supra-umbilical hernia sac | 0
    linear median incision along sub-umbilical linea alba | 0
    preperitoneal plane assessment | 0
    limited viscerolysis | 0
    abdominal wall defect corrected | 0
    rectus abdominis muscle plasty | 0
    Vicryl 1.0 stitches | 0
    umbilicus reconstruction using Santanelli technique | 0
    two Redon type surgical drains placed | 0
    weak peristalsis | 48
    resumption of intestinal flow | 48
    afebrile | 0
    good general conditions | 0
    deambulation started | 48
    bowels open for gas | 72
    bowels open for faeces | 72
    postoperative course uneventful | 0
    normal bowel function | 0
    drains removed | 96
    discharged | 96
    first follow-up | 96
    clean healing wound | 96
    deterged and dressed wound | 96
    four follow-up visits | 120
    stitches removed | 552
    fever episode | 696
    epigastric bulg | 696
    median epigastric bulg | 696
    xipho(umbilical region ballottement | 696
    erythema of overlying skin | 696
    pain during abdominal wall palpation | 696
    60 cc pus drained | 696
    cavity cleaned | 696
    subcutaneous abscess in epigastric region | 696
    purulent material collected | 696
    microbiological testing | 696
    Streptococcus anginosus positive | 696
    antibiotic therapy with Levoxacin 500 mg | 696
    persistent pain | 744
    xipho/umbilical bulge draining purulent exudate | 744
    dyspnoea after rinsing | 744
    chest X-ray showing sub-diaphragmatic free gas | 744
    abdominal CT scan confirming free endoperitoneal gas | 744
    intestinal perforation | 744
    exploratory laparotomy | 744
    plastic peritonitis | 744
    extended right and transverse colectomy | 744
    perforation located | 744
    abscessing mass located | 744
    ileal loops damaged | 744
    right monolateral salpingo-ovariectomy | 744
    temporary ileostomy | 744
    histological examination | 744
    resected small intestines | 744
    resected right colon | 744
    resected right ovary | 744
    resected right Fallopian tube | 744
    haemorrhagic serositis of distal ileum and caecum | 744
    ischaemic necrosis | 744
    ulceration in right colon | 744
    transferred to ICU | 744
    Metronidazole administered | 744
    Levofloxacin administered | 744
    Imipenem administered | 744
    Tigecicline administered | 744
    Fluconazole administered | 744
    ileostomy reversal surgery | 2016
    discharged after reversal | 2016
    