24 years old | 0
primigravida | 0
37 weeks of gestation | 0
referred to institute | 0
supplemental oxygen (Venturi mask) | 0
Rapid test diagnosis of Plasmodium falciparum malaria | 0
acute icteric leptospirosis | 0
microscopic agglutination test (MAT) titers for Leptospira ictero-haemorrhagiae | 0
high grade fever | -72
decreased urine output | -72
yellowish discolouration | -72
altered sensorium | -72
disoriented | 0
febrile | 0
icteric | 0
sub-conjunctival haemorrhages | 0
fine basal crepitations on auscultation | 0
intravenous artesunate | 0
ceftriaxone | 0
doxycycline capsules | 0
anaemia | 0
jaundice | 0
deranged liver function | 0
coagulopathy | 0
thrombocytopenia | 0
increased total leucocyte count | 0
elevated blood urea nitrogen | 0
serum creatinine | 0
singleton pregnancy | 0
adequate liquor | 0
umbilical artery systolic-diastolic ratio of 2:1 | 0
mild hepato-splenomegaly | 0
emergency caesarean delivery | 0
non-reassuring fetal heart rate | 0
aspiration prophylaxis | 0
high-risk consent | 0
rapid sequence intubation | 0
cricoid pressure | 0
thiopental | 0
succinylcholine | 0
right internal jugular vein cannulation | 0
left radial artery cannulation | 0
baseline serum glucose level normal | 0
isoflurane in N2O-O2 mixture | 0
atracurium | 0
delivery of 2.25 kg baby | 0
fentanyl administration | 0
oxytocin infusion | 0
Apgar score of 6 at 1 min | 0
Apgar score of 8 at 5 min | 0
cord blood pH of 7.28 | 0
base deficit of 5.4 | 0
cord blood sugar level of 50 mg/dl | 0
hypotension after placental separation | 0
packed red blood cells transfusion | 0
fresh frozen plasma transfusion | 0
platelets transfusion | 0
noradrenaline infusion | 0
mild acidosis | 0
normal electrolytes | 0
serum glucose normal | 0
shifted to ICU | 0
intubated state | 0
noradrenaline infusion continued | 0
ultrasound guided bilateral transverse abdominis plane block | 0
pulmonary haemorrhage on second postoperative day | 24
coagulopathy | 24
blood products transfusion | 24
fibre-optic bronchoscopy | 24
erythematous mucosa | 24
blood clots | 24
active oozing | 24
diffuse bleeding from distal airway | 24
broncho alveolar lavage | 24
Factor VIIa administration | 24
bleeding cessation | 24
reduction of inspired oxygen fraction (FiO2) | 24
bilateral non-homogeneous opacities on chest radiograph | 24
chest radiograph almost clear | 24
acute kidney injury | 24
severe hyperbilirubinemia | 24
haemolytic uremic syndrome | 24
high serum lactate dehydrogenase | 24
schistocytes in peripheral blood | 24
plasmapheresis | 24
dialysis | 24
computed tomography of the brain showing diffuse cerebral oedema | 24
cerebroprotective measures | 24
blood cultures negative | 24
urine cultures negative | 24
Weil-Felix test negative | 24
typhi dot negative | 24
dengue serology negative | 24
hepatitis viruses serology negative | 24
stress ulcer prevention | 24
deep vein thrombosis prophylaxis (pneumatic compression) | 24
glycemic control | 24
fever intensity reducing | 96
consciousness improved | 96
inotropic support tapered | 96
urine output improved | 96
liver function test improving trends | 96
coagulation parameters improving trends | 96
Pao2/Fio2 ratio improved | 96
extubation on sixth post-operative day | 144
shifted to wards | 144
discharged from hospital | 144
jaundice |; 0
