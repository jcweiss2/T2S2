71 years old | 0
female | 0
obese | 0
type 2 diabetes | 0
admitted to the hospital | 0
obstructive jaundice | 0
total bilirubin level 13.6 mg/dL | 0
abdominal ultrasound | 0
multiple gallbladder stones | 0
impacted stone in the cystic duct | 0
thickened gallbladder wall | 0
magnetic resonance cholangiopancreatography | 0
ERCP with biliary stent insertion | 0
cholangiography | 0
subhilar stenosis | 0
intrahepatic cholestasis | 0
early stent occlusion | 72
cholangitis | 72
antibiotic treatment with ceftriaxone and metronidazole | 72
discharged | 216
readmission | 504
fever | 504
cholangial sepsis | 504
hypotension | 504
renal failure | 504
CRP value 314 mg/dL | 504
computed tomography | 504
liver abscess | 504
percutaneous drainage | 504
blood culture | 504
Enterococcus faecalis | 504
Streptococcus anginosus | 504
liver abscess culture | 504
vancomycin-resistant Enterococcus faecium | 504
meropenem and linezolid treatment | 504
double pigtail plastic stent exchange | 504
intrahepatic biloma abscess | 504
elevated total bilirubin level 44 mg/dL | 504
prolonged systemic VRE sepsis | 1008
pleural effusions | 1008
articular effusions | 1008
central venous catheter infection | 1008
linezolid-resistant VRE | 1344
core genome multilocus sequence typing | 1344
G2576T mutation | 1344
antimicrobial treatment with meropenem and tigecycline | 1344
double-sided percutaneous biliary drainage | 1344
discharged | 1440
improvement in infection | 1440
re-admission | 1496
cholangial septic shock | 1496
emergency cholecystectomy | 1496
bile duct revision | 1496
t-tube insertion | 1496
histology | 1496
moderate differentiated adenocarcinoma | 1496
gallbladder cancer | 1496
death | 1500