60 years old | 0
male | 0
admitted to the hospital | 0
chronic alcoholic | 0
self-induced vomiting (5–6 episodes per day) | -72
cough | -72
expectoration | -72
hiccups | -72
altered behavior | -72
dizziness | -72
fall in washroom | -24
past history of admission for symptomatic hyponatremia | -264
serum sodium: 123 mEq L−1 | -264
serum potassium: 4.9 mEq L−1 | -264
managed with 3% hypertonic saline | -264
serum sodium was 129 mEq L−1 within 12 hours | -264
rate of correction maintained at 0.5 mEq L−1 per hour | -264
symptomatically improved | -264
discharged home on sixth day of hospital stay | -264
presented to neurology department after 10 days of discharge | 240
complain of imbalance | 240
slurred speech | 240
drowsiness | 240
fever | 240
cough | 240
systemic examination | 240
Glasgow Coma Scale E4V1M1 | 240
hypertonic bilateral upper and lower limbs | 240
hyperreflexia | 240
bilateral extensor plantar | 240
nystagmus | 240
restricted extraocular muscle movements | 240
shifted to ICU | 240
intubated | 240
antibiotics | 240
antimalarials | 240
stress ulcer prophylaxis | 240
deep venous thrombosis prophylaxis | 240
injection thiamine | 240
intravenous fluids | 240
differential diagnosis of CPM | 240
extrapontine myelinolysis | 240
subdural hemorrhage | 240
associated sepsis with delirium | 240
hepatic encephalopathy | 240
Wernicke–Korsakoff syndrome | 240
autoimmune encephalitis | 240
routine blood investigations within normal limits | 240
urine investigations within normal limits | 240
radiological investigations within normal limits | 240
MRI brain showing hyperintensities in central pons | 240
hyperintensities forming trident pattern in upper pons | 240
involvement of tegmentum of midbrain | 240
bilateral thalamic involvement | 240
parts of globus pallidus involvement | 240
supportive management | 240
tracheostomy on seventh day of ICU stay | 312
poor cough reflex | 312
absent gag reflex | 312
gradually weaned from ventilator | 312
put on T-piece | 312
multidisciplinary management | 312
neurology opinion | 312
ophthalmology opinion | 312
psychiatry opinion | 312
physical medicine rehabilitation opinion | 312
medicine opinion | 312
conscious oriented (GCS – E4VTM6) | 312
vitals stable | 312
rigidity persisted in all four limbs | 312
hyperreflexia persisted in all four limbs | 312
shifted from ICU | 312
followed up until discharge | 312
continuous cycles of physical rehabilitation | 312
able to walk with support over 2 months | 312
discharged | 312
