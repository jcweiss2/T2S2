47 years old | 0
man | 0
alcohol-induced dilated cardiomyopathy | 0
chronic atrial fibrillation | 0
admitted for New York Heart Association class IV dyspnea | 0
history of excess alcohol consumption | -175200
more than 100 g of alcohol daily | -175200
over 20 years | -175200
hospitalized 4 times in a 7-year period | -504
symptoms of heart failure | -504
presented with dyspnea | 0
presented with azotemia | 0
managed with continuous infusion of dobutamine | 0
managed with continuous infusion of milrinone | 0
managed with continuous renal replacement therapy | 0
experienced cardiac arrest | 792
ventricular fibrillation | 792
returned to spontaneous circulation | 792
transthoracic echocardiography showed decreased left ventricular systolic function | 0
tricuspid annular plane systolic excursion, 8.5 mm | 0
severe mitral regurgitation | 0
severe tricuspid regurgitation | 0
inferior vena cava was dilated | 0
diameter of 3.1 cm | 0
associated plethora | 0
right ventricular systolic pressure was 44.3 mm Hg | 0
severe cardiomegaly | 0
pericardial effusion | 0
could not lay supine | 0
right heart catheterization could not be performed | 0
serum creatinine level was 1.81 mg/dL | 0
estimated glomerular filtration rate was 40.4 mL/min/m2 | 0
total bilirubin level was 3.1 mg/dL | 0
recent alcohol abuser | 0
extensive discussion on further management of severe heart failure | 0
psychiatric evaluation | 0
psychologically dependent on alcohol | 0
physiologically dependent on alcohol | 0
wife and parents planned to provide psychosocial support | 0
accepted their plan | 0
agreed to proceed with left ventricular assist device (LVAD) insertion | 0
agreed to proceed with tricuspid annuloplasty | 0
severe right ventricular failure | 0
LVAD offered under the condition of remaining alcohol-free for at least 6 months | 0
possible later heart transplantation | 0
performed surgery | 1176
median sternotomy performed | 1176
cardiopulmonary bypass initiated | 1176
arterial cannulation into the ascending aorta | 1176
bicaval venous cannulation performed | 1176
without aortic cross-clamping | 1176
right atriotomy | 1176
beating heart tricuspid annuloplasty performed | 1176
Carpentier Edwards MC3 30-mm ring used | 1176
left ventricular apex sutured with a sewing ring | 1176
incised | 1176
fixed with an LVAD inflow cannula | 1176
driveline pulled out through left upper quadrant abdominal wall | 1176
double-tunnel technique used | 1176
outflow cannula anastomosed to the right side of the proximal ascending aorta | 1176
LVAD initiated | 1176
careful de-airing | 1176
successfully weaned from cardiopulmonary bypass | 1176
inotropic support with dobutamine [3 μg/kg/min] | 1176
inotropic support with milrinone [0.7 μg/kg/min] | 1176
LVAD flow increased to 4.5 L/min at 2,500 rpm | 1176
stable vital signs | 1176
transferred to the cardiovascular intensive care unit (ICU) | 1176
stable for a few hours | 1176
awoke | 1176
coughed | 1176
hypotension developed | 1176
tachycardia developed | 1176
inotrope infusion | 1176
nitric oxide inhalation | 1176
still unstable | 1176
mean arterial blood pressure (MBP) 40 mm Hg | 1176
high central venous pressure (CVP; range, 15–18 mm Hg) | 1176
low LVAD flow (2.5 L/min) | 1176
low pulmonary arterial pressure | 1176
systolic pulmonary arterial pressure 23 mm Hg | 1176
diastolic pulmonary arterial pressure 15 mm Hg | 1176
decided to perform emergent insertion of extracorporeal right ventricular assist device (RVAD) | 1176
veno-pulmonary artery extracorporeal life support | 1176
performed in ICU | 1176
avoid repeat sternotomy | 1176
percutaneous femoral venous cannulation | 1176
pulmonary artery cannulation via left anterior mini-thoracotomy | 1176
22F venous cannula inserted into femoral vein | 1176
Seldinger technique used | 1176
left anterior thoracotomy performed at second intercostal space | 1176
double purse-string suturing | 1176
return arterial cannulation (15F) placed in main pulmonary artery | 1176
extracorporeal RVAD initiated with flow of 4.4 L/min | 1176
LVAD flow increased to 4.7 L/min at 2,500 rpm | 1176
thoracotomy closed | 1176
maintaining stable LVAD flow | 1176
after RVAD implantation | 1176
inhaled nitric oxide tapered | 1176
stable hemodynamics | 1176
CVP of 8 mm Hg | 1176
MBP >60 mm Hg | 1176
heart rate 80–90/min | 1176
RVAD rpm and flow rates slowly decreased | 1176
spontaneous recovery of right ventricular systolic function | 1176
RVAD removed | 1584
general anesthesia in ICU | 1584
return cannulation into main pulmonary artery removed | 1584
redo thoracotomy using previous incision | 1584
venous cannulation removed from right femoral insertion site | 1584
transferred to general ward | 1752
resolution of lower leg pitting edema | 1752
rehabilitation therapy | 1752
discharged | 3096
noncompliant with medical therapy | 3096
readmitted for recurrent alcohol abuse | 3096
subsequent right ventricular failure | 3096
LVAD turned off due to irreversible septic encephalopathy | 6024
coma | 6024
impossible to get written informed consent | 6024
presented with azotemia |6 0
