47 years old| 0
female | 0
hypertension | 0
chronic kidney disease-5 | 0
thrice weekly hemodialysis | 0
cough | -672
expectoration | -672
breathlessness | -672
fever | -240
managed in outside facility | -168
amlodipine | -168
erythropoietin | -168
imipenem | -168
hemodialysis | -168
supportive care for CKD | -168
presentation | 0
conscious | 0
well-oriented | 0
heart rate 116 beats/min | 0
non-invasive blood pressure 108/66 mmHg | 0
temperature 100.2°F | 0
respiratory rate 34/min | 0
accessory muscles used | 0
bilateral normal vesicular breath sounds | 0
decreased air entry | 0
occasional coarse crepts | 0
right lower lobe consolidation/collapse | 0
pleural effusion | 0
blood cultures sterile | 0
urine cultures sterile | 0
managed in medical ICU | 0
non-invasive ventilation | 0
injection imipenem 500 mg BID | 0
received imipenem for 2 days prior to admission | -48
clinical deterioration on 3rd day of admission | 72
TLC 28,600/mm3 | 72
repeat blood cultures | 72
teicoplanin | 72
caspofungin | 72
provisional report of gram-negative coccobacilli | 96
Acinetobacter baumannii | 96
colistin 1 MU OD | 96
colistin loading dose 2 MU | 96
fever decrease | 168
TLC decrease | 168
caspofungin de-escalated | 168
imipenem stopped after 10 days | 240
off and on low-grade fever | 0
alternate day hemodialysis | 0
sudden onset facial twitchings | 384
circumoral twitchings | 384
neck twitchings | 384
seizures controlled with midazolam | 384
phenytoin 1 g IV | 384
phenytoin 100 mg BID | 384
another episode of seizures | 384
generalized tonic clonic seizures | 384
midazolam 1 mg + 1 mg IV bolus | 384
levirecetam 1 g IV | 384
levirecetam 500 mg BID | 384
no acute metabolic derangements | 384
normal liver profile | 384
normal neuroimaging | 384
normal electroencephalography | 384
normal nerve conduction velocity | 384
lumbar puncture | 384
clear CSF | 384
normal CSF pressure | 384
CSF glucose 56 mg/dl | 384
CSF proteins 37 | 384
CSF TLC nil | 384
imipenem stopped 1 week prior to seizures | 384
colistimethate considered causative agent | 384
colistin stopped | 384
blood cultures sterile after 48 h | 432
no recurrence of seizures | 432
antiepileptics tapered after 1 week | 432
shifted to ward | 792
discharged after 33 days | 792
