58 years old | 0
female | 0
Hispanic | 0
admitted to the hospital | 0
fever | -120
dizziness | -120
hypertension | -8760
denies dyspnea | 0
denies cough | 0
denies chills | 0
denies night sweats | 0
denies headache | 0
denies gastrointestinal symptoms | 0
no history of anorexia | 0
no history of weight loss | 0
born in the Dominican Republic | -524160
moved to New York City | -175680
denies use of tobacco | 0
denies use of alcohol | 0
denies use of recreational drugs | 0
febrile | 0
hypotensive | 0
cervical lymph nodes palpable | 0
bilateral rhonchi | 0
abdominal examination unremarkable | 0
neurological examination unremarkable | 0
cardiac examination unremarkable | 0
no organomegaly | 0
skin intact | 0
diffuse bilateral infiltrates on chest radiograph | 0
leukopenia | 0
thrombocytopenia | 0
elevated serum lactate dehydrogenase | 0
received IV fluids | 0
received ceftriaxone | 0
received azithromycin | 0
persistent fever | 0
blood cultures negative | 0
urine cultures negative | 0
respiratory cultures negative | 0
acid-fast bacilli stains negative | 0
antibiotics changed to IV piperacillin-tazobactam | 0
antibiotics changed to IV vancomycin | 0
transthoracic echocardiogram normal | 0
computed tomography of chest revealed bilateral infiltrates | 0
computed tomography of chest revealed mediastinal and subcarinal lymphadenopathy | 0
mild splenomegaly on CT of abdomen | 0
underwent flexible fiber optic bronchoscopy | 144
underwent bronchoalveolar lavage | 144
underwent transbronchial biopsies | 144
underwent endobronchial ultrasound transbronchial needle aspiration | 144
all cultures from FFB negative | 144
pathology from TBNA revealed T cell lymphoma | 144
CD4 positive | 144
CD3 positive | 144
CD43 positive | 144
BCL-2 positive | 144
CD20 negative | 144
CD10 negative | 144
CD79a negative | 144
PAX5 negative | 144
clinical condition deteriorated | 360
developed hypoxic respiratory failure | 360
required intubation and mechanical ventilation | 360
cervical lymph node excisional biopsy | 360
pathology of lymph node biopsy positive for peripheral T-cell lymphoma | 360
immunohistochemical stain results consistent with T cell lymphoma | 360
CD3 positive | 360
CD4 positive | 360
CD5 positive | 360
CD43 positive | 360
Ki67 positive | 360
CD20 negative | 360
CD79A negative | 360
CD7 negative | 360
CD15 negative | 360
bone marrow biopsy revealed hemophagocytic lymphocytic histiocytosis | 456
stains of bone marrow for AFB and fungal infection negative | 456
developed tumor lysis syndrome | 456
developed acute renal failure | 456
required hemodialysis | 456
required rasburicase | 456
cyclophosphamide started | 456
vincristine started | 456
patient died | 480
cultures for AFB from cervical lymph nodes positive | 480
Mycobacterium tuberculosis complex identified | 480
pathology stain demonstrated AFB | 480