36 years old | 0
female | 0
gravida 4 | 0
para 3 | 0
pregnant | 0
16 weeks and 1 day pregnant | 0
lower abdominal and flank pain | -24
vaginal spotting | -24
mild dysuria | -24
urinary frequency | -24
urgency | -24
no fever | -24
no chills | -24
no sick contacts | -24
referred to the emergency department | -24
arrived in the United States from Pakistan | -672
blood pressure of 103/70 mmHg | -24
heart rate of 133 bpm | -24
temperature of 99.9°F | -24
respiratory rate of 16 per minute | -24
oxygen saturation of 99% | -24
tachycardia | -24
suprapubic tenderness | -24
pelvic examination with slight bleeding | -24
no uterine tenderness | -24
leukocytosis of 16.1 K/μL | -24
88% polymorphonuclear leukocytes | -24
normal complete blood count | -24
normal chemistry panels | -24
normal urinalysis | -24
live intrauterine pregnancy | -24
estimated gestational age of 16 weeks and 0 days | -24
fetal heart rate of 182 beats per minute | -24
normal MRI of the abdomen | -24
no evidence of appendicitis | -24
received 4 liters of normal saline | -24
received 2 mg of morphine sulfate | -24
received 975 mg of acetaminophen | -24
heart rate improved to 100 bpm | -24
felt better | -24
discharged home | -24
returned to the ED with sudden onset of vaginal bleeding | 24
abdominal pain | 24
heart rate of 139 bpm | 24
blood pressure of 149/88 mmHg | 24
respiratory rate of 30 per minute | 24
oxygen saturation of 100% | 24
actively delivering the products of conception | 24
delivered an intact fetus and gestational sac | 24
received 800 mg of rectal misoprostol | 24
tympanic temperature of 105°F | 24
persistently tachycardic | 24
hemodynamically unstable | 24
blood pressure of 84/35 mmHg | 24
central intravenous access obtained | 24
given acetaminophen | 24
given intravenous normal saline | 24
given vancomycin | 24
given piperacillin/tazobactam | 24
working diagnosis of sepsis of unknown etiology | 24
venous pH of 7.22 | 24
anion gap of 21 | 24
lactate concentration of 10.8 mmol/L | 24
white blood cell count of 14.9 K/μL | 24
85% polymorphonuclear leukocytes | 24
normal MRI findings | 24
normal urinalysis findings | 24
no symptoms to suggest colitis | 24
no symptoms to suggest skin infection | 24
no symptoms to suggest other soft tissue infections | 24
given norepinephrine | 24
admitted to the medical intensive care unit | 24
received ampicillin | 24
received gentamycin | 24
received clindamycin | 24
suspected chorioamnionitis | 24
ultrasonogram suggestive of retained products of conception | 48
underwent dilatation and curettage | 48
removal of tissue debris | 48
discharged from the hospital | 96
blood cultures came back positive for H influenzae | 24
non–β-lactamase producing | 24
pathology report showed retroplacental hemorrhage | 48
placental abruption | 24
no histologic evidence of acute chorioamnionitis | 48