101 years old | 0
male | 0
Ashkenazi Jewish | 0
admitted to the hospital | 0
pulmonary oedema | 0
mechanical ventilation | 0
tracheostomy | 24
gram-negative bacteraemia | 168
sepsis | 168
haemodynamic instability | 168
oliguric | 840
acidemic | 840
rise in creatinine level | 840
abdominal aortic aneurysm | -8760
ischaemic heart disease | -8760
tricuspid regurgitation | -8760
pulmonary hypertension | -8760
congestive heart failure | -8760
pacemaker insertion | -8760
chronic kidney disease | -8760
diabetes | -8760
cardiorenal syndrome | -8760
intellectual capacity preserved | -8760
active rabbi and teacher | -8760
extremely frail | 840
unable to speak | 840
decreased level of consciousness | 840
uraemic encephalopathy | 840
haemodialysis | 840
cuffed, tunneled catheter | 840
dialysis initiated | 840
56 haemodialysis treatments | 840
death | 3360
acute on chronic renal failure | 840
poor functional status | 840
comorbidities | 840
advanced age | 840
multi organ failure | 840
preexisting CKD | 840
initiation of haemodialysis | 840
nursing home resident | -8760
uraemia | -8760
improved quality of life | -8760
improved mental status | -8760
decision to start haemodialysis | 840
aggressive treatments | 840
poor prognosis | 840
futile treatments | 840
empirically define futile treatments | 840
Renal Physicians Association guidelines | 840
American Society of Nephrology guidelines | 840
Shared Decision-Making | 840
initiation of and withdrawal from dialysis | 840
conflict resolution processes | 840
time limited trials of dialysis | 840
law in most jurisdictions | 840
Texas Advance Directive Act of 1999 | 840
Dying Patient Act of 2005 | 840
withhold life-sustaining treatments | 840
patient autonomy | 840
excessive suffering | 840
Ultra-Orthodox Judaism | 840
supreme sanctity of human life | 840
modest prolongation of life | 840
undue suffering | 840
excessive pain and suffering | 840
resource utilization | 840
treatment costs | 840
allocation of nursing and technician staff | 840
time in ICU | 840