47 years old|0
female|0
admitted to the oncology ward|0
low abdominal pain|-1440
nausea|-1440
vomiting|-1440
hyporexia|-1440
dehydration|-1440
weight loss|-1440
hypogastric mass|0
ascites|0
asymmetric edema in right calf|0
deep venous thrombosis (DVT)|0
Eastern Cooperative Oncology Group performance status (ECOG-PS) 3|0
anemia|0
hemoglobin 10.6 g/dL|0
normal electrolytes|0
ionic calcium|0
preserved renal function|0
preserved hepatic function|0
pelvic mass (21 × 11 × 16 cm) in right adnexal region|0
infiltration of left hepatic lobe|0
infiltration of peritoneum|0
multiple para-aortic lymph nodes|0
multiple iliac lymph nodes|0
bilateral pleural effusion|0
pleural fluid positive for neoplastic cells|0
ascitic fluid positive for neoplastic cells|0
image-guided biopsy of peritoneal nodule|0
poorly differentiated small-cell neoplasia|0
solid pattern|0
CD56 positive|0
vimentin positive|0
cytokeratins 35BH11 focally positive|0
WT1 negative|0
estrogen receptor negative|0
TTF-1 negative|0
inhibin negative|0
carcinoma with neuroendocrine differentiation|0
ovarian biopsy|0
emergency laparotomy|0
acute peritonitis|0
poorly differentiated small-cell neoplasia with extensive necrosis|0
CD99 focally positive|0
cytokeratin negative|0
S-100 negative|0
desmin negative|0
WT-1 negative|0
primitive neuroectodermal tumor (PNET) suspected|0
FLI-1 protein assay|0
peritoneal nodule FLI-1 focally positive|0
ovarian specimen FLI-1 focally positive|0
diagnosis of undifferentiated carcinoma with neuroendocrine differentiation|0
small-cell ovarian carcinoma (SCOC) hypercalcemic type|0
venous hydration|0
anticoagulation with low-molecular weight heparin|0
systemic chemotherapy with cisplatin and etoposide|0
cisplatin 80mg/m2 on day 1|0
etoposide 80mg/m2 on days 1, 2, & 3|0
significant reduction of abdominal mass|0
improvement of ECOG performance status to 2|0
serum uric acid 13.1 mg/dL|48
serum potassium 6.6 mEq/L|48
serum phosphate 9.7 mg/dL|48
tumor lysis syndrome (TLS) diagnosis|48
intravenous hydration with saline|48
second chemotherapy cycle|672
septic shock|1008
febrile neutropenia|1008
acute peritonitis|1008
admission to Intensive Care Unit|1008
broad-spectrum antibiotics|1008
emergency laparotomy|1008
no bowel perforation|1008
necrotic adnexal mass|1008
abscess resected|1008
death due to sepsis|1680
