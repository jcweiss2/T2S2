85 years old | 0
male | 0
type 2 diabetes mellitus | -672
hypertension | -672
dyslipidemia | -672
iron deficiency anemia | -672
chronic kidney disease | -672
dementia | -672
furosemide | -672
hydralazine | -672
β-blocker | -672
ferrous sulphate | -672
reduced oral intake | -168
recurrent vomiting | -168
decreased level of consciousness | -168
severely dehydrated | 0
hypotensive | 0
mildly tachypneic | 0
Glasgow coma scale of 11 | 0
melena | 0
leukocytosis | 0
low hemoglobin | 0
high C-reactive protein | 0
high urea | 0
acute kidney injury | 0
elevated lactate | 0
elevated procalcitonin | 0
urinary tract infection | 0
admitted to the intensive care unit | 0
severe sepsis | 0
hemoglobin dropped | 48
esophagogastroduodenoscopy | 48
hiatus hernia | 48
Hill's classification grade 4 | 48
sessile polyp | 48
Paris classification of 0-Is | 48
gastric pseudomelanosis | 48
duodenal pseudomelanosis | 48
histological examination | 48
intact lining epithelium | 48
brownish-black pigment-laden macrophages | 48
Perl's Prussian blue stain positive | 48
iron deposition | 48
hyperplastic duodenal polyp | 48
urosepsis managed with antibiotics | 48
kidney injury managed conservatively | 48
intravenous fluids | 48
supportive measures | 48
transferred to the wards | 120
renal function back to baseline | 120
septic markers improved | 120
discharged home | 288
full recovery | 288