27 years old | 0
male | 0
mitochondrial neurogastrointestinal encephalopathy disease | -672
percutaneous endoscopic gastrostomy | -672
total parenteral nutrition | -672
central catheter line | -672
jejunal diverticulosis | -672
pseudo-obstructions | -672
partial small bowel resection | -672
insulin-dependent type I diabetes mellitus | -672
admitted to the hospital | 0
fever | 0
vomiting | 0
abdominal pain | 0
core temperature of 38.5°C | 0
heart rate of 120 beat/min | 0
blood pressure of 120/70 mmHg | 0
rapid heart sounds | 0
no additional heart sounds or murmurs | 0
no abnormalities on lung auscultation | 0
mild abdominal tenderness | 0
marked redness around the central catheter line | 0
pussy secretion | 0
no stigmata of endocarditis | 0
leukocytosis | 0
WBC 20 K/uL | 0
C-reactive protein 25 mg/dL | 0
acute kidney injury | 0
creatinine 1.3 mg/dL | 0
urea 50 mg/dL | 0
diabetic ketoacidosis | 0
serum glucose level 420 mg/dL | 0
positive ketones in peripheral blood | 0
metabolic acidosis | 0
pH 7.2 | 0
pCO2 32 mmHg | 0
HCO3 11 mmHg | 0
regular sinus rhythm | 0
RR interval of 120 | 0
normal axis | 0
no PR or QT segment prolongation | 0
no changes in ST segments or T waves | 0
normal chest X-ray | 0
gastric distention | 0
no signs of obstruction or perforation | 0
central line-associated bloodstream infection | 0
central line removed | 0
blood cultures sent | 0
anti-staphylococcal antibiotic initiated | 0
hypoxemic respiratory failure | 24
intubated | 24
moved to the intensive care unit | 24
bilateral consolidations with hyperdensities | 24
marked bilateral consolidations | 24
hyperdensities in the apex and base of the right lung | 24
preserved function on TTE | 48
no obvious vegetations on TTE | 48
mild mitral and tricuspid regurgitations | 48
small mobile mass on the eustachian valve | 48
large 2×1.5 cm vegetation at the anterior leaflet of the mitral valve | 48
no echo-cardiographic evidence of an intra-atrial shunt | 48
refractory septic shock | 72
conservative approach with extended antibiotics regimen | 72
positive MSSA cultures | 96
hemodynamic and respiratory deterioration | 96
vasopressor support | 96
massive bilateral consolidations with cavitation | 120
septation on the right upper quadrant | 120
septic emboli | 120
large frontoparietal infarct | 120
middle cerebral artery occlusion | 120
ventilation-associated pneumonia | 144
disseminated intravascular coagulopathy | 144
death | 168