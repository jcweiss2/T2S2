32 years old | 0
male | 0
admitted to the emergency department | 0
beating | 0
multiple blunt trauma | 0
no penetrating injury | 0
Glasgow Coma Scale score 10 | 0
heart rate 95 | 0
blood pressure 120/80 mmHg | 0
loss of consciousness | 0
no nausea | 0
no vomiting | 0
pain on bilateral upper quadrants | 0
no abdominal tenderness | 0
no rebound tenderness | 0
no abdominal rigidity | 0
no hematuria | 0
leukocytosis 30,000×106/ml | 0
hemoglobin 14.8 g/dl | 0
AST 496 U/l | 0
ALT 940 U/l | 0
direct bilirubin 0.44 mg/dl | 0
total bilirubin 0.82 mg/dl | 0
computed tomography scan with IV contrast | 0
right parietal bone depression fracture | 0
free perihepatic fluid | 0
free perisplenic fluid | 0
splenic laceration suspected | 0
observation | 0
another abdominal CT scan | 4
cranial CT | 4
increased perihepatic fluid | 4
heterogeneous appearance at falciform ligament | 4
focal enlargement of duodenum | 4
mural thickening of duodenum | 4
initial diagnosis of bleeding from liver laceration | 4
neurosurgeons decided to operate | 4
postoperative follow-up in neurosurgical ICU | 4
decreased pain on abdomen | 24
leukocyte count decreased to 15,800×106/ml | 24
AST 2265 U/l | 24
ALT 2224 U/l | 24
Hgb 9.5 g/dl | 24
evaluated by general surgery team | 48
tachycardia | 48
tenderness on four quadrants of abdomen | 48
total bilirubin 24.63 mg/dl | 48
serum total bilirubin 8.69 mg/dl | 48
direct bilirubin 10.8 mg/dl | 48
serum direct bilirubin 5.7 mg/dl | 48
urea 48 mg/dl | 48
serum urea 39 mg/dl | 48
creatinine 0.93 mg/dl | 48
serum creatinine 1.08 mg/dl | 48
amylase 214 U/l | 48
serum amylase 310 U/l | 48
exploratory laparotomy | 48
intestines covered with bile | 48
free bile in abdomen | 48
no gastric perforation | 48
no intestinal perforation | 48
common hepatic duct fully transected | 48
cholecystectomy | 48
instability of patient | 48
inflammation on tissues | 48
decision to wait for hepaticojejunostomy | 48
drain placed to common hepatic duct | 48
multiple drains placed | 48
operation ended | 48
postoperative follow-up in general surgery ward | 48
abdominal drains removed day by day | 48
discharged postoperatively 10th day | 240
biliary drain changed for percutaneous drainage | 720
patient did not follow regular appointments | 720
continued with percutaneous drain | 720
accepted second operation | 8760
Roux-en-Y hepaticojejunostomy applied | 8760
discharged postoperatively 10th day | 8770
full recovery | 8770
blood pressure 120/80 mmHg |$[{'timestamp': 0, 'event': '32 years old'}, {'timestamp': 0, 'event': 'male'}, {'timestamp': 0, 'event': 'admitted to the emergency department'}, {'timestamp': 0, 'event': 'beating'}, {'timestamp': 0, 'event': 'multiple blunt trauma'}, {'timestamp': 0, 'event': 'no penetrating injury'}, {'timestamp': 0, 'event': 'Glasgow Coma Scale score 10'}, {'timestamp': 0, 'event': 'heart rate 95'}, {'timestamp': 0, 'event': 'blood pressure 120/80 mmHg'}, {'timestamp': 0, 'event': 'loss of consciousness'}, {'timestamp': 0, 'event': 'no nausea'}, {'timestamp': 0, 'event': 'no vomiting'}, {'timestamp': 0, 'event': 'pain on bilateral upper quadrants'}, {'timestamp': 0, 'event': 'no abdominal tenderness'}, {'timestamp': 0, 'event': 'no rebound tenderness'}, {'timestamp': 0, 'event': 'no abdominal rigidity'}, {'timestamp': 0, 'event': 'no hematuria'}, {'timestamp': 0, 'event': 'leukocytosis 30,000×106/ml'}, {'timestamp': 0, 'event': 'hemoglobin 14.8 g/dl'}, {'timestamp': 0, 'event': 'AST 496 U/l'}, {'timestamp': 0, 'event': 'ALT 940 U/l'}, {'timestamp': 0, 'event': 'direct bilirubin 0.44 mg/dl'}, {'timestamp': 0, 'event': 'total bilirubin 0.82 mg/dl'}, {'timestamp': 0, 'event': 'computed tomography scan with IV contrast'}, {'timestamp': 0, 'event': 'right parietal bone depression fracture'}, {'timestamp': 0, 'event': 'free perihepatic fluid'}, {'timestamp': 0, 'event': 'free perisplenic fluid'}, {'timestamp': 0, 'event': 'splenic laceration suspected'}, {'timestamp': 0, 'event': 'observation'}, {'timestamp': 4, 'event': 'another abdominal CT scan'}, {'timestamp': 4, 'event': 'cranial CT'}, {'timestamp': 4, 'event': 'increased perihepatic fluid'}, {'timestamp': 4, 'event': 'heterogeneous appearance at falciform ligament'}, {'timestamp': 4, 'event': 'focal enlargement of duodenum'}, {'timestamp': 4, 'event': 'mural thickening of duodenum'}, {'timestamp': 4, 'event': 'initial diagnosis of bleeding from liver laceration'}, {'timestamp': 4, 'event': 'neurosurgeons decided to operate'}, {'timestamp': 4, 'event': 'postoperative follow-up in neurosurgical ICU'}, {'timestamp': 24, 'event': 'decreased pain on abdomen'}, {'timestamp': 24, 'event': 'leukocyte count decreased to 15,800×106/ml'}, {'timestamp': 24, 'event': 'AST 2265 U/l'}, {'timestamp': 24, 'event': 'ALT 2224 U/l'}, {'timestamp': 24, 'event': 'Hgb 9.5 g/dl'}, {'timestamp': 48, 'event': 'evaluated by general surgery team'}, {'timestamp': 48, 'event': 'tachycardia'}, {'timestamp': 48, 'event': 'tenderness on four quadrants of abdomen'}, {'timestamp': 48, 'event': 'total bilirubin 24.63 mg/dl'}, {'timestamp': 48, 'event': 'serum total bilirubin 8.69 mg/dl'}, {'timestamp': 48, 'event': 'direct bilirubin 10.8 mg/dl'}, {'timestamp': 48, 'event': 'serum direct bilirubin 5.7 mg/dl'}, {'timestamp': 48, 'event': 'urea 48 mg/dl'}, {'timestamp': 48, 'event': 'serum urea 39 mg/dl'}, {'timestamp': 48, 'event': 'creatinine 0.93 mg/dl'}, {'timestamp': 48, 'event': 'serum creatinine 1.08 mg/dl'}, {'timestamp': 48, 'event': 'amylase 214 U/l'}, {'timestamp': 48, 'event': 'serum amylase 310 U/l'}, {'timestamp': 48, 'event': 'exploratory laparotomy'}, {'timestamp': 48, 'event': 'intestines covered with bile'}, {'timestamp': 48, 'event': 'free bile in abdomen'}, {'timestamp': 48, 'event': 'no gastric perforation'}, {'timestamp': 48, 'event': 'no intestinal perforation'}, {'timestamp': 48, 'event': 'common hepatic duct fully transected'}, {'timestamp': 48, 'event': 'cholecystectomy'}, {'timestamp': 48, 'event': 'instability of patient'}, {'timestamp': 48, 'event': 'inflammation on tissues'}, {'timestamp': 48, 'event': 'decision to wait for hepaticojejunostomy'}, {'timestamp': 48, 'event': 'drain placed to common hepatic duct'}, {'timestamp': 48, 'event': 'multiple drains placed'}, {'timestamp': 48, 'event': 'operation ended'}, {'timestamp': 48, 'event': 'postoperative follow-up in general surgery ward'}, {'timestamp': 48, 'event': 'abdominal drains removed day by day'}, {'timestamp': 240, 'event': 'discharged postoperatively 10th day'}, {'timestamp': 720, 'event': 'biliary drain changed for percutaneous drainage'}, {'timestamp': 720, 'event': 'patient did not follow regular appointments'}, {'timestamp': 720, 'event': 'continued with percutaneous drain'}, {'timestamp': 8760, 'event': 'accepted second operation'}, {'timestamp': 8760, 'event': 'Roux-en-Y hepaticojejunostomy applied'}, {'timestamp': 8770, 'event': 'discharged postoperatively 10th day'}, {'timestamp': 8770, 'event': 'full recovery'}]
no rebound tenderness |# 动态规划
