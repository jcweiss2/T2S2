2.980 Kg | 0
male | 0
born trans-vaginally | 0
40-week gestation | -2800
prolonged second stage of labour | -1
prolonged third stage of labour | -1
perinatal asphyxia | 0
non-invasive ventilation | 0
oxygen saturation 80% | 0
intubated | 0
Apgar score 4 | 0
Apgar score 7 | 5
Apgar score 10 | 10
transferred to NICU | 10
blood pressure 70/50 mm Hg | 10
heart rate 144 beats/min | 10
breathing rate 66/min | 10
respiratory distress | 48
afebrile | 48
tachypnic | 48
no history of aspiration | 48
no lethargy | 48
no rash | 48
blood pressure 52/38 mm Hg | 48
pulse rate 186/min | 48
S1 and S2 muffled | 48
lungs clear on auscultation | 48
low voltage QRS complex | 48
non-specific ST-T wave changes | 48
mild leucocytosis | 48
normal cardiac troponin | 48
normal myocardial enzymes | 48
halo sign on chest X-ray | 48
endotracheal tube in right main bronchus | 48
air bubbles in pericardial sac on echocardiography | 48
diastolic collapse of right atrium and right ventricular outflow tract | 48
cardiac tamponade | 48
normal bi-ventricular functions | 48
infection ruled out | 48
sepsis ruled out | 48
ARDS ruled out | 48
myocarditis ruled out | 48
pericardiocentesis planned | 48
intravenous fluid started | 48
ceftriaxone administered | 48
sub-costal area prepared | 48
skin infiltrated with xylocaine | 48
needle entered into pericardial cavity | 48
air bubbles in syringe | 48
guide wires inserted | 48
radial angiographic sheath inserted | 48
wire and dilator removed | 48
sheath left in situ | 48
air aspirated from underwater seal | 48
hemodynamic stability restored | 48
blood pressure rose to 66/42 mm Hg | 48
endotracheal tube repositioned | 48
repeated ECG showed minimal air on anterior cardiac surface | 72
pericardial sheath removed | 72
repeated chest X-ray showed complete resolution of PPC | 72
weaned off mechanical ventilation | 168
discharged | 240