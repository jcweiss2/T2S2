39 years old | 0
male | 0
admitted to the hospital | 0
temperature of 38°C | 0
abdominal pain | 0
7-day diarrhea | 0
tachycardia | 0
tachypnea | 0
leucocytosis | 0
raised serum transaminases | 0
inflammatory markers | 0
C-reactive protein level of 308 mg/l | 0
procalcitonin level of 39 ng/l | 0
multiple liver abscesses | 0
empirical antibiotic treatment with i.v. meropenem | 0
acute clinical deterioration | 1
transferred to surgical Intensive Care Unit (ICU) | 1
endotracheally intubated | 1
mechanical ventilation | 1
vasopressor support | 1
septic shock | 1
percutaneous CT-guide drainage of the liver abscesses | 2
micro-biological samples obtained | 2
liver aspirate revealed a positive visualization on the wet-mount slide of structures of 15–20 µm in diameter | 5
compatible with E. histolytica trophozoites | 5
genomic DNA isolated from clinical samples | 5
detection of Entamoeba histolytica DNA by real-time PCR (RT-PCT) | 5
i.v. metronidazole 750 mg 3 times daily | 5
oral paromomycin, 750 mg 3 times daily | 5
respiratory deterioration | 6
thoracoabdominal CT scan | 6
bilateral pleural effusion | 6
abscess in the right lower pulmonary lobe | 6
small disseminated intraabdominal abscesses | 6
amebic skin lesions on the chest and face | 10
RT- PCR for E. histolytica were positive in all samples obtained | 10
HIV serology and PCR for Acanthamoeba spp, Balamuthia mandrillaris, and Naegleria fowleri were negative | 10
neurological symptoms with aphasia and right-sided hemiplegia | 15
cranial CT scan | 15
multiple brain abscesses in left basal ganglia and in the right temporal lobe and right lenticular nucleus | 15
conservative management | 15
total of 10 weeks of i.v. metronidazole therapy | 15
neurological symptoms improved | 16
full recovery of language | 16
slight paresis in the right arm | 16
end-of-treatment CT scans showed residual liver and brain abscesses | 16
co-infection of liver abscesses by Staphylococcus epidermidis | 16
Clostridium difficile pseudomembranous colitis | 16
discharged after a 16-week stay in the surgical ICU | 16
stable and rehabilitating | 16
malnutrition | -672
alcohol abuse | -672
smoking | -672
pulmonary tuberculosis | -672
treated and cured | -672
amebiasis | -672 
Entamoeba histolytica infection | -672 
invasive amebiasis | 0 
intestinal amebiasis | 0 
extraintestinal amebiasis | 0 
liver abscess | 0 
peritoneal abscess | 6 
lung abscess | 6 
brain abscess | 15 
cutaneous amebiasis | 10 
amebic colitis | 5 
septic shock | 1 
respiratory failure | 6 
neurological symptoms | 15 
aphasia | 15 
right-sided hemiplegia | 15 
paresis in the right arm | 16 
disseminated intraabdominal abscesses | 6 
bilateral pleural effusion | 6 
amebic pleural effusions | 6 
Staphylococcus epidermidis co-infection | 16 
Clostridium difficile pseudomembranous colitis | 16 
HIV negative | 10 
Acanthamoeba spp negative | 10 
Balamuthia mandrillaris negative | 10 
Naegleria fowleri negative | 10 
RT-PCR positive for E. histolytica | 5 
microscopy positive for E. histolytica trophozoites | 5 
antigen detection in stool | 5 
serology | 10 
molecular analysis by RT-PCR | 5 
amebicidal tissue-active agent | 5 
luminal cysticidal agent | 5 
metronidazole | 5 
paromomycin | 5 
diloxanide | 5 
tinidazole | 5 
surgical drainage | 2 
antimicrobial treatment | 5 
conservative management | 15 
neurosurgery consultation | 15 
cranial CT scan | 15 
thoracoabdominal CT scan | 6 
abdominal CT scan | 0 
liver aspirate | 2 
blood samples | 10 
skin biopsy | 10 
bronchial aspirate | 10 
pleural drainage | 10 
stool samples | 5 
RT-PCR of liver aspirate | 5 
RT-PCR of stool | 5 
RT-PCR of pleural fluid | 10 
RT-PCR of blood | 10 
RT-PCR of skin biopsy | 10 
QIAamp DNA Mini Kit | 5 
real-time PCR (RT-PCT) | 5 
SSU rRNA gene | 5 
Gal/GalNAc lectin antigens | 5 
EhMIF (proinflammatory cytokine macrophage migration inhibitory factor) | 5 
interferon gamma (IFN-γ) | 5 
genetic susceptibility | 5 
immune status | 5 
young age | 5 
pregnancy | 5 
corticosteroid therapy | 5 
malnutrition | 5 
alcohol abuse | 5 
smoking | 5 
pulmonary tuberculosis | 5 
treated and cured | 5 
amebiasis diagnosis | 5 
differential diagnosis | 5 
pyogenic liver abscess | 5 
hepatoma | 5 
echinococcal cyst | 5 
liver abscess rupture | 6 
peritoneal involvement | 6 
pleural involvement | 6 
hematogenous spread | 6 
brain abscess formation | 15 
cerebral amebiasis | 15 
neurosurgical consultation | 15 
conservative management | 15 
antimicrobial treatment | 15 
metronidazole therapy | 15 
tinidazole therapy | 15 
diloxanide therapy | 15 
paromomycin therapy | 15 
luminal agent therapy | 15 
amebicidal tissue-active agent therapy | 15 
cysticidal agent therapy | 15 
surgical drainage | 2 
percutaneous CT-guide drainage | 2 
liver abscess drainage | 2 
brain abscess drainage | 15 
neurosurgery | 15 
craniotomy | 15 
antimicrobial therapy | 5 
antiparasitic therapy | 5 
supportive care | 5 
intensive care unit (ICU) | 1 
mechanical ventilation | 1 
vasopressor support | 1 
septic shock management | 1 
respiratory failure management | 6 
neurological symptoms management | 15 
aphasia management | 15 
right-sided hemiplegia management | 15 
paresis in the right arm management | 16 
disseminated intraabdominal abscesses management | 6 
bilateral pleural effusion management | 6 
amebic pleural effusions management | 6 
Staphylococcus epidermidis co-infection management | 16 
Clostridium difficile pseudomembranous colitis management | 16 
HIV management | 10 
Acanthamoeba spp management | 10 
Balamuthia mandrillaris management | 10 
Naegleria fowleri management | 10 
RT-PCR positive for E. histolytica management | 5 
microscopy positive for E. histolytica trophozoites management | 5 
antigen detection in stool management | 5 
serology management | 10 
molecular analysis by RT-PCR management | 5 
amebicidal tissue-active agent management | 5 
luminal cysticidal agent management | 5 
metronidazole management | 5 
paromomycin management | 5 
diloxanide management | 5 
tinidazole management | 5 
surgical drainage management | 2 
antimicrobial treatment management | 5 
conservative management management | 15 
neurosurgery consultation management | 15 
cranial CT scan management | 15 
thoracoabdominal CT scan management | 6 
abdominal CT scan management | 0 
liver aspirate management | 2 
blood samples management | 10 
skin biopsy management | 10 
bronchial aspirate management | 10 
pleural drainage management | 10 
stool samples management | 5 
RT-PCR of liver aspirate management | 5 
RT-PCR of stool management | 5 
RT-PCR of pleural fluid management | 10 
RT-PCR of blood management | 10 
RT-PCR of skin biopsy management | 10 
QIAamp DNA Mini Kit management | 5 
real-time PCR (RT-PCT) management | 5 
SSU rRNA gene management | 5 
Gal/GalNAc lectin antigens management | 5 
EhMIF (proinflammatory cytokine macrophage migration inhibitory factor) management | 5 
interferon gamma (IFN-γ) management | 5 
genetic susceptibility management | 5 
immune status management | 5 
young age management | 5 
pregnancy management | 5 
corticosteroid therapy management | 5 
malnutrition management | 5 
alcohol abuse management | 5 
smoking management | 5 
pulmonary tuberculosis management | 5 
treated and cured management | 5 
amebiasis diagnosis management | 5 
differential diagnosis management | 5 
pyogenic liver abscess management | 5 
hepatoma management | 5 
echinococcal cyst management | 5 
liver abscess rupture management | 6 
peritoneal involvement management | 6 
pleural involvement management | 6 
hematogenous spread management | 6 
brain abscess formation management | 15 
cerebral amebiasis management | 15 
neurosurgical consultation management | 15 
conservative management management | 15 
antimicrobial treatment management | 15 
metronidazole therapy management | 15 
tinidazole therapy management | 15 
diloxanide therapy management | 15 
paromomycin therapy management | 15 
luminal agent therapy management | 15 
amebicidal tissue-active agent therapy management | 15 
cysticidal agent therapy management | 15 
surgical drainage management | 2 
percutaneous CT-guide drainage management | 2 
liver abscess drainage management | 2 
brain abscess drainage management | 15 
neurosurgery management | 15 
craniotomy management | 15 
antimicrobial therapy management | 5 
antiparasitic therapy management | 5 
supportive care management | 5 
intensive care unit (ICU) management | 1 
mechanical ventilation management | 1 
vasopressor support management | 1 
septic shock management management | 1 
respiratory failure management management | 6 
neurological symptoms management management | 15 
aphasia management management | 15 
right-sided hemiplegia management management | 15 
paresis in the right arm management management | 16 
disseminated intraabdominal abscesses management management | 6 
bilateral pleural effusion management management | 6 
amebic pleural effusions management management | 6 
Staphylococcus epidermidis co-infection management management | 16 
Clostridium difficile pseudomembranous colitis management management | 16 
HIV management management | 10 
Acanthamoeba spp management management | 10 
Balamuthia mandrillaris management management | 10 
Naegleria fowleri management management | 10 
RT-PCR positive for E. histolytica management management | 5 
microscopy positive for E. histolytica trophozoites management management | 5 
antigen detection in stool management management | 5 
serology management management | 10 
molecular analysis by RT-PCR management management | 5 
amebicidal tissue-active agent management management | 5 
luminal cysticidal agent management management | 5 
metronidazole management management | 5 
paromomycin management management | 5 
diloxanide management management | 5 
tinidazole management management | 5 
surgical drainage management management | 2 
antimicrobial treatment management management | 5 
conservative management management management | 15 
neurosurgery consultation management management | 15 
cranial CT scan management management | 15 
thoracoabdominal CT scan management management | 6 
abdominal CT scan management management | 0 
liver aspirate management management | 2 
blood samples management management | 10 
skin biopsy management management | 10 
bronchial aspirate management management | 10 
pleural drainage management management | 10 
stool samples management management | 5 
RT-PCR of liver aspirate management management | 5 
RT-PCR of stool management management | 5 
RT-PCR of pleural fluid management management | 10 
RT-PCR of blood management management | 10 
RT-PCR of skin biopsy management management | 10 
QIAamp DNA Mini Kit management management | 5 
real-time PCR (RT-PCT) management management | 5 
SSU rRNA gene management management | 5 
Gal/GalNAc lectin antigens management management | 5 
EhMIF (proinflammatory cytokine macrophage migration inhibitory factor) management management | 5 
interferon gamma (IFN-γ) management management | 5 
genetic susceptibility management management | 5 
immune status management management | 5 
young age management management | 5 
pregnancy management management | 5 
corticosteroid therapy management management | 5 
malnutrition management management | 5 
alcohol abuse management management | 5 
smoking management management | 5 
pulmonary tuberculosis management management | 5 
treated and cured management management | 5 
amebiasis diagnosis management management | 5 
differential diagnosis management management | 5 
pyogenic liver abscess management management | 5 
hepatoma management management | 5 
echinococcal cyst management management | 5 
liver abscess rupture management management | 6 
peritoneal involvement management management | 6 
pleural involvement management management | 6 
hematogenous spread management management | 6 
brain abscess formation management management | 15 
cerebral amebiasis management management | 15 
neurosurgical consultation management management | 15 
conservative management management management | 15 
antimicrobial treatment management management | 15 
metronidazole therapy management management | 15 
tinidazole therapy management management | 15 
diloxanide therapy management management | 15 
paromomycin therapy management management | 15 
luminal agent therapy management management | 15 
amebicidal tissue-active agent therapy management management | 15 
cysticidal agent therapy management management | 15 
surgical drainage management management | 2 
percutaneous CT-guide drainage management management | 2 
liver abscess drainage management management | 2 
brain abscess drainage management management | 15 
neurosurgery management management | 15 
craniotomy management management | 15 
antimicrobial therapy management management | 5 
antiparasitic therapy management management | 5 
supportive care management management | 5 
intensive care unit (ICU) management management | 1 
mechanical ventilation management management | 1 
vasopressor support management management | 1 
septic shock management management management | 1 
respiratory failure management management management | 6 
neurological symptoms management management management | 15 
aphasia management management management | 15 
right-sided hemiplegia management management management | 15 
paresis in the right arm management management management | 16 
disseminated intraabdominal abscesses management management management | 6 
bilateral pleural effusion management management management | 6 
amebic pleural effusions management management management | 6 
Staphylococcus epidermidis co-infection management management management | 16 
Clostridium difficile pseudomembranous colitis management management management | 16 
HIV management management management | 10 
Acanthamoeba spp management management management | 10 
Balamuthia mandrillaris management management management | 10 
Naegleria fowleri management management management | 10 
RT-PCR positive for E. histolytica management management management | 5 
microscopy positive for E. histolytica trophozoites management management management | 5 
antigen detection in stool management management management | 5 
serology management management management | 10 
molecular analysis by RT-PCR management management management | 5 
amebicidal tissue-active agent management management management | 5 
luminal cysticidal agent management management management | 5 
metronidazole management management management | 5 
paromomycin management management management | 5 
diloxanide management management management | 5 
tinidazole management management management | 5 
surgical drainage management management management | 2 
antimicrobial treatment management management management | 5 
conservative management management management management | 15 
neurosurgery consultation management management management | 15 
cranial CT scan management management management | 15 
thoracoabdominal CT scan management management management | 6 
abdominal CT scan management management management | 0 
liver aspirate management management management | 2 
blood samples management management management | 10 
skin biopsy management management management | 10 
bronchial aspirate management management management | 10 
pleural drainage management management management | 10 
stool samples management management management | 5 
RT-PCR of liver aspirate management management management | 5 
RT-PCR of stool management management management | 5 
RT-PCR of pleural fluid management management management | 10 
RT-PCR of blood management management management | 10 
RT-PCR of skin biopsy management management management | 10 
QIAamp DNA Mini Kit management management management | 5 
real-time PCR (RT-PCT) management management management | 5 
SSU rRNA gene management management management | 5 
Gal/GalNAc lectin antigens management management management | 5 
EhMIF (proinflammatory cytokine macrophage migration inhibitory factor) management management management | 5 
interferon gamma (IFN-γ) management management management | 5 
genetic susceptibility management management management | 5 
immune status management management management | 5 
young age management management management | 5 
pregnancy management management management | 5 
corticosteroid therapy management management management | 5 
malnutrition management management management | 5 
alcohol abuse management management management | 5 
smoking management management management | 5 
pulmonary tuberculosis management management management | 5 
treated and cured management management management | 5 
amebiasis diagnosis management management management | 5 
differential diagnosis management management management | 5 
pyogenic liver abscess management management management | 5 
hepatoma management management management | 5 
echinococcal cyst management management management | 5 
liver abscess rupture management management management | 6 
peritoneal involvement management management management | 6 
pleural involvement management management management | 6 
hematogenous spread management management management | 6 
brain abscess formation management management management | 15 
cerebral amebiasis management management management | 15 
neurosurgical consultation management management management | 15 
conservative management management management management | 15 
antimicrobial treatment management management management | 15 
metronidazole therapy management management management | 15 
tinidazole therapy management management management | 15 
diloxanide therapy management management management | 15 
paromomycin therapy management management management | 15 
luminal agent therapy management management management | 15 
amebicidal tissue-active agent therapy management management management | 15 
cysticidal agent therapy management management management | 15 
surgical drainage management management management | 2 
percutaneous CT-guide drainage management management management | 2 
liver abscess drainage management management management | 2 
brain abscess drainage management management management | 15 
neurosurgery management management management | 15 
craniotomy management management management | 15 
antimicrobial therapy management management management | 5 
antiparasitic therapy management management management | 5 
supportive care management management management | 5 
intensive care unit (ICU) management management management | 1 
mechanical ventilation management management management | 1 
vasopressor support management management management | 1 
septic shock management management management management | 1 
respiratory failure management management management management | 6 
neurological symptoms management management management management | 15 
aphasia management management management management | 15 
right-sided hemiplegia management management management management | 15 
paresis in the right arm management management management management | 16 
disseminated intraabdominal abscesses management management management management | 6 
bilateral pleural effusion management management management management | 6 
amebic pleural effusions management management management management | 6 
Staphylococcus epidermidis co-infection management management management management | 16 
Clostridium difficile pseudomembranous colitis management management management management | 16 
HIV management management management management | 10 
Acanthamoeba spp management management management management | 10 
Balamuthia mandrillaris management management management management | 10 
Naegleria fowleri management management management management | 10 
RT-PCR positive for E. histolytica management management management management | 5 
microscopy positive for E. histolytica trophozoites management management management management | 5 
antigen detection in stool management management management management | 5 
serology management management management management | 10 
molecular analysis by RT-PCR management management management management | 5 
amebicidal tissue-active agent management management management management | 5 
luminal cysticidal agent management management management management | 5 
metronidazole management management management management | 5 
paromomycin management management management management | 5 
diloxanide management management management management | 5 
tinidazole management management management management | 5 
surgical drainage management management management management | 2 
antimicrobial treatment management management management management | 5 
conservative management management management management management | 15 
neurosurgery consultation management management management management | 15 
cranial CT scan management management management management | 15 
thoracoabdominal CT scan management management management management | 6 
abdominal CT scan management management management management | 0 
liver aspirate management management management management | 2 
blood samples management management management management | 10 
skin biopsy management management management management | 10 
bronchial aspirate management management management management | 10 
pleural drainage management management management management | 10 
stool samples management management management management | 5 
RT-PCR of liver aspirate management management management management | 5 
RT-PCR of stool management management management management | 5 
RT-PCR of pleural fluid management management management management | 10 
RT-PCR of blood management management management management | 10 
RT-PCR of skin biopsy management management management management | 10 
QIAamp DNA Mini Kit management management management management | 5 
real-time PCR (RT-PCT) management management management management | 5 
SSU rRNA gene management management management management | 5 
Gal/GalNAc lectin antigens management management management management | 5 
EhMIF (proinflammatory cytokine macrophage migration inhibitory factor) management management management management | 5 
interferon gamma (IFN-γ) management management management management | 5 
genetic susceptibility management management management management | 5 
immune status management management management management | 5 
young age management management management management | 5 
pregnancy management management management management | 5 
corticosteroid therapy management management management management | 5 
malnutrition management management management management | 5 
alcohol abuse management management management management | 5 
smoking management management management management | 5 
pulmonary tuberculosis management management management management | 5 
treated and cured management management management management | 5 
amebiasis diagnosis management management management management | 5 
differential diagnosis management management management management | 5 
pyogenic liver abscess management management management management | 5 
hepatoma management management management management | 5 
echinococcal cyst management management management management | 5 
liver abscess rupture management management management management | 6 
peritoneal involvement management management management management | 6 
pleural involvement management management management management | 6 
hematogenous spread management management management management | 6 
brain abscess formation management management management management | 15 
cerebral amebiasis management management management management | 15 
neurosurgical consultation management management management management | 15 
conservative management management management management management | 15 
antimicrobial treatment management management management management | 15 
metronidazole therapy management management management management | 15 
tinidazole therapy management management management management | 15 
diloxanide therapy management management management management | 15 
paromomycin therapy management management management management | 15 
luminal agent therapy management management management management | 15 
amebicidal tissue-active agent therapy management management management management | 15 
cysticidal agent therapy management management management management | 15 
surgical drainage management management management management | 2 
percutaneous CT-guide drainage management management management management | 2 
liver abscess drainage management management management management | 2 
brain abscess drainage management management management management | 15 
neurosurgery management management management management | 15 
craniotomy management management management management | 15 
antimicrobial therapy management management management management | 5 
antiparasitic therapy management management management management | 5 
supportive care management management management management | 5 
intensive care unit (ICU) management management management management | 1 
mechanical ventilation management management management management | 1 
vasopressor support management management management management | 1 
septic shock management management management management management | 1 
respiratory failure management management management management management | 6 
neurological symptoms management management management management management | 15 
aphasia management management management management management | 15 
right-sided hemiplegia management management management management management | 15 
paresis in the right arm management management management management management | 16 
disseminated intraabdominal abscesses management management management management management | 6 
bilateral pleural effusion management management management management management | 6 
amebic pleural effusions management management management management management | 6 
Staphylococcus epidermidis co-infection management management management management management | 16 
Clostridium difficile pseudomembranous colitis management management management management management | 16 
HIV management management management management management | 10 
Acanthamoeba spp management management management management management | 10 
Balamuthia mandrillaris management management management management management | 10 
Naegleria fowleri management management management management management | 10 
RT-PCR positive for E. histolytica management management management management management | 5 
microscopy positive for E. histolytica trophozoites management management management management management | 5 
antigen detection in stool management management management management management | 5 
serology management management management management management | 10 
molecular analysis by RT-PCR management management management management management | 5 
amebicidal tissue-active agent management management management management management | 5 
luminal cysticidal agent management management management management management | 5 
metronidazole management management management management management | 5 
paromomycin management management management management management | 5 
diloxanide management management management management management | 5 
tinidazole management management management management management | 5 
surgical drainage management management management management management | 2 
antimicrobial treatment management management management management management | 5 
conservative management management management management management management | 15 
neurosurgery consultation management management management management management | 15 
cranial CT scan management management management management management | 15 
thoracoabdominal CT scan management management management management management | 6 
abdominal CT scan management management management management management | 0 
liver aspirate management management management management management | 2 
blood samples management management management management management | 10 
skin biopsy management management management management management | 10 
bronchial aspirate management management management management management | 10 
pleural drainage management management management management management | 10 
stool samples management management management management management | 5 
RT-PCR of liver aspirate management management management management management | 5 
RT-PCR of stool management management management management management | 5 
RT-PCR of pleural fluid management management management management management | 10 
RT-PCR of blood management management management management management | 10 
RT-PCR of skin biopsy management management management management management | 10 
QIAamp DNA Mini Kit management management management management management | 5 
real-time PCR (RT-PCT) management management management management management | 5 
SSU rRNA gene management management management management management | 5 
Gal/GalNAc lectin antigens management management management management management | 5 
EhMIF (proinflammatory cytokine macrophage migration inhibitory factor) management management management management management | 5 
interferon gamma (IFN-γ) management management management management management | 5 
genetic susceptibility management management management management management | 5 
immune status management management management management management | 5 
young age management management management management management | 5 
pregnancy management management management management management | 5 
corticosteroid therapy management management management management management | 5 
malnutrition management management management management management | 5 
alcohol abuse management management management management management | 5 
smoking management management management management management | 5 
pulmonary tuberculosis management management management management management | 5 
treated and cured management management management management management | 5 
amebiasis diagnosis management management management management management | 5 
differential diagnosis management management management management management | 5 
pyogenic liver abscess management management management management management | 5 
hepatoma management management management management management | 5 
echinococcal cyst management management management management management | 5 
liver abscess rupture management management management management management | 6 
peritoneal involvement management management management management management | 6 
pleural involvement management management management management management | 6 
hematogenous spread management management management management management | 6 
brain abscess formation management management management management management | 15 
cerebral amebiasis management management management management management | 15 
neurosurgical consultation management management management management management | 15 
conservative management management management management management management | 15 
antimicrobial treatment management management management management management | 15 
metronidazole therapy management management management management management | 15 
tinidazole therapy management management management management management | 15 
diloxanide therapy management management management management management | 15 
paromomycin therapy management management management management management | 15 
luminal agent therapy management management management management management | 15 
amebicidal tissue-active agent therapy management management management management management | 15 
cysticidal agent therapy management management management management management | 15 
surgical drainage management management management management management | 2 
percutaneous CT-guide drainage management management management management management | 2 
liver abscess drainage management management management management management | 2 
brain abscess drainage management management management management management | 15 
neurosurgery management management management management management | 15 
craniotomy management management management management management | 15 
antimicrobial therapy management management management management management | 5 
antiparasitic therapy management management management management management | 5 
supportive care management management management management management | 5 
intensive care unit (ICU) management management management management management | 1 
mechanical ventilation management management management management management | 1 
vasopressor support management management management management management | 1 
septic shock management management management management management management | 1 
respiratory failure management management management management management management | 6 
neurological symptoms management management management management management management | 15 
aphasia management management management management management management | 15 
right-sided hemiplegia management management management management management management | 15 
paresis in the right arm management management management management management management | 16 
disseminated intraabdominal abscesses management management management management management management | 6 
bilateral pleural effusion management management management management management management | 6 
amebic pleural effusions management management management management management management | 6 
Staphylococcus epidermidis co-infection management management management management management management | 16 
Clostridium difficile pseudomembranous colitis management management management management management management | 16 
HIV management management management management management management | 10 
Acanthamoeba spp management management management management management management | 10 
Balamuthia mandrillaris management management management management management management | 10 
Naegleria fowleri management management management management management management | 10 
RT-PCR positive for E. histolytica management management management management management management | 5 
microscopy positive for E. histolytica trophozoites management management management management management management | 5 
antigen detection in stool management management management management management management | 5 
serology management management management management management management | 10 
molecular analysis by RT-PCR management management management management management management | 5 
amebicidal tissue-active agent management management management management management management | 5 
luminal cysticidal agent management management management management management management | 5 
metronidazole management management management management management management | 5 
paromomycin management management management management management management | 5 
diloxanide management management management management management management | 5 
tinidazole management management management management management management | 5 
surgical drainage management management management management management management | 2 
antimicrobial treatment management management management management management management | 5 
conservative management management management management management management management | 15 
neurosurgery consultation management management management management management management | 15 
cranial CT scan management management management management management management | 15 
thoracoabdominal CT scan management management management management management management | 6 
abdominal CT scan management management management management management management | 0 
liver aspirate management management management management management management | 2 
blood samples management management management management management management | 10 
skin biopsy management management management management management management | 10 
bronchial aspirate management management management management management management | 10 
pleural drainage management management management management management management | 10 
stool samples management management management management management management | 5 
RT-PCR of liver aspirate management management management management management management | 5 
RT-PCR of stool management management management management management management | 5 
RT-PCR of pleural fluid management management management management management management | 10 
RT-PCR of blood management management management management management management | 10 
RT-PCR of skin biopsy management management management management management management | 10 
QIAamp DNA Mini Kit management management management management management management | 5 
real-time PCR (RT-PCT) management management management management management management | 5 
SSU rRNA gene management management management management management management | 5 
Gal/GalNAc lectin antigens management management management management management management | 5 
EhMIF (proinflammatory cytokine macrophage migration inhibitory factor) management management management management management management | 5 
interferon gamma (IFN-γ) management management management management management management | 5 
genetic susceptibility management management management management management management | 5 
immune status management management management management management management | 5 
young age management management management management management management | 5 
