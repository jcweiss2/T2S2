34 years old | 0
female | 0
Japanese | 0
cough | -72
fever | -72
husband and son ill with COVID-19 | -72
nasopharyngeal swab for COVID-19 positive | -72
admitted to hospital for COVID-19 infection | 0
bilateral and peripheral ground-glass opacity | 0
moderate COVID-19 pneumonia | 0
intravenous remdesivir | 0
oral dexamethasone | 0
discharged from hospital | 240
chest pain | 240
ECG showed ST elevation | 240
inferior-wall acute myocardial infarction | 240
emergency coronary angiography | 240
embolic occlusion in left circumflex branch | 240
anticoagulation with heparin sodium | 240
right renal infarction | 240
acute multi-territory ischemic stroke | 240
fever | 240
blood culture positive for Gram-positive coccus | 240
tranthoracic echocardiography | 240
11-mm vegetation on posterior mitral valve leaflet | 240
native mitral valve IE | 240
intravenous vancomycin | 240
cefazolin | 240
transferred to university hospital | 240
clear consciousness level | 240
no apparent neurological deficit | 240
blood pressure 74/48 mmHg | 240
pulse 69 beats/minute | 240
body temperature 39.1℃ | 240
conjunctiva petechiae | 240
hemorrhagic spots on soft palate | 240
grade II/VI pansystolic murmur | 240
white blood cell count 20.9 K/μL | 240
C-reactive protein 10.12 mg/dL | 240
Troponin T 0.627 ng/mL | 240
NT-proBNP 4,041 pg/mL | 240
lactate 2.9 mmol/L | 240
chest X-ray showed no enlargement of cardiac silhouette | 240
sinus rhythm with heart rate of 70/min | 240
large and mobile vegetations on mitral posterior leaflet | 240
severe mitral regurgitation | 240
causative organism methicillin-susceptible Staphylococcus aureus | 240
optimal antimicrobial therapy | 240
surgical mitral valve replacement | 336
postoperative course uneventful | 336
discharged without complication | 600