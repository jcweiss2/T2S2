79 years old | 0
lady | 0
occipital headache | -48
nausea | -48
vomiting | -48
previous herpes zoster infection | -6720
hypertension | -6720
hyperlipidemia | -6720
labyrinthitis | -6720
Ramsay Hunt syndrome | -6720
hysterectomy | -6720
tonsillectomy | -6720
breast operation | -6720
cataract operation | -6720
ramipril | 0
bisoprolol | 0
atorvastatin | 0
clopidogrel | 0
aspirin | 0
zolpidem | 0
alfacalcidol | 0
calcium | 0
hyponatremia | 0
increased GGT | 0
bilirubin | 0
normal urinalysis | 0
normal CT brain | 0
mild pulmonary vascular congestion | 0
no chest pain | 0
no abdominal pain | 0
encephalitis | 0
antibiotics | 0
lumbar puncture | 96
herpes simplex virus 1 infection | 96
acyclovir | 96
nonspecific abdominal pain | 288
cholelithiasis | 288
conservative treatment | 288
pain localized to the right iliac fossa | 312
CT abdomen pelvis | 312
ischemia | 312
pneumatosis | 312
laparotomy | 432
bowel ischemia | 432
retrocaecal perforation | 432
terminal ileal band | 432
internal herniation | 432
gangrene | 432
extended right hemicolectomy | 432
Bogota bag | 432
re-look surgery | 456
no progression of ischemia | 456
ileostomy | 456
closure of abdomen | 456