57-year-old woman | 0  
    diabetes | 0  
    metformin | 0  
    vitamin D deficiency | 0  
    diagnosed with Ph+ CML in AP | -24  
    hepatosplenomegaly | -24  
    spleen 25 cm | -24  
    liver 22 cm | -24  
    imatinib | -24  
    hematological remission | -24  
    clinical resistance to imatinib | -24  
    imatinib dose increased to 600 mg/day | -24  
    pallor | -24  
    hepatosplenomegaly | -24  
    hemoglobin 7 g/dL | -24  
    platelet count 194,000/μL | -24  
    WBC count 26,000/μL | -24  
    0% basophils | -24  
    1% eosinophils | -24  
    10% blasts | -24  
    hypercellular BM (90% cellularity) | -24  
    11% blasts | -24  
    CD45 positive | -24  
    CD34 positive | -24  
    CD33 positive | -24  
    CD117 positive | -24  
    CD56 negative | -24  
    karyotype 47,XX,+7,t(9,22)(q34,q11.2) | -24  
    FISH BCR/ABL fusion signals 5% | -24  
    switched to dasatinib 100 mg/day | 0  
    minimal interruption of treatment | 0  
    GCSF | 0  
    blood product transfusions | 0  
    progressive shortness of breath | 168  
    lung infiltrates | 168  
    abdominal pain | 168  
    CT scan abdomen and pelvis | 168  
    mild hepatosplenomegaly | 168  
    portal venous hypertension | 168  
    small hypo-attenuated splenic lesion | 168  
    no lymphadenopathy | 168  
    bowels unremarkable | 168  
    complete cytogenetic remission | 432  
    Philadelphia chromosome disappearance | 432  
    trisomy 7 disappearance | 432  
    FISH negative | 432  
    BCRABL p210 not detectable | 432  
    JAK-2 V617F mutation negative | 432  
    severe headache | 432  
    nausea | 432  
    generalized tonic-clonic seizures | 432  
    brain MRI abnormal signal intensity | 432  
    contrast signal enhancement | 432  
    leptomeningeal infiltration | 432  
    CSF WBCs 130/μL | 432  
    51% blasts | 432  
    43% myeloblasts positive CD34, CD117, CD33 | 432  
    negative HLA-DR | 432  
    negative CD3 | 432  
    negative CD13 | 432  
    dasatinib | 432  
    TIT chemotherapy | 432  
    methotrexate 15 mg | 432  
    cytarabine 50 mg | 432  
    hydrocortisone 50 mg | 432  
    CSF clear after 5 rounds | 432  
    refused further TIT chemotherapy | 432  
    refused allo-SCT | 432  
    severe headache | 1680  
    second CNS relapse | 1680  
    brain MRI interval improvement | 1680  
    leukemic leptomeningeal infiltration resolution | 1680  
    new T2 hyperintensity | 1680  
    CSF blasts 52% | 1680  
    CD34 positive | 1680  
    CD117 positive | 1680  
    CD33 positive | 1680  
    CD13 positive | 1680  
    CD7 positive | 1680  
    whole-brain radiation therapy 30 Gy | 1680  
    dasatinib 100 mg/day | 1680  
    hepatosplenomegaly fluctuating | 1680  
    spleen size 18 cm | 1680  
    BM cellularity 50% | 1680  
    trilineage hematopoiesis | 1680  
    <1% blasts | 1680  
    cytogenetic analysis normal 46,XX | 1680  
    hypothyroidism | 2280  
    levothyroxine | 2280  
    minimal pleural effusion | 2280  
    diuretics | 2280  
    GCSF support | 2280  
    neutrophil count maintained | 2280  
    dasatinib decreased to 70 mg/day | 2280  
    dasatinib increased to 100 mg/day | 2832  
    dasatinib halted | 2832  
    diarrhea | 2832  
    edema | 2832  
    BCR-ABL transcripts undetectable | 2832  
    pegylated interferon%2a | 2832  
    doses 45-135 μg | 2832  
    hepatosplenomegaly resolved | 2832  
    unable to tolerate PegINF%2a | 2832  
    PegINF%2a discontinued | 2832  
    spleen growth | 2832  
    autoimmune disorder | 2832  
    joint pains | 2832  
    minimal left-sided pleural effusion | 2832  
    chronic diarrhea | 2832  
    lupus anticoagulant positive | 2832  
    ANA positive | 2832  
    anticardiolipin IgG positive | 2832  
    anticardiolipin IgM positive | 2832  
    B2GP1 positive | 2832  
    anti-dsDNA antibodies positive | 2832  
    refused prophylactic anticoagulation | 2832  
    referred to rheumatology | 2832  
    spleen size 17.1 cm | 2832  
    CML therapy on hold | 2832  
    deep molecular remission | 2832  
    BCR-ABL transcripts undetectable | 2832  
    bloody diarrhea | 2832  
    adenocarcinoma of rectum | 2832  
    invasion of uterus | 2832  
    septic shock | 2832  
    admitted to ICU | 2832  
    CT abdomen and pelvis | 2832  
    splenic infarct | 2832  
    moderate to massive ascites | 2832  
    omental thickening | 2832  
    peritoneal deposits | 2832  
    adnexal mass left 7.7x6 cm | 2832  
    adnexal mass right 6x6.7 cm | 2832  
    rectal mass infiltrated anal canal | 2832  
    nodules | 2832  
    inguinal lymph nodes increased | 2832  
    non-occlusive thrombosis left external iliac vein | 2832  
    common femoral vein thrombosis | 2832  
    bilateral pleural effusions | 2832  
    basilar atelectasis | 2832  
    traction bronchiectasis | 2832  
    pulmonary embolism | 2832  
    bilateral pulmonary nodules | 2832  
    unfit for chemotherapy | 2832  
    palliative supportive care | 2832  
    died | 2832  
    septic shock | 2832  
    cancer-related venous thromboembolism | 2832  
    possible autoimmune disorder | 2832  
    progressive adenocarcinoma of rectum | 2832  
    supportive therapy | 2832  
    treatment-free remission 18 months | 2832  
    