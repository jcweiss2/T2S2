48 years old | 0
female | 0
end-stage renal disease | -10080
hypertensive | -10080
maintenance hemodialysis | -432
elective robotic assisted laparoscopic renal transplantation | 0
living related donor | 0
preoperative hemodialysis | -24
standard monitoring | 0
balanced general anesthesia | 0
heart rate 94/min | 0
mean arterial pressure 103 mm of Hg | 0
SpO2 100% | 0
central venous pressure 12 cm of H2O | 0
core temperature 98.6°F | 0
arterial blood gas analysis | 0
lactate 1.9 mM/L | 0
volume controlled ventilation | 0
EtCO2 between 35 mm and 40 mm of Hg | 0
hemodynamic parameters deteriorated | 180
heart rate 122/min | 180
mean arterial pressure 72 mm of Hg | 180
central venous pressure 16 cm of H2O | 180
metabolic acidosis | 180
elevated lactate levels | 180
hyperglycemia | 180
elevated anion gap | 180
fall in hemoglobin | 180
blood sample for ketone bodies tested negative | 180
IV fluids | 180
packed red blood cells transfused | 180
noradrenaline infusion | 180
sodium bicarbonate infusion | 180
insulin infusion | 180
vascular anastomosis of the graft kidney | 180
allograft reperfused | 205
urine output established | 205
shifted to Intensive Care Unit | 420
elective ventilation | 420
continuous renal replacement therapy | 420
ABG analysis in ICU | 420
progressively increasing lactic acidosis | 420
hyperglycemia refractory to bicarbonate and insulin infusion | 420
average urine output 300 mL/h | 420
procalcitonin levels obtained | 420
procalcitonin level 14.6 ng/mL | 420
thiamine deficiency suspected | 420
empirical thiamine 300 mg administered intravenously | 420
ABG analysis after thiamine administration | 540
lactate and sugar levels decreased | 540
improvement in MAP | 540
bicarbonate infusion stopped | 540
insulin infusion stopped | 540
noradrenaline infusion stopped | 540
extubated | 630
thiamine injection 300 mg IV repeated | 630
ABG analysis after second thiamine injection | 720
lactic acidosis resolved | 720
shifted to posttransplant isolation ward | 840