57 years old | 0
male | 0
wine-grower | 0
heavy consumption of alcohol | 0
admitted to the hospital | 0
low back pain | -240
lumbar torsion | -240
loss of balance | -240
rough ground | -240
persistent and progressive lumbar pain | -240
slight fever | -72
dental pain | -240
untreated dental pain | -240
teeth 27 and 28 | -240
paravertebral painful muscular contracture | 0
lumbar spine | 0
no neurological deficit | 0
normal reflexes | 0
normal and symmetrical reflexes | 0
Lasègue and Bragard manoeuvres were negative | 0
systemic inflammatory syndrome | 0
erythrocyte sedimentation rate of 60 mm/hour | 0
C-reactive protein of 111 mg/L | 0
white cell count of 23 G/L | 0
91% of segmented neutrophils | 0
blood cultures were collected | 0
lumbar radiographs | 0
degenerative signs | 0
lumbar MRI | 0
epidural abscess | 0
posteriorly of the thecal sac | 0
L3-L4 and L4-L5 levels | 0
anteriorly at the L5-S1 level | 0
L5-S1 discopathy | 0
suspected psoas abscess | 0
emergency surgery | 0
posterior approach | 0
decompressive laminectomy | 0
right cross-over shape | 0
L3 to S1 | 0
no stabilisation | 0
two distinct collections | 0
microbiological studies | 0
thecal sac looked free of compression | 0
intravenous amoxicillin-clavulanic acid | 0
abscess cultures | 24
multisensitive Streptococcus mitis/oralis | 24
blood cultures were positive | 24
same pathogen | 24
became negative after 48 hours | 72
antibiotic treatment | 0
transoral echocardiography | 24
no evidence for endocarditis | 24
BARD 5f picc-line | 24
left basilic vein | 24
continuous intravenous antibiotic treatment | 24
empiric antibiotic treatment | 0
penicillin-G | 48
5M of units | 48
four times per day | 48
10 days | 48
minimum inhibitory concentration | 48
0.125 mg/L | 48
lumbar pain decreased | 24
no fever | 24
CRP decreased | 72
WCC became normal | 96
discharged from the hospital | 264
surgical wound healing well | 264
antibiotic treatment changed | 264
intravenous ceftriaxone | 264
2 g daily | 264
remaining 4 weeks | 264
infected teeth treated | 264
surgical avulsion | 264
teeth 27 and 28 | 264
asymptomatic | 432
CRP was 6 mg/L | 432
satisfactory wound healing | 432
lumbar MRI | 432
same collapse of the L5-S1 | 432
no sign of persistent or recurrent infection | 432
1-year follow-up | 876
no sign of persistent or recurrent abscess | 876
no evidence of spondylolisthesis | 876
peripheral inflammatory pannus resolved | 876