37 years old|0
man|0
no significant previous medical history|0
presented to the emergency department|0
fever|-96
vomiting|-24
loose stools|-24
abdominal cramps|-24
headache|-24
intermittent fever|-96
low grade fever|-96
generalized headache|-24
nonbilious vomiting|-24
tachycardia|0
mild tachypnea|0
blood pressure 100/70 mmHg|0
macular erythematous rash over both feet|0
Glasgow coma scale score 15|0
no neck stiffness|0
thrombocytopenia|0
high serum creatinine|0
high serum urea|0
high total bilirubin|0
high aspartate aminotransferase|0
high alanine aminotransferase|0
high C-reactive protein|0
chest X-rays bilateral haziness|0
started on empirical ceftriaxone|0
started IV fluids|0
provisionally diagnosed with acute gastroenteritis|0
acute kidney injury|0
admitted to the hospital|0
continued IV fluids|0
continued antibiotics|0
increased tachypnea|24
increased tachycardia|24
fever spike 38.3°C|24
hypoglycemia 2.9 mmol/L|24
worsening tachycardia|48
worsening tachypnea|48
hypotension|48
transferred to ICU|48
blood culture gram-negative bacilli|48
started piperacillin/tazobactam|48
intubated|48
ventilated due to respiratory distress|48
required vasopressors|72
required higher PEEP|72
blood culture positive for S. moniliforms|96
diagnosed with Rat Bite Fever|96
started intravenous penicillin G|96
weaned off ventilator|144
vasopressor tapered|144
improved renal functions|144
improved acidosis|144
extubated|144
discharged|240
no history of rat bite|0
rats present in house and workplace|0
frequently leaves food uncovered|0
no heart failure|240
no infective endocarditis|240
