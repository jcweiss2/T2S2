79 years old | 0
male | 0
admitted to the hospital | 0
increased shortness of breath | -96
pleuritic chest pain | -96
fevers | -96
non-productive cough | -96
Parkinson’s disease | 0
ischaemic heart disease | 0
hiatus hernia | 0
dysphagia | 0
tachycardic | 0
tachypnoeic | 0
hypotensive | 0
febrile | 0
reduced air entry in the right upper zone | 0
right basal crepitations | 0
aspiration pneumonia | 0
Acute Kidney Injury (AKI) stage 1 | 0
intravenous amoxicillin | 0
intravenous metronidazole | 0
intravenous fluids | 0
afebrile | 72
blood pressure 118/76 mmHg | 72
oxygen saturations 92% on 2 litres of oxygen per minute | 72
respiratory rate 20 breaths per minute | 72
CRP 297 | 72
WBC 8.0 | 72
improved renal function | 72
tachycardic | 96
tachypnoeic | 96
increasing oxygen requirements | 96
coarse crackles in the lung’s right lower zone | 96
intravenous piperacillin with tazobactam | 96
clarithromycin | 96
subcutaneous emphysema in the right hemithorax | 96
subcutaneous emphysema in the right neck | 96
subcutaneous emphysema in the right upper limb | 96
oxygen saturation 90% on 35% oxygen | 96
Type 1 Respiratory Failure | 96
stable blood pressure | 96
soft, non-tender abdomen | 96
no external signs of chest wall trauma | 96
extensive subcutaneous emphysema | 96
suspected pneumomediastinum | 96
urgent CT scan | 120
marked bilateral consolidation | 120
significant subcutaneous emphysema of the chest | 120
extensive pneumomediastinum | 120
right 2–3 mm anterior pneumothorax | 120
no pre-existing lung disease | 120
pneumomediastinum and subcutaneous emphysema secondary to severe pneumonia | 120
subcutaneous emphysema descended into his abdominal wall | 144
subcutaneous emphysema descended into his lower limbs | 144
clindamycin | 144
DNAR (Do Not Attempt Resuscitation) decision | 216
reviewed by the palliative care team | 216
died of septic shock | 216