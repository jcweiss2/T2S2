72 years old | 0
male | 0
admitted to the hospital | 0
history of hypertension | -8760
history of alcohol abuse | -8760
history of meningitis | -105120
acute change in mental status | -168
unsteady gait | -168
febrile | 0
tachycardic | 0
left band shift | 0
leukocytosis without elevated WBC | 0
WBC 6.2 × 103/µL | 0
nuchal rigidity | 0
altered mental status | 0
septic shock | 0
intravenous ceftriaxone | 0
intravenous vancomycin | 0
intravenous dexamethasone | 0
Streptococcus pneumoniae | 0
elevated total protein | 0
low albumin | 0
mild anemia | 0
elevated serum creatinine | 0
unprovoked pneumococcal infection | 0
multiple myeloma | 0
monoclonal gammopathy | 0
elevated IgG | 0
elevated β2-microglobulin | 0
hypercellular bone marrow | 0
monoclonal IgG lambda restricted plasma cells | 0
transferred to acute rehab | 168
neurological deficits | 168
fevers | 504
leukocytosis | 504
broad-spectrum antibiotics | 504
sepsis of unknown source | 504
Candida auris | 504
intravenous micafungin | 504
antifungal therapy | 504
induction chemotherapy | 672
CyBorD regimen | 672
cyclophosphamide | 672
bortezomib | 672
dexamethasone | 672
lenalidomide | 672
complete remission | 1344
recurrent infections | 1344