48 years old | 0
male | 0
admitted to the hospital | 0
generalised abdominal pains | -48
fever | -48
scanty urine | -48
painful irreducible right groin swelling | -120
absolute constipation | -120
vomiting | -120
reducible right groin swelling 11 years ago | -96288
ill-looking | 0
pale | 0
jaundiced | 0
dehydrated | 0
febrile (39.2°C) | 0
respiratory rate 25 breaths/min | 0
pulse rate 108 beats/min | 0
blood pressure 98/55 mmHg | 0
globally distended abdomen | 0
tense abdomen | 0
peritonism | 0
irreducible right inguinoscrotal swelling | 0
septic shock | 0
resuscitation with intravenous fluids | 0
intravenous ciprofloxacin 400 mg | 0
intravenous metronidazole 500 mg | 0
intranasal oxygen 4 L/min | 0
adrenaline administration | 0
blood transfusion 2 pints | 0
nasogastric tube insertion | 0
urethral catheter insertion | 0
optimal urine output >0.6 ml/kg/hour | 0
SPO2 94% | 0
blood pressure 115/70 mmHg | 0
pulse rate 86 bpm | 0
respiratory rate 22 cycles/min | 0
haemoglobin 7.4 g/dL | 0
leucocytosis 21×10^3 | 0
neutrophilia 83% | 0
decreased platelets 58×10^3 | 0
blood urea 11.2 mmol/L | 0
creatinine 162 μmol/L | 0
retroviral positive | 0
random blood sugar 6.1 mmol/L | 0
ASA score III | 0
informed consent for surgery | 0
general anaesthesia | 0
intubation | 0
extended midline incision | 0
free fluid with faecal matter | 0
herbal residue | 0
extensive exudate | 0
gangrenous perforated caecum | 0
mattered small bowel | 0
hernia sac containing redundant large bowel | 0
right hemicolectomy | 0
herniotomy | 0
nylon darn repair of posterior wall | 0
abdominal drain insertion | 0
peritoneum lavage | 0
post-operative blood transfusion | 24
continued intravenous antibiotics | 24
continued fluids | 24
analgesia | 24
intravenous KCL 50 mmol/day | 24
intravenous omeprazole 40 mg daily | 24
nil per oral | 24
graded oral intake after 72 hours | 72
oral medications | 72
several days to resume full feeds | 24
intravenous combined vitamins | 24
local formulated high carbohydrate diet | 24
weight loss 13.2 kg by week 4 | 672
exposed wound on day 2 | 48
cleaning with savlon | 48
normal saline irrigation | 48
povidone-iodine soaked gauze | 48
serosanguinous discharge | 48
offensive pus drainage by day 3 | 72
massive scrotal collection | 72
copious exudate | 72
daily wound cleaning | 72
cavity packed with povidone-iodine soaked gauze | 72
discharge subsided after 2 weeks | 336
daily dressing after 2 weeks | 336
granulation over nylon darn sutures at 5th week | 840
secondary suturing after 6th week | 1008
discharge after 8 weeks | 1344
parts of abdominal wound healed | 1344
continued wound dressing at primary facility | 1344
methylated spirit use | 1344
further investigations at Anti-Retroviral Clinic | 1344
no hernia recurrence 6 years after discharge | 52560
postoperative critical clinical events | 0
weight loss 13.2 kg within 2 weeks | 336
surgical site infection | 48
prolonged infection | 48
prolonged admission time | 48
extended antibiotics treatment | 48
extended dressing requirement | 48
perforated caecum | 0
soiled peritoneum | 0
major surgery (right hemicolectomy) | 0
retroviral status predisposing to infection | 0
nylon darn repair withstood infection | 0
granulation tissue over posterior wall repairs | 840
attempted closure of groin wound at 6th week | 1008
partially healed abdominal wound at discharge | 1344
HIV-associated lipodystrophy syndrome | -96288
rectus abdominis muscle separation | -96288
anterior abdominal wall hernias | -96288
risk factors for SSI | 0
advanced age | 0
ASA score > 2 | 0
immunosuppression | 0
emergency surgery | 0
low resource settings | 0
general anaesthesia use | 0
concurrent bilateral hernia repairs | 0
sliding hernia repairs | 0
viral load impact | 0
CD4 count impact | 0
increased risk of pneumonia | 0
increased mortality | 0
overall complications | 0
advanced disease consequences | 0
malnutrition | 0
infections | 0
hernia repair options | 0
open mesh repairs | 0
end-laparoscopic interventions | 0
Bassini method | 0
Shouldice method | 0
nylon darn repairs | 0
research on repair materials | 0
prolonged absorption duration | 0
improved tensile strength | 0
limited knots | 0
flexibility | 0
biocompatibility | 0
bacterial transmission prevention | 0
ideal material properties | 0
chemical impregnation | 0
poly-4-hydroxybutyrate use | 0
avoidance of porcine/human mesh | 0
bacteria resistance of nylon | 0
elasticity of nylon suture | 0
pore size maintenance | 0
purulent material escape | 0
minimal intersections and pull-outs | 0
successful management factors | 0
method of repair | 0
infected nylon darn maintained properties | 0
no hernia recurrence after 6 years | 52560
no prior lower urinary tract symptoms | -96288
no prior chronic cough | -96288
no prior chronic constipation | -96288
no prior co-morbidity | -96288
no diagnostic investigation | 0
no intensive care unit admission | 0
no mesh removal | 0
no advanced disease | 0
no chronic cough | -96288
no chronic constipation | -96288
no co-morbidity | -96288
no antiretroviral treatment | 0
no hernia recurrence | 52560
no evidence of hernia recurrence | 52560
no conflict of interest | 0
