22 years old | 0
male | 0
admitted to the hospital | 0
Crohn's colitis | -8760
fistulectomy | -8760
complex perianal fistula | -8760
severe weight loss | -8760
diarrhea | -8760
abdominal pain | -8760
recurrent perianal tenderness | -8760
mesalamine | -8760
herbal medicine | -8760
fistular openings | 0
subcutaneous abscess pockets | 0
severe tenderness | 0
mild fever | 0
complicated anal fistulas | 0
perianal abscesses | 0
multiple and diffuse aphthous ulcerations | 0
multifocal inflammatory wall thickening | 0
thick-walled abscess pockets | 0
subcutaneous small abscesses | 0
Crohn's disease activity index (CDAI) was 244 | 0
abscess drainage | 0
seton operation | 0
AZA administered | 0
high fever | 14
myalgia | 14
leukocytes were 180/μl | 14
hemoglobin was 6.6 g/dl | 14
platelets were 48,000/μl | 14
ESR was 55 mm/h | 14
CRP was 24.7 mg/l | 14
AZA discontinued | 14
pancytopenia | 14
septicemia | 14
human recombinant granulocyte colony-stimulating factor | 14
broad-spectrum antibiotic therapy | 14
fever subsided | 28
cell count fully recovered | 28
Escherichia coli found on blood culture | 28
TPMT was the wild type (*1/*1) | 28
frequency of bowel movements decreased | 28
perianal pain and oozing improved | 28
follow-up colonoscopy | 84
diffuse fibrotic scar | 84
gained 10 kg | 168
CDAI score = 114 | 168
clinical recurrence | 0