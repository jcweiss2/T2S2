fever | -72
chills | -72
pain in left leg | -72
cellulitis | -72
high-temperature spikes | -48
tachycardia | -48
tachypnea | -48
hypotensive | -48
encephalopathic | -48
admitted to ICU | 0
intravenous clindamycin | -72
intravenous benzylpenicillin | -72
levodopa / carbidopa | -72
rasagiline | -72
ropinirole | -72
trihexyphenidyl | -72
amantadine | -72
metformin | -72
glipizide | -72
intravenous linezolid | 24
intravenous piperacillin with tazobactam | 24
confused | 24
drowsy | 24
disoriented | 24
altered sensorium | 24
myoclonus | 24
tremors | 24
jerky movements | 24
no neck stiffness | 24
computed tomography of the brain | 24
cerebrospinal fluid analysis | 24
improving white blood cell counts | 24
better glycemic control | 24
sterile blood and pus cultures | 24
high temperature | 48
altered mental status | 48
myoclonus | 48
jerky movements | 48
tremors | 48
suspected serotonin syndrome | 48
stopped linezolid | 48
stopped rasagiline | 48
temperature settled | 56
heart rate normal | 72
sensorium improved | 72
tremors subsided | 72
shifted out of ICU | 96
started walking with support | 240
discharged from hospital | 240
added rasagiline | 240
stable and asymptomatic for serotonin syndrome | 240