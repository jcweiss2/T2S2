54 years old | 0
male | 0
chronic alcoholic | 0
COPD | 0
admitted to the hospital | 0
delirious state | 0
alcohol withdrawal syndrome | 0
deteriorated clinically | 24
high-grade fever | 24
continuous cough | 24
hypotension | 24
hypoxemia | 24
sepsis | 24
Type II respiratory failure | 24
neutrophilic leukocytosis | 24
anemia | 24
low RBC count | 24
high MCV | 24
high MCHC | 24
bandemia | 24
toxic granulation | 24
clumping of RBCs | 24
polychromatophilic cells | 24
nucleated RBCs | 24
high reticulocyte count | 24
hemoglobinemia | 24
raised lactate dehydrogenase | 24
mildly raised unconjugated bilirubin | 24
agglutination of blood | 24
autoagglutination | 24
atypical pneumonia | 24
bilateral pulmonary interstitial infiltrates | 24
cold agglutinin disease (CAD) | 24
discharged | 120
advice to avoid cold temperature | 120
COPD diagnosis | -8760
alcoholism diagnosis | -8760
admission to acute medical ward | 0
shifted to intensive care unit | 24
treated for sepsis | 24
treated for atypical pneumonia | 24
treated for alcohol withdrawal syndrome | 24
treated for COPD | 24
diagnosed with CAD | 24
Coomb's test negative | 24
autoagglutination test positive | 24 
chest X-ray | 24 
blood sampling | 24 
peripheral blood smear | 24 
biochemical tests | 24 
supravital stain | 24 
incubation at 37°C | 24 
refrigeration | 24 
warming of sample | 24 
analysis of report | 24 
reversal of agglutination | 24 
maintenance of pregnancy | -8760 
transfusion | -8760 
cross-matching | -8760 
in-line warmer | -8760 
severe hemolysis | -8760 
renal shutdown | -8760 
gangrene of fingers or toes | -8760 
patient consent | 0 
financial support | 0 
conflicts of interest | 0 
acknowledgment | 0