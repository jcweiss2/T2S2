82 years old | 0
woman | 0
arterial hypertension | -0
admitted to ICU | 0
septic shock | 0
heart rate 124/min | 0
blood pressure 80/45 mmHg | 0
no response after 1-L crystalloid fluid expansion | 0
polypnea 28 cycles/min | 0
no respiratory distress sign | 0
tense abdomen | 0
painful abdomen on palpation | 0
hyperlactatemia | 0
metabolic acidosis | 0
pH 7.21 | 0
PCO2 24 mmHg | 0
bicarbonate 14 mmol/L | 0
lactate 9 mmol/L | 0
liver abscess | 0
mechanical ventilation | 0
continuous norepinephrine infusion 8 mg/h | 0
piperacillin/tazobactam 4g daily | 0
gentamicin 480 mg | 0
emergency laparotomy | 0
liver abscess drainage | 0
crepitation of thoracic and cervical region | 0
subcutaneous emphysema | 0
massive subcutaneous emphysema | 0
pneumoperitoneum | 0
no SE during first physical examination | 0
no SE on first CT scan | 0
no upper airway injuries | 0
no pneumothorax | 0
suspected surgical complication | 0
second emergency laparotomy | 0
perforated transverse colon | 0
5 cm colon removed | 0
colostomy | 0
multiorgan failure | 0
death | 120
arterial hypertension | -8760
gentamicin 480 mg |;0
crepitation of thoracic and cervical region | 12
subcutaneous emphysema | 12
massive subcutaneous emphysema | 12
pneumoperitoneum | 12
suspected surgical complication | 24
second emergency laparotomy | 24
perforated transverse colon | 24
5 cm colon removed | 24
colostomy | 24
multiorgan failure | 120
- arterial hypertension | -8760 (assuming 1 year prior)
