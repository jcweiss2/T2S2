2 years old | 0
female | 0
born full term | -7300
spontaneous vaginal delivery | -7300
prolonged obstructive jaundice | -168
steatorrhea | -168
generalized itchiness | -168
ultrasound abdomen | -168
contrast-enhanced computed tomography (CT) scan | -168
choledochol cyst | -168
scheduled for portoenterostomy (KASAI procedure) | -168
scheduled for liver biopsy | -168
scheduled for on-table cholangiogram | -168
caudal epidural catheter insertion | 0
skin to space distance was 1.5 cm | 0
catheter advanced 10 cm | 0
minimal twisting | 0
measuring at approximately the T7 dermatome | 0
ultrasound guidance | 0
surgery | 0
extubated | 24
discharged back to ward | 24
epidural infusion functioning well | 24
pain well-controlled | 24
planned to remove epidural catheter | 48
resistance encountered while removing catheter | 48
catheter suddenly “fell off” | 48
end segment sheared off | 48
6 cm left inside space | 48
segment appeared to be twisted and crimped | 48
no remnant of catheter noted around skin area | 48
informed surgeon and patient's parents | 48
urgent MRI thoracolumbar | 48
non-contrast CT scan spine | 48
catheter tip retained from upper border of L4 vertebra | 48
retained catheter segment approximately 6 cm in length | 48
no other remnant of catheter noted | 48
persistent vomiting | 72
fever | 72
total white count increased | 72
no neurological deficit | 72
differential diagnosis includes pathology from laparotomy | 72
differential diagnosis includes sepsis | 72
differential diagnosis includes retained catheter tip | 72
CT brain urgent | 72
normal finding without mass effect or hydrocephalus | 72
repeated CT scan spine | 72
no catheter migration | 72
no other abnormal findings | 72
no focal swelling or collection | 72
fever subsided | 120
vomiting persists | 120
relaparotomy | 432
adhesions found | 432
adhesiolysis | 432
small bowel resection | 432
side-to-side anastomosis | 432
extubated well | 456
discharged home | 504
decided to let fragment remain in situ | 504
continue to follow-up patient | 504
patient's parents advised to report adverse symptoms | 504
patient remained asymptomatic | 8760
no symptoms of complication | 8760