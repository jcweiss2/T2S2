9-year-old | 0
boy | 0
presented to the emergency department | 0
abdominal pain | -12
abdominal pain worsened in the supile position | -12
two episodes of nonbilious vomiting | -12
no fever | 0
stool output via colostomy was normal | 0
spina bifida | 0
hydrocephalus | 0
imperforate anus | 0
scoliosis | 0
solitary kidney | 0
multiple urinary tract infections | 0
ventriculoperitoneal shunt | 0
colostomy | 0
titanium rib placement | 0
Monti procedure | -1680
Monti procedure performed 2½ months prior to ED visit | -1680
catheterization schedule every 3 hours from 6 AM to 9 PM | 0
always having a little blood with catheterization | 0
intermittent difficulty catheterizing the vesicostomy for 1 week | -168
catheter deviating to the right | -168
mild difficulty inserting the catheter | 0
good output | 0
heart rate 166 beats/min | 0
blood pressure 132/90 | 0
respiratory rate 25 breaths/min | 0
temperature 99.6 | 0
oxygen saturation 98% | 0
alert | 0
talkative | 0
comfortable in sitting position | 0
pain when placed supine | 0
abdominal distension in superior quadrants | 0
evaluation for tenderness and guarding difficult due to body habitus and sensory level at T10 | 0
white blood cell count 32.1 ×10³/mm³ | 0
77% neutrophils | 0
14% bands | 0
serum bicarbonate 12 mEq/L | 0
BUN 24 mg/dL | 0
Foley catheter initially obtained cloudy, blood-tinged fluid | 0
malodorous urine | 0
urine with 50–100 RBC/HPF | 0
urine with 50–100 WBC/HPF | 0
nitrite negative | 0
leukocyte esterase 3+ | 0
Foley catheter left in ileovesicostomy | 0
balloon inflated | 0
CT scan of abdomen and pelvis with IV contrast obtained | 24
ascitic fluid larger than expected | 24
no evidence of pseudocyst | 24
worsening hydronephrosis of solitary kidney | 24
CT cystogram performed | 24
urine extravasation into peritoneal cavity | 24
Foley catheter balloon outside bladder through perforation of continent ileovesicostomy | 24
infected urine causing peritonitis | 24
neurosurgery consulted | 24
urology consulted | 24
CT scan of brain requested | 24
cerebrospinal fluid clear | 24
head CT showed mild increase in ventricular size | 24
fracture in shunt tubing at postauricular level | 24
plans to externalize proximal portion of shunt | 24
remove indwelling shunt | 24
urology provided details of urologic procedure 10 weeks previously | -1680
bladder neck reconstruction | -1680
right ureteral implant | -1680
construction of Monti channel vesicostomy | -1680
bladder not augmented | 0
no appendix at time of reconstruction | 0
urologist planned endoscopy of Monti channel | 24
cystoscopy with further intervention | 24
received fluid bolus | 24
received cefepime in ED | 24
admitted to PICU | 24
worsening tachycardia | 24
diminished pulses | 24
compensated septic shock | 24
given vancomycin | 24
additional fluid bolus | 24
fluid resuscitation | 24
taken to surgery | 24
proximal shunt externalized | 24
incision on abdomen | 24
distal catheter removed | 24
distal peritoneal catheter externalized | 24
purulent material aspirated from peritoneal cavity | 24
endoscopy of catheterizable stoma revealed large posterior false passage | 24
catheter placed across stoma into bladder | 24
cystoscopy and cystogram after proper catheter placement | 24
no bladder perforation | 24
additional Foley catheter placed into bladder via native urethra | 24
dilation of bladder neck | 24
required mechanical ventilation | 48
low-dose norepinephrine for 24 hours | 48
urine culture grew Escherichia coli | 48
different sensitivities than culture 6 weeks previously | 48
all cultures of shunt and peritoneal fluid negative | 48
removal of retained fractured shunt catheter in supraclavicular region | 144
peritoneal catheter removed | 144
original shunt converted to ventriculocardiac shunt | 264
discharged after 14 days of intravenous antibiotics | 336
urethral catheter to gravity drainage | 336
vesicostomy catheters to gravity drainage | 336
Monti catheter left in place for 4 weeks | 336
cystoscopy performed for perceived difficulty in catheterization | 672
no stenosis | 672
no false passage | 672
catheterization difficulty | 1344
urinary retention | 1344
another cystoscopy revealed false passage | 1344
Monti revision for stenosis of channel at bladder junction | 4032
