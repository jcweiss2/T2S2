64 years old | 0
male | 0
hypertension | 0
type II diabetes mellitus | 0
admitted to the hospital | 0
left-sided hemiparesis | 0
right-sided facial deviation | 0
slurring of speech | 0
Broca's aphasia | 0
upper motor neuron (UMN) type VIIth cranial nerve (CN) palsy | 0
up-going plantar reflex on the left side | 0
power on the left upper limb 3/5 | 0
power on the left lower limb 4/5 | 0
Total Leukocytes Count 15.5 | 0
Neutrophil 65 | 0
Lymphocyte 28 | 0
Hemoglobin 14.8 | 0
Platelet Count 213 | 0
Urea 41 | 0
Creatinine 1.2 | 0
Sodium 140 | 0
Potassium 5.1 | 0
Bilirubin Total 1.1 | 0
Bilirubin Direct 0.4 | 0
Alkaline Phosphatase (ALP) 85 | 0
Alanine Transferase (ALT) 20 | 0
Aspartate Transferase (AST) 23 | 0
Prothrombin Time 13.1 | 0
International Normalized Ratio 1.0 | 0
HbA1C 13.9 | 0
Random Blood Glucose 331 | 0
infarction over the right hemisphere (temporo-parietal area) | 0
Ramipril 5 mg once daily | 0
Amlodipine 5 mg once daily | 0
Metformin 500 mg once daily | 0
Sitagliptin 100 mg once daily | 0
Empaglifozin 10 mg once daily | 0
Insulin 10 units subcutaneously once daily | 0
Aspirin 75 mg once daily | 0
Statins 10 mg once daily | 0
GRBS 186 | 24
GRBS 103 | 48
GRBS 117 | 72
GRBS 145 | 96
drowsy | 120
rapid breathing | 120
fall in Glasgow Coma scale (GCS) | 120
E3V4M5 | 120
GRBS 218 | 120
oxygen saturation 98% | 120
blood pressure 120/80 mmHg | 120
severe metabolic acidosis | 120
pH 7.124 | 120
HCO3 4.1 | 120
PaCO2 12.7 mm of Hg | 120
PaO2 90 mm of Hg | 120
Anion gap 25 | 120
Lactate 1.86 | 120
urine acetone positive | 120
Euglycemic DKA | 120
NaHCO3 50 mEq | 120
ABG analysis | 120
pH 7.214 | 120
HCO3 5.1 | 120
PCO2 13 | 120
PO2 116 | 120
Lactate 1.71 | 120
normal saline infusion | 120
NaHCO3 50 mEq | 120
piperacillin and tazobactam 4.5 gm thrice daily | 120
regular insulin infusion 2 units/hour | 120
empaglifozin stopped | 120
shifted to ICU | 120
ABG analysis | 144
bicarbonate level 13.4 mEq/L | 144
normal anion gap | 144
intubated and mechanically ventilated | 168
sepsis | 168
qSOFA score 2 | 168
blood pressure 110/80 mmHg | 168
respiratory rate 28 | 168
GCS 11/15 | 168
levofloxacin 750 mg once daily | 168
vancomycin 15 mg/kg/dose every 8 hours | 168
linezolid 600 mg every 12 hours | 168
colistin 300 mg loading dose | 168
colistin 150 mg twice daily | 168
spontaneous CPAP breathing trial | 312
passed the breathing trial | 312
shifted to HCU | 312
glycemic control target 110-180 mg/dl | 312
Insulin Glargine 10 units subcutaneous once daily | 312
Insulin Aspart 4 units subcutaneously before meal thrice daily | 312
stable in HCU | 312
normal vital parameters | 312
bed side mobilization | 312
chest/limb physiotherapy | 312
discharged from the hospital | 432