18 years old | 0\
male | 0\
Mayer Rokitansky-Küster-Hauser (MRKH) syndrome | 0\
congenital aplasia of the uterus and upper part of the vagina | 0\
normal secondary sex characteristics | 0\
female karyotype | 0\
primary amenorrhea | 0\
adolescence | -672\
diagnosed with MRKH syndrome | -672\
treatment options | -672\
creation of a functional neovagina | -672\
sigmoid vaginoplasty | -672\
safe procedure for vaginal agenesis | -672\
good cosmetic results | -672\
large lumen | -672\
thick walls resistant to trauma | -672\
adequate secretions for lubrification | -672\
not requiring prolonged dilatation | -672\
short recovery time | -672\
perforation of the neovagina | -672\
extremely rare | -672\
rare with only handful of cases reported | -672\
all cases occurred in transgender patients | -672\
27 years old | 0\
presented to the clinic | 0\
lower abdominal pain | 0\
bilateral pelvic pain | 0\
two weeks duration | 0\
denies routinely irrigating or dilating her neovagina | 0\
normally had penetrative sexual intercourse | 0\
every couple of weeks | 0\
life stressors | 0\
had not had intercourse in a few months | 0\
CT imaging of the abdomen | 0\
tubular, heterogenous, fluid-filled structure | 0\
extending from the pelvis to the lower abdomen | 0\
measuring 7.1 cm × 20 cm | 0\
blind ending | 0\
outpatient referral to the gynecologist | 0\
abdominal pain acutely worsened | 24\
presented to the local Emergency Department (ED) | 24\
diaphoresis | 24\
significant distress due to pain | 24\
unremarkable vitals | 24\
Complete blood count (CBC) | 24\
leukocytosis of 15.6 k/mm3 | 24\
absolute neutrophils of 9.8 k/mm3 | 24\
repeat abdominal CT | 24\
increasing inflammatory process in the pelvis | 24\
surrounding the reconstructed vagina | 24\
empiric intravenous (IV) piperacillin-tazobactam | 24\
transferred emergently to our children’s hospital | 24\
associated with her urologist | 24\
on arrival to our facility | 24\
hypotensive | 24\
tachycardic | 24\
afebrile | 24\
tachypneic | 24\
oxygen saturation of 95 % on room air | 24\
four IV fluid boluses | 24\
antimicrobials were empirically changed | 24\
IV ceftriaxone, IV vancomycin, and IV metronidazole | 24\
taken emergently to the operative room (OR) | 24\
exploratory laparotomy, cystoscopy, and vaginoscopy | 24\
intra-operatively | 24\
normal bladder and urethra | 24\
entirely obliterated introitus | 24\
diffuse intra-abdominal spillage of the mucus | 24\
perforated sigmoid neovagina | 24\
about one liter of purulent fluid was drained | 24\
three intrabdominal drains were placed | 24\
post-operatively | 24\
remained intubated requiring mechanical ventilation | 24\
in septic shock requiring three vasopressor agents | 24\
antimicrobials were transitioned | 24\
IV cefepime, IV vancomycin, and IV metronidazole | 24\
due to preliminary peritoneal culture growing gram-negative rods | 24\
blood cultures remained negative | 24\
peritoneal cultures finalized | 24\
Bacterioides thetaioaomicron, Bacteroides caccae, and Actinomyces species | 24\
antimicrobials were changed | 24\
IV piperacillin-tazobactam | 24\
day 7 of her hospitalization | 168\
weaned off vasopressors | 168\
extubated | 168\
day 8 | 168\
transferred to the general floor | 168\
Infectious Diseases team was consulted | 168\
antimicrobial management | 168\
additional susceptibilities for the Bacteroides species | 168\
were requested | 168\
pending | 168\
patient was discharged home | 168\
day 15 | 168\
abdominal wound vacuum | 168\
IV piperacillin-tazobactam for four weeks | 168\
plan for close follow-up | 168\
two weeks post-discharge | 168\
experienced generalized malaise | 168\
diffuse abdominal pain | 168\
readmitted with sepsis | 168\
laboratory data revealed | 168\
white blood count 13.2 k/cmm3 | 168\
absolute neutrophil count 9.5 k/cmm3 | 168\
d-dimer >5000 ng/mL DDU | 168\
lactate 0.9 mmol/L | 168\
CT of the chest, abdomen and pelvis | 168\
bilateral pleural effusions | 168\
loculated left pleural effusion | 168\
multiple new abdominal abscesses | 168\
largest next to the liver (15.6 cm) | 168\
transcutaneous drainage catheter in pelvis | 168\
open anterior midline wound with wound vacuum | 168\
due to hypoxemia | 168\
transferred to the intensive care unit (ICU) | 168\
IV piperacillin-tazobactam was continued | 168\
placement of a right perihepatic drain | 168\
aspiration of 20 mL of purulence | 168\
unsuccessful drainage of peri-splenic collection | 168\
blood cultures remained negative | 168\
interventional radiology was reconsulted | 168\
drained 350 mL of pus from the right perinephric abscess | 168\
90 mL of pus from her perisplenic abscess | 168\
broad-spectrum PCR was sent | 168\
on the drained fluid from the abscesses | 168\
positive for Gleimia europaea | 168\
Alistipes onderdonkil | 168\
Varibaculum timonense | 168\
Jonquetella anthropi | 168\
antimicrobials were narrowed | 168\
IV ampicillin-sulbactam | 168\
day 32 from the initial presentation | 192\
discharged | 192\
based on the susceptibilities from the original surgical cultures | 192\
broad-spectrum PCR from the fluid | 192\
positive for Gleimia europaea | 192\
Alistipes onderdonkil | 192\
Varibaculum timonense | 192\
Jonquetella anthropi | 192\
followed up at the adult infectious diseases clinic | 192\
continued on ampicillin-sulbactam | 192\
plans to reimage on day 60 | 192\
repeat CT abdomen | 192\
demonstrated decreased in the size of right and left sub-phrenic abscesses | 192\
transitioned from IV ampicillin-sulbactam | 192\
oral amoxicillin-clavulanate | 192\
several weeks | 192\
until complete resolution of the abscesses | 192\
day 60 | 240