31 years old | 0
female | 0
Aboriginal | 0
admitted to the hospital | 0
congenital bicuspid aortic valve | -6336
bicuspid aortic valve diagnosis | -6336
severe stenosis | -6336
severe regurgitation | -6336
aneurysm of the ascending aorta | -6336
aortic valve replacement | -2184
aortic root replacement | -2184
biventricular pacemaker insertion | -2184
type 2 diabetes mellitus | -2184
hypertension | -2184
smoking | -2184
suboptimal adherence to metformin | -2184
suboptimal adherence to bisoprolol | -2184
suboptimal adherence to aspirin | -2184
headaches | -168
fevers | -168
confusion | -168
seizures | -168
aeromedical retrieval | 24
meningoencephalitis treatment | 24
blood cultures positive for methicillin-resistant Staphylococcus aureus | 72
transoesophageal echocardiogram confirming aortic prosthetic valve endocarditis | 72
cardiac case conference | 144
medical treatment with flucloxacillin and rifampicin | 144
craniotomy and drainage of brain abscess | 360
brain abscess culture positive for S. aureus | 360
baseline positron emission tomography-fluorodeoxyglucose | 1008
para-valvular and peri-aortic abscess formation | 1080
bilateral pseudo-aneurysms | 1080
aeromedical transfer to interstate cardiothoracic surgery facility | 1200
redo-bioprosthetic aortic valve replacement | 1344
aortic root replacement | 1344
biventricular pacemaker explantation | 1344
biventricular pacemaker re-insertion | 1350
discharged against medical advice | 2112
lost to follow-up | 2112
presented to remote community clinic | 2760
commenced high-dose oral dicloxacillin and rifampicin | 2760
PET-FDG with no AVR or extra-cardiac uptake | 2976
CTCA showing two pseudo-aneurysms stable in size | 2976
CTCA showing two pseudo-aneurysms essentially unchanged | 4704
transthoracic echocardiogram showing normal bioprosthetic valve function | 10008
normocytic anaemia | 0
elevated C-reactive protein | 0
normal white cell count | 0
lumbar puncture results suggesting bacterial meningitis | 0
septic shock | 0
intensive care unit admission | 0
antibiotics rationalised to IV flucloxacillin | 0
treatment for hyperglycaemia | 0
treatment for anaemia | 0
red blood cell transfusion | 0
diuresis for biventricular heart failure | 0
electrocardiogram showing sinus rhythm with ventricular pacing | 0
electrocardiogram showing left bundle branch block | 0
cardiac imaging revealing a small mobile echodensity on the bioprosthetic AVR | 0
magnetic resonance imaging brain confirming multiple cerebral infarcts | 144
CT brain showing an evolving left frontal lobe cerebral abscess | 312
neurosurgical intervention with drainage of a 30 × 40 × 20 mm abscess | 312
repeat transthoracic echocardiogram unchanged | 312
rifampicin added for adjuvant biofilm activity | 312
discharged against medical advice from the ward | 312
interruptions to IV flucloxacillin and oral rifampicin | 312
fluorodeoxyglucose-positron emission tomography | 1008
follow-up TTE revealed new mild paravalvular aortic incompetence | 1080
transoesophageal echocardiogram demonstrating formation of two pseudo-aneurysms | 1080
CT coronary angiogram confirming para-valvular and peri-aortic abscess formation | 1080
bilateral pseudo-aneurysms | 1080
urgent transfer to interstate cardiac surgical centre | 1200
redo-bioprosthetic aortic valve replacement | 1344
aortic root replacement | 1344
biventricular pacemaker explantation | 1344
biventricular pacemaker re-insertion | 1350
planned for a further 6 weeks IV flucloxacillin and rifampicin post AVR | 1344
discharged against medical advice | 2112
lost to follow-up | 2112
presented to remote community clinic | 2760
commenced high-dose oral dicloxacillin and rifampicin | 2760
PET-FDG with no AVR or extra-cardiac uptake | 2976
CTCA showing two pseudo-aneurysms stable in size | 2976
CTCA showing two pseudo-aneurysms essentially unchanged | 4704
transthoracic echocardiogram showing normal bioprosthetic valve function | 10008