20 years old | 0
female | 0
primigravida | 0
admitted to the hospital | 0
breathing difficulty | 0
intubated | 0
respiratory distress | 0
transferred to critical care department | 0
no significant past medical history | 0
no genetic history | 0
no history of complications during pregnancy | 0
Glasgow coma scale (GCS) was E4M6Vt | 0
temperature was 101°F | 0
pulse was 122 beats/minute | 0
blood pressure was 118/78 mm Hg | 0
no rash | 0
bilateral crepitations | 0
bilateral infiltrates on chest X-ray | 0
poor left ventricle (LV) systolic function | 0
no right atrium (RA)/right ventricle (RV) dilatation | 0
treated for pneumonia | 0
treated for sepsis | 0
treated for acute kidney injury (AKI) | 0
treated for peripartum cardiomyopathy | 0
persistent high-grade fever | 24
gross muscle weakness | 120
involving all four limbs | 120
predominantly in proximal muscles | 120
dark colored urine | 120
positive urine myoglobin | 120
raised erythrocyte sedimentation rate (ESR) | 120
raised serum creatine phosphokinase (CPK) levels | 120
raised lactate dehydrogenase (LDH) levels | 120
normal thyroid function tests | 120
Systemic lupus erythematosus (SLE) ruled out | 120
negative antinuclear antibody (ANA) | 120
negative anti-dsDNA antibody | 120
rhabdomyolysis considered as differential diagnosis | 120
inflammatory myopathy suspected | 120
Magnetic resonance imaging (MRI) of cervical spine showed diffuse edema | 144
Electromyography (EMG) showed myopathic pattern | 144
muscle biopsy from the left thigh muscle showed inflammatory reaction | 144
Polymyositis diagnosed | 144
started on high dose of intravenous (IV) steroids | 144
tracheostomy performed | 240
liberated from mechanical ventilator | 456
decannulated | 456
bulbar weakness persisted | 456
intermittent cough | 456
intolerance to oral feeds | 456
retained secretions | 456
Videolaryngoscopy performed | 456
dysphagia due to cricopharyngeal muscle discordance | 456
continued to feed through Ryles tube | 456
improved gradually | 504
CPK levels decreased | 504
able to walk without support | 504
started to take oral feeds | 504
discharged on tapering dose of oral steroids | 504
followed up after 2 weeks | 720
followed up monthly | 720
prednisone dose tapered | 720
counseled to avoid conception for a year | 720
delivered a dead fetus | -96
pregnancy | -672
intrauterine fetal death | -96