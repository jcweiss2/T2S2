78 years old | 0
male | 0
presented to the emergency department | 0
dyspnea exacerbating | -240
shortness of breath | 0
cough | 0
anosmia | 0
myalgia | 0
hypertension | 0
Valsartan tablet 80 mg | 0
tachycardia | 0
normal core temperature | 0
tachypnea | 0
oxygen saturation 72% | 0
Glasgow Coma Scale 12 | 0
nasopharyngeal swab test positive | 0
plasma lactate 65 mg/dL | 0
albumin 2.5 g/L | 0
C-Reactive Protein 163 mg/L |:0
high sensitivity troponin 103 ng/ml | 0
creatine kinase myocardial band 66 IU/L | 0
chest CT diffuse bilateral ground-glass opacities | 0
mild pleural effusion | 0
cardiomegaly | 0
atrial fibrillation | 0
reduced left ventricular ejection fraction 15% | 0
high pulmonary arterial pressure 50 mmHg | 0
mildly enlarged LV | 0
moderate to severe LV dysfunction | 0
mild diastolic dysfunction grade 1 | 0
mild mitral valve regurgitation | 0
normal septal thickness | 0
intubated | 0
transferred to ICU | 0
USCOM low systemic vascular resistance | 0
low cardiac output | 0
low oxygen delivery | 0
cardiogenic shock | 0
septic shock | 0
Hydroxychloroquine 400 mg twice daily | 0
Hydroxychloroquine 200 mg twice daily | 0
Dexamethasone 16 mg daily | 0
Intravenous Immunoglobulin 10 g | 0
Ascorbic acid 1 g four times daily | 0
Melatonin 18 mg daily | 0
broad-spectrum antibiotics | 0
echocardiographic LVEF 25% | 600
PAP 38 mmHg | 600
moderate LV dysfunction | 600
right ventricular dilation | 600
LVEF 35% | 840
PAP 55 mmHg | 840
mild RV dilation | 840
respiratory distress improved | 840
LVEF 45% | 1008
PAP 45 mmHg | 1008
mild RV dilation | 1008
vasopressor | 0
amiodarone | 0
Midodrine | 0
hemodynamic parameters stable | 1008
wean mechanical ventilation | 1008
discharged from ICU | 1008
respiratory arrest | 1104
cardiopulmonary resuscitation | 1104
expired | 1104
