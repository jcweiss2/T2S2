20 years old | 0  
    male | 0  
    motor vehicle accident | 0  
    severe and diffuse trauma to the abdomen | 0  
    severe and diffuse trauma to the trunk | 0  
    severe and diffuse trauma to the extremities | 0  
    unstable vital signs | 0  
    flaccid paraplegia | 0  
    cord level at T10 | 0  
    complete loss of voluntary control over bowel function | 0  
    complete loss of voluntary control over bladder function | 0  
    FAST examination negative | 0  
    multiple rib fractures | 0  
    bilateral hemothoraces | 0  
    hemoperitoneum | 0  
    AAST grade 4 splenic injury | 0  
    left-sided renal injury | 0  
    left-sided adrenal injury | 0  
    right-sided scapular fracture | 0  
    transdiscal AO type C fracture | 0  
    bilateral facet subluxation of T11 over T12 | 0  
    pneumothoraces drained through chest tubes | 0  
    exploratory laparotomy | 0  
    splenectomy | 0  
    left retroperitoneal space packed | 0  
    large retroperitoneal hematoma | 0  
    kidney injury | 0  
    adrenal injury | 0  
    Damage Control surgery | 0  
    hemodynamic instability | 0  
    no other lesions identified | 0  
    transferred to Intensive Care Unit | 0  
    PAD 1 | 24  
    MRI of the spine | 24  
    subluxation of T11 over T12 | 24  
    rupture of the intervertebral disc | 24  
    rupture of the posterior longitudinal ligament | 24  
    9 mm-thick epidural hematoma overlying T11 | 24  
    medullary contusion at T11-T12 | 24  
    PAD 2 | 48  
    spinal surgery | 48  
    reduction of the subluxation | 48  
    trans-pedicular screw fixation from T9 to L2 | 48  
    intra-operative post-traumatic dural tear | 48  
    small leak of CSF | 48  
    no repair attempted | 48  
    PAD 3 | 72  
    second look laparotomy | 72  
    no bleeding observed | 72  
    persistence of the retroperitoneal hematoma | 72  
    small amount of turbid liquid identified | 72  
    no lesions found in small intestine | 72  
    no lesions found in colon | 72  
    intense back pain | 72  
    not responsive to opiates | 72  
    hallucinations | 72  
    agitated | 72  
    septic state | 72  
    thoracolumbar MRI | 72  
    thoraco-abdominal CT | 72  
    large bilateral paravertebral fluid collections | 72  
    large retroperitoneal fluid collections | 72  
    AAST grade 3 pancreatic injury | 72  
    retroperitoneal hematoma | 72  
    revision of the thoraco-lumbar wound | 72  
    CSF leak from circular dural breach | 72  
    fibrin sealant repair | 72  
    debridement of necrotic tissue | 72  
    drainage of purulent collections | 72  
    copious irrigation with normal saline | 72  
    tight closure of the facia | 72  
    tight closure of the subcutaneous tissue | 72  
    Penrose drains left in superficial layers | 72  
    retroperitoneal fluid collections evacuated | 72  
    percutaneous CT-guided drain placement | 72  
    blood cultures positive for Enterobacter cloacae | 72  
    paravertebral fluid collections positive for Enterobacter cloacae | 72  
    abdominal fluid collections positive for Enterobacter cloacae | 72  
    intravenous Meropenem | 72  
    paravertebral collections increased | 72  
    abdominal collections increased | 72  
    repeat cultures positive for Enterobacter cloacae | 72  
    paravertebral collections exteriorized through dorsal skin | 72  
    three new locations of exteriorization | 72  
    serum amylase high up to 3 times norm | 168  
    serum lipase high up to 3 times norm | 168  
    serum amylase returned to baseline | 168  
    serum lipase returned to baseline | 168  
    high amylase in dorsal spinal fluid collections | 168  
    high lipase in dorsal spinal fluid collections | 168  
    ERCP performed | 168  
    stent placement bridging defect of main duct | 168  
    reoperation for debridement | 168  
    drainage of recurrent paravertebral collection | 168  
    fibrin sealant reapplication | 168  
    total parenteral nutrition for 15 days | 168  
    subcutaneous somatostatin introduced | 168  
    proton pump inhibitors | 168  
    enteral feeding by naso-jejunal tube | 168  
    parenteral alimentation | 168  
    gradual oral feeding | 168  
    enteral intake weaned off | 168  
    parenteral intake weaned off | 168  
    general condition improvement | 168  
    progressive resolution of fluid collections | 168  
    drains removed | 168  
    transferred to rehabilitation facility | 1248  
    complete paraplegia | 1248  
    sensory level at T10 | 1248  
    antibiotic treatment for 7 months | 1248  
    complete resolution of spinal collections | 1248  
    complete resolution of retroperitoneal collections | 1248  
