66 years old | 0
male | 0
evaluated at the emergency department | 0
asthenia | -24
adynamia | -24
mild dyspnoea | -24
dry cough | -24
chills | -24
fever | -24
diaphoresis | -24
alteration of the consciousness state | -24
disorientation | -24
episodes of agitation | -24
great respiratory difficulty | -24
desaturation | -24
hypertensive nephropathy | -8760
polycystic kidney disease | -8760
renal transplantation | -8760
immunosuppressive treatment with tacrolimus | -8760
tacrolimus | -8760
prednisolone | -8760
azathioprine | -8760
chest x-ray performed | 0
consolidation in the middle third of the left pulmonary field | 0
shifted to the intensive care unit | 24
respiratory failure | 24
invasive mechanical ventilation support | 24
septic shock | 24
multiple organ failure syndrome | 24
neurological compromise | 24
progression to stupor | 24
presence of signs of systemic inflammatory response | 24
described pulmonary findings | 24
history of immunosuppression | 24
risk of infection by opportunistic germs | 24
empirical antibiotic treatment | 24
piperacillin/tazobactam | 24
vancomycin | 24
clarithromycin | 24
fluconazole | 24
oseltamivir | 24
assessed by the Department of Infectious Diseases | 48
rule out infection due to Histoplasma | 48
rule out infection due to Cryptococcus | 48
rule out infection due to Aspergillus | 48
urinary antigen testing for Histoplasma | 48
urinary antigen testing for Cryptococcus | 48
bronchoalveolar lavage galactomannan test | 48
tests were negative | 48
liposomal amphotericin B initiated | 96
suspicion of opportunistic fungal infection | 96
recent history of positive viral load for cytomegalovirus | 48
ganciclovir initiated | 48
viral load for cytomegalovirus undetectable | 384
reports of viral load for cytomegalovirus showed reactivity | 48
decreasing loads | 48
cytomegalovirus infection not considered the cause | 48
blood cultures | 48
oral tracheal secretion cultures for common aerobic germs | 48
cultures were negative | 48
suspending sedation | 48
patient persisted with an altered state of consciousness | 48
brain tomography performed | 48
intra-axial lesion with expansive behaviour | 48
ring enhancement | 48
associated vasogenic oedema | 48
right anterior subinsular vasogenic oedema | 48
lesions identified as foci of cerebritis | 48
open biopsy performed | 48
subcortical mass with lumpy consistency | 48
yellowish mass | 48
partially vascularised | 48
without cleavage planes | 48
suggestive of a secondary tumour | 48
no purulent material | 48
no signs of cerebritis | 48
samples taken for microbiological studies | 48
samples taken for histopathological studies | 48
histopathological studies not conclusive | 48
fresh examination of samples | 48
presence of large, irregular, septate and dematiaceous hyphae | 48
optimizing antifungal management | 48
amphotericin B | 48
voriconazole | 48
treatment extended for 42 days | 48
subsequent treatment with voriconazole for 6 months to 1 year | 48
patient's condition improved | 48
ventilation support discontinued | 48
alertness restored | 48
Sabouraud agar growth | 72
grey-white colonies | 72
colour turned to greenish black | 72
dark brown colour on the back of the colony | 72
strain sent for identification | 72
septate dematiaceous hyphae | 72
septate conidiophores | 72
microbiological typing concluded phaeohyphomycosis | 72
disseminated by Alternaria spp. | 72
MRI scan on day 5 | 120
collection on the surgical bed | 120
persistence of oedema in the right subinsular region | 120
excision of the lesion not radical | 120
optimise dematiaceous treatment | 120
inclusion of terbinafine treatment | 120
satisfactory progress | 120
no evidence of new neurological deficits | 120
subsequent CT scans showed no significant changes | 120
no progression of mycosis | 120
no other organs compromised | 120
patient dies | 2928
death cause other than fungal infection | 2928
