21 years old | 0
male | 0
allergic to cefuroxime | 0
allergic to metronidazole | 0
admitted to the hospital | 0
sore throat | -96
shortness of breath | -96
left tonsillitis | -96
septic shock | 0
transferred to the Intensive Care Unit | 0
fever | -96
poor oral intake | -96
low-grade temperature of 37.6°C | 0
bilateral lower zone infiltrates | 0
bilateral pleural effusion | 0
respiratory failure | 0
intubated | 0
doxycycline | 0
clindamycin | 0
vancomycin | 0
antibiotics upgraded to meropenem | 24
antibiotics upgraded to doxycycline | 24
throat swab negative | 24
urine culture negative | 24
sputum culture negative | 24
endotracheal aspirates for influenza negative | 24
endotracheal aspirates for other viruses negative | 24
blood culture yielded Fusobacterium necrophorum | 48
Fusobacterium necrophorum sensitive to metronidazole | 48
Fusobacterium necrophorum minimal inhibitory concentration of clindamycin 0.12 μg/mL | 48
meropenem alone | 48
persistent leukocytosis | 120
neck pain | 120
computed tomography of neck and thorax | 144
left internal jugular thrombophlebitis | 144
multiple cavitating lung nodules | 144
distal thromboembolism | 144
Lemierre's syndrome | 144
right internal jugular vein patent | 144
left brachiocephalic vein patent | 144
superior vena cava patent | 144
continue antibiotics | 144
no internal jugular vein ligation | 144
discharged to general ward | 168
intravenous amoxicillin-clavulanate | 168
antibiotic desensitization protocol | 168
satisfactory progress | 240
discharged home | 240
oral amoxicillin-clavulanate | 240
no anticoagulation | 240
follow-up with chest X-ray | 336
resolution of lung infiltrates | 336
antibiotic stopped | 432