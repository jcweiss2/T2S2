53 years old | 0
female | 0
Caucasian | 0
admitted to the hospital | 0
myeloablative allogeneic hematopoietic cell transplant | -7920
relapsing acute lymphoblastic leukaemia | -8760
CAR-T therapy | -264
cyclophosphamide | -264
fludarabine | -264
grade 1 CRS | -168
tocilizumab | -168
methylprednisolone | -168
levetiracetam | -168
fevers | -168
Escherichia coli bacteraemia | -168
admitted to the ward | -168
pancytopenia | -168
new fevers | -120
dyspnoea | -120
hypoxemia | -120
CT imaging of the chest | -120
consolidations in the right upper, right middle and left upper lobes | -120
vancomycin-resistant enterococcal bacteraemia | -120
foscarnet | -120
pentamidine | -120
isavuconazole | -120
levofloxacin | -120
meropenem | -120
linezolid | -120
restlessness | -96
agitation | -96
obtundation | -96
intubation | -96
ICU transfer | -96
basic metabolic panel | -96
mild elevation of the total bilirubin | -96
minor increased international normalised ratio | -96
normal kidney function | -96
blood urea nitrogen | -96
complete blood count | -96
pancytopenia | -96
encephalopathy workup | -96
thyroid-stimulating hormone | -96
vitamin B1 | -96
vitamin B12 | -96
electroencephalogram | -96
head CT | -96
lumbar puncture | -96
ammonia level | -96
391 µmol/L | -96
doxycycline | -72
lactulose | -72
methylprednisolone | -72
ICU day #1 | -72
bronchoscopy | -72
bronchoalveolar lavage | -72
bacterial, fungal and viral cultures | -72
PCR | -72
staining | -72
Ureaplasma PCR | -72
ammonia rose to 643 µmol/L | -48
electroencephalography | -48
epileptiform activity | -48
benzodiazepine infusion | -48
levetiracetam | -48
lacosamide | -48
propofol infusion | -48
pentobarbital | -48
status epilepticus | -48
CT imaging of the head | -48
mildly diminished gray–white differentiation | -48
cerebral oedema | -48
renal replacement therapy | -48
ammonia clearance | -48
meropenem | -48
ceftazidime/avibactam | -48
amphotericin B | -48
acyclovir | -48
genetics consult | -24
hyperammonemia | -24
inborn errors of metabolism | -24
urine organic acids | -24
urine orotic acid | -24
plasma amino acids | -24
plasma acylcarnitine levels | -24
dextrose | -24
levocarnitine | -24
arginine infusion | -24
sodium phenylbutyrate | -24
MRI of the brain | 0
diffuse worsening of the cerebral oedema | 0
Ureaplasma PCR | 0
levofloxacin | 0
withdraw care | 24
death | 24