61 years old | 0
male | 0
White | 0
admitted to the hospital | 0
long-standing arterial hypertension | -8760
severe heart failure | -8760
left ventricular ejection fraction of 30% | -8760
pharmacological treatment with carvedilol | -8760
pharmacological treatment with ivabradine | -8760
pharmacological treatment with losartan | -8760
stage IIIB chronic renal failure | -8760
no dialysis therapy | -8760
urinary symptoms | -8760
fever | -8760
diaphoresis | -8760
low back pain | -8760
hypotension | -8760
dyspnea | -8760
increased acute phase reactants | -8760
sepsis of urinary origin | -8760
hospitalization in the intensive care unit | -8760
multidisciplinary treatment | -8760
alterations in calcium behavior | -8760
severe hyperparathyroidism | -8760
functional adenoma in the lower left parathyroid | -8760
surgery for parathyroid adenoma | -8760
control of symptoms and levels of calcium and phosphorus | -8760
chest x-ray showed 2 lesions of tumor aspect with internal lytic areas | -24
lesions in the fourth right and eighth left costal arches | -24
first lesion measured 25 × 21 mm | -24
second lesion measured 77 × 54 mm | -24
growth toward the left pleural cavity | -24
physical examination | 0
thin patient with chronic disease | 0
deformity in the neck with anterior flexion | 0
severe dorsal kyphoscoliosis | 0
secondary asymmetry of the right ribcage | 0
retracted right ribcage | 0
decreased intercostal spaces | 0
increased dyspnea with the activities of daily life | 0
NYHA functional class III | 0
blood pressure 120/70 mm Hg | 0
heart rate 100 beats per minute | 0
breathing frequency 16 breaths per minute | 0
no cyanosis | 0
jugular engorgement at 90° | 0
no neck masses | 0
tachycardic rhythmic heart | 0
no murmurs or gallop | 0
decreased breath sounds at both lung bases | 0
abdomen without ascites or masses | 0
extremities with edema grade II | 0
no identifiable lesions in the chest wall | 0
blood work | 0
mild anemia of normal volumes | 0
spirometry showed a moderate restrictive ventilatory pattern | 0
no significant post-bronchodilator changes | 0
diffusing capacity of carbon monoxide in normal limits | 0
chronic kidney disease was stable | 0
thoracic computed tomography scan | 0
heterogeneous rounded lytic lesion | 0
sclerotic edges | 0
growth toward the pulmonary cavity | 0
expansive type | 0
displacement of pulmonary parenchyma | 0
severe dorsal kyphoscoliosis | 0
hospitalization in the intensive care unit for pre-surgical conditioning | -24
left ventricular ejection fraction of 30% | -24
cycle of intravenous levosimendan | -24
red blood cell transfusion | -24
resection of the left costal mass by thoracoscopy | 0
involvement of the eighth rib and soft tissues of the seventh to ninth left ribs | 0
no infiltration into the lung tissue or pleural cavity | 0
partial resection of the three ribs | 0
no pulmonary lobectomy | 0
difficult evolution in the immediate postsurgical period | 24
hemodynamic instability | 24
vasoactive support with norepinephrine | 24
prolonged mechanical ventilation | 24
need for a tracheostomy | 24
long-standing recovery process | 24
removal of vasoactive drugs | 168
invasive ventilatory support | 168
tracheostomy | 168
complete physical and respiratory rehabilitation | 168
pathology reported morphological findings compatible with ossifying lipoma | 168
histological sections showed a benign neoplastic lesion | 168
mature adipose tissue | 168
thin capsule of fibroconective tissue | 168
proliferation of thin bone trabeculae | 168
no Medullary stroma | 168
no other mesenchymal tissues within the mass | 168
discussion with the patient and his family | 168
no chemotherapeutic treatment or other specific oncological interventions | 168
benign nature of the mass | 168
post excisional curative potential | 168
frequent control with several medical specialties | 168
no evidence of recurrence of the lesions | 720