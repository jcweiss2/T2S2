46 years old | 0\
male | 0\
arterial hypertension | -672\
obesity | -672\
admitted to the hospital | 0\
fever | 0\
hypotension | 0\
asthenia | 0\
COVID-19 infection | -336\
rhinitis | -336\
mild cough | -336\
alert | 0\
oriented | 0\
cooperative | 0\
asthenic | 0\
blood pressure 85/55 mmHg | 0\
heart rate 120 bpm | 0\
arterial oxygen saturation 85% | 0\
body temperature 38.3 C° | 0\
femoral central venous catheter | 0\
sinus tachycardia | 0\
diffuse low voltages | 0\
absence of significant repolarization abnormalities | 0\
neutrophilic leukocytosis | 0\
C-reactive protein elevation | 0\
Procalcitonin elevation | 0\
elevated high sensitivity Troponin | 0\
elevated brain natriuretic peptide | 0\
elevated creatinine | 0\
elevated transaminases | 0\
elevated total bilirubin | 0\
COVID-19 IgM antibody test positive | 0\
normal left ventricular cavitary dimensions | 0\
diffuse LV parietal thickening | 0\
severely reduced LV global systolic function | 0\
grade II LV diastolic dysfunction | 0\
normal cavitary dimensions | 0\
reduced global right ventricular systolic function | 0\
dilated inferior vena cava | 0\
right ventricular systolic pressure 41 mmHg | 0\
absence of hemodynamically significant valvulopathy | 0\
slight pericardial effusion | 0\
blood cultures | 0\
broad-spectrum antibiotic therapy | 0\
crystalloid hydration | 0\
nasal cannula ventilatory therapy | 0\
norepinephrine | 0\
poor hemodynamic response | 0\
levosimendan | 0\
BP 100/60 mmHg | 12\
heart rate 110 bpm | 12\
BP 125/70 mmHg | 24\
heart rate 95 bpm | 24\
diuresis 1800 ml | 24\
improvement of systolic performance indices | 12\
improvement of systolic performance indices | 24\
LV EF 66% | 24\
dP/dT ratio 1275 mmHg/sec | 24\
TAPSE 23 mm | 24\
tricuspid S-wave velocity at TDI 11.2 cm/sec | 24\
SVi 27 ml/m2 | 24\
CI 2.5 l/min/m2 | 24\
LV diastolic function normal | 24\
IVC diameter 18 mm | 24\
IVC collapse 100% | 24\
RVSP 28 mmHg | 24\
cardiac magnetic resonance imaging | 24\
endomyocardial biopsy | 48\
lymphocytic myocarditis | 48\
coronary arteriography | 48\
normal coronary circulation | 48\
discharged | 504\
TTE normal findings | 744\
TTE normal findings | 1008