70 years old | 0
    male | 0
    admitted to the intensive care unit | 0
    bullous pemphigoid | 0
    sepsis | 0
    fundus fluorescein angiography | -1440
    senile macular degeneration | -1440
    fluorescein extravasation | -1440
    pruritus | -1440
    erythema | -1440
    essential hypertension | 0
    glaucoma | 0
    senile macular degeneration | 0
    oral metoprolol 50 mg | 0
    oral aspirin 100 mg | 0
    brimonidine tartrate 0.2% | 0
    allergy to human albumin solution | -131400
    bypass surgery | -131400
    erythematous patches on scalp | 0
    erythematous patches on chest | 0
    erythematous patches on anogenital region | 0
    vesicles | 0
    tense bullae | 0
    daily oral methylprednisolone 48 mg | 0
    topical clobetasol dipropionate 0.05% cream | 0
    topical 4% urea lotion | 0
    relative eosinophilia | 0
    punch biopsies | 0
    subepidermal blistering | 0
    dermal infiltrates of mononuclear cells | 0
    dermal infiltrates of eosinophils | 0
    focal areas of collagen flame figures | 0
    direct immunofluorescence linear reactivity for C3c | 0
    direct immunofluorescence linear reactivity for IgG | 0
    salt extraction testing consistent with bullous pemphigoid | 0
    regression of lesions | 144
    daily oral azathioprine 150 mg | 144
    resolution of all lesions | 144
    discharged | 144
    oral methylprednisolone 40 mg | 144
    topical 4% urea lotion | 144
    oral azathioprine 150 mg daily | 144
    admitted to the ICU | 720
    sepsis secondary to urinary tract infection | 720
    decreased immune response | 720
    died from cardiac failure | 984
    