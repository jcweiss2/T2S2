61 years old | 0
African-Canadian | 0
woman | 0
admitted to the hospital | 0
fever | 0
dyspnea | 0
pneumonia | 0
chronic kidney disease | -168
previous pyoderma gangrenosum | -168
left above-knee amputation | -168
diabetes mellitus | -168
hypertension | -168
osteoarthritis | -168
sarcoidosis | -168
deteriorated kidney function | -168
permanent hemodialysis catheter insertion | -168
hemodialysis started | -168
discharged | -168
presented with diarrhea | -168
presented with vomiting | -168
blood pressure 157/79 mm Hg | 0
heart rate 97 beats per minute | 0
respiratory rate 20 breaths per minute | 0
temperature 38.3°C | 0
oxygen saturation 98% on room air | 0
purulent discharge around catheter exit site | 0
redness around catheter exit site |5 0
induration along the tunnel | 0
redness along the tunnel | 0
tenderness along the tunnel | 0
admitted with dialysis catheter tunnel infection diagnosis | 0
central blood samples sent for cultures | 0
peripheral blood samples sent for cultures | 0
swab from purulent discharge around catheter exit site sent for cultures | 0
received intravenous cloxacillin 2 g every 6 hours | 0
received vancomycin 15 mg/kg bolus | 0
subsequent vancomycin doses targeting 15 to 20 mg/L trough levels | 0
catheter removed | 0
catheter tip sent for culture | 0
transthoracic echocardiogram showed no valvular vegetations | 0
continued high-grade fever | 168
leukocytosis | 168
swelling at catheter tunnel exit site expanded | 168
ulcerated with multiple points of purulent discharge over 5 cm × 5 cm area | 168
small collection at clavicle lanced | 168
1 to 2 mL pus expressed | 168
new painful nodular lesion developed on abdominal wall | 168
lesion at site of subcutaneous low-molecular-weight heparin injections | 168
ulcerated | 168
blood cultures repeated multiple times | 168
negative blood cultures | 168
negative catheter tip culture | 168
negative swab from exit site | 168
negative pus from clavicular collection | 168
negative swabs from abdominal ulcer | 168
stool enteric cultures negative | 168
clostridium difficile toxin negative | 168
urine culture negative | 168
surgical review requested | 168
lesions deemed too small for incision and drainage | 168
antibiotic coverage broadened on third day | 72
intravenous piperacillin/tazobactam 2.25 g every 8 hours | 72
vancomycin continued | 72
clinical diagnosis of pyoderma gangrenosum entertained on seventh day | 168
consultation with rheumatology | 168
decision to avoid biopsy | 168
insertion of new dialysis line deferred | 168
diuretics maximized | 168
stable without dialysis for 11 days | 168
initiation of steroids delayed | 168
concerns of ongoing infection | 168
not taking maintenance steroids for sarcoid | 168
developed hemodynamic instability on eighth day | 192
blood pressure 94/39 mm Hg | 192
acute alteration of mental status | 192
C-reactive protein 335 mg/L | 192
leukocyte count 28.7 × 109/L | 192
normal serum lactate | 192
resuscitated with intravenous fluids | 192
transferred to intensive care unit | 192
computed tomography of chest, abdomen, and pelvis with intravenous contrast | 192
left lower lobe consolidation | 192
mediastinal lymphadenopathy | 192
no other pathology | 192
treated with intravenous hydrocortisone 50 mg every 6 hours | 192
antibiotics continued unchanged | 192
no hemodynamic or ventilatory support required | 192
fever resolved within 2 days of steroid initiation | 216
pain at lesion sites markedly improved | 216
new tunneled dialysis line inserted | 216
hemodialysis resumed | 216
intravenous hydrocortisone changed to oral prednisone 50 mg/day | 216
piperacillin/tazobactam stopped | 216
vancomycin continued for total of 4 weeks | 216
discharged after 4 weeks of hospitalization | 672
discharge medications included oral prednisone 50 mg daily | 672
discharge medications included hydroxychloroquine 200 mg twice a day | 672
skin ulceration continued to improve | 1344
ulcers almost completely healed after 2 months | 1344
