69 years old | 0
male | 0
admitted to the hospital | 0
coronary artery disease | -672
aspirin | -672
hypertension | -672
type 2 diabetes mellitus | -672
fever | -168
malaise | -168
shortness of breath | -168
temperature of 103.1 °F | 0
pulse of 106 beats per minute | 0
respiratory rate of 18 per minute | 0
blood pressure of 142/70 mm Hg | 0
saturation of 89% on room air | 0
decreased breath sounds bilaterally at base with crepitations | 0
hemoglobin 12.7 g/dL | 0
white blood cell count of 4.5 × 103 | 0
platelet count of 164 × 103 | 0
neutrophil 76.4% | 0
lymphocyte 14.9% | 0
absolute lymphocytes 0.7 | 0
C-reactive protein (CRP) 12.07 mg/dL | 0
D-dimer 570 ng/mL | 0
influenza A and B serology was negative | 0
COVID-19 RT-PCR was positive | 0
bilateral infiltrates at the lung bases | 0
hydroxychloroquine | 0
azithromycin | 0
supplemental oxygen with nasal cannula | 0
prophylactic enoxaparin | 0
worsening of bilateral infiltrates | 24
optiflow (100% FiO2 at 55 L/min) | 24
elevated D-dimer to 1,763 ng/mL | 48
therapeutic enoxaparin | 48
abdominal pain | 480
hypovolemic shock | 480
hemoglobin level of 8.9 g/dL | 480
computed tomography (CT) scan of the abdomen and pelvis | 480
hemorrhage along entire length of right psoas muscle | 480
transferred to intensive care unit (ICU) | 480
resuscitated with 2 L intravenous fluid | 480
3 units of packed red blood cells (PRBC) | 480
vasopressors | 480
post-transfusion hemoglobin of 6.6 g/dL | 480
two more units of PRBC | 480
1 unit of fresh frozen plasma | 480
arterial embolization | 480
left common femoral artery accessed | 480
abdominal aortogram | 480
subtle extravasation from branches of the right L3 and L4 lumbar arteries | 480
selectively catheterized with a 5 French Mickelson catheter | 480
high flow microcatheter placed | 480
active extravasation identified | 480
Embosphere particles administered | 480
microcoils placed | 480
no active contrast extravasation identified | 480
one more unit of PRBC | 480
hemoglobin stabilized to 7.9 g/dL | 480
vasopressor requirement decreased | 480
vasopressor requirement discontinued | 480
repeat CT scan showed decreased size of hematoma | 504
weaned off optiflow | 504
transferred to the medical floors | 504