70 years old | 0
male | 0
admitted to the ICU | 0
BP | 0
sepsis | 0
fundus fluorescein angiography | -144
senile macular degeneration | -144
fluorescein extravasation | -144
pruritus | -144
erythema | -144
essential hypertension | 0
glaucoma | 0
senile macular degeneration | 0
oral metoprolol | 0
oral aspirin | 0
brimonidine tartrate | 0
allergy to human albumin solution | -13140
bypass surgery | -13140
erythematous patches | 0
vesicles | 0
tense bullae | 0
methylprednisolone | 0
clobetasol dipropionate | 0
topical 4% urea lotion | 0
relative eosinophilia | 0
punch biopsies | 0
subepidermal blistering | 0
dermal infiltrates | 0
eosinophils | 0
collagen flame figures | 0
direct immunofluorescence | 0
linear reactivity for C3c | 0
linear reactivity for IgG | 0
salt extraction testing | 0
regression of lesions | 144
oral azathioprine | 144
resolution of lesions | 240
discharged | 240
sepsis secondary to urinary tract infection | 720
decreased immune response | 720
cardiac failure | 888
died | 888