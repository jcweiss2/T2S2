17 years old | 0
male | 0
admitted to the hospital | 0
shortness of breath | -2
pleuritic chest pain | -2
dry cough | -720
fatigue | -720
weight loss | -720
fever | -24
chills | -24
pleuritic chest pain worsened | -2
shortness of breath worsened | -2
cardiac tamponade | 6
pericardiocentesis | 6
pus-like fluid drained | 6
intravenous ceftriaxone | 0
Mycobacterium tuberculosis polymerase chain reaction (TB PCR) test positive | 24
isoniazid | 24
rifampin | 24
ethambutol | 24
pyrazinamide | 24
pyridoxine | 24
yeast growth in pericardial fluid culture | 72
intravenous fluconazole | 72
Candida parapsilosis identified | 96
fever persisted | 96
gram-positive bacterium growth in pericardial fluid culture | 96
vancomycin | 96
ciprofloxacin | 96
pneumopericardium | 168
vancomycin and ciprofloxacin switched to vancomycin and ertapenem | 168
Peptostreptococcus asaccharolyticus identified | 216
Streptococcus anginosus identified | 216
Methicillin-sensitive Staphylococcus aureus identified | 216
Prevotella oralis identified | 216
pericardiectomy | 240
pus and inflammatory material observed | 240
irrigation with suction and removal of septations | 240
pericardial tissue biopsy | 240
acute and chronic inflammation with liquefactive necrosis | 240
discharged | 720
oral antifungal | 720
antibiotic | 720
anti-TB medication | 720
amoxicillin/clavulanic acid stopped | 2160
fluconazole stopped | 4320
anti-TB medication continued | 4320
returned to normal activity | 4320
heart rate around 70 beats/min | 4320
echocardiography showed no cardiac relaxation abnormality | 4320
ejection fraction minimally decreased | 4320