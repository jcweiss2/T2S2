67 years old | 0
    male | 0
    cardiogenic cerebral infarction | -672
    visited hospital | 0
    chills | 0
    right chest pain | 0
    daily exercise | -672
    no tobacco use | -672
    no excessive alcohol use | -672
    no subsequent comorbidities of cerebral infarction | -672
    body temperature 36.4°C | 0
    blood pressure 82/66 mmHg | 0
    pulse rate 110/min | 0
    oxygen saturation 90% | 0
    respiratory rate 30 breaths/min | 0
    right coarse crackles | 0
    white blood cell count 9500/μl | 0
    neutrophils 7695/μl | 0
    platelets 165,000/μl | 0
    C-reactive protein 2.59 mg/dl | 0
    chest radiograph right S2-infiltrate | 0
    chest computed tomography right S2-infiltrate | 0
    systemic blood pressure declined to 60 mmHg | 2
    oxygen saturation decreased to 70% | 2
    transferred to ICU | 2
    mechanical ventilation support | 2
    oxygenation not fully recovered | 2
    bronchoscopy large amount of bleeding (>1000 ml) | 2
    right upper bronchus bleeding | 2
    B6 segments obstruction | 2
    repetitive chest radiograph complete opacification right hemithorax | 2
    repetitive chest CT complete opacification right hemithorax | 2
    veno8-venous ECMO introduced | 2
    P. aeruginosa identified bronchial secretion | 2
    P. aeruginosa identified blood | 2
    meropenem | 2
    ciprofloxacin | 2
    withdrawal of v-v ECMO | 336
    abscess formation right lung | 336
    P. aeruginosa empyema | 336
    purulent sputum | 336
    minor bleeding right lung | 336
    right pneumonectomy | 336
    pleural lavage | 336
    discharged from ICU | 2208
    home whirlpool bath use | -672
    P. aeruginosa in whirlpool bathtub | -672
    exoS gene-positive P. aeruginosa | -672
    virulent P. aeruginosa strain exposure | -672
    fulminant pneumonia | 0
    sepsis recovery | 336
    vital signs improved | 336
    unaffected left lung competent | 336
    surgical intervention | 336
    infection resolution | 2208
    patient's wife no pneumonia | -672
    wife immunocompromised | -672
    wife no jet bath use | -672
    bathroom dry and clean | -672
    black mud emitted jet system | -672
    genomic analysis P. aeruginosa | 336
    MLST ST-900 | 336
    drug resistance genes | 336
    virulent factor exoS | 336
    life-threatening pneumonia | 0
    surgical resection therapeutic option | 336
    contaminated aerosol inhalation | -672
    severe bacterial pneumonia | 0
    intensive management | 2
    antimicrobial therapy | 2
    lung abscess prolonged | 336
    purulent sputum damage left lung | 336
    right lung resection | 336
    sepsis resolved | 336
    P. aeruginosa infection resolved | 2208
    discharge | 2208
    