34 years old | 0
female | 0
gravid 2 | 0
para 1 | 0
previous uncomplicated normal vaginal delivery | 0
ITP | 0
anemia | 0
suspected hypoplastic anemia | 0
received blood transfusion | 0
on iron supplement | 0
denies smoking | 0
denies alcohol intake | 0
admitted to hospital | 0
threatened preterm labor | 0
delivery plan | 0
low hemoglobin level | 0
low platelet count | 0
hematologist ordered 2 units of blood | 0
IVIG at a dose of 0.5 g/kg/day for 4 days | 0
hemoglobin level increased | -6
hemoglobin level dropped | 0
platelet count remained | 0
Hgb 8.6 g/dl | -24
platelet 25 × 10^3/μl | -24
diagnosis of intrauterine growth retardation | -24
counseled regarding mode of delivery | -24
avoidance of operative vaginal delivery | -24
opted for an elective cesarean section | -24
scheduled at 36 weeks of gestation | -24
no amniocentesis | -24
RCOG guideline recommends antenatal corticosteroids | -24
dexamethasone tablets administered orally | -12
last dose completed | -3.5
baby girl born | 0
born at 36 weeks of gestation | 0
weight 2235 g | 0
1-min Apgar score 9 | 0
5-min Apgar score 10 | 0
mild grunting | 1
incubator care with supplemental oxygen | 1
admitted to neonatal ward | 6
mild respiratory distress | 6
mild grunting and retraction | 6
oxygen saturation 94-95% | 6
respiratory rate 64/min | 6
temperature 36.6 °C | 6
heart rate 148/min | 6
blood pressure 65/35 mmHg | 6
suspected to have Transient Tachypnea of Newborn | 6
nasal cannula 2 L flow/min in room air | 6
weaned and discontinued on the third day | 72
neonatal jaundice | 48
phototherapy for two days | 48
feeding started | 48
gradually increased to full feed | 72
discharged home | 96
chest X-ray showed features suggestive of TTN | 24
complete blood counts and serum electrolytes were normal | 8
blood culture was negative | 8