32 years old | 0
    male | 0
    pneumonia | 0
    sepsis | 0
    shifted to intensive care unit (ICU) | 0
    replaced PVC ETT with Portex Blue Line SACETT™ | 0
    sudden desaturation | 48
    audible leak around ETT | 48
    ventilator disconnection alarm | 48
    decreased expiratory tidal volume | 48
    pilot balloon deflated | 48
    inability to inflate pilot balloon | 48
    suspected ETT cuff rupture | 48
    exchanged ETT over tube exchange catheter | 48
    inflation line disconnection found | 48
    adhesive tape fixation of inflation line | 48
    evaluation of possible causes | 48
    ruled out patient pulling inflation line | 48
    intact inflation line length | 48
    no stretching features | 48
    suspected adhesive tape issue | 48
    insertion sites at 21 and 22 cm marks | 48
    ETT fixation at oral level | 48
    suggestion to move insertion sites above 24 cm | 48
    possible manufacturing defect | 48
    inadequate bonding solvent use | 48
    lack of standards for inflation line attachment | 48
    recommendation for peruse test | 48
    <|eot_id|>
    