57 years old | 0
male | 0
diagnosed with lepromatous leprosy | -672
treatment with rifampicin/clofazimine/dapsone | -672
abdominal distension | 0
constipation | 0
vomiting | 0
10-kg weight loss | 0
peripheral lymphadenopathy | 0
distended abdomen | 0
positive shifting dullness | 0
computed tomography scan of abdomen | 0
mural thickening of terminal ileum | 0
enlarged mesenteric lymph nodes | 0
mesenteric fat stranding | 0
intra-abdominal free fluid | 0
abdominal paracentesis | 0
atypically large lymphocytes | 0
flow cytometry | 0
abnormal CD4/CD8 double-negative T-cell population | 0
cervical lymph node biopsy | 0
high-grade peripheral T-cell lymphoma | 0
bone marrow examination | 0
stage IV lymphoma | 0
started on dexamethasone | 0
transfer to ICU | 0
severe sepsis | 0
antibiotics and antifungals | 0
ICU care | 24
transfer to national cancer center | 168
commenced on EPOCH chemotherapy | 168
CNS prophylaxis | 168
complete metabolic remission | 672
febrile neutropenia episodes | 336
recurrent bacteremia | 336
generalized weakness | 0
decreased power in muscles | 0
neurological team involvement | 0
neurophysiological electromyogram/nerve conduction study | 0
repetitive nerve stimulation | 0
presynaptic neuromuscular junction disorder | 0
VGCC antibodies requested | 0
started on intravenous immunoglobulins | 0
significant improvement of motor function | 24
planned for autologous bone marrow transplant | 0
re-admitted to medical ICU | 0
severe sepsis and multiorgan failure | 0
passed away | 4320