77 years old | 0
male | 0
benign prostatic hyperplasia | 0
nocturia | 0
increased frequency | 0
hypertension | 0
fatty liver | 0
hemiparesis | -2160
acute infarction of the basal ganglia | -2160
cilostazol | -336
discontinued cilostazol | -336
no history of general anesthesia | 0
no family history of MH | 0
normal laboratory tests | 0
normal chest X-ray examination | 0
normal electrocardiography | 0
normal pulmonary function testing | 0
ejection fraction of 60.4% | 0
mild to moderate aortic regurgitation | 0
mild aortic stenosis | 0
mild concentric left ventricular hypertrophy | 0
antihypertensive medication stopped | -12
stable vital signs | -12
general anesthesia induced | 0
propofol administered | 0
rocuronium administered | 0
remifentanil administered | 0
laryngeal mask airway insertion | 0
sevoflurane administered | 0
mechanical ventilation | 0
constant tidal volume of 400 mL | 0
respiratory rate of 12 breaths/minute | 0
blood pressure 114/63 mmHg | 0
heart rate 60 beats/minute | 0
oxygen saturation 99% | 0
EtCO2 30 mmHg | 0
bispectral index 30 | 0
total anesthesia time 85 minutes | 0
vital signs before end of anesthesia | 85
blood pressure 180/90 mmHg | 85
heart rate 89 beats/minute | 85
body temperature 37.8°C | 85
oxygen saturation 99% | 85
EtCO2 31 mmHg | 85
shivering | 95
severe anxiety | 95
pethidine administered | 95
fentanyl administered | 95
mental status deteriorated | 95
masseter muscle rigidity | 95
muscle rigidity of both arms | 95
sudden hyperventilation | 95
oxygen mask | 95
blood pressure 220/168 mmHg | 95
heart rate 134 beats/minute | 95
respiratory rate 30 breaths/minute | 95
body temperature 38.1°C | 95
oxygen saturation 98% | 95
suspected MH | 105
increased body temperature | 105
worsening masseter muscle rigidity | 105
MH clinical classification score 53 points | 105
diagnosis of MH | 105
aggressive cooling | 105
esmolol administered | 105
arterial blood gas analysis | 105
compensated metabolic acidosis | 105
pH 7.35 | 105
PaCO2 33 mmHg | 105
PaO2 79 mmHg | 105
bicarbonate 18.2 mmol/L | 105
follow-up biochemical tests | 105
increased CPK | 105
increased LDH | 105
increased myoglobin | 105
dantrolene sodium administered | 115
body temperature decreased | 115
systemic muscle rigidity disappeared | 115
entry into intensive care unit | 120
consciousness restored | 120
no remnant muscle rigidity | 120
general weakness | 120
stable respiratory pattern | 120
body temperature maintained | 120
urinalysis | 120
myoglobinuria not confirmed | 120
mild fever | 144
pulmonary edema | 144
white blood cell count 28,700/µL | 144
hemoglobin concentration 10.3 g/dL | 144
hematocrit 31% | 144
platelet count 74,000/µL | 144
C-reactive protein concentration 10.51 mg/dL | 144
arterial blood gas analysis | 144
pH 7.48 | 144
PaCO2 28 mmHg | 144
PaO2 66 mmHg | 144
bicarbonate concentration 20.9 mmol/L | 144
oxygen saturation 94% | 144
antibiotics started | 144
body temperature varied | 168
renal function testing | 168
improvement in blood urea nitrogen concentration | 168
improvement in creatinine concentration | 168
sanguineous urine | 168
oral diet started | 288
Klebsiella pneumoniae identified | 288
transferred to general ward | 432
discharged | 576
explanation of treatment history | 576
informed of MH recurrence risk | 576