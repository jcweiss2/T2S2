44 years old | 0
male | 0
admitted to the hospital | 0
DWD | -64800
mild acne | -51600
seborrheic distribution | -51600
summertime exacerbations | -51600
systemic retinoids | -64800
sepsis | -14400
Kaposi varicelliform eruption | -14400
local infection episodes | -14400
Staphylococcus aureus | -14400
Morganella morganii | -14400
atypical Mycobacterium cutaneous infection | -7200
widespread erythema | -720
hypertrophic warty keratotic papules | -720
plaques | -720
cysts | -720
nodules | -720
giant comedones | -720
macerations of the skin | -720
severe fetor | -720
leoninelike facies | -720
diffuse palmo-plantar keratoderma | -720
extreme cachexia | -720
tachycardia | -720
keratotic plugs | -720
dyskeratosis | -720
corps ronds | -720
grains | -720
suprabasal clefts | -720
anemia | -720
leukocytosis | -720
hypoalbuminemia | -720
skin cultures positive for S aureus | -720
skin cultures positive for M morganii | -720
skin cultures positive for Streptococcus group G | -720
blood cultures positive for S aureus | -720
fungal infection excluded | -720
HIV serology negative | -720
polymerase chain reaction test results for herpes simplex type 1 and 2 and varicella zoster negative | -720
blood absorption indexes low | -720
neutrophil phagocytosis normal | -720
chemotaxis normal | -720
super oxide production normal | -720
flow cytometry test results unremarkable | -720
computed tomography enterography normal | -720
spinal radiographs normal | -720
chest radiographs normal | -720
transthoracic cardiac echo test normal | -720
genetic test for the 3-base deletion in exon 2 of leucine negative | -720
intravenous broad-spectrum antibiotics | -720
high-dose oral isotretinoin | -720
topical keratolytic therapy | -720
discharged from the department | 0
severe sepsis | 8760
severe hypoglycemia | 8760
widespread erythema | 8760
died | 8762