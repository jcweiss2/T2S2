77 years old | 0
male | 0
admitted to the hospital | 0
unstable angina | -67200
coronary stent insertion | -67200
Sigmart (nicorandil 5 mg) | -67200
aspirin (enteric coated tab, 100 mg) | -67200
Almarl (arotinolol 5 mg) | -67200
Herben (diltiazem 30 mg) | -67200
normal chest X-ray | -24
left ventricular ejection fraction of 61% | -24
grade 2 diastolic dysfunction | -24
mild aortic regurgitation | -24
trivial mitral regurgitation | -24
tricuspid regurgitation | -24
normal blood urea nitrogen/creatinine (BUN/Cr) of 11.0/0.8 mg/dL | -24
low hemoglobin of 11.9 g/dL | -24
aspirin stopped 7 days before surgery | -168
no medication administered on the morning of surgery | -24
blood pressure (BP) of 144/79 mmHg | -24
heart rate (HR) of 68 beats/min | -24
SpO2 of 97% | -24
bupivacaine (0.5%, 10 mg) injected into the subarachnoid space at T10 | -24
intravenous dexmedetomidine infused (0.5 μg/kg/min for first 10 min, then at 0.4-0.6 μg/kg/min) | -24
pneumatic thigh tourniquet applied intraoperatively at 300 mmHg for 100 min | -24
total anesthesia time of 2 hours and 10 minutes | -24
600 mL of crystalloid administered | -24
150 mL of urine collected | -24
estimated blood loss of 90 mL | -24
BP of 100-130/50-70 mmHg | -24
HR of 45-55 beats/min | -24
SpO2 of 97%-99% | -24
BP of 97/55 mmHg | 0
HR of 41 beats/min | 0
SpO2 of 100% | 0
BP of 95-100/55-60 mmHg | 24
HR of 40-45 beats/min | 24
SpO2 of 98%-100% | 24
90 mL of urine | 24
70 mL of blood drained | 24
400 mL of crystalloid administered | 24
intravenous patient-controlled analgesia (AutoFuser) | 24
1 mg fentanyl | 24
baseline infusion rate of 2 mL/h | 24
bolus demand dose of 2 mL | 24
lock-out time of 15 min | 24
antibiotics (Refosporen, 1 g and cefazedone sodium 1 g) injected bid | 24
severe pain on the right thigh | 24
overnight shivering | 24
Tridol Injection (tramadol hydrochloride 50 mg/mL) injected | 24
drowsy mental state | 24
Glasgow coma scale score of 8/15 (M5/V2/E1) | 24
BP of 110/70 mmHg | 24
HR of 122 beats/min | 24
body temperature of 37.9 °C | 24
SpO2 of 86%-90% | 24
normal electrocardiogram | 24
right thigh stiff and dark brown | 24
no swelling | 24
surgical site unaffected | 24
distal extremity unaffected | 24
dark colored urine | 24
urine output every 8 h after operation of 100 mL, 220 mL, 250 mL | 24
total urine output of 570 mL/d | 24
CK increased to 2763 IU/L | 24
CK-MB elevated to 13.26 ng/mL | 24
AST elevated | 24
BUN/Cr elevated | 24
normal troponin-I at 0.100 ng/mL | 24
prolonged coagulation battery | 24
thrombocytopenia | 24
high fibrinogen degradation product | 24
high D-dimer | 24
progressive deterioration of DIC | 24
continued deterioration of laboratory parameters in ICU | 48
mild small vessel disease on brain MRI | 24
no notable hemorrhage | 24
no infarction | 24
serum myoglobin of 1027 ng/mL | 24
urine myoglobin of 25.3 ng/mL | 24
red blood cell count of 100/high powered field (HPF) | 24
tourniquet-induced rhabdomyolysis diagnosed | 24
AKI (AKIN criteria stage 1) | 24
DIC | 24
BP dropped to 88/62 mmHg | 24
norepinephrine (0.5-1 μg/kg/min) infused | 24
admitted to ICU | 24
arterial line placed in left radial artery | 24
central line secured in right internal jugular vein | 24
nephrologist consulted | 24
fluid treatment of 5 L/d prescribed | 24
dialysis scheduled | 24
fluid loading with normal saline at 400 mL/h for 2 h | 24
fluid decreased to 250 mL/h | 24
Lasix (furosemide, 20 mg injection) administered | 24
sodium bicarbonate (40 mL injection of 8.4%) administered | 24
urine output of 110 mL for first 3 h | 24
urine output of 600 mL for next 4 h | 24
Denogan (propacetamol hydrochloride 1 g injection) administered | 24
mental status restored to alert | 24
BP of 90-110/60-70 mmHg | 24
HR of 104 beats/min | 24
body temperature of 36.2 °C | 24
SpO2 of 98% on room air | 24
body temperature elevated to 38.0 °C | 24
BP and HR dropped suddenly | 24
cardiac arrest | 24
cardiopulmonary resuscitation performed for 1 h | 24
resuscitation stopped | 24
patient expired | 24
