69 years old | 0  
    male | 0  
    generalized abdominal pain | -192  
    bilious vomiting | -192  
    obstipation | -96  
    diabetes | 0  
    chronic alcoholism | 0  
    tachycardia | 0  
    abdominal distension | 0  
    generalized tenderness | 0  
    leucocytosis | 0  
    ultrasonography findings | 0  
    CECT findings | 0  
    Rigler's triad | 0  
    exploratory laparotomy | 0  
    gallstone impacted in ileum | 0  
    enterotomy | 0  
    cholecystoduodenal fistula | 0  
    chronic cholecystitis | 0  
    reactive lymphadenitis | 0  
    full diet started | 120  
    suture line healthy | 192  
    left abdominal drain removed | 192  
    right abdominal drain removed | 216  
    respiratory infection | 288  
    shock | 288  
    acute kidney injury | 288  
    intubated | 288  
    ventilated | 288  
    blood transfusions | 288  
    intravenous antibiotics | 288  
    inotropic support | 288  
    electrolyte corrections | 288  
    pneumonia | 504  
    sepsis | 504  
    death | 504