59 years old | 0
male | 0
visited Karachi, Pakistan | -48
began to have a persistent fever | -48
seen in the clinic | -46
prescribed antipyretics | -46
antipyretics failed to improve his fever | -44
continuous, nonprojective vomiting | -44
headaches | -44
no apparent contact with sick individuals | -48
no history of upper respiratory tract infection (URTI) symptoms | -48
no ear problems | -48
no animal contact | -48
no swimming in any local river streams or bathing ponds | -48
admitted to the emergency department | 0
cerebrospinal fluid (CSF) sample was taken | 0
neurology team assessed him | 0
awake, confused and agitated | 0
became drowsy | 1
barely responsive to painful stimuli | 1
no longer protecting his airway | 1
intubated | 1
admitted to the intensive care unit | 1
impression of septic shock secondary to a primary central nervous system infection | 1
laboratory investigations | 1
radiological imaging of the brain | 1
computed tomography (CT) brain angiogram | 1
no evidence of acute intracranial insult | 1
computed tomography angiography (CTA) | 1
no significant stenosis or focal occlusion | 1
CT of the brain without contrast | 1
new onset of diffuse brain oedema | 1
moderate diffuse narrowing of the CSF spaces | 1
scattered hyperattenuating foci in the subarachnoid spaces | 1
leptomeningeal process | 1
infectious disease team was consulted | 2
antimicrobial treatment | 2
physical examination | 2
coma | 2
fixed dilated pupils | 2
vital signs were stable on inotropic support | 2
other examinations were within normal limits | 2
broad antimicrobial coverage of community-acquired meningitis | 2
lumbar puncture | 2
cultures remained negative | 2
CSF sample was preserved for metagenomics-based diagnosis | 2
clinical condition worsened | 4
antimicrobial treatment regimen was modified | 4
technetium-99 m HMPO brain perfusion scan | 72
brain death | 72
passed away | 216
metagenomics-based analytical protocols | 216
retrospective metagenomic sequencing | 216
primary amoebic meningoencephalitis (PAM) | 216
N. fowleri as the aetiological agent | 216
metagenomic next generation sequencing (mNGS)-based protocol | 216
draft assembly of the first N. fowleri clinical isolate genome | 216
Karachi-NF001 | 216