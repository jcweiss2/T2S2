18 years old | 0
male | 0
parkinsonism | -720
diabetes | -720
levodopa | -720
carbidopa | -720
ropinirole | -720
trihexyphenidyl | -720
amantadine | -720
metformin | -720
glipizide | -720
cellulitis | -72
clindamycin | -72
benzylpenicillin | -72
admitted to the hospital | 0
high-temperature spikes | 0
tachycardia | 0
tachypnea | 0
hypotensive | 0
encephalopathic | 0
shifted to ICU | 0
linezolid | 0
piperacillin | 0
tazobactam | 0
inotropic supports | 0
stopped oral hypoglycemic agents | 0
switched to insulin | 0
confused | 0
drowsy | 0
disoriented | 0
altered sensorium | 0
myoclonus | 0
tremors | 0
jerky movements | 0
Computed tomography of the brain | 0
cerebrospinal fluid analysis | 0
improving white blood cell counts | 0
better glycemic control | 0
no other abnormalities | 0
blood and pus cultures | 0
high temperature | 24
altered mental status | 24
myoclonus | 24
jerky movements | 24
tremors | 24
stopped rasagiline | 24
stopped linezolid | 24
temperature settled | 32
normal heart rate | 48
improved sensorium | 48
tremors subsided | 48
shifted out of the ICU | 96
started walking with support | 120
discharged from the hospital | 120
anti-parkinsonism drugs | 120
rasagiline | 120