67 years old | 0
female | 0
admitted to the hospital | 0
fever | -96
chills | -96
cough | -96
dyspnea | -96
diabetes mellitus | -6720
temperature 38.9°C | 0
mildly icteric | 0
bilateral rhonchi | 0
crepitations | 0
no tenderness over the right hypochondrial region | 0
raised white blood cell count | 0
neutrophils 90.2% | 0
hemoglobin level 11.0 g/dL | 0
platelet count 81,000/μL | 0
aspartate aminotransferase level 86 units/L | 0
alanine aminotransferase 78 units/L | 0
bilirubin level high | 0
blood glucose high | 0
acute kidney injury | 0
blood urea nitrogen 24 mg/dL | 0
creatinine 1.7 mg/dL | 0
SPE | 0
multiple peripheral nodules in both lungs | 0
wedge-shaped peripheral lesions | 0
bilateral pleural effusions | 0
mass within the liver | 0
mild tricuspid regurgitation | 0
no vegetations on the heart valves | 0
intravenous imipenem | 0
fever worsened | 24
chills worsened | 24
dyspnea worsened | 24
contrast-enhanced abdominal CT | 24
large liver abscess | 24
no evidence of gas formation | 24
pneumocardia | 24
air within the right ventricle | 24
supine Trendelenburg position | 24
100% oxygen | 24
telemetry unit | 24
liver abscess drained | 48
ultrasonographic guidance | 48
antibiotic treatment continued | 48
symptoms improved | 48
transthoracic echocardiography | 48
no evidence of air within the heart | 48
blood cultures yielded K pneumoniae | 48
pus culture from the liver abscess yielded K pneumoniae | 48
discharged | 600
full recovery | 600
follow-up at 10 months | 7440