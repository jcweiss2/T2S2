39 years old | 0
male | 0
African American | 0
admitted to the emergency department | 0
painful rash | -336
swelling of his eyelids and lips | -336
rash involving his face, scalp, torso, and perianal area | -336
pain moving his bowels | -336
passing bright red blood per rectum | -336
diagnosed with HIV | -336
not compliant with antiretroviral therapy | -336
anal receptive intercourse with men | -336
fever | 0
coalescing vesiculopustular patches | 0
nasal bridge, eyebrows, and scalp were ulcerated | 0
coalescing lesion with crusting and purulent discharge surrounded his anus | 0
rectal exam was refused | 0
electrolytes, blood urea nitrogen, and creatinine were normal | 0
hemoglobin was 5.4 g/dL | 0
leukocytes 5.32 × 10^3/uL | 0
neutrophils 49.1% | 0
lymphocytes 24.1% | 0
eosinophils 2.1% | 0
monocytes 11.5% | 0
basophils 0.4% | 0
absolute CD4 count was 29 cells/uL | 0
liver tests were normal | 0
rectal tissue swab for MPX DNA PCR was positive | 0
HIV viral load was 90,000 | 0
anal, rectal, and oral swab for chlamydia and gonorrhea were negative | 0
IgM for Herpes Simplex 1 and 2, and Herpes 8 were negative | 0
human papilloma virus was not assessed | 0
abdominal computed tomography showed marked circumferential thickening of the rectum | 0
near obliteration of the lumen | 0
pericolonic mesenteric stranding | 0
perianal fistulas extending from the distal rectum to the medial gluteal cleft | 0
started on oral immunotherapy with tecovirimat | 0
started on antiretroviral therapy with Biktarvy | 0
offered MPX vaccine but declined | 0
given polyethylene glycol for constipation | 0
given parenteral opiates for pain | 0
changed to tramadol and gabapentin for pain | 0
transfused two units of blood | 0
discharged to a respite home for recovery | 24
started on AIDS prophylaxis therapies including Bactrim and Azithromycin | 24
readmitted with continued facial swelling, rectal pain, and spreading of his rash | 48
spiking fevers | 48
secondarily infected with Salmonella, Covid19, and MRSA | 48
started on intravenous TPOXX | 48
given smallpox immunoglobulin | 48
commenced on methylprednisolone | 48
developed acute hypoxemic respiratory failure | 72
required intensive care unit admission | 72
commenced on vasopressors | 72
developed cardiac arrest | 96
expired from overwhelming sepsis with multiorgan failure | 120