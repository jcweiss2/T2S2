26 years old | 0
African American | 0
female | 0
hospitalization for possible rheumatic fever | -72
pyrexia | -72
polyserositis | -72
cardiac tamponade | -72
pericardial drainage | -72
pericarditis | -72
abdominal pain | 0
nausea | 0
vomiting | 0
diarrhea | 0
recently quit smoking | -24
family history of mild hypertension | 0
colchicine | 0
lisinopril | 0
omeprazole | 0
pantoprazole | 0
ranitidine | 0
tramadol | 0
penicillin G | 0
albuterol | 0
tachycardia | 0
systolic murmur | 0
severe leukocytosis | 0
low hemoglobin | 0
low serum albumin | 0
normal serum creatinine | 0
proteinuria | 0
severe abdominal and pelvic pain | 0
colitis | 0
mild ascites | 0
sepsis | 0
Clostridium difficile colitis | 0
intravenous metronidazole | 0
intravenous fluids | 0
oral vancomycin | 0
admitted to the transitional intensive care unit | 0
nephrology consultation | 96
oliguric acute tubular necrosis | 96
vasculitis | 96
increased serum creatinine | 96
increased leukocyte count | 96
decreased platelet count | 96
stable hemoglobin | 96
percutaneous renal biopsy | 96
new-onset anemia | 96
hemolytic anemia | 96
schistocytes | 96
elevated lactate dehydrogenase | 96
thrombotic thrombocytopenic purpura | 96
high-dose steroids | 96
daily plasma exchange | 96
ADAMTS13 level | 120
inconclusive ADAMTS13 level | 120
transferred | 312
continued daily plasma exchange | 312
dialysis | 312
mycophenolate mofetil | 312
seizure disorder | 312
levetiracetam | 312
vision loss | 312
bilateral retinal damage | 312
disc, macular, and retinal hemorrhages | 312
vitreous hemorrhage | 312
blindness | 312
discharged | 312
outpatient dialysis | 312
outpatient plasma exchange | 312
follow-up with retinal specialist | 312
bilateral central artery and vein occlusion | 312
eculizumab | 576
improved renal indices | 576
little interdialytic weight gain | 576
increased urinary output | 576
discontinued hemodialysis | 720
discontinued plasma exchange | 720
hypertensive emergency | 912
altered mental status | 912
shortened eculizumab dosing schedule | 912
improved sight | 1092
improved functional status | 1092
walked without assistance | 1092
continued eculizumab | 1092
normal platelet count | 1092
normal hemoglobin | 1092
normal lactate dehydrogenase | 1092
stable serum creatinine | 1092