26 years old | 0
male | 0
admitted to the hospital | 0
spontaneous labor | 0
spontaneous rupture of membranes | -8
respiratory distress | -5
grunting | -5
lethargic | -5
hypoglycemic | -5
blood glucose: 26 mg/dL | -5
oxygen initiated via nasal cannula | -5
intravenous access obtained | -5
ampicillin administration | -5
gentamicin administration | -5
chest X-ray revealed bibasilar infiltrates | -5
severe leukopenia | -5
white blood cell count: 2.3 × 10e9/L | -5
NICU referral | -5
transport team intubated | -5
fluid resuscitation started | -5
progressive respiratory failure | -5
poor perfusion | -5
lactic metabolic acidosis | 0
severe neutropenia | 0
absolute neutrophil count: 500 × 10e9/L | 0
thrombocytopenia | 0
platelet count 111 × 10e9/L | 0
chest radiograph revealed infiltrates | 8
blood culture grew gram-negative rods | 12
lumbar puncture | 12
urinary catheterization | 12
tracheal aspiration | 12
cerebrospinal fluid analysis | 12
normal white blood cell count (17 cells/µL) | 12
elevated red blood cell count (258 cells/µL) | 12
normal protein | 12
normal glucose concentrations | 12
negative Gram's stain | 12
unremarkable urinalysis | 12
tracheal aspirate showed few gram-negative rods | 12
fewer than 25 polymorphonuclear cells | 12
persistent pulmonary hypertension | 0
progressive septic shock | 0
hypotension | 0
poor perfusion | 0
infectious diseases consultation obtained | 0
antibiotics broadened to meropenem | 0
multiple vasoactive medications | 0
inhaled nitric oxide | 0
blood culture revealed P. multocida | 24
tracheal culture revealed P. multocida | 24
cerebral spinal fluid culture negative | 24
urine culture negative | 24
subsequent blood cultures negative | 24
multiple pets in parents' home | 0
maternal vaginal culture positive for P. multocida | 0
molecular diagnostic studies performed | 24
MALDI-TOF mass spectrometry identification | 24
16S rRNA gene sequencing performed | 24
sequences matched P. multocida subspecies septica | 24
maternal vaginal colonization related to pet exposure | 0
mother treated with amoxicillin-clavulanic acid | 24
infant ventilator support weaned | 120
cardiovascular support weaned | 120
hemodynamically stable | 120
respiratory support discontinued | 120
neutropenia resolved | 120
thrombocytopenia worsened | 120
platelet nadir 36 × 10e9/L | 120
transfusion administered | 120
C-reactive protein peak 174 mg/L | 60
antibiotic therapy narrowed to ceftazidime | 168
gentamicin used for synergy | 168
completed 14-day antibiotic course | 336
discharged | 408
infancy without noted morbidities | 408
