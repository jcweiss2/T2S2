21 years old | 0
male | 0
admitted to the hospital | 0
protracted febrile urinary tract infection | -72
no significant medical history | 0
normal physical examination on admission | 0
mild thrombocytopenia | 0
elevated liver enzymes | 0
primary EBV infection | 0
MRI of the kidneys revealed no abnormalities | 0
splenomegaly |*0
multiple smallest inconclusive hepatic lesions | 0
inconclusive MRI of the liver | 0
antibiotic therapy stopped immediately | 0
paracetamol replaced by metamizole | 0
no causative microorganism in urine culture | 0
no causative microorganism in blood culture | 0
liver function decreased dramatically | 96
acute liver failure | 96
acute renal failure | 96
leucopenia | 96
thrombopenia | 96
significantly elevated ferritin level | 96
beginning of severe immune dysregulation | 96
transferred to University Hospital Vienna | 96
genital lesions suggestive of HSV infection | 96
intravenous acyclovir started immediately | 96
patient's condition rapidly deteriorated | 96
multiorgan failure | 96
died | 144
EBV DNA detected by PCR | 120
primary EBV infection confirmed by serology | 120
VCA IgM antibodies detected | 120
VCA IgG antibodies of low avidity detected | 120
HSV1 PCR highly positive | 120
HSV IgG antibody seroconversion confirmed primary HSV1 infection | 120
postmortem analysis of tissues by PCR revealed HSV1 and EBV DNA | 144
high concentrations of HSV1 DNA in liver and spleen tissues | 144
EBV DNA concentration in liver and spleen tissues | 144
histopathology of liver samples displayed HSV hepatitis | 144
confluent necroses in geographical pattern | 144
mixed reactive inflammatory infiltrate | 144
polymorph nuclear leucocytes | 144
hepatocytes with typical nuclear inclusions | 144
immunoperoxidase staining confirmed HSV1 hepatitis | 144
EBV-hepatitis features found | 144
EBV LMP1 detected by alkaline phosphatase staining | 144
EBV DNA extracted from liver tissue | 144
trapping of erythrocytes in portal macrophages | 144
activated Kupffer cells showed erythrophagocytosis | 144
consistent with SHLH | 144
five diagnostic criteria fulfilled | 144
elevated sCD25 level in serum sample | 144
sixth diagnostic criterion fulfilled | 144
multiorgan failure due to SHLH | 144
primary EBV infection | 144
primary HSV1 infection | 144
no mucocutaneous lesions initially | 0
delay in diagnosis and treatment | 0
no bone marrow or spleen histopathology | 144
