57 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
menopausal | 0 | 0 | Factual
admitted to the gynecological emergency unit | 0 | 0 | Factual
left lower quadrant abdominal pain | -1008 | 0 | Factual
pelvic heaviness | -1008 | 0 | Factual
urinary frequency | -1008 | 0 | Factual
past history of 5 miscarriages | 0 | 0 | Factual
tubal ligation | 0 | 0 | Factual
active smoker | 0 | 0 | Factual
no medication | 0 | 0 | Factual
large and painful mass | 0 | 0 | Factual
pelvic MRI | 0 | 0 | Factual
mass measuring 18 × 17 × 12 cm | 0 | 0 | Factual
no lymphadenopathy | 0 | 0 | Factual
no ascites | 0 | 0 | Factual
no peritoneal implants | 0 | 0 | Factual
uterus and adnexa were normal | 0 | 0 | Factual
serum tumor markers were negative | 0 | 0 | Factual
surgical pelvic exploration | -672 | -672 | Factual
30-centimeter mass of the left broad ligament | -672 | -672 | Factual
no ascites | -672 | -672 | Factual
no peritoneal carcinomatosis | -672 | -672 | Factual
uterus and right adnexa were normal | -672 | -672 | Factual
total hysterectomy with adnexectomy | -672 | -672 | Factual
removal of the mass | -672 | -672 | Factual
definitive histological diagnosis was leiomyosarcoma | -672 | -672 | Factual
isolated fever | 48 | 48 | Factual
major inflammatory syndrome | 48 | 48 | Factual
leukocytes 15,000/μL | 48 | 48 | Factual
C-reactive protein 317 mg/dL | 48 | 48 | Factual
contrast-enhanced computed tomography scan | 48 | 48 | Factual
bilobed air and fluid collection | 48 | 48 | Factual
abscess | 48 | 48 | Factual
blood pressure dropped | 48 | 48 | Factual
vasopressor therapy | 48 | 120 | Factual
noradrenaline | 48 | 120 | Factual
emergency revision surgery | 72 | 72 | Factual
peritoneal cavity exploration | 72 | 72 | Factual
moderately abundant non-purulent serosanginous peritoneal fluid | 72 | 72 | Factual
adhesions to the Douglas pouch | 72 | 72 | Factual
peritonitis | 72 | 72 | Factual
antibacterial treatment with piperacillin/tazobactam and gentamicin | 72 | 168 | Factual
extubated | 96 | 96 | Factual
hemodynamic support with noradrenaline | 96 | 120 | Factual
transferred to the intensive care unit | 96 | 96 | Factual
clinically improved | 120 | 168 | Factual
noradrenaline requirement decreased | 120 | 120 | Factual
discontinuation of noradrenaline | 120 | 120 | Factual
decrease in inflammatory markers | 120 | 168 | Factual
microbiological analysis of the peritoneal fluid | 120 | 120 | Factual
Gardnerella vaginalis | 120 | 120 | Factual
discontinuation of gentamicin | 120 | 120 | Factual
addition of metronidazole | 120 | 168 | Factual
Atopobium vaginae | 144 | 144 | Factual
antibacterial susceptibility testing | 144 | 144 | Factual
Gardnerella vaginalis resistant to metronidazole | 144 | 144 | Factual
Gardnerella vaginalis susceptible to penicillin G | 144 | 144 | Factual
Atopobium vaginae susceptible to metronidazole | 144 | 144 | Factual
piperacillin/tazobactam active against both bacteria | 144 | 144 | Factual
final diagnosis was an early postoperative peritonitis-induced septic shock | 168 | 168 | Factual
discharged from the intensive care unit | 168 | 168 | Factual
antibacterial therapy stopped | 168 | 168 | Factual