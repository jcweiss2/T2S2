53 years old | 0
male | 0
admitted to the emergency department | 0
complained of four-month progressive fatigue | -672
pain of his legs | -168
weakness of his legs | -168
taking diclofenac | -672
no fever | 0
no weight loss | 0
no night sweats | 0
spastic paraparesis | 0
sensitive level at the eight thoracic medullar segment | 0
pale | 0
gingival hemorrhage | 0
ecchymosis of the left thigh | 0
hepatomegaly | 0
spinal magnetic resonance imaging | 0
posterolateral extradural mass | 0
medullar compression | 0
anemia | 0
thrombocytopenia | 0
white blood count of 7.5 x 10^9/L | 0
absolute promyelocyte count of 4.8 | 0
blast count of 1.3 | 0
fibrinogen below normal limits | 0
international normalized ratio of 1.86 | 0
partial thromboplastin time within normal limits | 0
electrolytes within normal range | 0
hepatic and renal functions within normal range | 0
uric acid elevated | 0
lactate dehydrogenase elevated | 0
bone marrow biopsy | 0
hypercellularity | 0
massive infiltration of promyelocytes | 0
palisades of Auer rods | 0
diagnosis of APL | 0
qualitative polymerase chain reaction for the PML-RARα gene positive | 0
cytogenetic examination identified a t(15;17)(q22q21) abnormality | 0
ATRA therapy initiated | 0
daunorubicin initiated | 48
ATRA syndrome | 24
febrile neutropenia | 24
dexamethasone | 24
ceftazidime | 24
amikacin | 24
deterioration in the weakness of his legs | 72
lost bladder sphincter control | 72
radiotherapy for the extradural lesion | 120
nephrotic syndrome | 168
ATRA interrupted | 168
hematological remission of APL | 240
persistence of the extradural mass | 240
respiratory distress | 336
hypotension | 336
shock | 336
pneumonia | 336
vancomycin | 336
imipenem | 336
intensive care with ventilation support | 336
died of sepsis | 408