72 years old | 0
    male | 0
    dermatomyositis | -40320
    pancytopenic | -3360
    methotrexate therapy | -3360
    aplastic anemia | -3360
    bone marrow biopsy | -3360
    hypocellularity | -3360
    neutropenic fever | -720
    second hospitalization | -720
    neutropenic fever | -720
    ATG therapy considered | 0
    hypersensitivity testing | 0
    equine ATG ID test | 0
    wheal and flare reaction | 0
    respiratory distress absence | 0
    generalized urticaria absence | 0
    systemic symptoms absence | 0
    prednisone use | -720
    white blood cell count 500 | 0
    lymphocytes 400 | 0
    epicutaneous skin test | 120
    nonreactive epicutaneous test | 120
    histamine control positive | 120
    saline control nonreactive | 120
    white blood cell count 200 | 0
    lymphocytes 200 | 0
    horse dander testing | 120
    horse dander negative | 120
    informed consent | 0
    desensitization regimen | 0
    prednisone 40 mg daily | 0
    intensive care transfer | 0
    emergency medications available | 0
    resuscitation equipment available | 0
    premedication diphenhydramine | 0
    premedication ranitidine | 0
    premedication acetaminophen | 0
    premedication methylprednisolone | 0
    ranitidine every 8 hours | 0
    acetaminophen for fever prevention | 0
    ID desensitization doses | 0
    subcutaneous desensitization doses | 0
    intravenous desensitization doses | 0
    no localized reaction | 0
    no systemic reaction | 0
    premedication before dose 12 | 0
    full therapeutic dosing | 24
    continuous ATG infusion | 24
    fungal septicemia | 672
    death | 672

    