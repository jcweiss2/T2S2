43 years old | 0
female | 0
productive cough | -240
diarrhoea | -240
vomiting | -240
end-stage renal failure | -10080
crescentic IgA nephropathy | -10080
live related renal transplant | -10920
chronic transplant glomerulopathy | -10920
poor transplant function | 0
estimated glomerular filtration rate 15 mL/min | 0
tacrolimus | 0
mycophenolate mofetil | 0
sodium bicarbonate | 0
atenolol | 0
ramipril | 0
methoxy polyethylene glycol-epoetin beta | 0
severe hyponatraemia | 0
serum sodium 102 mmol/L | 0
acute-on-chronic kidney injury | 0
bilateral consolidation | 0
no fluid overload | 0
septic screen | 0
atypical respiratory serology | 0
antibiotics | 0
community-acquired pneumonia | 0
intensive care unit | 0
CVVHD | 0
protocol for sodium concentration adjustment | 0
sodium concentration adjustment | 0
serum sodium 100 mmol/L | 0
potassium 5.3 mmol/L | 0
creatinine 416 μmol/L | 0
urea 39.4 mmol/L | 0
magnesium N/A | 0
bicarbonate N/A | 0
chloride N/A | 0
phosphate 1.94 mmol/L | 0
eGFR N/A | 0
CRP 83.7 mg/L | 0
serum osmolality 248 mOsm/kg | 0
urine osmolality 246 mOsm/kg | 0
TSH N/A | 0
confusion | 72
agitation | 72
intubation | 72
lumbar puncture | 72
CT brain | 72
cerebrospinal fluid analysis | 72
no meningism | 72
no encephalitis | 72
serum sodium 116 mmol/L | 72
tacrolimus level 32 μg/L | 72
sepsis | 72
renal failure | 72
extubation | 96
normal cognitive function | 96
normal neurological function | 96
transfer to renal unit | 144
serum sodium 135 mmol/L | 144
dialysis dependent | 144
discharge from hospital | 240