44 years old | 0
male | 0
chronic hepatitis B virus carrier | 0
normal liver function | 0
admitted to the local hospital | 0
seven-day history of dry cough | -168
seven-day history of shortness of breath | -168
seven-day history of hypodynamia | -168
three days prior to admission experienced frequent coughing | -72
three days prior to admission experienced yellow-white sputum | -72
three days prior to admission experienced high fever (38.9°C) | -72
20-year history of smoking | -175200
approximately twenty cigarettes daily | -175200
denied recent exposure to sick animals | 0
denied visiting to farms | 0
temperature of 38.7°C | 0
heart rate of 134/min | 0
respiratory rate of 24/min | 0
blood pressure of 124/70 mmHg | 0
fine crackles in the left lung | 0
chest computed tomography (CT) scan demonstrated patchy high-density shadows with blurred margins | 0
pan-lobar pneumonia | 0
slightly elevated leucocyte count (10.77 × 109/L) | 0
elevated D-dimer (31.21 mg/L) | 0
elevated glucose levels (9.93 mmol/L) | 0
elevated blood urea nitrogen (27.57 mmol/L) | 0
elevated creatinine (576 umol/L) | 0
elevated C reactive protein (>200 mg/L) | 0
elevated procalcitonin (PCT) (36.33 ug/L) | 0
elevated alanine aminotransferase (107 IU/L) | 0
elevated aspartate aminotransferase (401 IU/L) | 0
elevated lactic dehydrogenase (2119 IU/L) | 0
elevated creatine kinase (4620 IU/L) | 0
elevated serum total bilirubin (67.1 umol/L) | 0
decreased serum albumin (25.8 g/L) | 0
decreased serum sodium levels (128 mmol/L) | 0
arterial blood gas analysis showed normal pH (7.45) | 0
normal PaO2 (71.3mmHg) | 0
normal blood lactate (1.5mmol/L) | 0
decreased PaCO2 (25.5mmHg) | 0
decreased PO2/FiO2 (216.1mmHg) | 0
samples collected for culture | 0
no pathogenic bacteria, fungi, or viruses found | 0
acid-fast staining of sputum negative | 0
diagnosed with pneumonia | 0
empiric treatment initiated with meropenem | 0
empiric treatment initiated with moxifloxacin | 0
respiratory status deteriorated after 6 hours | 6
delirium observed after 6 hours | 6
intubation and ventilator required | 6
transferred to ICU of local hospital | 6
repeated blood-gas analysis | 6
pH level 7.23 | 6
PaCO2 34mmHg | 6
PaO2 193.5mmHg | 6
PO2/FiO2 193.5mmHg | 6
blood lactate 1.3mmol/L | 6
transferred to our hospital | 6
experienced hypoxemia during transportation | 6
SpO2 60%-70% | 6
hemorrhagic fluid gushed out from tracheal tube | 6
wet and dry rales in both lungs | 6
arterial blood-gas analysis | 6
pH 7.29 | 6
PaCO2 30.4mmHg | 6
PaO2 73.7mmHg | 6
PO2/FiO2 73.7mmHg | 6
blood lactate 2.3mmol/L | 6
developed ARDS | 6
lung-protective ventilation administered | 6
deep sedation administered | 6
analgesia administered | 6
paralysis using neuromuscular blocker | 6
continuous renal replacement therapy administered | 6
prone-position ventilation administered | 6
condition worsened on second day after intubation | 30
increased bilateral pulmonary infiltrates | 30
leucocyte count increased (19.54 × 109/L) | 30
PCT levels increased (83.26 ug/L) | 30
ventilatory parameters high | 30
