65 years old | 0
male | 0
admitted to the hospital | 0
shortness of breath | -96
fever | -96
dry cough | -96
fatigue | -96
breath sounds reduced | 0
oxygen saturation 93% | 0
bilateral peripheral ground-glass attenuation | 0
patchy consolidation | 0
lung involvement 60%-70% | 0
SARS-CoV-2 RT-PCR test positive | 0
increased temperature | 0
saturation with free breathing decreased to 90% | 0
white cell count 7.93 х 109/ L | 0
hemoglobin 159 g/l | 0
platelet count 468 х 109/l | 0
Westergren ESR 41 mm/h | 0
interleukine 6 102 pg/ml | 0
С-reactive protein 142 mg/l | 0
ferritin 939.92 μg/ml | 0
D-dimer 609 ng/ml | 0
procalcitonin 0.11 ng/ml | 0
treatment with dexamethason | 0
treatment with heparin | 0
treatment with tocilizumab | 0
treatment with acetylcysteine | 0
treatment with pantoprazole | 0
treatment with nadroparin calcium | 0
oxygen supplementation | 0
air and pleural effusion in the right pleural cavity | 360
collapse of the right lung | 360
thoracentesis | 360
thoracostomy | 360
evacuation of 1400 ml of yellowish opaque liquid | 360
linezolid therapy | 360
imipenem/cilastatin therapy | 360
oxygen supplementation with flow rate of 8-10 l/min | 360
daily drainage volume 300-1000 ml | 360
pleural effusion with gas bubbles | 432
focal area of subpleural infiltration | 432
central cavity of destruction | 432
air layer up to 47 mm | 432
radiological signs of left side hydropneumothorax | 432
pleural fluid analysis | 432
exudative lymphocytic-rich effusion | 432
Acinetobacter baumannii in pleural fluid | 432
Pseudomonas aeruginosa in pleural fluid | 432
Klebsiella pneumonia in urine culture | 432
negative SARS-CoV-2 RT-PCR test | 504
needle thoracocentesis | 504
new pleural drainage | 504
air and creamy purulent mass aspirated | 504
serofibrinous hemorrhagic fluid drawn | 504
chest CT showed air and pleural effusion | 504
diagnosis of pleural empyema | 504
transfer to Surgical Department | 504
right pleural space irrigated with antiseptic solutions | 504
lung expansion by continuous vacuum aspiration | 504
encapsulated pleural effusion | 576
ultrasound-guided puncture | 576
new drainage of pleural cavity | 576
4-week antibiotic therapy | 672
discharged from hospital | 672
oxygen saturation 97% | 672
chest CT showed small amount of fluid | 672
lab test scores normal | 672
С-reactive protein 11.7 mg/l | 672
procalcitonin < 0.1 ng/ml | 672