20 years old | 0
male | 0
motor vehicle accident | -1
severe and diffuse trauma to the abdomen, trunk and extremities | -1
unstable vital signs | -1
flaccid paraplegia | -1
complete loss of voluntary control over bowel and bladder function | -1
FAST examination was negative | 0
multiple rib fractures | 0
bilateral hemothoraces | 0
hemoperitoneum | 0
AAST grade 4 splenic injury | 0
left-sided renal and adrenal injury | 0
right-sided scapular fracture | 0
transdiscal AO type C fracture | 0
bilateral facet subluxation of T11 over T12 | 0
pneumothoraces were drained through chest tubes | 0
exploratory laparotomy | 0
splenectomy | 0
left retroperitoneal space was packed | 0
“Damage Control” type surgery | 0
MRI of the spine | 24
subluxation of T11 over T12 | 24
rupture of the intervertebral disc | 24
rupture of the posterior longitudinal ligament | 24
9 mm-thick epidural hematoma | 24
medullary contusion at the level of T11–T12 | 24
spinal surgery | 48
reduction of the subluxation | 48
trans-pedicular screw fixation from T9 to L2 | 48
intra-operative post-traumatic dural tear | 48
small leak of CSF | 48
planned second look laparotomy | 72
depacking | 72
no bleeding | 72
persistence of the retroperitoneal hematoma | 72
small amount of turbid liquid | 72
intense back pain | 96
hallucinations | 96
agitated | 96
septic state | 96
thoracolumbar MRI | 96
thoraco-abdominal CT | 96
large bilateral para-vertebral and retroperitoneal fluid collections | 96
AAST grade 3 pancreatic injury | 96
revision of the thoraco-lumbar wound | 120
CSF leak from a circular dural breach | 120
breached area was repaired with a fibrin sealant | 120
debridement of necrotic tissue | 120
drainage of newly purulent collections | 120
copious irrigation with normal saline | 120
tight closure of the facia and subcutaneous tissue | 120
two Penrose drains were left in the superficial layers | 120
retroperitoneal fluid collections were evacuated | 120
blood cultures, paravertebral and abdominal fluid collections were positive for Enterobacter cloacae | 120
intravenous antibiotic treatment with Meropenem | 120
paravertebral and abdominal collections increased | 144
repeat cultures remained positive for Enterobacter cloacae | 144
paravertebral collections exteriorized through the dorsal skin | 144
serum amylase and lipase were measured high | -1
high levels of amylase and lipase were found in the dorsal spinal fluid collections | 168
ERCP was performed | 168
placement of a stent bridging the defect of the main duct | 168
total parenteral nutrition | 0
subcutanous somatostatine | 0
progressive enteral feeding by naso-jejunal tube | 168
patient could be orally fed | 240
enteral and parenteral nutritional intake could be weaned off | 240
patient's general condition slowly improved | 240
drains were removed | 1248
patient transferred to a rehabilitation facility | 1248
neurologic status of complete paraplegia | 1248
sensory level at T10 | 1248
antibiotic treatment was given for a total of 7 months | 0
CT showed complete resolution of the collections | 2016