Here is the table of events and timestamps:

10 years old | 0
male | 0
pre-term | -33.5
Russell-Silver syndrome | -6
proteinuria | -6
hypoalbuminemia | -6
nephrotic syndrome | -6
high-dose steroid | -6
calcineurin inhibitor | -6
renal function deteriorated | -6
right renal vein thrombosis | -3
pulmonary embolism | -3
anticoagulants | -3
persistent pulmonary hypertension | -3
sildenafil | -3
kidney transplantation | 0
immunosuppression | 0
prednisolone | 0
mycophenolate mofetil | 0
tacrolimus | 0
MMF discontinued | 70
steroid tapered | 70
pneumocystis pneumonia | 90
mechanical ventilation | 90
intravenous sulfamethoxazole/trimethoprim | 90
hematuria | 135
dysuria | 135
BUN 24 mg/dL | 135
creatinine 0.56 mg/dL | 135
C-reactive protein 0.42 mg/dL | 135
red blood cell count > 100/HPF | 135
white blood cell count > 100/HPF | 135
urine culture negative | 135
BK virus negative | 135
JC virus positive | 135
adenovirus positive | 135
hemodialysis | 135
hydration | 135
pain control | 135
hematuria persisted | 142
dysuria persisted | 142
RBC count > 100/HPF | 142
WBC count 1-4/HPF | 142
immunopression maintained | 142
fever | 159
general weakness | 159
chest tightness | 159
mild cough | 159
hematuria | 159
BUN 175 mg/dL | 159
creatinine 8.29 mg/dL | 159
C-reactive protein 30.23 mg/dL | 159
piperacillin/tazobactam | 159
sputum culture negative | 159
blood culture negative | 159
urine culture negative | 159
adenovirus real-time PCR positive | 159
CMV antigen positive | 159
immunopression reduction | 159
ganciclovir | 159
renal allograft biopsy | 159
diffuse necrotizing granulomatous tubulointerstitial nephritis | 159
CD3 negative | 159
C4d negative | 159
JC virus PCR positive | 159
CMV PCR positive | 159
granulocyte colony-stimulating factor | 159
immunoglobulin | 159
transfusion | 159
hemodialysis | 159
cidiocvir | 167
renal impairment dose | 167
hemodialysis | 167
cidiocvir | 170
renal impairment dose | 170
hemodialysis | 170
cidiocvir | 173
renal impairment dose | 173
hemodialysis | 173
cidiocvir | 176
renal impairment dose | 176
hemodialysis | 176
cidiocvir | 179
renal impairment dose | 179
hemodialysis | 179
cidiocvir | 182
renal impairment dose | 182
hemodialysis | 182
cidiocvir | 185
renal impairment dose | 185
hemodialysis | 185
cidiocvir | 188
renal impairment dose | 188
hemodialysis | 188
cidiocvir | 191
renal impairment dose | 191
hemodialysis | 191
cidiocvir | 194
renal impairment dose | 194
hemodialysis | 194
cidiocvir | 197
renal impairment dose | 197
hemodialysis | 197
cidiocvir | 200
renal impairment dose | 200
hemodialysis | 200
cidiocvir | 203
renal impairment dose | 203
hemodialysis | 203
cidiocvir | 206
renal impairment dose | 206
hemodialysis | 206
cidiocvir | 209
renal impairment dose | 209
hemodialysis | 209
cidiocvir | 212
renal impairment dose | 212
hemodialysis | 212
cidiocvir | 215
renal impairment dose | 215
hemodialysis | 215
generalized tonic-clonic seizure | 215
vancomycin | 215
meropenem | 215
acyclovir | 215
death | 215