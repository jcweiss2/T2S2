23 years old | 0
female | 0
Caucasian | 0
admitted to the hospital | 0
nonverbal acoustic hallucinations | -240
insomnia | -240
psychomotor slowing | 0
cerebral MRI normal | 0
CSF 73 leukocytes/μL | 0
isolated oligoclonal bands | 0
slightly increased lactate | 0
NMDAR antibodies in serum and CSF positive | 0
ovarian teratoma not detected | 0
methylprednisolone administered | 0
immunoglobulins administered | 0
oral prednisolone administered | 0
condition worsened | 24
dyskinesias | 24
dysautonomia | 24
respiratory insufficiency | 24
analgosedation and artificial ventilation | 24
multidrug analgosedation | 24
propofol administered | 24
midazolam administered | 24
esketamine administered | 24
sufentanil administered | 24
alpha-2 receptor agonists administered | 24
4-hydroxybutyrate administered | 24
drug-induced hepatotoxicity | 48
transaminases 36-fold of normal | 48
switched to isoflurane | 48
rituximab administered | 72
immunoadsorption | 72
dyskinesias reappeared | 120
isoflurane concentration increased | 120
MRI showed symmetrical striatal and dentate nuclei T2-weighted hyperintensities | 168
mesiotemporal atrophy | 168
CSF lactate increased | 168
CSF neurofilament light chain levels increased | 168
suspecting adverse reaction to isoflurane | 168
IV analgosedation reinstated | 168
arterial hypertension reappeared | 192
MRI showed posterior reversible encephalopathy syndrome | 216
striatal and dentate nucleus hyperintensities dissolved | 216
patient became alert and adequately oriented | 2160
severe flaccid tetraparesis | 2160
hypoesthesias | 2160
critical illness polyneuropathy/myopathy | 2160
minimal cognitive impairment | 4320
cerebellar ataxia | 4320
MRI showed reversible forebrain atrophy | 4320
cerebellar atrophy | 4320
cerebellar ataxia showed mild improvement | 8640