25 years old| 0  
    male| 0  
    referred to ICU for evaluation and treatment of unexplained shock syndrome| 0  
    recent asymptomatic COVID-19 infection| -672  
    no history of smoking, alcohol, or drug use| 0  
    no exposure to infectious or toxic agents| 0  
    recreational exercise| 0  
    double BNT162b2 vaccinated| -648  
    last vaccine dose nine months before admission| -648  
    presented to general practitioner with fever (>39°C)| -96  
    abdominal pain| -96  
    vomiting| -96  
    diarrhoea| -96  
    elevated Erythrocyte Sedimentation Rate| -96  
    elevated C-Reactive Protein (CRP)| -96  
    normal white blood cell count| -96  
    normal chest radiography| -96  
    prescribed amoxicillin/clavulanic acid| -96  
    switched to cefuroxime| -96  
    diffuse erythematous and maculopapular rash| -96  
    worsening clinical condition| 0  
    presented to emergency department| 0  
    ill patient with dyspnoea| 0  
    diffuse abdominal pain| 0  
    normal heart-lung auscultation| 0  
    rash persisted| 0  
    bilateral conjunctivitis| 0  
    no other mucosal lesions| 0  
    blood pressure 141/80 mmHg| 0  
    pulse 110 bpm| 0  
    temperature 37.8°C| 0  
    oxygen saturation 98% without supplemental oxygen| 0  
    sinus tachycardia on ECG| 0  
    new diffuse PR-depression on ECG| 0  
    neutrophilia| 0  
    thrombocytopenia| 0  
    lymphopenia| 0  
    high ferritin| 0  
    high D-dimer| 0  
    CRP doubling since GP visit| 0  
    increased serum creatinine| 0  
    increased gamma-glutamyl transferase| 0  
    increased alkaline phosphatase| 0  
    increased total bilirubin| 0  
    thoraco-abdominal CT performed| 0  
    suspected intra-abdominal sepsis| 0  
    uncomplicated ileocaecal inflammation| 0  
    mesenteric lymphadenopathy| 0  
    splenomegaly| 0  
    normal lung parenchyma| 0  
    discrete pericardial effusion| 0  
    transthoracic echocardiography (TTE) showed normal cardiac morphology and function| 0  
    no significant pericardial effusion on TTE| 0  
    blood, sputum, stool, and urine cultures incubated| 0  
    switched to intravenous ciprofloxacin and metronidazole| 0  
    developed hypotension over next two days| 48  
    high anion gap metabolic acidosis due to lactic acid accumulation| 48  
    necessitating fluid resuscitation| 48  
    necessitating norepinephrine| 48  
    developed type 1 respiratory insufficiency| 48  
    treated with High Flow Nasal Oxygen| 48  
    sedation| 48  
    intubation| 48  
    mechanical ventilation| 48  
    further clinical deterioration| 96  
    repeated thoraco-abdominal CT| 96  
    terminal ileitis| 96  
    diffuse colitis| 96  
    increased lymphadenopathy| 96  
    hepatosplenomegaly| 96  
    new ascites| 96  
    bilateral pleural effusions| 96  
    failure of shock resolution| 96  
    persistent inflammation| 96  
    antimicrobial escalation to meropenem and vancomycin| 96  
    persistent suspicion for intra-abdominal septic shock| 96  
    no etiological explanation on repeat imaging| 96  
    exploratory laparoscopy performed| 96  
    moderate clear ascites| 96  
    no signs of infection| 96  
    ascites recovered for culture| 96  
    unexplained shock with increasing vasopressor doses| 96  
    worsening peripheral perfusion| 96  
    increasing lactate| 96  
    repeat TTE performed| 96  
    mildly dilated left ventricle| 96  
    moderately decreased ejection fraction| 96  
    anteroseptal akinesia| 96  
    hypokinesia of other segments| 96  
    6 mm circumferential pericardial effusion| 96  
    no tamponade physiology| 96  
    new chest radiograph showed cardiomegaly| 96  
    bilateral pleural effusions| 96  
    pulmonary edema| 96  
    high sensitive troponin T elevated up to 288 ng/L| 96  
    NT-pro-BNP 28,770 pg/mL| 96  
    suspected myocarditis| 96  
    suspected cardiogenic shock| 96  
    dobutamine started| 96  
    levosimendan started| 96  
    cardiac MRI (CMR) performed| 96  
    moderately dilated left ventricle| 96  
    moderately reduced systolic function| 96  
    non-ischemic myocardial injury| 96  
    increased myocardial extracellular volume by T1-mapping| 96  
    focal myocardial edema in anterior and apicolateral segments on T2-weighted images| 96  
    no focal myocardial late gadolinium enhancement| 96  
    fulfilled 2018 Lake Louise criteria for myocarditis| 96  
    pericardial inflammation| 96  
    pericardial effusion| 96  
    pericardial thickening| 96  
    pericardial gadolinium enhancement| 96  
    retrospective CT evaluation confirmed normal coronary arteries| 96  
    no arrhythmia| 96  
    negative cultures| 96  
    negative auto-immune serology| 96  
    negative viral serology| 96  
    persistently high SARS-CoV-2 viral load| 96  
    presence of anti-N IgG| 96  
    diagnosed with MIS-A| 96  
    suggestive rash| 96  
    conjunctivitis| 96  
    gastro-intestinal symptoms| 96  
    thrombocytopenia| 96  
    fever| 96  
    major inflammation| 96  
    shock| 96  
    severe myocarditis| 96  
    cardiac failure| 96  
    lack of any other explanation| 96  
    intravenous immunoglobulins (IVIGs) administered| 96  
    pulse corticosteroids started| 96  
    patient improved| 120  
    weaned off ventilatory support| 120  
    weaned off inotropic support| 120  
    weaned off vasopressor support| 120  
    antibiotics discontinued| 144  
    regression of PR depression on ECG| 120  
    TTE showed improved anteroseptal contractility| 120  
    increased LVEF| 120  
    regressed pericardial effusion| 120  
    corticosteroids continued orally| 120  
    slowly tapered over six weeks| 120  
    proton pump inhibitor associated| 120  
    calcium/vitamin D supplements associated| 120  
    heart failure therapy started| 120  
    bisoprolol 2.5 mg| 120  
    lisinopril 10 mg daily| 120  
    left ventricular function improved rapidly| 120  
    lisinopril not escalated to valsartan-sacubitril| 120  
    no mineralocorticoid receptor antagonist associated| 120  
    low-dose aspirin associated| 120  
    asymptomatic at ambulatory follow-up| 168  
    no inflammation at ambulatory follow-up| 168  
    resting ECG normal| 168  
    TTE showed lower septum and posterior wall thicknesses| 168  
    normalisation of left ventricular diameters| 168  
    normalisation of systolic function| 168  
    heart failure therapy to be discontinued in future| 168  
    low dose aspirin to be discontinued in future| 168  

<|eot_id|>