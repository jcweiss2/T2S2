36 years old | 0
female | 0
admitted to the Emergency Department | 0
sudden loss of consciousness | 0
head trauma | 0
falling from her own height | -72
loss of strength in the lower extremities | -72
impaired ambulation | -72
sudden-onset disabling holocranial headache | -336
aggressive behavior | -336
vertigo | -336
no fever | -336
no malaise | -336
somatoform disorder diagnosis | -72
depressive episode diagnosis | -72
major depression | -13104
no adherence to medical treatment | -13104
two previous suicide attempts | -13104
recumbent patient | 0
Glasgow coma score of 11 | 0
no focal neurologic deficits | 0
no meningeal signs | 0
aware of her environment | 0
mutism | 0
no verbal contact | 0
no eye contact | 0
hydrated integumentary system | 0
no integumentary alterations | 0
horizontal nystagmus | 0
oculogyric crises | 0
no head and neck alterations | 0
stereotyped movements in all four extremities | 0
normal plantar reflexes | 0
normal deep tendon reflexes | 0
mass in the right axillary line | 0
blood pressure 94/60 mm Hg | 0
heart rate 77 bpm | 0
respiratory rate 20 rpm | 0
temperature 36.5°C | 0
body-weight 60 kg |%23420
