62 years old | 0
female | 0
Saudi | 0
admitted to King Khalid University Hospital | 0
elective laparoscopic sigmoid resection | 0
complicated and uncomplicated attacks of diverticulitis | -672
increase in urea | 0
increase in creatinine | 0
increase in potassium | 0
increase in white blood cells (WBCs) | 0
decrease in red blood cells (RBCs) | 0
decrease in hemoglobin | 0
decrease in hematocrit | 0
decrease in bicarbonate | 0
diagnosed with diverticulosis | 0
diverticula in the sigmoid and distal descending colon | 0
spiked a fever | 72
temperature of 38.9°C | 72
septic screening | 72
diagnosed with urinary tract infection | 72
antibiotics started | 72
low hemoglobin | 72
blood transfusion | 72
hypotensive | 72
blood pressure 85/52 mmHg | 72
oxygen saturation 94% | 72
pulse rate 110/min | 72
transfusion stopped | 72
hydrocortisone started | 72
transferred to surgical intensive care unit (SICU) | 72
dopamine given | 72
transfusion of 1 unit of packed RBCs | 72
transferred back to general ward | 144
follow-up WBC count 12.7 | 144
blood culture showed Escherichia coli | 144
urine culture showed Klebsiella pneumonia | 144
antibiotic changed | 144
complained of abdominal pain | 168
abdominal distention | 168
WBC 13.8 | 168
computed tomography (CT) showed air bubbles in abdominal cavity | 168
air bubbles in retroperitoneal with extension into mediastinum | 168
evidence of bowel air at serosal surface of gallbladder and omentum | 168
anastomotic leakage (AL) | 168
diagnostic laparoscopy | 168
laparoscopic Hartmann's sigmoid resection | 168
transferred to SICU postoperatively | 168
intubated | 168
started on inotrope | 168
CT scan showed no drainable intra-abdominal collection | 240
discharged | 240