21 years old | 0  
    male | 0  
    allergic to cefuroxime | 0  
    allergic to metronidazole | 0  
    sore throat | -96  
    shortness of breath | -96  
    left tonsillitis | -96  
    septic shock | -96  
    fever | -96  
    poor oral intake | -96  
    febrile | -96  
    low-grade temperature | -96  
    bilateral lower zone infiltrates | -96  
    bilateral pleural effusion | -96  
    respiratory failure | -96  
    intubation | -96  
    doxycycline | -96  
    clindamycin | -96  
    vancomycin | -96  
    clinical deterioration | 0  
    meropenem | 0  
    doxycycline continued | 0  
    throat swab negative | 0  
    urine culture negative | 0  
    sputum culture negative | 0  
    endotracheal aspirates negative | 0  
    blood culture positive for Fusobacterium necrophorum | 168  
    persistent leukocytosis | 168  
    neck pain | 168  
    CT neck | 168  
    CT thorax | 168  
    left internal jugular thrombophlebitis | 168  
    multiple cavitating lung nodules | 168  
    diagnosis of Lemierre's syndrome | 168  
    antibiotics continued | 168  
    intravenous amoxicillin-clavulanate | 168  
    discharged to general ward | 168  
    oral amoxicillin-clavulanate | 168  
    resolution of lung infiltrates | 168  
    antibiotic stopped | 672  
    no anticoagulation | 0  
    discharge home | 168  
    satisfactory progress | 168  
