67 years old | 0
male | 0
multiple cerebrovascular events | -672
myocardial infarction | -672
hypertension | -672
30 pack-year smoking history | -672
dull 5/10 sacral pain | -24
pelvic magnetic resonance imaging (MRI) examination | -24
large, well circumscribed, heterogeneously enhancing mass through the mid body of the sacrum | -24
core biopsy | -24
sacral chordoma | -24
preoperative external beam radiation | -168
sacrectomy | 0
abdominoperineal resection | 0
colostomy | 0
pelvic and perineal defect | 0
reconstructed using a right VRAM flap | 0
admission to the intensive care unit | 0
transferred to the orthopedic surgery unit | 120
regular flap checks | 120
flap consistently well perfused | 120
fever | 312
tachycardia | 312
abdominal discomfort | 312
increase in white blood cell count | 312
septic workup | 312
flap demonstrated signs of both venous and arterial insufficiency | 312
computed tomography of the pelvis | 312
markedly distended bladder | 312
bilateral hydronephrosis | 312
deep inferior epigastric pedicle occluded | 312
bladder decompressed | 312
improvement in the patient's clinical status | 312
perfusion to the flap did not improve | 312
total flap loss | 312
debridement of the VRAM flap | 504
thrombosis of the deep inferior epigastric pedicle | 504
flap debridement | 504
bilateral advancement flaps elevated for closure | 504
discharged from hospital | 960
wound completely healed | 1440