male | 0
newborn | 0
38 weeks and 6 days of gestational age | 0
3410 g | 0
Apgar score of 10/10/10 | 0
vaginal delivery | 0
oxytocin-induced labor | -672
uneventful cephalic presentation | -672
mother 31 years old | -672
gravida 5 | -672
para 4 | -672
previously healthy | -672
normal prenatal consultations | -672
follow-up | -672
immunity for rubella | -672
immunity for toxoplasmosis | -672
serologies for hepatitis B negative | -672
serologies for hepatitis C negative | -672
serologies for syphilis negative | -672
serologies for HIV negative | -672
blood type B+ | -672
evaluation for irregular blood group antibodies negative | -672
respiratory failure | 27
respiratory frequency of 98 respiratory movements per minute | 27
intense respiratory labor | 27
intercostal and subcostal retractions | 27
tachycardia | 27
pulse rate of 170 beats per minute | 27
capillary refill time of 7 seconds | 27
room air oximetry of 85% | 27
small amplitude arterial pulses | 27
mechanical ventilatory support | 27
umbilical vein catheterization | 27
fluid resuscitation | 27
administration of vasoactive drugs | 27
septic shock | 27
metabolic acidosis | 27
hypotension | 27
upper limbs systolic pressure higher than lower limbs | 27
echodopplercardiogram | 27
left ventricle hypoplasia | 27
prostaglandin infusion | 27
patency of ductus arteriosus | 27
adequate retrograde shunt to aortic arch and coronary arteries | 27
situs solitus | 27
hypoplastic aortic arch | 27
retrograde blood flow | 27
systemic and pulmonary venous drainage preserved | 27
mitral valve hypoplasia | 27
no communication between left ventricle and aortic arch | 27
aortic valve atresia | 27
ductus arteriosus patent | 27
bidirectional flow | 27
heart enlarged | 27
right chambers hypokinesia | 27
left ventricle normal size and thickness | 27
left ventricle hypokinetic | 27
left-to-right flow | 27
restrictive atrial septal defect | 27
interventricular communication | 27
pericardium normal | 27
death | 72
cardiogenic shock | 72
multiple organ failure | 72
congenital heart disease | 72
anasarca | 72
cyanosis of lower limbs and scrotum | 72
red-wine-stained skin | 72
focal areas of desquamation | 72
lungs congestion | 72
pulmonary parenchyma in alveolar stage of development | 72
diffuse congestion of capillaries | 72
areas of hemorrhage | 72
scales in alveolar lumen | 72
numerous neutrophils in alveolar lumen | 72
alveolar hemorrhage | 72
liver enlarged | 72
diffuse congestion | 72
preserved portal tracts | 72
severely congested and dilated hepatic sinusoids | 72
foci of necrosis in hepatic lobule | 72
hepatic extra medullary hematopoiesis | 72
spleen congested | 72
enlarged | 72
congestion of red pulp | 72
kidneys congested | 72
diffuse congestion of cortex and medulla | 72
acute tubular necrosis | 72
absence of nephrogenic zone | 72