57 years old | 0
male | 0
admitted to the hospital | 0
diarrhea | -1080
weight loss | -1080
intermittent fever | -1080
right loin pain | -1080
intermittent abdominal pain | -1080
small volume diarrhea | -1080
3–4 episodes/day | -1080
weight loss of 8 kg | -1080
over 8 months | -1080
denied fever | 0
denied vomiting | 0
denied cough | 0
denied urinary symptoms | 0
recurrent infections | -1080
history of tuberculosis | -1080
tuberculosis contact | -1080
denied exposure to cattle | 0
denied exposure to pets | 0
reported consumption of cooked food mostly | 0
reported no food intolerance | 0
lives in rural South India | -1080
walks barefooted in his farm | -1080
consumes alcohol daily | -1080
denied intravenous (IV) drug abuse | 0
denied high-risk sexual behavior | 0
not on steroids | 0
not on immunosuppressive drugs | 0
married | 0
two children | 0
family members healthy | 0
bank manager | 0
cachexia | 0
hypotension | 0
blood pressure 80/60 | 0
dry tongue | 0
sunken eyes | 0
oral candida | 0
perioral vitiligo | 0
generalized macular erythematous | 0
purpuric lesion over trunk and abdomen | 0
nonmigratory lesions | 0
right loin tenderness | 0
bilateral wheezes | 0
no neck stiffness | 0
normal cardiac examination | 0
chronic diarrhea syndrome | 0
possible sepsis | 0
admitted to medical Intensive Care Unit | 0
ertapenem | 0
flucanozole | 0
Gram-negative sepsis | 0
probable gut origin sepsis | 0
oral/esophageal candidiasis | 0
neutrophilic leucocytosis | 0
low protein | 0
low albumin (4.8/2.2 g/dl) | 0
macrocytic anemia | 0
low mg | 0
low K | 0
low B12 | 0
low folate | 0
normal cortisol | 0
stool sent for GI pathogen multiplex PCR panel | 0
no pathogens (FilmArray, bio’Merieux) | 0
stabilization of BP | 0
contrast CT of chest and abdomen | 0
ground glass opacities in lung | 0
ileocaecal thickening | 0
upper GI endoscopy | 0
biopsy | 0
antral gastritis | 0
colonoscopy | 0
colonoscopy biopsy | 0
small ulcers throughout colon | 0
blood culture grew Klebsiella pneumoniae | 0
extended-spectrum beta-lactamases producer | 0
stool routine initial sample revealed pinworms | 0
duodenal mucosa biopsy revealed Strongyloides larval forms | 0
colonic biopsy revealed chronic colitis | 0
no granuloma | 0
no Strongyloides in colonic biopsy | 0
repeat stool for Strongyloides positive for adult worms | 24
Strongyloides hyperinfection | 24
started on ivermectin | 24
diarrhea settled | 24
encephalopathy | 24
switched to meropenem | 24
meningitic dose | 24
brain imaging normal | 24
cerebral spinal fluid (CSF) analysis | 24
CSF cell count of 1200 | 24
CSF protein-213 | 24
CSF sugar-40 | 24
no organisms on Gram stain | 24
CSF multiplex PCR revealed Klebsiella | 24
CSF culture grew Enterococcus faecium | 48
resistant to penicillin | 48
sensitive to vancomycin | 48
improved with meropenem and vancomycin | 48
repeat stool routine revealed persistent Strongyloides worms | 48
albendazole 400 mg twice daily added | 48
skin lesions suggestive of larva migrans | 48
autoimmune workup negative | 48
HIV 1 and 2 antibody negative | 48
CD4 1270 | 48
low IgG | 48
low IgM | 48
low IgE | 48
normal IgA | 48
no thymoma | 48
no lymph node enlargements | 48
peripheral smear no abnormal cells | 48
common variable immunodeficiency considered | 48
HTLV serology negative | 48
CD19 and CD20 negative | 48
antiendomysial antibody negative | 48
tissue transglutaminase antibody negative | 48
persistent Strongyloides in repeat stool | 48
low Ig level | 48
IVIg 400 mg/kg | 48
low Ig due to low globulins | 48
cleared stool of Strongyloides | 48
improved remarkably | 48
