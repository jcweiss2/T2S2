73 years old | 0  
    male | 0  
    presented with altered mental status | -168  
    presented with decreased appetite | -168  
    presented with poor oral intake | -168  
    hepatocellular carcinoma | -2892  
    history of alcohol use | -2892  
    congestive heart failure | -2892  
    coronary artery disease | -2892  
    chronic kidney disease | -2892  
    previous occupation as a floor maker | -2892  
    alcohol abuse | -2892  
    cigarette smoking | -2892  
    stopped alcohol 20 years prior | -175200  
    stopped cigarettes 40 years prior | -350400  
    afebrile | 0  
    hypotensive | 0  
    hypoxic | 0  
    mild right upper quadrant tenderness | 0  
    shock | 0  
    admitted to ICU | 0  
    elevated liver transaminases | 0  
    blood cultures obtained | 0  
    started empiric antibiotics | 0  
    chest X-ray unremarkable | 0  
    urinalysis unremarkable | 0  
    CT abdomen showed increased metastases | 0  
    diagnosed with hepatocellular carcinoma | -2892  
    imaging at diagnosis showed left liver mass | -2892  
    biopsy showed moderately differentiated HCC | -2892  
    recent MI | -2892  
    deemed poor surgical candidate | -2892  
    TACE performed | -2892  
    second TACE required | -2892  
    post-TACE admission for chest pain | -2892  
    post-TACE sepsis | -2892  
    CT post-TACE showed embolized mass and hypodensities | -2892  
    presented current admission | 0  
    CT on admission showed liver abscesses | 0  
    Raoultella planticola in blood cultures | 0  
    intermediate ampicillin sensitivity | 0  
    antibiotics narrowed to ceftriaxone and metronidazole | 0  
    drains placed on day 4 | 96  
    drain fluid with elevated WBC | 96  
    no culture growth | 96  
    repeat imaging showed abscess decrease | 96  
    clinical improvement | 96  
    discharged on IV ceftriaxone | 96  
    discharged on oral metronidazole | 96  
    readmitted during therapy | 672  
    worsening lesions | 672  
    decompensation | 672  
    comfort-based care | 672  
    expired | 672  
    <|eot_id|>
    