seventy years old | 0
Kuwaiti | 0
female | 0
admitted to the hospital | 0
uncontrolled Diabetes Mellitus | -672
irregular treatment with Lantus | -672
Lantus 20 units once daily | -672
uncompliant to Lantus | -672
uncompliant to follow up | -672
infrequent blood sugar monitoring | -672
chronic renal disease | -672
hypertensive | -672
Zestril 10 mg once daily | -672
Zestoretic 20 one tab daily | -672
Norvasc 5 mg once daily | -672
pacemaker | -672
anticoagulants | -672
gradual progressive left deep ear pain | -24
ear pain started to be bearable | -24
ear pain became very severe | -12
gradual decrease in hearing on the left ear | -24
facial asymmetry | -24
no tinnitus | 0
no discharge | 0
no itching | 0
first time to experience this complaint | 0
conscious | 0
oriented | 0
alert | 0
febrile | 0
vital signs stable | 0
edematous left ear | 0
very painful on touch | 0
tympanic membrane not visible | 0
ear pack inserted in the left external canal | 0
polypoidal mass in the inferior-posterior part of the left external canal | 12
biopsy of the mass | 12
inflammatory mass | 12
facial nerve exam showed slight weakness | 0
facial palsy | 0
hypoglossal nerve palsy | 0
nasopharyngeal scope showed mild bulging | 0
mild mucosal thickening of the left sphenoidal sinus | 0
admitted as a case of left malignant otitis externa | 0
IV Tazocin | 0
Fortum | 0
baseline investigations | 0
COVID19 nasopharyngeal swab | 0
sudden slurred speech | 24
urgent Computerized tomography of ear and skull base | 24
urgent neurology consultation | 24
left nasopharyngeal heterogonous enhanced soft tissue mass lesion | 24
bone erosion and destruction of related part of skull base | 24
suspected jugular thrombosis | 24
opacity of left middle ear and mastoid | 24
mild mucosal thickening of the left sphenoidal sinus | 24
surgical debridement of the diseased tissues | 48
biopsy of nasopharynx and left ear mass | 48
histopathology result reported as fungal hyphae | 48
IV Tazocin and Fortum discontinued | 48
liposomal amphotericin b started | 48
insulin to control blood sugar | 48
Eliquis administered | 48
hypothermia | 72
AKI | 72
hyponatremia | 72
liposomal amphotericin b stopped | 72
Posaconazole syrup started | 72
septic shock | 96
shifted to intensive care unit | 96
levophid infusion | 96
died | 120