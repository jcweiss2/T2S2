19 years old|0
male|0
intermittent fever|-240
progressive shortness of breath|-240
methicillin-susceptible Staphylococcus aureus infection|0
broad-spectrum antibiotics administration|0
Sievers type I bicuspid aortic valve|0
moderate aortic insufficiency|0
vegetation on ventricular side of aortic leaflet|0
vegetation on A2 segment of mitral valve|0
mitral valve perforation|0
moderate mitral regurgitation|0
aortomitral pseudoaneurysm|0
positive Doppler flow|0
paradoxical expansion|0
multiple foci of septic emboli|0
small localized subarachnoid hemorrhage|0
3-cm aneurysm in right pre-central sulcus|0
urgent cardiac surgery|0
bioprosthetic valve implantation|0
cardiac exposure via sternotomy|0
aorta cannulation|0
cavae cannulation|0
cardiopulmonary bypass initiation|0
del Nido cardioplegia|0
aortic valve excision|0
aortomitral aneurysm debridement|0
left atriotomy|0
anterior mitral leaflet vegetation excision|0
bovine pericardial patch repair|0
antibiotic solution irrigation|0
25-mm Freestyle porcine aortic root prosthesis implantation|0
inversion of prosthesis|0
placement in left ventricular outflow tract|0
alignment of right coronary ostia|0
commissural sutures|0
suture prosthetic rim to aortic annulus|0
noncoronary cusp reconstruction|0
bovine pericardial strip|0
aortomitral defect obliteration|0
prosthesis eversion|0
coronary ostia reimplantation|0
distal graft to ascending aorta anastomosis|0
normal functioning aortic root prosthesis|0
mild central leak in mitral valve|0
successful aortomitral defect repair|0
separation from cardiopulmonary bypass|0
no rhythm abnormalities|0
uneventful postoperative ICU stay|24
excised tissue microbiology negative|24
intravenous flucloxacillin administration|24
discharge after antibiotic completion|168
no neurologic deficits at discharge|168
completely well at 6 weeks follow-up|1008
