52 years old|0
man|0
emergency department visit|0
diffuse vesicular skin rash over the trunk|-24
contact with co-workers diagnosed as varicella infection|-96
headache|-24
sore throat|-24
nausea|-24
denied prior history of chicken pox|0
immunosuppressants|-43800
methotrexate|-43800
azathioprine|-43800
prednisolone|-43800
cutaneous leukocytoclastic vasculitis|-43800
vesicle Tzank smear|0
multinucleated giant cells|0
herpes virus infection|0
white blood cell count 4100/uL|0
hemoglobin 14.8 gm/dL|0
platelets 134000/uL|0
serum creatinine 0.62 mg/dL|0
Aspartate transaminase 782 U/L|0
Alanine transaminase 603 U/L|0
total bilirubin 0.4 mg/dL|0
prothrombin time 12.6 s|0
C reactive protein 1.45 mg/L|0
varicella zoster|0
hepatitis|0
oral famciclovir 500 mg three times per day|0
immunosuppressive drugs discontinued|0
discharged|0
outpatient clinics follow up arranged|0
emergency department visit again|48
general malaise|48
nausea|48
acute ill looking|48
alert (E4V5M6)|48
temperature 36.2 °C|48
blood pressure 54/46 mmHg|48
pulse rate 102 beats/minute|48
respiratory rate 20 cycles/min|48
white blood cell 12700/uL|48
hemoglobin 15.4 g/dL|48
platelets 61000/uL|48
prothrombin time 35.7 s|48
activated partial thromboplastin time 44.5 s|48
fibrinogen <50 mg/dL|48
AST 8989 U/L|48
ALT 6048 U/L|48
total bilirubin 2.0 mg/dL|48
indirect total bilirubin 1.5 mg/dL|48
serum creatinine 2.99 mg/dL|48
blood arterial gas analysis PH 7.31|48
CO2 23 mmHg|48
O2 83 mmHg|48
HCO3 15.1 mm/L|48
nasal cannula oxygen flow 5 L/min|48
negative Hepatitis B surface antigen (HbsAg)|48
negative antibodies against hepatitis C (anti-HCV)|48
negative anti-hepatitis A IgM antibody|48
negative Epstein-Barr virus (EBV) viral capsid antigen IgM|48
negative EBV IgG|48
negative serum Cytomegalovirus (CMV) IgM|48
negative CMV IgG|48
negative CMV pp65 antigen test|48
negative serum Herpes simplex virus IgM|48
negative HSV IgG|48
negative serum HSV DNA PCR|48
positive VZV PCR|48
vesicular base viral isolation VZV|48
serum viral isolation VZV|48
negative VZV IgM|48
negative VZV IgG|48
admitted to intensive care unit|48
septic shock|48
multiple organ failure|48
disseminated intravascular coagulopathy|48
aggressive fluid resuscitation|48
broad-spectrum empirical antibiotics|48
glycopeptide|48
carbapenem|48
blood transfusion|48
correcting anemia|48
correcting coagulopathy|48
intravenous acyclovir|48
severe VZV infection|48
clinical condition deteriorated rapidly|48
intubated|48
comatose consciousness (E2M2V1)|48
dyspnea|48
profound shock|48
brain CT not done|48
lumbar puncture not considered|48
absence of meningeal sign|48
lactate acidosis|48
expired|72
