43 years old | 0
man | 0
presented to the hospital | 0
cough | -168
high fever | -168
anosmia | -168
nasopharyngeal PCR swab taken | 0
SARS-CoV-2 positive | 0
gout | 0
hypertension | 0
chronic kidney disease (CKD-3, eGFR 55) | 0
unprovoked lower limb venous thromboembolism (VTE) | 0
lupus anticoagulant (LAC) positive in 2017 | -8760
declined anticoagulation | -8760
B2-glycoprotein IgG negative | -8760
anti-cardiolipin IgM negative | -8760
homocysteine normal | -8760
anti-thrombin III normal | -8760
protein C levels normal | -8760
admitted to intensive care | 0
intubation required | 24
respiratory failure | 24
commencement of dual vasopressors | 24
refractory shock | 24
norepinephrine max 0.28 mcg/kg/min on day 2 | 48
norepinephrine stopped by day 9 | 216
vasopressin max 0.03 units/min on day 2 | 48
vasopressin stopped on day 3 | 72
continuous renal replacement therapy | 24
COVID-19 acute respiratory distress syndrome (H-type CARDS) | 24
prone-positioning required | 24
paralysis required | 24
progression towards refractory shock | 24
rapidly deteriorating CARDS | 24
high-grade fever | 24
multidisciplinary COVID-19 team review | 24
cytokine release syndrome (CRS) considered | 24
interleukin-6 (IL-6) level >1000 pg/mL | 24
D-dimer 8.56 mcg/mL | 24
ferritin 8109 ng/mL | 24
lactate dehydrogenase 2111 U/L | 24
aspartate transaminase 1896 U/L | 24
H-score 146 | 24
tocilizumab administered | 48
hydrocortisone administered (days 2-5) | 48
no other targeted COVID-19 intervention | 48
heparin infusion started | 48
heparin continued until day 17 | 408
overt lower gastrointestinal (GI) bleeding | 408
high-volume diarrhoea | 336
rectal tube insertion | 336
CT mesenteric angiogram (CTMA) on day 17 | 408
arterial blush in the caecum | 408
thickening of the terminal ileum | 408
embolisation of the culprit branch | 408
bleeding continued on day 18 | 432
repeated CTMA | 432
active bleeding in the ascending colon | 432
second embolisation performed | 432
continued bleeding | 432
significant blood transfusion required | 432
colonoscopy on day 20 | 480
endostasis attempted | 480
erythematous friable ileal mucosa | 480
luminal bleeding | 480
colitis of the caecum | 480
ascending colon colitis | 480
large ulcerations | 480
failure of endostasis | 480
right-sided hemicolectomy | 480
segmental resection of the terminal ileum | 480
gross examination showed extensive ulceration of the terminal ileum | 480
thickened dusky wall | 480
fat encroachment | 480
mesenteric stranding | 480
caecum showed three deep linear circumferential ulcers | 480
bowel wall perforation | 480
microscopic examination revealed extensive ulceration of the terminal ileum | 480
deep fissuring ulceration of the caecum | 480
perforation | 480
irregular, branching, disordered crypts | 480
regenerative changes | 480
no thrombi within large vessels | 480
smaller vessels with fibrin microthrombi | 480
low overall thrombus burden | 480
no ischaemic changes | 480
no severe ischaemic colitis | 480
no transmural lymphoid aggregates | 480
no viral inclusions | 480
no granulomas | 480
no parasites | 480
no vasculitic changes | 480
heparin infusion stopped on day 17 | 408
vasopressors stopped by day 9 | 216
hydrocortisone prescribed for 3 days | 48
no non-steroidal anti-inflammatory drugs prescribed | 0
superimposed infective cause excluded | 0
HIV screening negative | 0
Clostridium difficile testing negative | 0
tissue bacterial culture light growth of multidrug-resistant Pseudomonas | 480
Candida glabrata light growth | 480
acid-fast smears negative | 480
molecular testing for tuberculosis negative | 480
PCR tests varicella-zoster virus negative | 480
cytomegalovirus IgM negative | 480
blood PCR for cytomegalovirus negative | 480
histological analysis for viral inclusions negative | 480
stool PCR for SARS-CoV-2 negative | 480
stoma swab PCR for SARS-CoV-2 negative | 480
