22 years old | 0
    male | 0
    admitted to intensive care unit (ICU) | 0
    fever | -240
    cough | -192
    sputum production | -192
    respiratory distress | -24
    altered sensorium | -24
    no history of hospitalization within past 1 year | -8760
    altered sensorium | 0
    tachycardic | 0
    tachypnea | 0
    hypotensive | 0
    heart rate-130/min | 0
    blood pressure-90/60 mm Hg | 0
    hypoxemia | 0
    right lower lobe consolidation | 0
    haemoglobin-9.3 g% | 0
    white blood cell (WBC) count-3,500/cu.mm | 0
    platelets-80,000/cu.mm |DISCUSSIONSince the 1990s, CA-MRSA has emerged as a major cause of skin and soft-tissue infections.[1] Centers for Disease Control and Prevention has epidemiologically defined, CA-MRSA specimens as those recovered no more than 48 h after hospitalization and from a patient without a history of hospitalization, surgery, dialysis, residence in the long-term-care facility within the past 12 months, prior MRSA infection or indwelling devices.[2]Staphylococcal pneumonia is clinically defined by the signs of lower respiratory tract infection (e.g. cough, expectoration and chest pain) and pulmonary infiltrates on chest radiograph that were not attributable to other causes, coinciding with isolation of S. aureus as the only potential pathogen by at least one of the following procedures: (1) Puncture of a pleural effusion or lung abscess, (2) culture of BAL fluid (≥103 CFU/ml), Wimberg brushing (≥102 CFU/ml) or protected tracheal aspiration (≥105 CFU/ml); and (3) blood culture yielding the same S. aureus strain as that found in tracheal secretions.[3]This entity is common in children, but rarely reported in adults. This is the first reported case of CA-MRSA from Indian subcontinent. This disease affects the young, with 80% of patients in previous reports being younger than 50 years.[1] Severe leucopenia appears to be characteristic of CA-MRSA pneumonia, with WBC counts less than 2500/cu.mm seen in 63% (5/8) cases at presentation. Our case was a young male who met the CDC epidemiologic criteria for CA-MRSA. His initial WBC counts were 3500/cu mm as explainable from previous reports that leucopenia is an ominous prognostic factor in these patients, due to affinity of Panton-Valentine leukocidin (PVL) for neutrophils leading to their lysis. It is speculated that WBC count is an inverse biomarker of the PVL burden.[4]Hemoptysis is a common finding. Presenting vital signs are severe, reflecting incipient or frank septic shock. Cavitary pulmonary infiltrates may be seen on chest radiograph or chest computed tomography. Patient presented with hypoxemia and shock. Patient lacked hemoptysis, typical of most prior case reports, also bronchoscopy showed no hemorrhage. However, computed tomography revealed diffuse cavitations and necrosis. Clinical factors associated with fatal outcome are need for artificial ventilation, inotrope support, airway bleeding, ARDS, leucopenia, low platelet count.[3] Approximately, 50% of mortality is described in the literature.[1]The Staphylococcus isolate was resistant to penicillinase-resistant penicillins, but sensitive to macrolides, quinolones, linezolid, clindamycin and vancomycin. This sensitivity pattern is characteristic of CA-MRSA and distinct from that of hospital-acquired MRSA, which typically exhibits resistance to numerous agents other than penicillinase-resistant penicillins.[4] Therapeutic options in case of severe CA-MRSA infections are vancomycin and linezolid.[5] In less severe infections, clindamycin, trimethoprim — sulphamethoxazole (TMP — SMX) and doxycycline are therapeutic options. The majority of strains remain susceptible to TMP — SMX, but more than 30% of isolates are resistant to clindamycin and doxycycline. Fluoroquinolone are not recommended because resistance to these agents develops rapidly.[5]Commercially available intravenous immune globulin, which has in vitro activity against PVL, is another treatment alternative that was not used.[4] By the time, the diagnosis of necrotizing pneumonia is made, the pathology achieved by CA-MRSA and PVL is advanced and it may be difficult to neutralize the organism and its virulence factor. In absence of microbiological data, other etiology for necrotizing lesions on chest imaging includes Klebsiella pneumonia, Pseudomonas eruginosa, Nocardia, Actinomyces and anaerobes.[4] The ability to predict etiology of pneumonia from clinical signs is limited; in the presence of shock, leucopenia and severe hypoxemia suspicion for MRSA should be kept high. Early diagnosis and intervention may be critical in improving outcomes of necrotizing pneumonia due to CA-MRSA.We recommend considering CA-MRSA among pathogens that cause community-acquired pneumonia, in patients presenting to casualty with shock, hypoxemia and leucopenia.Source of Support: NilConflict of Interest: None declared
    <|eot_id|><|start_header_id|>assistant<|end_header_id|>
    22 years old | 0
    male | 0
    admitted to intensive care unit (ICU) | 0
    fever | -240
    cough | -192
    sputum production | -192
    respiratory distress | -24
    altered sensorium | -24
    no history of hospitalization within past 1 year | -8760
    altered sensorium | 0
    tachycardic | 0
    tachypnea | 0
    hypotensive | 0
    heart rate-130/min | 0
    blood pressure-90/60 mm Hg | 0
    hypoxemia | 0
    right lower lobe consolidation | 0
    haemoglobin-9.3 g% | 0
    white blood cell (WBC) count-3,500/cu.mm | 0
    platelets-80,000/cu.mm | 0
    serum creatinine-1.8 mg/dl | 0
    normal liver function test | 0
    normal general blood picture | 0
    intubated | 0
    mechanical ventilation | 0
    bronchoalveolar lavage (BAL) | 0
    blood samples sent for culture and sensitivity testing | 0
    provisional diagnosis of acute febrile illness | 0
    pneumonia | 0
    septic shock | 0
    started on piperacillin-tazobactum | 0
    vancomycin | 0
    antimalarials | 0
    tests for malaria | 0
    tests for leptospirosis | 0
    tests for dengue | 0
    tests for typhoid | 0
    all tropical infective profile tests negative | 0
    PaO2/FiO2 ratios 100 | 0
    ventilated as per acute respiratory distress syndrome (ARDS) net protocol | 0
    prone ventilation | 0
    blood cultures positive for MRSA | 0
    BAL cultures positive for MRSA | 0
    i.v. vancomycin added | 0
    PaO2/FiO2 ratios improved (P/F > 300) | 168
    extubated | 168
    continuing hypoxia | 168
    respiratory rate of 28-30/min | 168
    computed tomography pulmonary angiogram | 96
    high resolution computed tomography chest | 96
    patchy consolidation with cavity in lateral basal segment of right lower lobe | 96
    pulmonary angiogram normal | 96
    continued on vancomycin for 3 weeks | 168
    respiratory rate settled | 672
    discharged after 28 days of ICU stay | 672
    diffuse consolidation with air bronchograms | 96
    consolidation and areas of cavitation | 96
    right-sided pleural effusion | 96
    no hemoptysis | 0
    bronchoscopy showed no hemorrhage | 0
    diffuse cavitations and necrosis | 96
    MRSA resistant to penicillinase-resistant penicillins | 0
    MRSA sensitive to macrolides | 0
    MRSA sensitive to quinolones | 0
    MRSA sensitive to linezolid | 0
    MRSA sensitive to clindamycin | 0
    MRSA sensitive to vancomycin | 0
    leucopenia | 0
    low platelet count | 0
    septic shock | 0
    severe hypoxemia | 0
    cavitary pulmonary infiltrates | 96
    no airway bleeding | 0
    ARDS | 0
    inotrope support | 0
    artificial ventilation | 0
    leucopenia | 0
    low platelet count | 0
    severe leucopenia | 0
    WBC counts less than 2500/cu.mm | 0
    leucopenia as ominous prognostic factor | 0
    Panton-Valentine leukocidin (PVL) affinity for neutrophils leading to lysis | 0
    WBC count as inverse biomarker of PVL burden | 0
    no prior MRSA infection | -8760
    no indwelling devices | -8760
    CA-MRSA pneumonia | 0
    necrotizing pneumonia | 0
    multiorgan failure | 0
    shock | 0
    hypoxemia | 0
    leucopenia | 0
    severe hypoxemia | 0
    leucopenia | 0
    shock | 0
    cavitary pulmonary infiltrates | 96
    no pulmonary embolism | 96
    patchy consolidation | 96
    cavity in right lower lobe | 96
    right-sided pleural effusion | 96
    no Klebsiella pneumonia | 0
    no Pseudomonas aeruginosa | 0
    no Nocardia | 0
    no Actinomyces | 0
    no anaerobes | 0
    community-acquired pneumonia | 0
    CA-MRSA | 0
    <|eot_id|>