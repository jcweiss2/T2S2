76 years old | 0
female | 0
renal transplant | 0
admitted to ICU | 0
coma | 0
respiratory distress | 0
methylprednisolone | 0
tacrolimus | 0
mycophenolate mofetil | 0
candesartan | 0
arterial hypertension | 0
serum creatinine concentration 1.70 mg/dl | 0
estimated glomerular filtration rate 28 ml/min/1.73 m2 | 0
HBV reactivation | -432
HBV DNA copies/ml 109 | -432
dyspnea | -288
bilateral lung infiltrates | -288
CMV pneumonia | -288
quantitative CMV PCR 3130 copies/ml | -288
intravenous sodium ganciclovir | -288
ganciclovir 200 mg | -288
ganciclovir 400 mg | -276
white blood cell count 5080/mm3 | -288
white blood cell count 3430/mm3 | -276
renal function deterioration | -276
creatinine 2.67 mg/dl | -276
estimated GFR 17 ml/min/1.73 m2 | -276
hip fracture | -276
orthopedic surgery | -276
epidural anesthesia | -276
altered consciousness | -12
respiratory distress | -12
arterial blood gas analysis | -12
pH 6.79 | -12
pCO2 54 mm Hg | -12
bicarbonate 8 mmol/l | -12
lactate 20 mmol/l | -12
intubation | -12
mechanical ventilation | -12
intravenous sodium bicarbonate | -12
thiamine supplementation | -12
continuous venovenous hemofiltration | -12
arterial pH 7.31 | -6
central venous oxygen saturation 61.5% | -6
echocardiography | -6
left ventricular function preserved | -6
arterial lactate 27 mmol/l | -6
pyruvate 0.6 mmol/l | -6
L/P molar ratio 45 | -6
hypoglycemia | -6
dextrose 30% | -6
biological signs of ketogenesis | -6
urinary excretion of 3-hydroxybutyrate 256.2 mmol/mol creatinine | -6
dicarboxylic acids | -6
ganciclovir discontinued | 0
rhabomyolysis | 12
vasoplegia | 12
blood cultures sterile | 12
abdominal CT | 12
no bowel ischemia | 12
hyperlactatemia | 12
liver tests moderately disturbed | 12
ammonia level 109 μg/dl | 12
encephalopathy | 12
brain CT normal | 12
fatality | 14
hospital day 14 | 14