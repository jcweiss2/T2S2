65 years old | 0
    female | 0
    stage IIIA lung cancer | -16200
    abdominal pain | 0
    pancreatic head lesion | 0
    smoking history of greater than 40 pack years | 0
    hypertension | 0
    hypothyroidism | 0
    dyslipidemia | 0
    spiculated suprahilar 4.5 × 2.6 cm right upper lobe nodule | -16200
    multiple sub-centimeter left lung nodules | -16200
    lung-RADS 4X | -16200
    augmented activity in the RUL mass | -16200
    NSCLC | -16200
    adenocarcinoma | -16200
    lymph node sampling negative for nodal involvement | -16200
    T4N0M0 | -16200
    Program death ligand-1 expression 15% | -15840
    encasement of the pulmonary artery | -16200
    encasement of the superior vena cava | -16200
    7 rounds of carboplatin and paclitaxel | -16200
    8 rounds of radiation therapy | -16200
    decrease in the RUL mass from 4.5 × 2.6 cm to 3.5 × 2.1 cm | -14160
    adjuvant immunotherapy with durvalumab | -14160
    3 rounds of durvalumab | -14160
    pneumonitis | -14160
    steroid taper | -14160
    increase in the RUL mass to 5.0 × 2.8 cm | -14160
    increase in the RUL mass to 6.5 × 2.2 cm | -14160
    respiratory symptom management | -14160
    radiation oncology clinic follow-up | -14160
    hematology-oncology clinic follow-up | -14160
    thoracic, abdominal, and pelvic CT scan | -14160
    stable lung nodules | -14160
    radiation fibrosis | -14160
    epigastric pain | -840
    constipation | -840
    loss of appetite | -840
    weight loss | -840
    abdominal and pelvic CT scan showing pancreatic head mass | -840
    pancreatic ductal dilatation to 7 mm | -840
    endoscopic ultrasound-guided biopsy of the pancreatic head mass | -840
    tumor cells with nuclear pleomorphism | -840
    prominent nucleoli | -840
    irregular nuclear contours | -840
    coarse chromatin | -840
    CK7 positivity | -840
    TTF-1 positivity | -840
    Napsin-A positivity | -840
    negative for CDX-2 | -840
    negative for KOC | -840
    negative for synaptophysin | -840
    mixed Smad-4 staining pattern | -840
    morphologically similar to original lung adenocarcinoma | -840
    lung adenocarcinoma metastasized to the pancreas | -840
    AST 35 U/L | -840
    ALT 23 U/L | -840
    ALP 74 U/L | -840
    total bilirubin 0.5 mg/dL | -840
    direct bilirubin 0.2 mg/dL | -840
    CA 19.9 22.5 U/mL | -840
    PET/CT scan showing FDGC-avid pancreatic head mass | -840
    SUV max of 13.3 | -840
    increased uptake in the porta hepatis | -840
    SUV max of 4.2 | -840
    no other regions of metastases | -840
    no lymphadenopathy | -840
    brain MRI scan negative for intracranial metastasis | -840
    palliative radiation therapy to the pancreatic mass | 0
    combination chemotherapy with carboplatin and pemetrexed | 0
    3 cycles of chemotherapy | 720
    admitted for generalized weakness | 720
    dyspnea at rest | 720
    electrolyte derangements | 720
    acute anemia with hemoglobin 6.9 g/dL | 720
    transfusion | 720
    new 9 mm left lower lobe nodule | 720
    decreased metabolic activity in the pancreatic mass | 1080
    metabolic activity in the new left lower lobe nodule | 1080
    uncertainty regarding treatment continuation | 1080
    no further treatments | 1080
    saturating at 87% on 3 L oxygen | 2160
    use of accessory muscles | 2160
    blood pressure 84/70 | 2160
    heart rate 138 | 2160
    increased dyspnea | 2160
    cough | 2160
    generalized weakness | 2160
    right lung consolidation | 2160
    loculated pleural effusion | 2160
    acute hypoxic respiratory failure | 2160
    sepsis secondary to pneumonia | 2160
    vancomycin | 2160
    azithromycin | 2160
    cefepime | 2160
    oxygen supplementation | 2160
    altered mentation | 2160
    worsening hypoxemia | 2160
    vasopressor support | 2160
    bilevel-positive airway pressure | 2160
    transition to inpatient hospice care | 2160
    passed peacefully under comfort measures | 2160