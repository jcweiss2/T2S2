41 years old | 0
male | 0
unconscious | -240
multiple trauma | -240
admitted to the hospital | 0
respiratory failure | -240
sepsis | -240
hypotension | -240
vasopressors | -240
hematemesis | -240
drop of hemoglobin | -240
transfusions of packed red blood cells | -240
upper endoscopy | -240
large cratered ulcer | -240
visible bleeding vessel | -240
epinephrine injection | -240
bipolar cautery | -240
hemostasis | -240
vasopressor requirements decreased | -216
hemoglobin 8.5 g/dL | -216
hypotensive | -192
hemoglobin 5.8 g/dL | -192
computed tomography angiogram | -192
selective arteriograms | -192
extravasation of contrast | -192
coil embolization | -192
active bleeding | -192
salvage surgery | -192
laparotomy | -192
duodenotomy | -192
suture ligation | -192
repeat endoscopy | -168
new large ulcer | -168
spurting vessel | -168
epinephrine injection | -168
thermocoagulation | -168
oozing from the ulcer | -168
placement of hemostatic clips | -168
endoscopic sutures | -168
OverStitch endoscopic suture system | -168
interrupted suture | -168
running suture | -168
hemostasis | -168
discharge to subacute rehabilitation | 240
hemoglobin 8.1 g/dL | 240
negative Helicobacter pylori serology | 240
follow-up telephone call | 8760
no further gastrointestinal bleeding | 8760