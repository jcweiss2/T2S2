66 years old | 0\
male | 0\
admitted to the hospital | 0\
intermittent high-grade fever | -72\
generalized dull-aching abdominal pain | -72\
passing turbid urine | -240\
decrease in urine output | -240\
swelling of both feet | -240\
treated with intravenous medications | -168\
type II diabetes mellitus | -2628\
conscious | 0\
afebrile | 0\
tachycardic | 0\
heart rate of 136/min | 0\
blood pressure was 110/70 mmHg | 0\
renal angle tenderness bilaterally | 0\
high total leukocyte counts | 0\
left shift | 0\
elevated urea | 0\
elevated creatinine levels | 0\
pyuria | 0\
leukocyte esterase positivity | 0\
prolonged activated partial thromboplastin time | 0\
enlarged kidneys | 0\
bilateral renal abscesses | 0\
emergency ultrasound-guided drainage of renal abscesses | 24\
transfusion of blood products | 24\
coagulopathy | 24\
initiated on intravenous meropenem | 0\
pus smear from renal abscesses showed septate fungal hyphae | 24\
initiated on intravenous voriconazole | 24\
initiated on intravenous amphotericin B | 24\
cultures from both renal abscesses revealed growth of Aspergillus fumigatus | 48\
worsening renal function | 48\
acute pulmonary edema | 48\
hyperkalemia | 48\
metabolic acidosis | 48\
initiated on hemodialysis | 48\
initiated on noninvasive ventilation | 48\
sudden cardiac arrest | 216\
aspiration | 216\
succumbed to his illness | 216