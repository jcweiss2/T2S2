80 years old | 0
male | 0
admitted to the hospital | 0
peripheral artery disease | 0
hypertension | 0
end stage renal disease | 0
on peritoneal dialysis | 0
hypotension | 0
denies chest pain | 0
denies shortness of breath | 0
denies fever | 0
denies cough | 0
denies palpitation | 0
denies nausea | 0
denies vomiting | 0
denies abdominal pain | 0
denies changes in urinary or bowel habits | 0
blood pressure 63/29 | 0
pulse 72/min | 0
temperature 97.2 F | 0
WBC count 16.5 K/UL | 0
Hgb 14.3 GM/DL | 0
PLT 115 K | 0
Creatinine 12.59 MG/DL | 0
BUN 56 MG/DL | 0
Sodium 133 MMOL/L | 0
Potassium 5.4 MMOL/L | 0
BNP 143 PG/ML | 0
Troponin 0.05 NG/ML | 0
ST segment elevation in lead V3, V4 and V5 | 1
Q wave in lead II, III and AVF | 1
diagnosis of acute ST elevation MI | 1
oral aspirin 325 mg | 1
clopidogrel 300 mg | 1
atorvastatin 80 mg | 1
heparin 3500 units/kg | 1
emergent cardiac catheterization | 1
coronary angiography | 1
chronic total right coronary artery occlusion | 1
collaterals from left | 1
patent left coronary arteries | 1
left ventriculography | 1
wall motion abnormalities | 1
mid to apical akinesis | 1
basal hyperkinesis | 1
transferred to ICU | 1
levophed pressure support | 1
CK-MB 11.6 ng/ml | 4
Troponin 2.10 | 4
resolution of ST elevation in anterior leads | 6
broad spectrum antibiotics | 6
vancomycin | 6
Zosyn | 6
leukocytosis | 6
hypotension | 6
septic shock | 6
cardiogenic shock | 6
transthoracic echocardiography | 12
left ventricular ejection fraction 25-30% | 12
elevated left ventricular end diastolic pressure | 12
akinesis of left and right ventricle | 12
except in the basal region | 12
repeat echocardiogram | 24
sessile LV thrombus | 24
akinesis of both left and right ventricles | 24
except in the basal region | 24
anticoagulation with heparin | 24
died | 72
biventricular takotsubo cardiomyopathy | 0
LV thrombus | 24