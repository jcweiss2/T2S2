38 years old | 0
male | 0
admitted to the hospital | 0
chondrosarcoma | -672
involving the right second to fifth ribs | -672
extension into the anterior chest wall | -672
mild compressive atelectasis | -672
wide local excision of the lesion | 0
anterior chest wall defect | 0
missing ribs | 0
exposed cardiopulmonary structures | 0
rib cage reconstruction | 0
double-folded polypropylene mesh | 0
anchored using No. 1 prolene | 0
soft tissue reconstruction | 0
free anterolateral thigh flap (ALT) | 0
nipple areola complex (NAC) harvested | 0
free graft from the excised specimen | 0
secured to the flap with a bolster dressing | 0
intraoperative hemodynamic instability | 0
endotracheal tube | 0
noradrenaline | 0
injection vasopressin | 48
hemodynamic instability worsened | 48
spontaneous breathing trials (SBT) | 24
unsuccessful weaning from ventilator support | 24
pneumothorax detected | 24
chest tube inserted | 24
echocardiogram | 24
normal left ventricular ejection fraction | 24
antibiotics escalated | 48
blood culture came negative | 48
afebrile | 48
vacuum dressing applied | 120
polyurethane sponge and film at −125 mm Hg | 120
improvement in breathing mechanics | 120
reduced requirement of positive end expiratory pressure (PEEP) | 144
better tolerance of SBT and pressure support ventilation (PSV) | 144
extubated | 192
transitioned to high-flow nasal cannula | 192
shifted out of ICU | 240
removal of vacuum dressing | 264
flap, suture line, and free NAC graft were healthy | 264
discharged | 264
NPWT stopped | 360
minimal residual paradoxical breathing | 360
no discomfort in breathing | 360