2 years old | 0
male | 0
father had fever and exanthema | -720
father's disease remained undiagnosed | -720
contact with two dogs | 0
normal weight at birth | 0
breastfeed for six months | 0
vaccination was up to date | 0
fever | -72
nimesulide and amoxicilin | -72
pallor | -69
leucopenia | -66
anemia | -66
thrombocytopenia | -66
admission | 0
hypoalbuminemia | 2
high liver enzymes | 2
prolongation of coagulation times | 2
hyponatremia | 2
elevation of the C reactive protein | 2
enlarged lymph nodes | 2
hepatomegaly | 2
splenomegaly | 2
erythematous, macular, non-itching rash | 2
left inguinal adenopathy | 2
coughs | 2
bone marrow aspiration | 2
activated lymphocytes | 2
cytopenia | 7
anemia | 7
deep neutropenia | 7
thrombocytopenia | 7
hemorrhagic syndrome | 7
multiple transfusions | 7
liver failure | 14
incoagulable prothrombin time | 14
persistent hypoalbuminemia | 14
lactate dehydrogenase peaked | 14
serological tests for HIV, Epstein-Barr virus, Hepatitis A, B and C virus, Toxoplasma gondii, cytomegalovirus, rubella virus, herpes simplex, Treponema pallidum | 14
Weil-Felix reactions | 14
bone marrow biopsy | 14
cellularity of 70% | 14
inverted myeloid-erythroid ratio | 14
myeloid hypoplasia | 14
erythroid series hyperplasia | 14
megakaryocytic series | 14
histiocytes with hemophagocytosis | 14
lymph node biopsy | 14
ganglionic sinus partially infiltrated by histiocytic cells | 14
loss of architecture | 14
hyperplasic lymphoid follicle | 14
immunohistochemistry for Langerhans cells histiocytosis | 14
doxycycline | 21
remission of fever | 23
improvement of the general condition | 23
new fever peaks | 25
jaundice | 25
asthenia | 25
increased triglycerides | 25
persistence of cytopenia | 25
low fibrinogen levels | 25
Leptospira interrogans infection ruled out | 25
diagnosis of hemophagocytic lymphohistiocytosis | 25
steroids management | 25
methylprednisolone | 25
DNA extraction | 25
nested polymerase chain reaction for the 17-kDA gene of Rickettsia spp. | 25
in-house indirect immunofluorescence assay for IgM and IgG against Rickettsia rickettsii and Rickettsia typhi | 25
seroconversion | 32
hemorrhagic syndrome | 28
persistence of low fibrinogen levels | 28
petechiae | 28
gingivorrhagia | 28
admission to the Pediatric intensive care unit | 28
neurological and respiratory deterioration | 28
antimicrobial management | 28
Meropenem | 28
vancomycin | 28
amphotericin B | 28
nosocomial sepsis suspected | 28
doxycycline suspended | 28
dexamethasone | 33
poor response | 33
abdominal ultrasound | 33
diffuse hepatic and kidney damage | 33
altered cortex-marrow relationship | 33
hyperechoic pattern | 33
ascites | 33
urine output decreased | 38
neurological and hemodynamic sudden worsening | 38
mechanical ventilation | 38
vasopressor drugs | 38
alveolar diffuse hemorrhage | 38
anuria | 38
death | 41
post-mortem histopathological test | 41
lymph node biopsy | 41
immunohistochemistry | 41
positive result for Rickettsia | 41