53 years old | 0
man | 0
arterial hypertension | 0
dyslipidemia | 0
previous myocardial infarction | 0
coronary bypass surgery | -58560
admitted to the emergency department | 0
mild COVID-19 | -240
severe and sharp abdominal pain | -48
abdominal pain located in the epigastrium | -48
abdominal pain worsening in intensity | -24
fever | -48
no nausea | 0
no vomit | 0
no abnormal bowel movements | 0
no other respiratory symptoms | 0
no urinary complaints | 0
febrile | 0
stable patient | 0
blood pressure 125/82 mmHg | 0
heart rate 89 bpm | 0
normal cardiopulmonary auscultation | 0
abdomen non-distended | 0
tender mass in the epigastrium | 0
localized guarding | 0
hypoactive bowel sounds | 0
non-metallic bowel sounds | 0
no abdominal hernias | 0
normal white blood cell count | 0
segmented neutrophils 72.9% | 0
hemoglobin 13.80 g/dl | 0
d-dimer 0.94 μg/ml | 0
normal hepatobiliopancreatic parameters | 0
normal cardiac parameters | 0
normal renal parameters | 0
normal urinalysis | 0
normal arterial-blood gas test | 0
computed tomography scan with intravenous contrast | 0
short segment of small bowel with inflammatory signs | 0
localized free peritoneal fluid | 0
residual ground-glass opacities related to COVID-19 | 0
ruled out cholecystitis | 0
ruled out pancreatitis | 0
ruled out perforation of hollow viscus | 0
diagnostic exploratory laparotomy | 0
therapeutic exploratory laparotomy | 0
suppurative Meckel’s diverticulitis | 0
local abscess | 0
drainage | 0
segmental ileal resection | 0
primary anastomosis | 0
intravenous antibiotics | 0
no further rises in temperature | 0
no complications | 144
discharged | 144
active inflammation | 0
gangrenous Meckel’s diverticulum | 0
