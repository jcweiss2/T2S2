50 years old | 0
    male | 0
    admitted to the hospital | 0
    perianal swelling | 0
    discomfort | 0
    anal pain | -144
    discomfort | -144
    no obvious cause | -144
    no abdominal pain | -144
    no bleeding during defecation | -144
    visited local hospital | -48
    pain | -48
    diagnosed perianal abscess | -48
    incision and drainage | -48
    perianal swelling not subsided | -24
    spread to base of scrotum | -24
    local incision showed yellowish gray necrotic tissue | -24
    fishy odor | -24
    high fever | -24
    body temperature 38.2 °C | 0
    respiratory rate 21 breaths/min | 0
    heart rate 81 beats/min | 0
    blood pressure 105/69 mmHg | 0
    dysuresia | 0
    denied underlying diseases | 0
    no type 2 diabetes | 0
    no malignancy | 0
    no other common diseases | 0
    entire anal margin swollen | 0
    skin red and black | 0
    previous incision on posterior anal margin with yellow-white frothy secretions | 0
    severe pain | 0
    skin sides and base of scrotum tender and warm | 0
    crepitus when palpating left pubic symphysis | 0
    white cell count 14.29 × 109/L | 0
    neutrophils 85.10% | 0
    lymphocytes 6.70% | 0
    monocytes 8.00% | 0
    eosinophils 0.10% | 0
    hemoglobin 123.00 g/L | 0
    hematocrit 34.90% | 0
    platelet count 135.00 × 109/L | 0
    C-reactive protein 126.40 mg/L | 0
    sodium 140.40 mmol/L | 0
    potassium 3.50 mmol/L | 0
    chloride 101.20 mmol/L | 0
    calcium 2.11 mmol/L | 0
    urea nitrogen 7.08 mmol/L | 0
    creatinine 81.30 μmol/L | 0
    glucose 7.02 mmol/L | 0
    alanine aminotransferase 35.00 U/L | 0
    aspartate aminotransferase 35.00 U/L | 0
    albumin 33.70 g/L | 0
    D-dimer 7.30 mg/L | 0
    lower abdominal and pelvic CT scan showing gas in tissue | 0
    urine retention | 0
    multiple lymph nodes inguinal area | 0
    diagnosed perianal and perineal necrotizing fasciitis | 0
    aggravated by inadequate drainage | 0
    surgery under spinal anesthesia | 0
    urethra catheter surgery | 0
    lithotomy position | 0
    defect in anal gland near posterior dentate line | 0
    primary opening | 0
    previous wound connected | 0
    internal opening resource of infection | 0
    cryptoglandular infection | 0
    main incision excised and debrided | 0
    probe and clamp used to explore infection area | 0
    scissors and diathotomy used to remove necrotic tissues | 0
    multiple incisions performed | 0
    rubber catheters as loose setons | 0
    incision outside bilateral symphysis pubis | 0
    21 loose rubber setons | 0
    scrotum skin kept intact | 0
    transferred to intensive care unit | 0
    fourth-generation cephalosporin | 0
    metronidazole | 0
    human blood albumin | 0
    vitamins | 0
    lipids | 0
    daily laboratory examination | 0
    wound cleaned and changed daily | 0
    surgical area rinsed with hydrogen peroxide and oxygenate | 0
    necrotic tissue trimmed | 0
    rubber setons removed after no pus | 0
    necrotic perineal skin completely removed | 72
    CT scan showed loose setons | 72
    small amount of gas shadow | 72
    catheter drainage | 72
    final drainage incision at right groin and pubic symphysis | 72
    perianal MRI | 168
    stable laboratory results | 168
    transferred to general ward | 168
    antibiotic treatment stopped | 168
    nutrition support continued | 168
    daily dressing changes | 168
    clinically improved | 336
    discharged | 336
    outpatient follow-up once a week | 336
    wounds healed at 3 weeks post-discharge | 504
    perianal morphology retained | 504
    anorectal manometry results recovered | 504
    cured | 504
    satisfied with treatment | 504

    <|eot_id|>
    