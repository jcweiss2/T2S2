16-year-old | 0
boy | 0
admitted to a local hospital | 0
history of severe fatigue | -168
CT revealed large anterior mediastinal tumor | 0
hepatosplenomegaly | 0
multiple lymph node swelling | 0
diagnosed with T-lymphoblastic lymphoma | 0
treated with multiple cytotoxic agents | 0
refractory to initial treatment | -168
transferred to our hospital | 0
Eastern Cooperative Oncology Group performance status 1 | 0
vital signs within normal range | 0
physical examination detected mild hepatosplenomegaly | 0
electrocardiogram showed normal sinus rhythm | 0
normal range of voltage of R waves at V5 lead | 0
serum brain natriuretic peptide concentration 17.2 pg/mL | 0
transthoracic echocardiography showed 59.8% LVEF | 0
no wall motion asynergy | 0
no valvular dysfunction | 0
therapeutic courses before allo-HCT | 0
induction phase | 0
PR | 0
CPA 750 mg/m2 | 0
DXR 50 mg/m2 | 0
VCR 2 mg/body | 0
PSL 60 mg/m2 | 0
LD-asp 6000 U/m2 | 0
IT | 0
consolidation phase | 0
SD | 0
THP-ADR 25 mg/m2 | 0
Ara-C 75 mg/m2 | 0
6-MP 50 mg/m2 | 0
sanctuary phase | 0
PD | 0
MTX 3000 mg/m2 | 0
re-induction phase | 0
PSL 90 mg/m2 | 0
DNR 50 mg/m2 | 0
LD-asp 5000 U/body | 0
ETP 100 mg/m2 | 0
bridging to conditioning | 0
DXR 40 mg/m2 | 0
CPA 500 mg/m2 | 0
RT 20 Gy/10 fr | 0
conditioning regimen | 0
ETP 15 mg/kg | -240
CPA 60 mg/kg | -240
TBI 12 Gy/6 fr | -240
cord blood cell transplantation | 0
continuous intravenous tacrolimus administered | 0
no infectious diseases detected in pre-conditioning period | -96
fever 38.6°C | -96
treated with meropenem | -96
fever resolved | -96
high fever | 48
septic shock caused by Gram-positive cocci | 72
administered vancomycin | 72
transferred to ICU | 72
treated with circulatory assisting agents | 72
respiratory condition worsened | 144
required mechanical ventilation | 144
LVEF rapidly decreased to 10.3% | 144
AHF diagnosed | 144
TTE suggested left ventricular wall thickness | 144
ECG showed decrease in voltage of R waves at V5 lead | 144
increase in dobutamine dose | 144
addiction to milrinone | 144
heart rate up to 160 per minute | 144
body temperature 38-41°C | 144
treated with 1.2 mg/kg/day methylprednisolone | 288
fever did not subside | 288
serum BNP concentration increased to 2764 pg/mL | 384
serum troponin I concentration 2018 pg/mL | 624
CAD placement considered | 624
CAD use not considered | 624
LVEF maintained at 10% to 25% | 624
dobutamine 5 γ | 624
milrinone 0.45 γ | 624
heart failure progressing from acute to chronic phase | 624
start treatment for chronic heart failure | 624
dose reduction of dobutalone not allowed | 624
treated with ivabradine 5 mg/day | 624
heart rate decreased | 672
blood pressure maintained | 672
BNP level decreased | 672
reduce dose of circulatory assisting agents | 672
carvedilol 1.25 mg/day added | 768
doses of ivabradine and carvedilol increased | 768
dobutamine and milrinone decreased | 768
ceased administration of dobutamine and milrinone | 1416
discharged from ICU | 1416
withdrawn from ventilator | 2040
engraftment recognized | 456
neutrophils engraftment | 456
red blood cells engraftment | 960
platelets engraftment | 1248
grade 3 acute graft-versus-host disease | 888
treated with 2 mg/kg/day mPSL | 888
serum troponin I concentration decreased to 530 pg/mL | 840
LVEF improved to 45.7% | 3432
ECG improvements in voltage of R waves at V5 lead | 3432
died of relapsed lymphoma | 4032
