65 years old | 0\
male | 0\
admitted to the hospital | 0\
shortness of breath | -96\
fever | -96\
dry cough | -96\
fatigue | -96\
breath sounds were reduced in the lower segments of the lungs | 0\
oxygen saturation (SpO2) was 93% | 0\
bilateral peripheral ground-glass attenuation and patchy consolidation | 0\
lung involvement was 60%-70% | 0\
nasopharyngeal SARS-CoV-2 RT-PCR test was positive | 0\
increased temperature | 0\
saturation with free breathing decreased to 90% | 0\
white cell count: 7.93 х 109/ L | 0\
hemoglobin 159 g/l | 0\
platelet count: 468 × 109/l | 0\
Westergren ESR 41 mm/h | 0\
interleukine 6 102 pg/ml | 0\
С-reactive protein 142 mg/l | 0\
ferritin 939.92 μg/ml | 0\
D-dimer 609 ng/ml | 0\
procalcitonin 0,11 ng/ml | 0\
treatment of SARS-CoV-2 infection included dexamethason | 0\
treatment of SARS-CoV-2 infection included heparin | 0\
treatment of SARS-CoV-2 infection included tocilizumab | 0\
treatment of SARS-CoV-2 infection included acetylcysteine | 0\
treatment of SARS-CoV-2 infection included pantoprazole | 0\
treatment of SARS-CoV-2 infection included nadroparin calcium | 0\
oxygen supplementation through the simple face mask with a flow rate of 4 l/min | 0\
air and pleural effusion in the right pleural cavity with collapse of the right lung | 360\
thoracentesis and thoracostomy in the 6th intercostal space on the mid-axillary line | 360\
1400 ml of a yellowish opaque liquid was evacuated from the pleural cavity | 360\
linezolid and imipenem/cilastatin therapy was initiated | 360\
oxygen supplementation through the simple face mask with flow rate of 8-10 l/min | 360\
pleural effusion with gas bubbles extended along the posterior and inferior walls of the right hemithorax | 432\
right lung was reduced in volume by half | 432\
focal area of subpleural infiltration with a central cavity of destruction up to 6.5 mm in diameter | 432\
air layer up to 47 mm of anteroposterior thickness was revealed along the anterior chest wall | 432\
radiological sings of the left side hydropneumothorax | 432\
pleural fluid analysis confirmed an exudative lymphocytic-rich effusion | 432\
gram-negative bacteria as Acinetobacter baumannii and Pseudomonas aeruginosa were cultured | 432\
urine culture was positive for Klebsiella pneumonia | 432\
needle thoracocentesis and new pleural drainage in the second intercostal space on the midclavicular line | 504\
air and creamy purulent mass have been aspirated | 504\
200 to 800 ml of serofibrinous hemorrhagic fluid was drawn daily through 2 drainage tubes | 504\
diagnosis of pleural empyema was confirmed | 576\
transferred to the Surgical Department | 576\
right pleural space was daily irrigated with antiseptic solutions | 576\
lung expansion was achieved by continuous vacuum aspiration technique | 576\
encapsulated pleural effusion located in the upper anterior area of the right hemithorax | 736\
ultrasound-guided puncture of this effusion was performed | 736\
new drainage of the pleural cavity was installed | 736\
4-week antibiotic therapy | 736\
discharged from the hospital | 1008\
oxygen saturation (SpO2) was 97% on room air | 1008\
chest CT after chest tube removing showed the presence of a small amount of fluid in the right pleural cavity | 1008\
lab test scores came back to normal range | 1008\
level of С-reactive protein was 11.7 mg/l | 1008\
procalcitonin − < 0,1 ng/ml | 1008