29 years old | 0
male | 0
cardiogenic shock | -168
biventricular failure | -168
ejection fraction 5–10% | -168
myopericarditis | -168
constrictive physiology | -168
PICC line placed | -168
milrinone | -168
septic shock | 0
fever | 0
chills | 0
tachycardia | 0
hypotension | 0
PICC line removed | 0
vancomycin | 0
piperacillin/tazobactam | 0
vasopressor support | 0
Chryseobacterium indologenes | 48
ciprofloxacin | 48
piperacillin/tazobactam | 48
pericardiectomy | 240
discharged | 336
follow-up | 744
NYHA Class I | 744
no evidence of recurrent infection | 744
biventricular failure | -168
non-ischaemic cardiomyopathy | -168
myopericarditis | -168
constrictive pericarditis | -168
NYHA Class II symptoms | -168
home milrinone | -168
fevers/chills | 0
fatigue | -168
dyspnoea on exertion | -168
cardiomegaly | -168
dilated right atrium | -168
passive hepatic congestion | -168
right ventricular failure | -168
pericardial calcification | -168
atrial flutter with rapid ventricular response | -168
radiofrequency ablation | -168
inotrope therapy | -168
furosemide | -168
losartan | -168
metoprolol succinate | -168
milrinone | -168
spironolactone | -168
tachycardia | 0
fever | 0
hypotension | 0
elevated lactate level | 0
septic shock | 0
catheter-related bloodstream infection | 0
pericardiectomy | 240
dense areas of adhesions | 240
calcium | 240
adhesions taken down | 240
complete removal of the pericardium | 240
left ventricular EF increased | 288
right ventricular systolic dysfunction improved | 288
inotrope independent | 336
guideline-directed medical therapy for heart failure with reduced EF | 336
furosemide | 336
metoprolol succinate | 336
sacubitril-valsartan | 336