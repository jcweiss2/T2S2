74 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
hypertension | 0 | 0 | Factual
diabetes mellitus | 0 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
intermittent subjective fever | -96 | 0 | Factual
rigors | -96 | 0 | Factual
generalized headache | -96 | 0 | Factual
altered mentation | -96 | 0 | Factual
body malaise | -96 | 0 | Factual
nausea | -96 | 0 | Factual
vomiting | -96 | 0 | Factual
no history of loss of consciousness | 0 | 0 | Negated
no abdominal pain | 0 | 0 | Negated
no change in stool habits/urine color | 0 | 0 | Negated
no recent trauma or falls | 0 | 0 | Negated
febrile | 0 | 0 | Factual
tachypneic | 0 | 0 | Factual
disoriented | 0 | 0 | Factual
good nutritional status | 0 | 0 | Factual
not jaundiced | 0 | 0 | Negated
not cyanosed | 0 | 0 | Negated
pulse rate of 103 beats/min | 0 | 0 | Factual
respiratory rate of 23 breaths/min | 0 | 0 | Factual
blood pressure of 96/60 mmHg | 0 | 0 | Factual
saturating at 98% on room air | 0 | 0 | Factual
normal vesicular breath sounds | 0 | 0 | Factual
normal abdominal examination | 0 | 0 | Factual
IV resuscitation | 0 | 0 | Factual
analgesia | 0 | 0 | Factual
WBC of 8.2 × 103/μL | 0 | 0 | Factual
hemoglobin of 11.5 g/dL | 0 | 0 | Factual
thrombocytopenia of 46,000/mm3 | 0 | 0 | Factual
elevated creatinine 117 μmol/L | 0 | 0 | Factual
BUN 10.5 mmol/L | 0 | 0 | Factual
slightly low sodium of 131 mmol/L | 0 | 0 | Factual
normal serum electrolytes | 0 | 0 | Factual
normal liver profile | 0 | 0 | Factual
normal coagulation profile | 0 | 0 | Factual
normal chest X-ray | 0 | 0 | Factual
P. falciparum with high parasitemia | 0 | 0 | Factual
admitted to the ICU | 0 | 0 | Factual
intravenous artesunate-based regimen | 0 | 72 | Factual
supportive measures | 0 | 72 | Factual
improvement in clinical status | 72 | 72 | Factual
improvement in lab parameters | 72 | 72 | Factual
shifted to the general ward | 72 | 72 | Factual
acute abdomen | 120 | 120 | Factual
progressive abdominal pain | 120 | 120 | Factual
nausea | 120 | 120 | Factual
non-bilious vomiting | 120 | 120 | Factual
anxious | 120 | 120 | Factual
afebrile | 120 | 120 | Factual
diaphoretic | 120 | 120 | Factual
tachycardic | 120 | 120 | Factual
tachypneic | 120 | 120 | Factual
hypotensive | 120 | 120 | Factual
saturating well on room air | 120 | 120 | Factual
distended abdomen | 120 | 120 | Factual
tender on superficial palpation | 120 | 120 | Factual
inaudible bowel sounds | 120 | 120 | Factual
low Hb of 7.1 g/dL | 120 | 120 | Factual
hypoechoic nodular cystic area | 120 | 120 | Factual
splenomegaly | 120 | 120 | Factual
hyperdense intrasplenic hematoma | 120 | 120 | Factual
hypodense subcapsular hematoma | 120 | 120 | Factual
splenic laceration | 120 | 120 | Factual
intraperitoneal free fluid | 120 | 120 | Factual
grade 3 splenic injury | 120 | 120 | Factual
blood products mobilized | 120 | 120 | Factual
adequate resuscitation | 120 | 120 | Factual
explorative laparotomy | 120 | 120 | Factual
splenectomy | 120 | 120 | Factual
2.5 L of frank blood evacuated | 120 | 120 | Factual
enlarged spleen | 120 | 120 | Factual
long laceration on the upper pole | 120 | 120 | Factual
uneventful postoperative period | 120 | 168 | Factual
discharged home | 168 | 168 | Factual
fully recovered | 168 | 168 | Factual
scheduled clinic visits | 168 | 168 | Factual