57 years old | 0
male | 0
lepromatous leprosy | -1440
skin biopsy | -1440
rifampicin | -1440
clofazimine | -1440
dapsone | -1440
abdominal distension | -1440
constipation | -1440
vomiting | -1440
10-kg weight loss | -1440
admitted to the hospital | 0
vital stability | 0
peripheral lymphadenopathy | 0
distended abdomen | 0
positive shifting dullness | 0
computed tomography scan abdomen | 0
mural thickening of terminal ileum | 0
enlarged mesenteric lymph nodes | 0
mesenteric fat stranding | 0
intra-abdominal free fluid | 0
abdominal granulomatous infection | 0
neoplastic process | 0
abdominal paracentesis | 0
atypically large lymphocytes | 0
high-grade lymphoma | 0
flow cytometry | 0
abnormal CD4/CD8 double-negative T-cell population (38%) | 0
multiple phenotypic aberrancies | 0
cervical lymph node biopsy | 0
high-grade peripheral T-cell lymphoma (PTCL) | 0
NHL subtype | 0
bone marrow examination | 0
no involvement of T-cell NHL | 0
stage IV lymphoma | 0
dexamethasone | 0
tumor-lysis syndrome precautions | 0
clinical deterioration | 0
transfer to medical ICU | 0
severe sepsis | 0
antibiotics | 0
antifungals | 0
ICU care for 1 week | 168
transfer to national cancer center | 168
EPOCH chemotherapy protocol | 168
etoposide | 168
prednisone | 168
vincristine sulfate (oncovin) | 168
cyclophosphamide | 168
doxorubicin hydrochloride (hydroxydaunorubicin) | 168
six cycles | 168
CNS prophylaxis (intrathecal methotrexate) | 168
assessment after four cycles | 672
complete metabolic remission | 672
positron emission tomography/computed tomography | 672
multiple febrile neutropenia episodes | 672
recurrent bacteremia | 672
generalized weakness | 672
no sensory changes | 672
no clear fatigability | 672
decreased power in proximal and distal muscles (3/5) | 672
no other abnormalities | 672
previous history of ICU admission | 672
neurotoxic drug use | 672
malignancy | 672
differential diagnosis | 672
critical illness myopathy-neuropathy | 672
toxic neuropathy | 672
paraneoplastic syndrome | 672
neurophysiological electromyogram/nerve conduction study | 672
normal distal latencies | 672
normal compound muscle action potential | 672
normal conduction velocities | 672
normal F waves | 672
sensory nerve studies | 672
normal onset latencies | 672
normal sensory nerve action potential amplitude | 672
needle electromyogram | 672
proximal muscles | 672
distal muscles | 672
lower limbs | 672
upper limbs | 672
normal insertional activity | 672
no spontaneous activity | 672
normal motor unit action potential | 672
poor recruitment effects | 672
repetitive nerve stimulation (30–40 Hz) | 672
significant incremental response | 672
presynaptic neuromuscular junction disorder | 672
likely LEMS | 672
VGCC antibodies requested | 672
technical issues preventing VGCC antibodies test | 672
intravenous immunoglobulins for 5 days | 672
significant improvement of motor function | 672
ambulate afterward | 672
dramatic response to treatment | 672
planned autologous bone marrow transplant | 672
sepsis | 672
immunocompromised state | 672
re-admission to medical ICU | 672
severe sepsis | 672
multiorgan failure | 672
passed away | 4320
remission status maintained | 4320
