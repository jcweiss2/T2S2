63 years old | 0
male | 0
smoking | -6720
DVT | -12
rivaroxaban | -12
dyspnea | -8
pulmonary thromboembolism | -8
splenic infarctions | -8
renal infarctions | -8
cerebral and cerebellar areas | -8
nystagmus | -6
ataxia | -6
dysmetria | -6
adiadochokinesia | -6
lung cancer | -6
locally advanced non-small cell lung cancer | -6
large-cell carcinoma of the lung | -6
diplopia | -4
gait impairment | -4
substernal chest pain | -3
dyspnea | -3
sinus tachycardia | -3
ST segment elevation | -3
elevated serum troponin I | -3
reduced left ventricular ejection fraction | -3
mobile mass on the anterior leaflet of mitral valve | -3
moderate aortic insufficiency | -3
acute pulmonary edema | -2
respiratory failure | -2
coronary angiography | -2
reduced flow of the recurrent branch of the descending artery | -2
embolus | -2
aspirin | -2
β-blockers | -2
LMWH | -2
petechiae on the skin of the lower limbs | -2
abdominal pain | -1
loss of blood in the stool | -1
occlusion of a distal branch of the superior mesenteric artery | -1
thinning of the corresponding ileal loop | -1
bowel infarction | -1
emergency segmental ileo-cecal resection | -1
TEE | 0
mobile echogenic mass on the atrial surface of the anterior leaflet of the mitral valve | 0
moderate aortic insufficiency | 0
reduced LVEF | 0
coma | 2
multi-organ failure | 4
death | 70
admitted to the hospital | -8
discharged | -4
hospitalization | -4
NBTE | -3
PFO | -6
TTE | -6
cardio embolic origin of the brain lesions | -6
transesophageal echocardiogram | -4
Pembrolizumab therapy | -2
anticancer therapy | -2
anticoagulant therapy | -2
LMWH treatment | -2
fondaparinux | -2
edoxaban | -2
aspirin and β-blockers | -2
linezolid | -2
daptomycin | -2
piperacillin/tazobactam | -2
noninvasive ventilation | -2
coronary angiography | -2
emergency segmental ileo-cecal resection | -1
histological diagnosis of bowel infarction | -1
brain CT scan | 2
increased number and dimension of the bi-hemispheric infarct lesions | 2
novel ischemic events | 2
systemic embolisms | 2
cardiac vegetations | 2
aseptic thrombi | 2
valvular surface | 2
aortic and mitral valves | 2
embolization events | 2
spleen | 2
kidneys | 2
brain | 2
mesenteric | 2
coronary arterial circulation | 2
TTE | 2
TEE | 2
NBTE diagnosis | 2
anticoagulant therapy | 2
surgical intervention | 2
unfractionated heparin | 2
LMWH | 2
vitamin K antagonists | 2
fondaparinux | 2
direct oral anticoagulants | 2
rivaroxaban | 2
edoxaban | 2
bleeding events | 2
Pembrolizumab | 2
tyrosine kinase inhibitors | 2
immunotherapy agents | 2
pro-thrombotic effects | 2
cancer | 2
NBTE | 2
systemic embolisms | 2
sterile cardiac vegetations | 2
anticoagulant therapy | 2
anticancer therapy | 2
survival | 2
complications | 2