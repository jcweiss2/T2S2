3 years old | 0
female | 0
admitted to the hospital | 0
intermittent fever | -144
drowsiness | -24
nodding spasm | -8760
seizures | -336
electroencephalogram | -336
video-EEG | -336
myoclonic seizures | -336
epilepsy | -336
myoclonia | -336
sodium valproate | -336
discharged | -336
readmitted | 0
jaundice | 0
anuria | 0
hepatomegaly | 0
pharyngeal congestion | 0
low and dull cardiac sounds | 0
abdominal ultrasound | 0
hepatic failure | 0
acute kidney injury | 0
disseminated intravascular coagulation | 0
hemophagocytic syndrome | 0
pulmonary hemorrhage | 36
respiratory failure | 36
mechanical ventilation | 36
genomic DNA extraction | 0
molecular genetic analysis | 0
plasma exchange | 0
hemodialysis | 0
immunosupportive therapy | 0
component transfusion | 0
organ protection | 0
sodium valproate discontinued | 0
death | 168
NEXMIF variant | 0
whole exome sequencing | 720
mitochondrial DNA sequencing | 720
Sanger-sequencing analysis | 720
informed consent | 0
publication of case report | 0