74 years old | 0
man | 0
type 2 diabetes mellitus | -192
vague abdominal pain | -168
lower back pain | -168
leukocytosis | 0
white blood cell count of 25 × 10^9/L | 0
left shift | 0
dyspepsia | -672
upper gastrointestinal discomfort | -672
sore throat | -336
oral antibiotics | -336
magnetic resonance imaging | -168
computed tomography scan | 0
infrarenal aortic aneurysm rupture | 0
infectious etiology | 0
transferred to emergency department | 0
vancomycin | 3
piperacillin-tazobactam | 3
blood culturing | 3
hemodynamic stability | 0
autogenous NAIS reconstruction | 5
deep vein imaging | 5
two-team approach | 5
right femoral vein harvesting | 5
circumferential dissection | 5
infrarenal aortic clamp placement | 5
aorta debridement | 5
periaortic tissue debridement | 5
common iliac arteries debridement | 5
retroperitoneal tissues debridement | 5
femoral vein graft anastomosis | 5
omental flap | 5
thigh wound irrigation | 5
biphasic Doppler signals | 5
extubation | 72
intensive care unit stay | 168
lower extremity elevation | 168
compressive bandage wrapping | 168
thigh-high compression stockings | 168
group A streptococcus | 0
negative blood cultures | 72
transthoracic echocardiography | 72
intravenous ceftriaxone | 72
minimal stranding | 168
prolonged ileus | 408
discharged home | 408
thigh-high stockings | 408
aspirin | 408
intravenous antibiotics | 408
infectious disease follow-up | 720
oral amoxicillin | 720
vascular surgery follow-up | 720
afebrile | 720
well-healed incisions | 720
neurovascular examination | 720
stable imaging findings | 720
amoxicillin discontinuation | 720
ultrasound examination | 1752
CT angiography | 3504
annual follow-up | 3504
