58 years old | 0
female | 0
admitted to the emergency department | 0
lumbar back pain | -504
numbness in lower left leg and foot | -504
gait disorder | -120
urine incontinence | -120
bowel incontinence | -120
fever | -24
weight loss | -504
septic profile | 0
body temperature 38.8°C | 0
decreased strength in left leg | 0
strength MRC 3/5 in iliopsoas | 0
strength MRC 4/5 in tibialis anterior | 0
strength MRC 4+/5 in gastrocnemius | 0
normal sensation in saddle area | 0
normal sensation in perianal area | 0
normal anal sphincter tone | 0
positive Lasègue sign on left side | 0
leukocytosis | 0
elevated C-reactive protein level | 0
urine retention 1300 ml | 0
high-grade fever 40.9°C | 12
antibiotic therapy started | 12
Amoxicillin/Clavulanate | 12
transferred to intensive care unit | 12
MRI of spinal canal | 24
fistula from sigmoid colon to presacral abscess | 24
abscess expanded into spinal canal | 24
sacral osteomyelitis | 24
diffuse meningeal staining of conus medullaris and cauda equina | 24
chest/abdominal CT scan | 24
pleural fluid on both sides | 24
multiple fluid and air collections | 24
air in spinal canal and back muscles | 24
Hartmann's procedure | 48
multiple intra-abdominal abscesses drained | 48
intra-abdominal drains placed | 48
broad-spectrum antibiotics | 48
therapeutic heparin | 48
thrombus in left iliac vein | 48
extubated | 72
transferred to gastrointestinal surgery ward | 96
stoma production started | 96
neurological symptoms did not resolve | 96
discharged to primary care center | 336
enrolled in intensive rehabilitation program | 336