48 years old | 0
female | 0
diabetes | -720
coronary artery disease | -720
psoriasis | -720
acute onset of diffuse abdominal pain | -48
tachycardic | -48
heart rate of 130 | -48
hypotensive | -48
blood pressure of 78/45 | -48
afebrile | -48
alert and oriented to person, place and time | -48
resuscitated in the emergency department | -24
intravenous fluids | -24
normal WBC level of 8.3 thou/mcL | -24
acidotic | -24
pH of 7.29 | -24
lactic acid level of 3.5 mmol/l | -24
free air below the right hemidiaphragm | -24
distended abdomen | -24
tenderness | -24
guarding | -24
signs of peritonitis | -24
exploratory laparotomy | 0
repair of perforated viscus | 0
CT scan | 0
ruptured splenic abscess | 0
pneumoperitoneum | 0
increasingly confused | 12
worsening sepsis | 12
laparoscopic splenectomy | 12
converted to laparotomy with splenectomy | 12
gross contamination of the abdomen | 12
abdominal compartment copiously irrigated | 12
abdomen closed | 12
antibiotics | 12
intensive care unit | 12
post-operative care | 12
splenic abscess grew Prevotella intermedia | 24
blood cultures were negative | 24
transesophageal echocardiogram | 48
negative for any masses, thrombus or vegetation | 48
panorex | 48
negative | 48
tooth pain | -168
discharge | 240
splenectomy vaccinations | 336