38 years old | 0
male | 0
diagnosed with primary sclerosing cholangitis | -26304
no inflammatory bowel disease | -26304
ursodeoxycholic acid therapy | -26304
developed three episodes of bacterial cholangitis | -4320
last episode requiring intensive care unit admission | -4320
magnetic resonance cholangiography revealing mucosal irregularities | -4320
test of immunoglobulin type G4 serum level normal | -4320
carbohydrate antigen 19-9 level within normal limits | -4320
listed for liver transplantation | -4320
developed persistent pruritus | -2016
jaundice lasting for 3 months | -2016
fourth episode of bacterial cholangitis | -2016
Escherichia coli bacteremia in two prior episodes | -4320
Enterococcus fecalis in recent episode | -2016
fecal microbiota transplantation considered | -2016
donor screening completed | -2016
fecal microbiota transplantation performed weekly for 4 weeks | 0
antibiotics withheld during FMT | 0
ursodeoxycholic acid continued | 0
afebrile after third FMT | 168
anicteric after fourth FMT | 268
pruritus worsened for 6 weeks | 168
pruritus decreased to tolerable levels | 1008
liver function improvements observed | 0
circulating bile acids improved | 0
Proteobacteria decreased | 0
Bacteroidetes and Actinobacteria increased | 0
Enterobacter decreased | 0
Catenibacterium decreased | 0
Dialister decreased | 0
Clostridium emerged | 0
Veillonella emerged | 0
Fecalibacterium absent post-FMT | 0
Oscillopsira absent post-FMT |)
