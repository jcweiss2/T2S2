86 years old | 0
female | 0
anorexia | -72
vomiting | -72
incarcerated femoral hernia | -72
severe pain | -72
redness | -72
palpable bulge | -72
past appendectomy | -0
white blood cell count of 17.1 × 10^9/L | -72
C-reactive protein levels at 6.13 mg/dL | -72
abdominal computed tomography (CT) | -72
right incarcerated femoral hernia | -72
small bowel obstruction | -72
laparoscopic repair of an incarcerated femoral hernia | 0
incarcerated ileum perforation | 0
necrotic ileum resection | 0
right femoral hernia repair | 0
McVay procedure | 0
postoperative intensive care | 0
septic shock | 0
disseminated intravascular coagulation | 0
discharged | 720
umbilical incisional hernia | 2160
laparoscopic incisional hernia repair | 2160
multiple small white nodules | 2160
peritoneal wash cytology | 2160
frozen sections | 2160
multinucleated giant cell | 2160
foreign body | 2160
inflammatory cells | 2160
fibrosis | 2160
granulomatous formations | 2160
laparoscopic intraperitoneal onlay mesh repair | 2160
hernia orifice closure | 2160
postoperative clinical course | 2160
chest-to-abdominal enhanced CT | 3024
gastrointestinal and colon endoscopy | 3024
no malignancy | 3024
no recurrence of hernia | 3024
follow-up | 5040