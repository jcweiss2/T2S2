44 years old | 0 | 0 
female | 0 | 0 
admitted to the emergency department | 0 | 0 
left groin and inner thigh redness | -72 | 0 
left groin and inner thigh pain | -72 | 0 
left groin and inner thigh swelling | -72 | 0 
fever | -72 | 0 
chills | -72 | 0 
vomiting | -72 | 0 
treated with intravenous vancomycin | -24 | -24 
discharged from urgent care | -24 | -24 
afebrile | 0 | 0 
normotensive | 0 | 0 
tachycardia | 0 | 0 
mild tachypnea | 0 | 0 
left inner thigh and groin induration | 0 | 0 
morbidly obese | 0 | 0 
lactate 3.5 mmol/L | 0 | 0 
WBC 18.2 × 103 per mm3 | 0 | 0 
hemoglobin 12.3 g/dL | 0 | 0 
sodium 136 mmol/dL | 0 | 0 
glucose 225 mg/dL | 0 | 0 
creatinine 1.8 mg/dL | 0 | 0 
laboratory risk indicator for necrotizing fasciitis (LRINEC) score of 6 | 0 | 0 
bedside ultrasound performed | 0 | 0 
subcutaneous thickening | 0 | 0 
air | 0 | 0 
fascial fluid | 0 | 0 
started on intravenous vancomycin and piperacillin/tazobactam | 0 | 0 
surgery consulted | 0 | 0 
operative debridement of the left groin and perineum | 0 | 0 
excision of 15 cm × 23 cm of tissue | 0 | 0 
extensive washout | 0 | 0 
admitted to the surgical intensive care unit | 0 | 0 
septic shock | 0 | 0 
requiring vasopressors | 0 | 0 
requiring ventilator | 0 | 0 
repeat washouts with minor debridements | 0 | 72 
lactate normalization | 72 | 72 
down-trending WBC to 13.5 × 103 per mm3 | 72 | 72 
extubated | 120 | 120 
transferred to a step-down unit | 120 | 120 
plastic surgery consulted | 120 | 120 
wound vacuum-assisted closure (V.A.C.) device placed | 216 | 216 
transferred to the plastic surgery service | 216 | 216 
discharged home with a wound V.A.C. | 672 | 672 
skin graft | 672 | 672 
recovering well | 672 | 672