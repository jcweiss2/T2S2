20 years old | 0
female | 0
G1P1001 | 0
admitted to the hospital | 0
cough | -72
shortness of breath | -72
amenorrhea | -720
morning sickness | -120
evaluation for pulmonary embolism | 0
infectious etiologies | 0
Influenza A negative | 0
Influenza B negative | 0
SARS-CoV-2 negative | 0
beta-HCG 900,000 mIU/mL | 0
adnexal mass | 0
bilateral diffuse pulmonary nodules | 0
intubated | 0
hypoxemia | 0
empiric antibiotics | 0
septic shock | 0
transferred to hospital | 0
ECMO cannulation | 0
right ventricular failure | 0
tricuspid regurgitation | 0
dilated right ventricle | 0
systolic dysfunction | 0
intra-atrial septal bowing | 0
dual-lumen percutaneous right ventricular assist device | 0
ECMO circuit | 0
dilation and curettage | 0
heparin infusion | 0
vasopressors | 0
beta-HCG 917,929 mIU/mL | 0
induction chemotherapy | 12
cisplatin | 12
etoposide | 12
WHO score 14 | 0
extubated | 48
ECMO circuit complication | 48
oxygenator failure | 48
tachycardia | 48
hypoxia | 48
hypotension | 48
vasopressor support | 48
circuit exchange | 48
reintubation avoided | 48
final pathology | 0
no chorionic villi | 0
no fetal parts | 0
no implantation site | 0
no neoplasm | 0
gestational type endometrium | 0
breakdown | 0
CT-guided biopsy | 144
pelvic mass | 144
corpus luteum cyst | 144
oncologic plan | 0
EMA-CO chemotherapy | 0
thrombocytopenia | 120
neutropenia | 120
delayed chemotherapy | 120
magnetic resonance imaging | 120
brain negative for metastatic lesions | 120
respiratory status improved | 120
decannulated from ECMO | 240
clot on cannula | 240
tricuspid valve echodensity | 240
tumor | 240
thrombus | 240
vegetation | 240
beta-HCG 60,862 mIU/mL | 240
transferred out of ICU | 288
platelet counts improved | 288
ANC improved | 288
cycle 2 induction chemotherapy | 384
cycle 2 induction chemotherapy | 384
echocardiogram | 384
tricuspid valve echodensity | 384
enoxaparin | 384
respiratory status stable | 384
discharged home | 432
cycle 1 day 1 EMA-CO | 720
etoposide | 720
methotrexate | 720
dactinomycin | 720
cyclophosphamide | 744
vincristine | 744
filgrastim | 744
beta-HCG normalized | 1008
EMA-CO cycles | 1008
surveillance | 1008