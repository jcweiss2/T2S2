40 years old | 0
male | 0
admitted to the emergency department | 0
odynophagia | -168
dry cough | -168
exertional dyspnea | -168
fever | -168
arthralgias | -168
fatigue | -168
poorly controlled diabetes | 0
glycosylated hemoglobin 10.8 % | 0
insulin treatment with 44 IU of glargine | 0
insulin treatment with 16 UI of lispro | 0
body mass index of 28.3 kg/m² | 0
heart rate 110 beats per minute | 0
24 breaths per minute | 0
oxygen saturation of 82% at ambiance | 0
right lung rales | 0
no cyanosis | 0
no lower limb edema | 0
no direct contact with a coronavirus case | 0
arterial gases showed moderate oxygen impairment (PAFI 190) | 0
supplemental oxygen required | 0
normal blood count | 0
increased CRP | 0
right basal ground glass opacity on chest x-ray | 0
positive RT-PCR COVID-19 | 0
adenovirus isolated in respiratory viral panel | 0
increased lactate dehydrogenase | 0
markedly elevated ferritin | 0
positive D-dimer adjusted by age | 0
ground-glass opacities with multilobar involvement on chest tomography | 0
increased dyspnea | 144
tachypnea | 144
desaturation | 144
transferred to intensive care unit | 144
management with ampicillin-sulbactam | 144
management with clarithromycin | 144
hydroxychloroquine 200 mg twice daily | 144
corrected Qt interval monitored | 144
hypotension | 144
hypoxemia | 144
mechanical ventilation started | 144
norepinephrine started | 144
septic shock | 144
acute respiratory distress syndrome (ARDS) | 144
pronation required | 144
neuromuscular relaxation cycles required | 144
Klebsiella oxytoca isolated on blood cultures | 144
antibiotic escalation to cefepime | 144
10-day treatment completed | 144
successful extubation | 432
transferred to general floor | 432
symptoms resolved | 432
second RT-PCR SARS Cov2 negative | 432
discharged | 480
supplemental oxygen requirement at home | 480
no gastrointestinal symptoms | 0
no history of smoking | 0
no history of alcohol consumption | 0
