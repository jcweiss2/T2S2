55 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
nonalcoholic steatohepatitis | -672 | 0 | Factual
alpha 1 antitrypsin deficiency | -672 | 0 | Factual
orthotopic liver transplant | 0 | 0 | Factual
incarcerated inguinal hernia | -168 | -168 | Factual
hernia repair | -168 | -168 | Factual
cytomegalovirus viremia | -168 | -168 | Factual
valganciclovir | -168 | 0 | Factual
mycophenolate mofetil | 0 | 0 | Factual
tacrolimus | 0 | 0 | Factual
prednisone | 0 | 0 | Factual
encephalopathy | -48 | 0 | Factual
increasing home oxygen requirements | -48 | 0 | Factual
oxygen saturation <92% | -48 | 0 | Factual
sparse speech | 0 | 0 | Factual
disorientation | 0 | 0 | Factual
nonfocal neurologic examination | 0 | 0 | Factual
white blood cell count 9.3 × 10^9/L | 0 | 0 | Factual
creatinine 2.12 mg/dL | 0 | 0 | Factual
blood urea nitrogen 53 mg/dL | 0 | 0 | Factual
synthetic liver function normal | 0 | 0 | Factual
arterial ammonia 204 µmol/L | 0 | 0 | Factual
induction dosing of intravenous ganciclovir | 0 | 0 | Factual
empiric antibiotic coverage | 0 | 0 | Factual
vancomycin | 0 | 0 | Factual
meropenem | 0 | 0 | Factual
micafungin | 0 | 0 | Factual
intravenous micronutrient supplementation | 0 | 0 | Factual
B1 supplementation | 0 | 0 | Factual
B6 supplementation | 0 | 0 | Factual
levocarnitine supplementation | 0 | 0 | Factual
lumbar puncture | 0 | 0 | Factual
encapsulated yeast suspicious for Cryptococcus | 0 | 0 | Factual
liposomal amphotericin B | 0 | 0 | Factual
flucytosine | 0 | 0 | Factual
continuous renal replacement therapy (CRRT) | 0 | 0 | Factual
rifaximin | 0 | 0 | Factual
zinc | 0 | 0 | Factual
lactulose | 0 | 0 | Factual
ammonia level 692 µmol/L | 12 | 24 | Factual
neurological deterioration | 12 | 24 | Factual
mechanical ventilation | 24 | 24 | Factual
empiric intravenous doxycycline | 24 | 24 | Factual
urine and bronchial aspirate for Mycoplasma and Ureaplasma PCR | 24 | 24 | Factual
ammonia level <100 µmol/L | 48 | 48 | Factual
Cryptococcal serum and cerebrospinal fluid (CSF) antigen titers positive | 48 | 48 | Factual
cultures from bronchoalveolar lavage, CSF, and blood revealed cryptococcal growth | 48 | 48 | Factual
repeat lumbar punctures | 48 | 0 | Factual
opening pressures greater than 45 cmH2O | 48 | 0 | Factual
large volume drainage | 48 | 0 | Factual
thrombocytopenia | 48 | 0 | Factual
tracheostomy | 0 | 0 | Factual
hydrocephalus | 0 | 0 | Factual
oliguric renal failure | 0 | 0 | Factual
splenic infarcts with necrosis | 0 | 0 | Factual
splenectomy | 0 | 0 | Factual
sepsis | 0 | 0 | Factual
duodenal leak | 0 | 0 | Factual
failure to thrive | 0 | 0 | Factual
comfort care in hospice | 0 | 0 | Factual
urea cycle disorder screening studies | 0 | 0 | Factual
low urine orotic level | 0 | 0 | Factual
normal serum citrulline and arginine level | 0 | 0 | Factual