50 years old | 0
male | 0
hospitalized | 0
dry cough | -96
chills | -96
fever | -96
back pain | -96
cough | -96
no gastrointestinal symptoms | -96
acetaminophen | -96
carbocysteine | -96
symptoms did not improve | -96
referred to our hospital | -96
previous 20-pack-year smoker | 0
no alcohol consumption | 0
lived in an over 40-year-old house | 0
contaminated shower use presumed | 0
worked in a bar | 0
rainy season | 0
no use of humidifier | 0
no use of air conditioner | 0
no recent travel to spa | 0
no recent travel to other countries | 0
maintenance hemodialysis for three years | 0
diabetic kidney disease | 0
percutaneous coronary intervention eight years earlier | 0
angina pectoris eight years earlier | 0
congestive heart failure | 0
beta blockers | 0
angiotensin receptor blockers | 0
echocardiography four months earlier | -2880
ejection fraction 33% four months earlier | -2880
diffuse hypokinesis four months earlier | -2880
echocardiography on admission | 0
ejection fraction 30% | 0
no significant change from previous examination | 0
no history of gastrointestinal disorders | 0
no family history of diabetes | 0
no family history of hemodialysis | 0
no family history of immunodeficiency | 0
body temperature 38.9°C | 0
blood pressure 131/97 mmHg | 0
heart rate 117 per minute | 0
respiratory rate 18 per minute | 0
arterial oxygen saturation 96% | 0
intact consciousness | 0
left pulmonary rales | 0
bilateral lower leg edema | 0
no xerostomia | 0
elevated leukocyte count | 0
markedly elevated C-reactive protein | 0
severe liver function abnormalities | 0
elevated creatine kinase | 0
moderate hypoxemia | 0
electrocardiogram tachycardia | 0
no specific ST elevation | 0
chest radiograph lobular infiltrates left lower lung | 0
mild heart enlargement | 0
no significant pleural effusion | 0
CT lobar consolidation left lower lobe | 0
chronic liver injury | 0
fatty liver | 0
bacterial pneumonia diagnosis | 0
severe liver dysfunction diagnosis | 0
good general condition | 0
no dyspnea necessitating oxygen | 0
A-DROP score <1 | 0
quick Sequential Organ Failure Assessment score 0 | 0
piperacillin/tazobactam started | 0
immunodeficient expected | 0
laboratory results worsened next day | 24
negative blood cultures | 24
sputum culture oral microflora | 24
sputum serous components | 24
consideration of Legionnaires' disease | 24
oral azithromycin started day 1 | 24
consciousness deterioration | 34
systolic blood pressure deterioration | 34
septic shock diagnosis | 34
noradrenaline infusion started | 34
bradycardia day 2 | 48
cardiac arrest day 2 | 48
cardiopulmonary resuscitation | 48
defibrillation attempts | 48
adrenaline bolus doses | 48
return of spontaneous circulation | 48
transfer to ICU | 48
hydrocortisone phosphate started | 48
gamma globulin started | 48
CRRT started day 3 | 72
noradrenaline dose reduced | 72
blood pressure improved | 72
azithromycin changed to levofloxacin day 3 | 72
blood pressure drop day 5 | 120
CRRT discontinued | 120
death | 120
Legionella pneumophila serotype 1 detected postmortem | 120
autopsy lobar pneumonia | 120
hepatic lobular central congestion | 120
shock liver | 120
Legionnaires' disease confirmed | 120
