newborn female | 0 | 0 | Factual
24 weeks + 3 days | 0 | 0 | Factual
breech presentation | 0 | 0 | Factual
cord prolapse | 0 | 0 | Factual
birth weight of 645 g | 0 | 0 | Factual
HIV negative mother | 0 | 0 | Factual
Apgar score of 4 | 0 | 0 | Factual
Apgar score of 8 | 5 | 5 | Factual
mechanical ventilation | 0 | 216 | Factual
central umbilical catheters | 0 | 216 | Factual
total parenteral nutrition | 0 | 216 | Factual
empiric antibiotics | 0 | 216 | Factual
skin sensors | 0 | 216 | Factual
late-onset sepsis | -216 | -216 | Factual
Escherichia coli bacteremia | -216 | -216 | Factual
cefepime | -216 | -96 | Factual
adhesive patch removal | -192 | -192 | Factual
skin abrasion | -192 | -192 | Factual
erythema | -168 | -168 | Factual
induration | -168 | -168 | Factual
plaque with necrotic center | -168 | -168 | Factual
ulcer | -144 | -144 | Factual
subcutaneous cell tissue extension | -144 | -144 | Factual
necrotic area progression | -144 | -144 | Factual
intensive treatment | -144 | -72 | Factual
wound care team | -144 | -72 | Factual
healings | -144 | -72 | Factual
hydrating dermal wound dressings | -144 | -72 | Factual
sodium alginate | -144 | -72 | Factual
carboxymethylcellulose | -144 | -72 | Factual
hydrocolloids | -144 | -72 | Factual
thermic instability | -72 | -72 | Factual
metabolic acidosis | -72 | -72 | Factual
hyperglycemia | -72 | -72 | Factual
hypotension | -72 | -72 | Factual
clinical deterioration | -72 | -72 | Factual
cutaneous mucormicosis suspicion | -72 | -72 | Possible
skin biopsy | -72 | -72 | Factual
empiric antifungal treatment | -72 | -36 | Factual
liposomal amphotericin B | -72 | -36 | Factual
fungal biomarkers | -72 | -72 | Negated
serum galactomannan | -72 | -72 | Negated
1,3 beta-D-glucan | -72 | -72 | Negated
refractory shock | -36 | -36 | Factual
renal failure | -36 | -36 | Factual
death | 0 | 0 | Factual
Rhizopus spp. | -72 | -72 | Factual
Rhizopus arrhizus | -72 | -72 | Factual
broad aseptate hyphae | -72 | -72 | Factual
right angle branching | -72 | -72 | Factual
MALDI-TOF MS | -72 | -72 | Factual
PCR | -72 | -72 | Factual
panfungal PCR | -72 | -72 | Factual
sequencing | -72 | -72 | Factual
fungal blood cultures | -216 | -216 | Negated
necrotic eschar | -144 | -144 | Factual
skin abscesses | -144 | -144 | Possible
surgical debridement | -36 | -36 | Negated
anti-fungal treatment | -72 | -36 | Factual
L-AmB | -72 | -36 | Factual