55 years old | 0\
male | 0\
nonalcoholic steatohepatitis | -672\
alpha 1 antitrypsin deficiency | -672\
orthotopic liver transplant | 0\
incarcerated inguinal hernia | 24\
repaired incarcerated inguinal hernia | 48\
cytomegalovirus (CMV) viremia | 168\
treated with valganciclovir | 168\
discharged | 336\
immunosuppression of mycophenolate mofetil | 336\
immunosuppression of tacrolimus | 336\
immunosuppression of prednisone | 336\
encephalopathy | 336\
increasing home oxygen requirements | 336\
required 4L nasal cannula | 336\
oxygen saturation >92% | 336\
sparse speech | 336\
disorientation | 336\
nonfocal neurologic examination | 336\
white blood cell count was 9.3 × 109/L | 336\
creatinine 2.12 mg/dL | 336\
blood urea nitrogen of 53 mg/dL | 336\
arterial ammonia was unusually elevated at 204 µmol/L | 336\
induction dosing of intravenous ganciclovir | 336\
empiric antibiotic coverage with vancomycin | 336\
empiric antibiotic coverage with meropenem | 336\
empiric antibiotic coverage with micafungin | 336\
intravenous micronutrient supplementation for B1 | 336\
intravenous micronutrient supplementation for B6 | 336\
intravenous micronutrient supplementation for levocarnitine | 336\
lumbar puncture | 336\
opening pressure of 8 cmH2O | 336\
Gram stain revealed encapsulated yeast suspicious for Cryptococcus | 336\
liposomal amphotericin B | 336\
flucytosine | 336\
continuous renal replacement therapy (CRRT) | 336\
rifaximin | 336\
zinc | 336\
lactulose | 336\
ammonia proceeded to unexpectedly climb to 692 µmol/L | 360\
neurological deterioration | 360\
mechanical ventilation | 360\
empiric intravenous doxycycline | 360\
urine and bronchial aspirate was obtained for Mycoplasma and Ureaplasma polymerase chain reaction (PCR) | 360\
ammonia levels had fallen to <100 µmol/L | 384\
Cryptococcal serum and cerebrospinal fluid (CSF) antigen titers both returned positive at >1:2560 | 384\
cultures from bronchoalveolar lavage, CSF, and blood all revealed cryptococcal growth | 384\
repeat lumbar punctures revealed opening pressures greater than 45 cmH2O | 432\
large volume drainage every 48 hours | 432\
thrombocytopenia | 432\
nadir of 16 × 103/µL | 432\
mental status transiently improved | 432\
unable to wean from mechanical ventilation | 432\
tracheostomy | 432\
persistent hydrocephalus | 432\
oliguric renal failure | 432\
progressive splenic infarcts with necrosis | 432\
splenectomy | 432\
sepsis | 432\
duodenal leak | 432\
persisting renal failure | 432\
failure to thrive | 432\
moved to comfort care in hospice | 432\
urea cycle disorder screening studies eventually returned | 432\
low urine orotic level | 432\
normal serum citrulline and arginine level | 432