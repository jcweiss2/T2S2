18 years old | 0
male | 0
admitted to the hospital | 0
abdominal discomfort | -24
nausea | -24
vomiting | -24
fever | -24
vaginal discharge | -24
obstetric ultrasound | -24
abdominal pain | -6
nausea | -6
vomiting | -6
tachycardia | -6
diffuse abdominal pain | -6
guarding on the right quadrants | -6
neutrophilia | 0
low prothrombinemia | 0
acute renal failure | 0
high procalcitonin | 0
c-reactive protein | 0
moderate fluid in all quadrants | 0
good foetal vitality | 0
hypotension | 0
general abdominal guarding | 0
hyperlacticaemia | 0
hypokalaemia | 0
hyperglycaemia | 0
septic shock | 0
abdominal source | 0
exploratory laparotomy | 0
generalised purulent peritonitis | 0
perforated acute appendicitis | 0
pus | 0
multiple interloop abscesses | 0
retrosplenic abscess | 0
subfrenic abscess | 0
pelvic abscess | 0
retrouterine abscess | 0
appendicectomy | 0
thorough abdominal washing | 0
laparostomy | 0
vasopressor therapy | 0
dialysis | 0
intravenous piperacillin-tazobactam | 0
laparostomy revision | 24
bowel oedema | 24
distention | 24
mild intraabdominal soiling | 24
further peritoneal lavage | 24
new laparostomy | 24
progressive closure technique | 24
surgical revision | 96
abdominal cavity primary closed | 96
amoxicillin with clavulanic acid | 96
obstetric follow-up | 96
elective caesarean section | 168
healthy child | 168
ventral hernia | 168
3 months post-partum follow-up | 168