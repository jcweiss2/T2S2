42 years old | 0 | 0 
female | 0 | 0 
granular dystrophy | 0 | 0 
DALK | 0 | 0 
big bubble technique | 0 | 0 
8 mm recipient stromal flap partially dissected | 0 | 0 
air injected into the substance of the remaining stroma | 0 | 0 
donor button cut 8.25 mm | 0 | 0 
DM peeled off | 0 | 0 
donor button placed over the recipient DM | 0 | 0 
donor button sutured with recipient rim | 0 | 0 
age of donor cornea 36 years | 0 | 0 
in situ cornea excision | 0 | 0 
surgery gone well | 0 | 0 
whitish infiltrates along the graft-host junction | -24 | 24 
severe anterior chamber reaction | -24 | 24 
postoperative keratitis | -24 | 24 
graft removed | 24 | 24 
graft replaced by another stromal graft | 24 | 24 
corneal scrapings sent for microbiology | 24 | 24 
host DM clear and intact | 24 | 24 
topical vancomycin started | 27 | 48 
topical ceftazidime started | 27 | 48 
Gram-stain showed Gram-negative Bacilli | 48 | 48 
infiltrates along the entire graft host junction | 48 | 72 
hypopyon | 48 | 72 
topical antibiotics increased to half hourly | 72 | 72 
corneal scrapings revealed Klebsiella pneumoniae | 72 | 72 
Klebsiella pneumoniae resistant to multiple antibiotics | 72 | 72 
imipenem drops started | 96 | 120 
infiltration extended toward center of graft | 120 | 120 
hypopyon persisted | 120 | 120 
therapeutic penetrating keratoplasty | 168 | 168 
infiltrates observed in host DM | 168 | 168 
graft clear without infiltrates or hypopyon | 192 | 192 
imipenem continued | 192 | 192 
gatifloxacin drops added | 192 | 240 
prednisolone drops added | 240 | 240 
unaided vision 6/60 | 1008 | 1008 
vision improved to 6/18 with pin hole | 1008 | 1008 
graft clear | 1008 | 1008 
anterior segment quiet | 1008 | 1008 
intraocular pressure normal | 1008 | 1008 
pathogen eradicated | 1008 | 1008