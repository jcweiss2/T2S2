34 years old | 0
female | 0
gravida 4 | 0
para 3 | 0
presented to the Obstetric Department | 0
labor induction | 0
suspected macrosomic fetus | 0
39th gestational week | 0
medical history unremarkable | 0
periodic depression | -672
whiplash | -672
overweight | -672
BMI 34 | -672
entered the active phase of labor | 6
amniotomy | -6
oxytocin | 6
spontaneous birth | 10
male infant | 10
Apgar score 7 | 10
Apgar score 10 | 15
discharged | 4
readmitted to the hospital | 24
complaining of pain | 24
complaining of chills | 24
hypotension | 24
tachycardia | 24
fever | 24
oliguria | 24
generalized abdominal tenderness | 24
peritoneal signs | 24
enlarged uterus | 24
abdominal ultrasound examination | 24
transvaginal ultrasound examination | 24
empty uterus | 24
no intraabdominal fluid | 24
culture samples collected | 24
intravenous antibiotic therapy | 24
metronidazole | 24
cefuroxime | 24
elevated CRP | 24
elevated creatinine | 24
normal white blood cell counts | 24
normal hemoglobin | 24
normal platelets | 24
abdominal CT-scan | 32
enlarged uterus | 32
ascites | 32
transferred to the ICU | 32
circulatory instability | 32
tentative diagnosis severe puerperal endometritis | 32
manual exploration of the uterus | 38
progressive elevation of CRP | 38
leucocytosis | 38
antibiotic therapy changed | 38
meropenem | 38
fulminate circulatory shock | 40
fluid resuscitation | 40
vasopressor therapy | 40
cardiac arrest | 40
basic cardiopulmonary resuscitation | 40
intravenous adrenaline | 40
transthoracic echocardiography | 40
right ventricular heart failure | 40
left ventricular heart failure | 40
low ejection fraction | 40
transferred to the TICU | 40
invasive cardiopulmonary support | 40
cardiac failure reversed | 64
kidney function improved | 64
urine sample | 24
culture from vagina | 24
Group A streptococcus | 24
blood cultures negative | 24
allergy toward penicillin | 24
meropenem and metronidazole continued | 24
returned to the regional ICU | 168
stable condition | 168
intubated | 168
sedated | 168
circulatory unstable | 168
temperature increased | 168
active cooling | 168
CVVHDF | 168
new CT scan | 168
suspicion of necrosis in the uterus | 168
thrombosis in the right uterine artery | 168
explorative laparotomy | 168
total abdominal hysterectomy | 168
necrotic uterus | 168
enlarged uterus | 168
thromboembolus in the right uterine artery | 168
extensive acute necrotizing inflammation | 168
septic thromboemboli | 168
intensive care management | 168
respiratory assistance | 168
dialysis | 168
altered consciousness | 168
paralysis of all four extremities | 168
absent tendon reflexes | 168
preserved eye movements | 168
preserved oculus reflex | 168
MRI-scan | 168
EEG | 168
lumbar puncture | 168
Critical Illness Polyneuropathy | 168
transferred to a highly specialized department | 168
neurorehabilitation | 168
condition slowly improving | 336