63 years old| 0  
    man | 0  
    presented to the emergency department| 0  
    midepigastric pain | -72  
    intolerance to oral intake | -72  
    denied hematemesis | 0  
    denied hematochezia | 0  
    denied other gastrointestinal symptoms | 0  
    physical examination | 0  
    mild midepigastric tenderness | 0  
    computed tomography scan | 0  
    fluid collection | 0  
    thickened duodenum wall | 0  
    infrarenal saccular abdominal aortic aneurysm | 0  
    no evidence of free air | 0  
    esophagogastroduodenoscopy | 0  
    abnormal mucosa | 0  
    possible mass | 0  
    perforation of the third portion of the duodenum | 0  
    taken to the operating room | 0  
    gross contamination from intestinal fluid | 0  
    perforation of the posterior medial aspect of the second portion of the duodenum | 0  
    retroperitoneal space adjacent to the infrarenal aorta | 0  
    saccular mycotic aortic aneurysm | 0  
    aortic wall inflammation | 0  
    thinning representing impending rupture | 0  
    intraoperative hemodynamic stability | 0  
    pancreaticoduodenectomy | 0  
    open abdominal aortic aneurysm repair | 0  
    rifampin-soaked Dacron graft | 0  
    omental wrap | 0  
    staged Whipple reconstruction | 48  
    final pathologic examination | 0  
    moderately differentiated pancreatic ductal adenocarcinoma | 0  
    extension through the duodenum wall | 0  
    lymph node positive | 0  
    margins uninvolved | 0  
    Cooper triad for aortoenteric fistula | 0  
    upper gastrointestinal bleeding | 0  
    abdominal pain | 0  
    palpable abdominal mass | 0  
    primary aortoenteric fistula due to pancreatic cancer | 0  
    prolonged postoperative course | 0  
    intractable intra-abdominal sepsis | 0  
    died | 2880  
    
    <|eot_id|>
    
    63 years old|0
    man|0
    presented to the emergency department|0
    midepigastric pain|-72
    intolerance to oral intake|-72
    denied hematemesis|0
    denied hematochezia|0
    denied other gastrointestinal symptoms|0
    physical examination|0
    mild midepigastric tenderness|0
    computed tomography scan|0
    fluid collection|0
    thickened duodenum wall|0
    infrarenal saccular abdominal aortic aneurysm|0
    no evidence of free air|0
    esophagogastroduodenoscopy|0
    abnormal mucosa|0
    possible mass|0
    perforation of the third portion of the duodenum|0
    taken to the operating room|0
    gross contamination from intestinal fluid|0
    perforation of the posterior medial aspect of the second portion of the duodenum|0
    retroperitoneal space adjacent to the infrarenal aorta|0
    saccular mycotic aortic aneurysm|0
    aortic wall inflammation|0
    thinning representing impending rupture|0
    intraoperative hemodynamic stability|0
    pancreaticoduodenectomy|0
    open abdominal aortic aneurysm repair|0
    rifampin-soaked Dacron graft|0
    omental wrap|0
    staged Whipple reconstruction|48
    final pathologic examination|0
    moderately differentiated pancreatic ductal adenocarcinoma|0
    extension through the duodenum wall|0
    lymph node positive|0
    margins uninvolved|0
    Cooper triad for aortoenteric fistula|0
    upper gastrointestinal bleeding|0
    abdominal pain|0
    palpable abdominal mass|0
    primary aortoenteric fistula due to pancreatic cancer|0
    prolonged postoperative course|0
    intractable intra-abdominal sepsis|0
    died|2880