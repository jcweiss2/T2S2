67 years old | 0
female | 0
plasma cell leukemia | -8760
multiple myeloma | -8760
treatment for malignancy | -8760
generalized tiredness | -24
altered sensorium | -24
patent airway | 0
bilateral crackles at the lung base | 0
respiratory rate 30 cycles/min | 0
Spo2 70% in room air | 0
feeble peripheral pulses | 0
un-recordable blood pressure | 0
heart rate 120 bpm | 0
responding to verbal stimulus | 0
normal finger stick glucose levels | 0
pale | 0
jugular venous distension | 0
bilateral pitting pedal edema | 0
muffled heart sounds | 0
no focal deficits | 0
bilaterally equal pupils | 0
secure large bore intravenous lines | 0
IV fluid resuscitation | 0
vasopressor support | 1
inotrope support | 1
intubation | 2
continuous cardiac monitoring | 2
supplemental oxygen | 2
bedside goal-directed ECHO | 2
massive pericardial effusion | 2
right ventricular collapse | 2
plethoric IVC | 2
emergency pericardiocentesis | 3
pericardial fluid aspirated | 3
active aspiration | 3
250 ml of fluid aspirated | 3
heart globally expanded | 4
pericardial drain placement | 6
transfer to intensive care team | 6
cardiac tamponade | 0 
BECK’s triad | 0 
RUSH protocol | 2 
ultrasound guidance | 3 
central venous catheter | 3 
PHASED ARRAY probe | 3 
local anesthetic | 3 
trocar needle | 3 
pericardial sac punctured | 3 
3-way stopcock valve | 3 
syringe | 3 
pericardiocentesis | 3 
discharge from ED | -24 
admitted to ED | 0 
discharge from hospital | 48 
admitted to hospital | 0 
pericardial effusion | -24 
multiple myeloma diagnosis | -8760 
pericardial effusion diagnosis | 2 
cardiac tamponade diagnosis | 2 
ultrasound | 2 
pericardiocentesis procedure | 3 
pericardial fluid analysis | 4 
pericardial drain | 6 
intensive care | 6 
ventilator support | 2 
oxygen therapy | 2 
vasopressor | 1 
inotrope | 1 
IV fluid | 0 
pericardiocentesis guidance | 3 
ultrasound guidance | 3 
sub-xiphoid view | 3 
pericardial sac | 3 
pericardial fluid | 3 
right ventricle | 2 
inferior vena cava | 2 
heart rate monitoring | 2 
blood pressure monitoring | 2 
oxygen saturation monitoring | 2 
respiratory rate monitoring | 0 
pericardial effusion treatment | 3 
cardiac tamponade treatment | 3 
multiple myeloma treatment | -8760 
plasma cell leukemia treatment | -8760 
pericardiocentesis complication | 6 
pericardial drain complication | 6 
intensive care complication | 6 
ventilator complication | 6 
oxygen therapy complication | 6 
vasopressor complication | 6 
inotrope complication | 6 
IV fluid complication | 6 
pericardiocentesis outcome | 6 
pericardial effusion outcome | 6 
cardiac tamponade outcome | 6 
multiple myeloma outcome | 48 
plasma cell leukemia outcome | 48 
patient outcome | 48 
discharge | 48 
death | -1 
survival | 48 
recovery | 48 
relapse | -1 
remission | 48 
pericardial effusion recurrence | -1 
cardiac tamponade recurrence | -1 
multiple myeloma recurrence | -1 
plasma cell leukemia recurrence | -1 
pericardiocentesis recurrence | -1 
pericardial drain recurrence | -1 
intensive care recurrence | -1 
ventilator recurrence | -1 
oxygen therapy recurrence | -1 
vasopressor recurrence | -1 
inotrope recurrence | -1 
IV fluid recurrence | -1 
pericardiocentesis readmission | -1 
pericardial effusion readmission | -1 
cardiac tamponade readmission | -1 
multiple myeloma readmission | -1 
plasma cell leukemia readmission | -1 
intensive care readmission | -1 
ventilator readmission | -1 
oxygen therapy readmission | -1 
vasopressor readmission | -1 
inotrope readmission | -1 
IV fluid readmission | -1 
pericardiocentesis follow-up | 48 
pericardial effusion follow-up | 48 
cardiac tamponade follow-up | 48 
multiple myeloma follow-up | 48 
plasma cell leukemia follow-up | 48 
intensive care follow-up | 48 
ventilator follow-up | 48 
oxygen therapy follow-up | 48 
vasopressor follow-up | 48 
inotrope follow-up | 48 
IV fluid follow-up | 48 
pericardiocentesis aftercare | 48 
pericardial effusion aftercare | 48 
cardiac tamponade aftercare | 48 
multiple myeloma aftercare | 48 
plasma cell leukemia aftercare | 48 
intensive care aftercare | 48 
ventilator aftercare | 48 
oxygen therapy aftercare | 48 
vasopressor aftercare | 48 
inotrope aftercare | 48 
IV fluid aftercare | 48 
pericardiocentesis rehabilitation | 48 
pericardial effusion rehabilitation | 48 
cardiac tamponade rehabilitation | 48 
multiple myeloma rehabilitation | 48 
plasma cell leukemia rehabilitation | 48 
intensive care rehabilitation | 48 
ventilator rehabilitation | 48 
oxygen therapy rehabilitation | 48 
vasopressor rehabilitation | 48 
inotrope rehabilitation | 48 
IV fluid rehabilitation | 48 
pericardiocentesis therapy | 3 
pericardial effusion therapy | 3 
cardiac tamponade therapy | 3 
multiple myeloma therapy | -8760 
plasma cell leukemia therapy | -8760 
intensive care therapy | 6 
ventilator therapy | 2 
oxygen therapy | 2 
vasopressor therapy | 1 
inotrope therapy | 1 
IV fluid therapy | 0 
pericardiocentesis medication | 3 
pericardial effusion medication | 3 
cardiac tamponade medication | 3 
multiple myeloma medication | -8760 
plasma cell leukemia medication | -8760 
intensive care medication | 6 
ventilator medication | 2 
oxygen medication | 2 
vasopressor medication | 1 
inotrope medication | 1 
IV fluid medication | 0 
pericardiocentesis treatment outcome | 6 
pericardial effusion treatment outcome | 6 
cardiac tamponade treatment outcome | 6 
multiple myeloma treatment outcome | 48 
plasma cell leukemia treatment outcome | 48 
intensive care treatment outcome | 6 
ventilator treatment outcome | 6 
oxygen therapy treatment outcome | 6 
vasopressor treatment outcome | 6 
inotrope treatment outcome | 6 
IV fluid treatment outcome | 6 
pericardiocentesis prognosis | 48 
pericardial effusion prognosis | 48 
cardiac tamponade prognosis | 48 
multiple myeloma prognosis | 48 
plasma cell leukemia prognosis | 48 
intensive care prognosis | 48 
ventilator prognosis | 48 
oxygen therapy prognosis | 48 
vasopressor prognosis | 48 
inotrope prognosis | 48 
IV fluid prognosis | 48 
pericardiocentesis survival rate | 48 
pericardial effusion survival rate | 48 
cardiac tamponade survival rate | 48 
multiple myeloma survival rate | 48 
plasma cell leukemia survival rate | 48 
intensive care survival rate | 48 
ventilator survival rate | 48 
oxygen therapy survival rate | 48 
vasopressor survival rate | 48 
inotrope survival rate | 48 
IV fluid survival rate | 48 
pericardiocentesis life expectancy | 48 
pericardial effusion life expectancy | 48 
cardiac tamponade life expectancy | 48 
multiple myeloma life expectancy | 48 
plasma cell leukemia life expectancy | 48 
intensive care life expectancy | 48 
ventilator life expectancy | 48 
oxygen therapy life expectancy | 48 
vasopressor life expectancy | 48 
inotrope life expectancy | 48 
IV fluid life expectancy | 48 
pericardiocentesis quality of life | 48 
pericardial effusion quality of life | 48 
cardiac tamponade quality of life | 48 
multiple myeloma quality of life | 48 
plasma cell leukemia quality of life | 48 
intensive care quality of life | 48 
ventilator quality of life | 48 
oxygen therapy quality of life | 48 
vasopressor quality of life | 48 
inotrope quality of life | 48 
IV fluid quality of life | 48 
pericardiocentesis patient outcome | 48 
pericardial effusion patient outcome | 48 
cardiac tamponade patient outcome | 48 
multiple myeloma patient outcome | 48 
plasma cell leukemia patient outcome | 48 
intensive care patient outcome | 48 
ventilator patient outcome | 48 
oxygen therapy patient outcome | 48 
vasopressor patient outcome | 48 
inotrope patient outcome | 48 
IV fluid patient outcome | 48 
pericardiocentesis patient survival | 48 
pericardial effusion patient survival | 48 
cardiac tamponade patient survival | 48 
multiple myeloma patient survival | 48 
plasma cell leukemia patient survival | 48 
intensive care patient survival | 48 
ventilator patient survival | 48 
oxygen therapy patient survival | 48 
vasopressor patient survival | 48 
inotrope patient survival | 48 
IV fluid patient survival | 48 
pericardiocentesis patient recovery | 48 
pericardial effusion patient recovery | 48 
cardiac tamponade patient recovery | 48 
multiple myeloma patient recovery | 48 
plasma cell leukemia patient recovery | 48 
intensive care patient recovery | 48 
ventilator patient recovery | 48 
oxygen therapy patient recovery | 48 
vasopressor patient recovery | 48 
inotrope patient recovery | 48 
IV fluid patient recovery | 48 
pericardiocentesis patient rehabilitation | 48 
pericardial effusion patient rehabilitation | 48 
cardiac tamponade patient rehabilitation | 48 
multiple myeloma patient rehabilitation | 48 
plasma cell leukemia patient rehabilitation | 48 
intensive care patient rehabilitation | 48 
ventilator patient rehabilitation | 48 
oxygen therapy patient rehabilitation | 48 
vasopressor patient rehabilitation | 48 
inotrope patient rehabilitation | 48 
IV fluid patient rehabilitation | 48 
pericardiocentesis patient aftercare | 48 
pericardial effusion patient aftercare | 48 
cardiac tamponade patient aftercare | 48 
multiple myeloma patient aftercare | 48 
plasma cell leukemia patient aftercare | 48 
intensive care patient aftercare | 48 
ventilator patient aftercare | 48 
oxygen therapy patient aftercare | 48 
vasopressor patient aftercare | 48 
inotrope patient aftercare | 48 
IV fluid patient aftercare | 48 
pericardiocentesis patient follow-up | 48 
pericardial effusion patient follow-up | 48 
cardiac tamponade patient follow-up | 48 
multiple myeloma patient follow-up | 48 
plasma cell leukemia patient follow-up | 48 
intensive care patient follow-up | 48 
ventilator patient follow-up | 48 
oxygen therapy patient follow-up | 48 
vasopressor patient follow-up | 48 
inotrope patient follow-up | 48 
IV fluid patient follow-up | 48 
pericardiocentesis patient therapy | 3 
pericardial effusion patient therapy | 3 
cardiac tamponade patient therapy | 3 
multiple myeloma patient therapy | -8760 
plasma cell leukemia patient therapy | -8760 
intensive care patient therapy | 6 
ventilator patient therapy | 2 
oxygen therapy patient therapy | 2 
vasopressor patient therapy | 1 
inotrope patient therapy | 1 
IV fluid patient therapy | 0 
pericardiocentesis patient medication | 3 
pericardial effusion patient medication | 3 
cardiac tamponade patient medication | 3 
multiple myeloma patient medication | -8760 
plasma cell leukemia patient medication | -8760 
intensive care patient medication | 6 
ventilator patient medication | 2 
oxygen therapy patient medication | 2 
vasopressor patient medication | 1 
inotrope patient medication | 1 
IV fluid patient medication | 0 
pericardiocentesis patient treatment outcome | 6 
pericardial effusion patient treatment outcome | 6 
cardiac tamponade patient treatment outcome | 6 
multiple myeloma patient treatment outcome | 48 
plasma cell leukemia patient treatment outcome | 48 
intensive care patient treatment outcome | 6 
ventilator patient treatment outcome | 6 
oxygen therapy patient treatment outcome | 6 
vasopressor patient treatment outcome | 6 
inotrope patient treatment outcome | 6 
IV fluid patient treatment outcome | 6 
pericardiocentesis patient prognosis | 48 
pericardial effusion patient prognosis | 48 
cardiac tamponade patient prognosis | 48 
multiple myeloma patient prognosis | 48 
plasma cell leukemia patient prognosis | 48 
intensive care patient prognosis | 48 
ventilator patient prognosis | 48 
oxygen therapy patient prognosis | 48 
vasopressor patient prognosis | 48 
inotrope patient prognosis | 48 
IV fluid patient prognosis | 48 
pericardiocentesis patient survival rate | 48 
pericardial effusion patient survival rate | 48 
cardiac tamponade patient survival rate | 48 
multiple myeloma patient survival rate | 48 
plasma cell leukemia patient survival rate | 48 
intensive care patient survival rate | 48 
ventilator patient survival rate | 48 
oxygen therapy patient survival rate | 48 
vasopressor patient survival rate | 48 
inotrope patient survival rate | 48 
IV fluid patient survival rate | 48 
pericardiocentesis patient life expectancy | 48 
pericardial effusion patient life expectancy | 48 
cardiac tamponade patient life expectancy | 48 
multiple myeloma patient life expectancy | 48 
plasma cell leukemia patient life expectancy | 48 
intensive care patient life expectancy | 48 
ventilator patient life expectancy | 48 
oxygen therapy patient life expectancy | 48 
vasopressor patient life expectancy | 48 
inotrope patient life expectancy | 48 
IV fluid patient life expectancy | 48 
pericardiocentesis patient quality of life | 48 
pericardial effusion patient quality of life | 48 
cardiac tamponade patient quality of life | 48 
multiple myeloma patient quality of life | 48 
plasma cell leukemia patient quality of life | 48 
intensive care patient quality of life | 48 
ventilator patient quality of life | 48 
oxygen therapy patient quality of life | 48 
vasopressor patient quality of life | 48 
inotrope patient quality of life | 48 
IV fluid patient quality of life | 48 
pericardiocentesis patient outcome | 48 
pericardial effusion patient outcome | 48 
cardiac tamponade patient outcome | 48 
multiple myeloma patient outcome | 48 
plasma cell leukemia patient outcome | 48 
intensive care patient outcome | 48 
ventilator patient outcome | 48 
oxygen therapy patient outcome | 48 
vasopressor patient outcome | 48 
inotrope patient outcome | 48 
IV fluid patient outcome | 48 
pericardiocentesis patient survival | 48 
pericardial effusion patient survival | 48 
cardiac tamponade patient survival | 48 
multiple myeloma patient survival | 48 
plasma cell leukemia patient survival | 48 
intensive care patient survival | 48 
ventilator patient survival | 48 
oxygen therapy patient survival | 48 
vasopressor patient survival | 48 
inotrope patient survival | 48 
IV fluid patient survival | 48 
pericardiocentesis patient recovery | 48 
pericardial effusion patient recovery | 48 
cardiac tamponade patient recovery | 48 
multiple myeloma patient recovery | 48 
plasma cell leukemia patient recovery | 48 
intensive care patient recovery | 48 
ventilator patient recovery | 48 
oxygen therapy patient recovery | 48 
vasopressor patient recovery | 48 
inotrope patient recovery | 48 
IV fluid patient recovery | 48 
pericardiocentesis patient rehabilitation | 48 
pericardial effusion patient rehabilitation | 48 
cardiac tamponade patient rehabilitation | 48 
multiple myeloma patient rehabilitation | 48 
plasma cell leukemia patient rehabilitation | 48 
intensive care patient rehabilitation | 48 
ventilator patient rehabilitation | 48 
oxygen therapy patient rehabilitation | 48 
vasopressor patient rehabilitation | 48 
inotrope patient rehabilitation | 48 
IV fluid patient rehabilitation | 48 
pericardiocentesis patient aftercare | 48 
pericardial effusion patient aftercare | 48 
cardiac tamponade patient aftercare | 48 
multiple myeloma patient aftercare | 48 
plasma cell leukemia patient aftercare | 48 
intensive care patient aftercare | 48 
ventilator patient aftercare | 48 
oxygen therapy patient aftercare | 48 
vasopressor patient aftercare | 48 
inotrope patient aftercare | 48 
IV fluid patient aftercare | 48 
pericardiocentesis patient follow-up | 48 
pericardial effusion patient follow-up | 48 
cardiac tamponade patient follow-up | 48 
multiple myeloma patient follow-up | 48 
plasma cell leukemia patient follow-up | 48 
intensive care patient follow-up | 48 
ventilator patient follow-up | 48 
oxygen therapy patient follow-up | 48 
vasopressor patient follow-up | 48 
inotrope patient follow-up | 48 
IV fluid patient follow-up | 48 
pericardiocentesis patient therapy | 3 
pericardial effusion patient therapy | 3 
cardiac tamponade patient therapy | 3 
multiple myeloma patient therapy | -8760 
plasma cell leukemia patient therapy | -8760 
intensive care patient therapy | 6 
ventilator patient therapy | 2 
oxygen therapy patient therapy | 2 
vasopressor patient therapy | 1 
inotrope patient therapy | 1 
IV fluid patient therapy | 0 
pericardiocentesis patient medication | 3 
pericardial effusion patient medication | 3 
cardiac tamponade patient medication | 3 
multiple myeloma patient medication | -8760 
plasma cell leukemia patient medication | -8760 
intensive care patient medication | 6 
ventilator patient medication | 2 
oxygen therapy patient medication | 2 
vasopressor patient medication | 1 
inotrope patient medication | 1 
IV fluid patient medication | 0 
pericardiocentesis patient treatment outcome | 6 
pericardial effusion patient treatment outcome | 6 
cardiac tamponade patient treatment outcome | 6 
multiple myeloma patient treatment outcome | 48 
plasma cell leukemia patient treatment outcome | 48 
intensive care patient treatment outcome | 6 
ventilator patient treatment outcome | 6 
oxygen therapy patient treatment outcome | 6 
vasopressor patient treatment outcome | 6 
inotrope patient treatment outcome | 6 
IV fluid patient treatment outcome | 6 
pericardiocentesis patient prognosis | 48 
pericardial effusion patient prognosis | 48 
cardiac tamponade patient prognosis | 48 
multiple myeloma patient prognosis | 48 
plasma cell leukemia patient prognosis | 48 
intensive care patient prognosis | 48 
ventilator patient prognosis | 48 
oxygen therapy patient prognosis | 48 
vasopressor patient prognosis | 48 
inotrope patient prognosis | 48 
IV fluid patient prognosis | 48 
pericardiocentesis patient survival rate | 48 
pericardial effusion patient survival rate | 48 
cardiac tamponade patient survival rate | 48 
multiple myeloma patient survival rate | 48 
plasma cell leukemia patient survival rate | 48 
intensive care patient survival rate | 48 
ventilator patient survival rate | 48 
oxygen therapy patient survival rate | 48 
vasopressor patient survival rate | 48 
inotrope patient survival rate | 48 
IV fluid patient survival rate | 48 
pericardiocentesis patient life expectancy | 48 
pericardial effusion patient life expectancy | 48 
cardiac tamponade patient life expectancy | 48 
multiple myeloma patient life expectancy | 48 
plasma cell leukemia patient life expectancy | 48 
intensive care patient life expectancy | 48 
ventilator patient life expectancy | 48 
oxygen therapy patient life expectancy | 48 
vasopressor patient life expectancy | 48 
inotrope patient life expectancy | 48 
IV fluid patient life expectancy | 48 
pericardiocentesis patient quality of life | 48 
pericardial effusion patient quality of life | 48 
cardiac tamponade patient quality of life | 48 
multiple myeloma patient quality of life | 48 
plasma cell leukemia patient quality of life | 48 
intensive care patient quality of life | 48 
ventilator patient quality of life | 48 
oxygen therapy patient quality of life | 48 
vasopressor patient quality of life | 48 
inotrope patient quality of life | 48 
IV fluid patient quality of life | 48 
pericardiocentesis patient outcome | 48 
pericardial effusion patient outcome | 48 
cardiac tamponade patient outcome | 48 
multiple myeloma patient outcome | 48 
plasma cell leukemia patient outcome | 48 
intensive care patient outcome | 48 
ventilator patient outcome | 48 
oxygen therapy patient outcome | 48 
vasopressor patient outcome | 48 
inotrope patient outcome | 48 
IV fluid patient outcome | 48 
pericardiocentesis patient survival | 48 
pericardial effusion patient survival | 48 
cardiac tamponade patient survival | 48 
multiple myeloma patient survival | 48 
plasma cell leukemia patient survival | 48 
intensive care patient survival | 48 
ventilator patient survival | 48 
oxygen therapy patient survival | 48 
vasopressor patient survival | 48 
inotrope patient survival | 48 
IV fluid patient survival | 48 
pericardiocentesis patient recovery | 48 
pericardial effusion patient recovery | 48 
cardiac tamponade patient recovery | 48 
multiple myeloma patient recovery | 48 
plasma cell leukemia patient recovery | 48 
intensive care patient recovery | 48 
ventilator patient recovery | 48 
oxygen therapy patient recovery | 48 
vasopressor patient recovery | 48 
inotrope patient recovery | 48 
IV fluid patient recovery | 48 
pericardiocentesis patient rehabilitation | 48 
pericardial effusion patient rehabilitation | 48 
cardiac tamponade patient rehabilitation | 48 
multiple myeloma patient rehabilitation | 48 
plasma cell leukemia patient rehabilitation | 48 
intensive care patient rehabilitation | 48 
ventilator patient rehabilitation | 48 
oxygen therapy patient rehabilitation | 48 
vasopressor patient rehabilitation | 48 
inotrope patient rehabilitation | 48 
IV fluid patient rehabilitation | 48 
pericardiocentesis patient aftercare | 48 
pericardial effusion patient aftercare | 48 
cardiac tamponade patient aftercare | 48 
multiple myeloma patient aftercare | 48 
plasma cell leukemia patient aftercare | 48 
intensive care patient aftercare | 48 
ventilator patient aftercare | 48 
oxygen therapy patient aftercare | 48 
vasopressor patient aftercare | 48 
inotrope patient aftercare | 48 
IV fluid patient aftercare | 48 
pericardiocentesis patient follow-up | 48 
pericardial effusion patient follow-up | 48 
cardiac tamponade patient follow-up | 48 
multiple myeloma patient follow-up | 48 
plasma cell leukemia patient follow-up | 48 
intensive care patient follow-up | 48 
ventilator patient follow-up | 48 
oxygen therapy patient follow-up | 48 
vasopressor patient follow-up | 48 
inotrope patient follow-up | 48 
IV fluid patient follow-up | 48 
pericardiocentesis patient therapy | 3 
pericardial effusion patient therapy | 3 
cardiac tamponade patient therapy | 3 
multiple myeloma patient therapy | -8760 
plasma cell leukemia patient therapy | -8760 
intensive care patient therapy | 6 
ventilator patient therapy | 2 
oxygen therapy patient therapy | 2 
vasopressor patient therapy | 1 
inotrope patient therapy | 1 
IV fluid patient therapy | 0 
pericardiocentesis patient medication | 3 
pericardial effusion patient medication | 3 
cardiac tamponade patient medication | 3 
multiple myeloma patient medication | -8760 
plasma cell leukemia patient medication | -8760 
intensive care patient medication | 6 
ventilator patient medication | 2 
oxygen therapy patient medication | 2 
vasopressor patient medication | 1 
inotrope patient medication | 1 
IV fluid patient medication | 0 
pericardiocentesis patient treatment outcome | 6 
pericardial effusion patient treatment outcome | 6 
cardiac tamponade patient treatment outcome | 6 
multiple myeloma patient treatment outcome | 48 
plasma cell leukemia patient treatment outcome | 48 
intensive care patient treatment outcome | 6 
ventilator patient treatment outcome | 6 
oxygen therapy patient treatment outcome | 6 
vasopressor patient treatment outcome | 6 
inotrope patient treatment outcome | 6 
IV fluid patient treatment outcome | 6 
pericardiocentesis patient prognosis | 48 
pericardial effusion patient prognosis | 48 
cardiac tamponade patient prognosis | 48 
multiple myeloma patient prognosis | 48 
plasma cell leukemia patient prognosis | 48 
intensive care patient prognosis | 48 
ventilator patient prognosis | 48 
oxygen therapy patient prognosis | 48 
vasopressor patient prognosis | 48 
inotrope patient prognosis | 48 
IV fluid patient prognosis | 48 
pericardiocentesis patient survival rate | 48 
pericardial effusion patient survival rate | 48 
cardiac tamponade patient survival rate | 48 
multiple myeloma patient survival rate | 48 
plasma cell leukemia patient survival rate | 48 
intensive care patient survival rate | 48 
ventilator patient survival rate | 48 
oxygen therapy patient survival rate | 48 
vasopressor patient survival rate | 48 
inotrope patient survival rate | 48 
IV fluid patient survival rate | 48 
pericardiocentesis patient life expectancy | 48 
pericardial effusion patient life expectancy | 48 
cardiac tamponade patient life expectancy | 48 
multiple myeloma patient life expectancy | 48 
plasma cell leukemia patient life expectancy | 48 
intensive care patient life expectancy | 48 
ventilator patient life expectancy | 48 
oxygen therapy patient life expectancy | 48 
vasopressor patient life expectancy | 48 
inotrope patient life expectancy | 48 
IV fluid patient life expectancy | 48 
pericardiocentesis patient quality of life | 48 
pericardial effusion patient quality of life | 48 
cardiac tamponade patient quality of life | 48 
multiple myeloma patient quality of life | 48 
plasma cell leukemia patient quality of life | 48 
intensive care patient quality of life | 48 
ventilator patient quality of life | 48 
oxygen therapy patient quality of life | 48 
vasopressor patient quality of life | 48 
inotrope patient quality of life | 48 
IV fluid patient quality of life | 48 
pericardiocentesis patient outcome | 48 
pericardial effusion patient outcome | 48 
cardiac tamponade patient outcome | 48 
multiple myeloma patient outcome | 48 
plasma cell leukemia patient outcome | 48 
intensive care patient outcome | 48 
ventilator patient outcome | 48 
oxygen therapy patient outcome | 48 
vasopressor patient outcome | 48 
inotrope patient outcome | 48 
IV fluid patient outcome | 48 
pericardiocentesis patient survival | 48 
pericardial effusion patient survival | 48 
cardiac tamponade patient survival | 48 
multiple myeloma patient survival | 48 
plasma cell leukemia patient survival | 48 
intensive care patient survival | 48 
ventilator patient survival | 48 
oxygen therapy patient survival | 48 
vasopressor patient survival | 48 
inotrope patient survival | 48 
IV fluid patient survival | 48 
pericardiocentesis patient recovery | 48 
pericardial effusion patient recovery | 48 
cardiac tamponade patient recovery | 48 
multiple myeloma patient recovery | 48 
plasma cell leukemia patient recovery | 48 
intensive care patient recovery | 48 
ventilator patient recovery | 48 
oxygen therapy patient recovery | 48 
vasopressor patient recovery | 48 
inotrope patient recovery | 48 
IV fluid patient recovery | 48 
pericardiocentesis patient rehabilitation | 48 
pericardial effusion patient rehabilitation | 48 
cardiac tamponade patient rehabilitation | 48 
multiple myeloma patient rehabilitation | 48 
plasma cell leukemia patient rehabilitation | 48 
intensive care patient rehabilitation | 48 
ventilator patient rehabilitation | 48 
oxygen therapy patient rehabilitation | 48 
vasopressor patient rehabilitation | 48 
inotrope patient rehabilitation | 48 
IV fluid patient rehabilitation | 48 
pericardiocentesis patient aftercare | 48 
pericardial effusion patient aftercare | 48 
cardiac tamponade patient aftercare | 48 
multiple myeloma patient aftercare | 48 
plasma cell leukemia patient aftercare | 48 
intensive care patient aftercare | 48 
ventilator patient aftercare | 48 
oxygen therapy patient aftercare | 48 
vasopressor patient aftercare | 48 
inotrope patient aftercare | 48 
IV fluid patient aftercare | 48 
pericardiocentesis patient follow-up | 48 
pericardial effusion patient follow-up | 48 
cardiac tamponade patient follow-up | 48 
multiple myeloma patient follow-up | 48 
plasma cell leukemia patient follow-up | 48 
intensive care patient follow-up | 48 
ventilator patient follow-up | 48 
oxygen therapy patient follow-up | 48 
vasopressor patient follow-up | 48 
inotrope patient follow-up | 48 
IV fluid patient follow-up | 48 
pericardiocentesis patient therapy | 3 
pericardial effusion patient therapy | 3 
cardiac tamponade patient therapy | 3 
multiple myeloma patient therapy | -8760 
plasma cell leukemia patient therapy | -8760 
intensive care patient therapy | 6 
ventilator patient therapy | 2 
oxygen therapy patient therapy | 2 
vasopressor patient therapy | 1 
inotrope patient therapy | 1 
IV fluid patient therapy | 0 
pericardiocentesis patient medication | 3 
pericardial effusion patient medication | 3 
cardiac tamponade patient medication | 3 
multiple myeloma patient medication | -8760 
plasma cell leukemia patient medication | -8760 
intensive care patient medication | 6 
ventilator patient medication | 2 
oxygen therapy patient medication | 2 
vasopressor patient medication | 1 
inotrope patient medication | 1 
IV fluid patient medication | 0 
pericardiocentesis patient treatment outcome | 6 
pericardial effusion patient treatment outcome | 6 
cardiac tamponade patient treatment outcome | 6 
multiple myeloma patient treatment outcome | 48 
plasma cell leukemia patient treatment outcome | 48 
intensive care patient treatment outcome | 6 
ventilator patient treatment outcome | 6 
oxygen therapy patient treatment outcome | 6 
vasopressor patient treatment outcome | 6 
inotrope patient treatment outcome | 6 
IV fluid patient treatment outcome | 6 
pericardiocentesis patient prognosis | 48 
pericardial effusion patient prognosis | 48 
cardiac tamponade patient prognosis | 48 
multiple myeloma patient prognosis | 48 
plasma cell leukemia patient prognosis | 48 
intensive care patient prognosis | 48 
ventilator patient prognosis | 48 
oxygen therapy patient prognosis | 48 
vasopressor patient prognosis | 48 
inotrope patient prognosis | 48 
IV fluid patient prognosis | 48 
pericardiocentesis patient survival rate | 48 
pericardial effusion patient survival rate | 48 
cardiac tamponade patient survival rate | 48 
multiple myeloma patient survival rate | 48 
plasma cell leukemia patient survival rate | 48 
intensive care patient survival rate | 48 
ventilator patient survival rate | 48 
oxygen therapy patient survival rate | 48 
vasopressor patient survival rate | 48 
inotrope patient survival rate | 48 
IV fluid patient survival rate | 48 
pericardiocentesis patient life expectancy | 48 
pericardial effusion patient life expectancy | 48 
cardiac tamponade patient life expectancy | 48 
multiple myeloma patient life expectancy | 48 
plasma cell leukemia patient life expectancy | 48 
intensive care patient life expectancy | 48 
ventilator patient life expectancy | 48 
oxygen therapy patient life expectancy | 48 
vasopressor patient life expectancy | 48 
inotrope