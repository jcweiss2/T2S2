37 years old | 0
male | 0
healthcare worker | 0
fever | -672
diarrhoea | -672
lethargy | -672
symptoms subsided | -552
recurrence of fever | -120
recurrence of diarrhoea | -120
dizziness | 0
admitted to the emergency department | 0
clinical shock | 0
blood pressure 75/50 | 0
heart rate 120 beats per minute | 0
febrile 39°C | 0
tachypnoeic >30 breaths per minute | 0
oxygen saturation 97% | 0
raised jugular venous pressure | 0
coarse crepitations | 0
global moderate-to-severe left ventricular systolic dysfunction | 0
transferred to critical care | 0
milrinone commenced | 0
noradrenaline commenced | 0
worsening myocardial function | 24
ejection fraction 25% | 24
intravenous immunoglobulin administered | 24
hydrocortisone commenced | 24
anticoagulation with heparin | 24
high-dose vitamin B & C initiated | 24
leucocytosis 36 × 10^9/L | 0
lymphopenia 0.6 × 10^9/L | 0
elevated troponin 490 ng/L | 0
brain natriuretic peptide >35,000 ng/L | 0
ferritin 8681 µg/L | 0
D-dimer 2782 ng/mL | 0
acute kidney injury | 0
creatinine 130 µmol/L | 0
coagulopathy INR 1.5 | 0
transaminitis ALT 538 U/L | 0
procalcitonin 14.78 µg/L | 0
negative blood cultures | 0
negative urine cultures | 0
negative stool cultures | 0
negative nasopharyngeal swab Day 1 | 0
negative nasopharyngeal swab Day 3 | 72
negative nasopharyngeal swab Day 5 | 120
negative influenza test | 0
negative HIV test | 0
normal serum autoimmune panel | 0
sinus tachycardia | 0
bilateral lower lobe consolidation | 0
small pleural effusions | 0
linezolid commenced | 0
clarithromycin commenced | 0
piperacillin-tazobactam commenced | 0
worsening biventricular function | 72
LVEF reduction to 21% | 72
right ventricular function worsening | 72
LV wall thickening | 72
bi-atrial dilatation | 72
increased pulmonary artery systolic pressures | 72
LVEF improvement to 29% | 120
prednisolone substituted for hydrocortisone | 168
rapid recovery in myocardial function | 168
troponin 108 ng/L | 264
radiological improvement in cardiac function | 264
CMR evidence of myocarditis | 264
LV wall thickening | 264
inhomogeneity of T1/T2 mapping | 264
patchy non-infarct pattern late gadolinium enhancement | 264
LVEF 70% | 264
normalization of RV volumes | 264
SARS-CoV-2 IgG positive | 312
ACE inhibitor commenced | 288
beta-blocker commenced | 288
mineralocorticoid receptor antagonist commenced | 288
discharged | 336
prednisolone 40 mg | 336
troponin normalization | 456
BNP normalization | 456
absence of dizziness | 456
improved exercise tolerance | 456
repeat CMR significant improvement | 696
patchy late gadolinium enhancement | 696
normal biventricular size | 696
normal systolic function | 696
prednisolone weaning reduced by 1 mg every 3 weeks | 4992
prednisolone 4 mg | 4992
beta-blocker continued | 4992
ACE inhibitor continued | 4992
MRA continued | 4992
