90 years old | 0
    female | 0
    presented to the emergency department | 0
    hematemesis (five episodes) | 0
    low back pain | -672
    taking nonsteroidal anti-inflammatory medications | -672
    hypertension | 0
    stable vitals | 0
    unremarkable physical examination | 0
    urgent esophagogastroduodenoscopy (OGD) | 0
    Mallory Weiss tear in the esophagus | 0
    Forrest 1a ulcer on the anterior wall of the first to second part of the duodenum | 0
    hemoclips deployed to the duodenal ulcer | 0
    hemostasis (OGD) | 0
    intravenous proton pump inhibitor | 0
    hemodynamic instability (three days later) | 72
    drop in hemoglobin (9.0 to 6.5 g/dL) | 72
    second OGD | 72
    slow active bleeding from vessel at site of intact clips | 72
    additional hemoclips and adrenaline injection | 72
    hemostasis (second OGD) | 72
    melena (twelve days later) | 288
    repeat OGD | 288
    friable tissue | 288
    active bleeding at site of previous duodenal ulcer | 288
    three hemoclips deployed | 288
    CT mesenteric angiogram | 288
    no evidence of bleeding from the gastrointestinal tract | 288
    no signs of pancreatitis | 288
    refractory UGI bleeding | 288
    referred to Interventional Radiology | 288
    embolize the GDA | 288
    super selective angiograms of the GDA, SPDA, and IPDA | 288
    no active contrast extravasation | 288
    no pseudoaneurysm | 288
    embolization of the GDA using microcoils | 288
    no gel foam or particles used | 288
    completion angiograms | 288
    no contrast opacification of the GDA | 288
    sudden onset of severe epigastric pain | 288
    hematemesis (post embolization) | 288
    remained hemodynamically stable | 288
    urgent OGD (post embolization) | 288
    fresh blood in the esophagus | 288
    large blood clot in the gastric antrum extending to the pylorus | 288
    blood in the duodenum | 288
    increased serum amylase (716 U/L) | 288
    increased serum lipase (>600 U/L) | 288
    normal liver enzymes | 288
    exploratory laparotomy with pyloromyoduodenotomy | 288
    gastrojejunal bypass | 288
    edematous pancreas | 288
    generalized bruising | 288
    fat saponification on the surface | 288
    hemorrhagic pancreatitis | 288
    recovery in surgical intensive care unit | 288
    high dependency unit | 288
    pseudomonas septicemia | 288
    atrial fibrillation | 288
    CT scan (1 week later) | 384
    acute focal pancreatitis | 384
    loculated peripancreatic collection extending into the lesser sac | 384
    failed to recover | 384
    died from multiorgan failure | 384
    