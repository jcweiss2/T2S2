47 years old | 0
female | 0
poorly controlled type 1 diabetes mellitus (T1DM) | -1464
heart failure with a mildly reduced ejection fraction of 47% | -1464
mild severe acute coronavirus respiratory virus-2 (SARS-COV-2) | -1464
left lower extremity deep vein thrombosis | -1464
presented with altered mental status | 0
presented with a burning sensation of her left hand | 0
cachectic | 0
alert to self | 0
appeared comfortable | 0
blood pressure of 104/65 mmHg | 0
pulse of 88 beats/min | 0
respiratory rate of 20 breaths/min | 0
oxygen saturation of 99% on room air | 0
wet gangrene of the left fourth digit | 0
leukocytosis | 0
white blood cell count of 15 ×10(9)/L | 0
acute kidney injury | 0
creatinine of 6.63 mg/dl | 0
diabetic ketoacidosis (DKA) | 0
glucose of 746 mg/dl | 0
anion gap of 30 | 0
X-ray of the left hand revealed atrophy of the fourth digit with subcutaneous gas | 0
CT scan of the brain was unremarkable | 0
CT scan of the abdomen and pelvis revealed consolidative and reticular opacities in the right lower lung | 0
CT scan of the chest showed a cavitary right lower lobe lesion with possible reversed halo sign | 0
started on vancomycin | 0
started on piperacillin-tazobactam | 0
started on clindamycin | 0
admitted to the intensive care unit (ICU) | 0
management of DKA | 0
sepsis from suspected pulmonary and skin/soft tissue infections | 0
resolution of DKA on hospital day 2 | 48
taken to the operating room for amputation of her left fourth digit | 48
concern for a necrotizing hand infection from a gas-producing organism | 48
no viable tissue observed throughout the hand | 48
left wrist disarticulation | 48
worsening leukocytosis | 72
white blood cell count peaked at 54,320 | 72
antimicrobial coverage broadened to vancomycin | 72
antimicrobial coverage broadened to meropenem | 72
antimicrobial coverage broadened to doxycycline | 72
addition of liposomal amphotericin B on hospital day 3 | 72
concern for underlying invasive fungal infection (IFI) | 72
pending surgical pathology results | 72
pending infectious studies (bacterial, fungal, and mycobacterial cultures) | 72
pending autoimmune laboratory panel | 72
bronchoscopy performed | 72
infiltrates of the right middle and lower lobe | 72
diffuse necrotic tissue past the right lower lobe bronchus with fibrinous clot | 72
concerning for IFI | 72
thoracic surgery consulted | 72
right lower lobectomy performed | 72
surgical source control through a posterolateral thoracotomy | 72
posaconazole added to anti-fungal regimen | 72
evaluation for dissemination of IFI | 72
bilateral frontal lobe punctate infarcts on MRI of the brain | 72
1.6 centimeter right atrial vegetation | 72
patent foramen ovale (PFO) on TEE | 72
urgent AngioVac extraction of the right atrial vegetation | 72
elevated risk of right-to-left embolization through PFO | 72
intraoperatively noted small vegetation not seen on pre-operative TEE | 72
suspected embolized vegetation | 72
no tissue obtained for culture or pathology | 72
bronchoalveolar lavage cytologic specimen demonstrated pauciseptate hyphae of a zygomycete | 72
right lower lobe surgical specimen demonstrated pauciseptate hyphae of a zygomycete | 72
left hand surgical specimen demonstrated pauciseptate hyphae of a zygomycete | 72
cultures grew a Rhizopus species | 72
hyphae present within vessels | 72
hyphae around nerves | 72
transferred to the general medicine floor | 72
re-admitted to the ICU for hypothermia | 144
re-admitted to the ICU for hypotension requiring vasopressor support | 144
prolonged hospital course complicated by acute metabolic encephalopathy | 144
bilateral pleural effusions managed with percutaneous drains | 144
acute kidney injury | 144
mixed transaminitis thought secondary to antifungal medications | 144
poor prognosis of disseminated mucormycosis | 144
progressive renal dysfunction | 144
progressive hepatic dysfunction | 144
family decided to discontinue further treatment | 144
transitioned to comfort care | 144
passed away | 144
