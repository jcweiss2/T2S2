36 years old | 0
    woman | 0
    presented to emergency room | 0
    34 weeks of gestation | 0
    worsening dyspnea | -48
    severe vomiting | -48
    poor oral intake | -48
    bronchial asthma diagnosed | -168000
    age 15 years | -168000
    experienced 2 episodes of near-fatal asthma | -168000
    misperception regarding effects of asthma medications during pregnancy | -672
    stopped taking asthma medication since becoming pregnant | -672
    increased asthma attack frequency | -168
    frequent use of rescue medication | -168
    denied smoking history | 0
    denied alcohol consumption | 0
    denied illicit drug usage | 0
    outpatient labor surveillance | -672
    glucose tolerance testing | -672
    no abnormalities | -672
    clear consciousness | 0
    agitated | 0
    tachypnea | 0
    inspiratory wheezing | 0
    expiratory wheezing | 0
    Kussmaul breathing | 0
    pulse 138 beats/min | 0
    respiratory rate 25 breaths/min | 0
    blood pressure 126/78 mm Hg | 0
    temperature 37°C | 0
    height 1.65 m | 0
    weight 72.2 kg | 0
    arterial blood gas analysis | 0
    mixed respiratory alkalosis | 0
    metabolic acidosis | 0
    no hypoxia | 0
    supplemental oxygen | 0
    high-dose short-acting beta-agonist | 0
    ipratropium via nebulizer | 0
    intravenous steroids | 0
    condition deteriorated | 0
    high respiratory rate | 0
    accessory muscle use | 0
    intubated | 2
    admitted to ER | 0
    prevented maternal fatigue | 0
    deterioration of oxygenation | 0
    postintubation ventilator settings | 2
    pressure-control ventilation mode | 2
    pressure level 18 cm H2O | 2
    respiratory rate 15 breaths/min | 2
    PEEP 5 cm H2O | 2
    FiO2 80% | 2
    Ti 1 s | 2
    hydrated with 0.9% saline | 2
    severe vomiting | -48
    fetal viability monitored | 0
    cardiotocography | 0
    blood tests | 0
    elevated C-reactive protein | 0
    leucocyte count 15.85 × 109/L | 0
    normal renal function | 0
    normal liver function | 0
    normal creatinine kinase | 0
    random capillary blood glucose 152 mg/dL | 0
    normal glycosylated hemoglobin | 0
    urinalysis | 0
    2+ acetone | 0
    no glycosuria | 0
    no proteinuria | 0
    admitted to ICU | 8
    intubation | 2
    initial management in ER | 0
    adjusted ventilator settings | 8
    pressure-support ventilation | 8
    pressure level 16 cm H2O | 8
    PEEP 8 cm H2O | 8
    FiO2 50% | 8
    administered inhaled short-acting beta-agonist | 8
    inhaled corticosteroid | 8
    intravenous magnesium sulfate | 8
    breathless | 8
    deep breathing | 8
    labored breathing | 8
    dynamic hyperinflation | 8
    intrinsic end-expiratory pressure | 8
    adjusted ventilator settings to lower tidal volumes | 8
    tidal volumes 6–8 mL/kg | 8
    ideal body weight 55.8 kg | 8
    sedated with propofol | 8
    rapid respiratory rates | 8
    intermittent high tidal volume | 8
    high minute ventilation | 8
    partial sedation | 8
    no response to high-dose propofol | 8
    labored breathing | 8
    chest radiography | 8
    subcutaneous emphysema | 8
    suspected pneumomediastinum | 8
    follow-up arterial blood gas analysis | 29
    decreased bicarbonate levels | 29
    increased anion gap | 29
    respiratory compensation | 29
    worsening metabolic acidosis | 29
    labored breathing | 29
    deep breathing | 29
    difficult to control asthma | 29
    lactic acidosis unlikely | 29
    normal serum lactate | 29
    sepsis work-up | 29
    no infection | 29
    serum ketone levels 3.7 mmol/L | 29
    pH 7.216 | 29
    bicarbonate 11.6 mmol/L | 29
    high anion gap metabolic acidosis | 29
    diagnosed starvation ketoacidosis | 29
    vomiting | 29
    stress during third trimester | 29
    hydrated with D5NS | 29
    partially resolved ketoacidosis | 29
    aggressive treatment for asthma attack | 29
    concern for beta-agonist and corticosteroid effects | 29
    high-dose propofol adverse effects | 29
    emergency caesarean section | 29
    general anesthesia | 29
    betamethasone administered | 29
    prevented fetal respiratory distress syndrome | 29
    delivered 2.3 kg girl | 29
    umbilical cord arterial pH 7.143 | 29
    Apgar score 9 | 29
    intensive care for newborn | 29
    extubated | 49
    post-delivery | 29
    rapid resolution of metabolic derangement | 29
    panendoscopy | 29
    superficial gastritis | 29
    mother discharged | 49
    baby discharged | 49
    favorable outcome | 49
    ketoacidosis induced by short-term starvation | 29
    near-fatal asthma attack | 29
    nondiabetic | 0
    pregnant | 0
    third trimester | 0
    placenta-derived hormones contribution | 29
    fuel homeostasis during starvation | 29
    stress during pregnancy | 29
    pharmacological effects | 29
    acidosis reversal via caesarean delivery | 29
    favorable outcome | 49
    life-threatening events | 0
    acidosis | 0
    asthma | 0
    conflicting treatments | 0
    emergency caesarean section delivery | 29
    ketoacidosis and asthma resolved | 49
    uncontrolled asthma | 29
    high anion gap metabolic derangement | 29
    GOLD MARK mnemonic | 29
    glycols excluded | 29
    5-oxoproline excluded | 29
    lactate excluded | 29
    methanol excluded | 29
    aspirin excluded | 29
    renal failure excluded | 29
    rhabdomyolysis excluded | 29
    ketoacidosis diagnosis | 29
    previously healthy | 0
    nonalcoholic | 0
    nondiabetic | 0
    no ketogenic diet | 0
    no long-term fasting | 0
    no previous ketoacidosis episodes | 0
    normal blood glucose | 0
    normal glycosylated hemoglobin | 0
    metabolic alkalosis from vomiting | -48
    respiratory alkalosis | 0
    short-term fasting | -48
    insulinopenia | 29
    insulin resistance | 29
    accelerated starvation | 29
    third trimester | 0
    lipid metabolism adaptation | 29
    placenta-derived hormones | 29
    cortisol | 29
    glucagon | 29
    gluconeogenesis | 29
    glycogenolysis | 29
    ketogenesis | 29
    increased glucose counter-regulatory hormones | 29
    pharmacological effects | 29
    beta# 网络拓扑结构

## 网络结构图
![网络结构图](NetworkTopology.png)

## 网络结构说明
网络结构中存在四个服务器，两个服务器位于内网，两个位于公网。其中，公网的服务器有两个：一个用于运行主程序（如网站服务），另一个用于代理服务器；内网的两台服务器，一台用于数据库，另一台用于缓存。

## 访问流程说明
用户通过访问代理服务器来获取服务。代理服务器作为入口，将请求分发到内网的主程序服务器。主程序在处理请求时，根据需要会访问缓存服务器或数据库服务器。这种结构确保了主程序服务器不直接暴露于公网，提高了安全性。同时，代理服务器还可能承担负载均衡和流量管理的职责。