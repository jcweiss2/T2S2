72 years old | 0
male | 0
right-hand dominant | 0
retired mechanic | 0
admitted to the hospital | 0
left shoulder remote rotator cuff injury | -672
adhesive capsulitis | -672
aneurysmal dilation of the ascending aorta | -672
mild aortic insufficiency | -672
crush injury to the left forearm and hand | -672
rib fractures | -672
pneumohemothorax | -672
acute treatment of injuries | -672
transferred to home hospital | -668
admitted to the intensive care unit | -668
symptoms of sepsis | -668
left upper extremity appeared to be infected | -668
imaging and surgical exploration | -668
preoperative x-ray | -668
surgery | -664
postoperative day 5 | -660
second surgery | -660
extensive debridement and lavage | -660
deep infection | -660
flexor carpi radialis nonviable | -660
hand intrinsic muscles nonviable | -660
long flexors nonviable | -660
extensors nonviable | -660
wound packed | -660
surgery ended | -660
discussion of limb salvage versus amputation | -660
postoperative day 7 | -657
transradial below-elbow amputation | -657
postoperative day 19 | -649
debridement of the amputation site | -649
split-thickness skin grafting | -649
recovered well | -649
discharged home | -645
referral for prosthetic fitting and training | -645
rehabilitation and prosthetic fitting impaired by PLP | -645
PLP | -645
intense sensation of flexion and cramping of digits 1 to 3 | -645
short-term trials of medication | -645
avoid long-term daily medication use | -645
nonpharmacological management | -645
multiple modifications to the socket | -645
desensitization therapy | -645
compressive stump covers | -645
mirror therapy | -645
discontinuation of prosthesis use | -645
gabapentin | -645
pregabalin | -645
tramadol | -645
hydromorphone | -645
xylocaine injections | -645
x-ray of the residual limb | -624
heterotopic ossification | -624
median nerve | -624
local HO in close anatomical proximity to the median nerve | -624
management options reviewed | -624
daily bisphosphonates | -624
analgesic effects | -624
patient refused long-term daily treatments | -624
calcitonin | -624
possible treatment option for PLP | -624
possible aid in HO management | -624
two-week trial of intranasal calcitonin | -624
extension to four weeks | -624
one month follow-up | -592
significant reduction in PLP | -592
discontinued all other scheduled and as-needed analgesic medication | -592
not returned to using the prosthesis | -592
three-month follow-up | -564
pain at a minimum | -564
repeat x-ray | -564
no progression of HO | -564
six-month follow-up | -536
returned to prosthesis use | -536
18-month follow-up | -468
minimal phantom pain | -468
continued prosthesis use | -468
no desire to pursue surgical management with HO excision | -468