52 years old | 0
male | 0
goiter | -504
neck pain | -168
dysphagia | -168
difficulty breathing | -168
thyroidectomy | -504
post-operative hematoma | -504
Jackson-Pratt wound drain placement | -504
neck enlargement | 0
neck tenderness | 0
normal PT | 0
normal INR | 0
normal PTT | 0
normal fibrinogen | 0
neck hematoma (CT scan) | 0
hematoma evacuation (otolaryngology) | 0
desmopressin (DDAVP) administration | 0
cessation of bleeding | 0
discharge | 0
severe oral mucosal bleeding (post-dental) | 12960
ICU admission | 12960
red blood cell transfusion | 12960
platelet transfusion | 12960
fresh frozen plasma transfusion | 12960
DDAVP administration | 12960
Humate-P administration | 12960
aminocaproic acid administration | 12960
surgical packing | 12960
bleeding control | 12960
normal PTT | 12960
normal Factor II | 12960
normal Factor V | 12960
normal Factor VII | 12960
normal Factor VIII | 12960
normal Factor IX | 12960
normal Factor X | 12960
normal Factor XI | 12960
normal Factor XII | 12960
normal Von Willebrand Factor antigen | 12960
normal Von Willebrand activity | 12960
normal platelet function assay | 12960
prolonged PT (13.9s) | 12960
elevated INR (1.3) | 12960
PT mixing study corrected | 12960
definitive diagnosis not established | 12960
bleeding diathesis education | 12960
aminocaproic acid taper | 12960
hematology follow-up | 12960
failure to follow-up (socio-financial) | 12960
abdominal pain | 21600
distention | 21600
massive hepatosplenomegaly | 21600
no liver disease history | 21600
no alcohol abuse | 21600
coagulopathy workup initiated | 21600
elevated PT | 21600
PT mixing study corrected | 21600
Factor VII deficiency (29%) | 21600
transjugular liver biopsy planned | 21600
recombinant factor VIIa (rFVIIa) prophylaxis | 21600
vitamin K prophylaxis | 21600
liver biopsy (Congo red stain) | 21600
AL (kappa) amyloid deposition | 21600
readmission for biopsy site bleeding | 21600
bleeding control (rFVIIa, vitamin K) | 21600
readmission for abdominal pain | 21600
retroperitoneal hematoma | 21600
ICU admission | 21600
FFP transfusion | 21600
cryoprecipitate transfusion | 21600
aminocaproic acid infusion | 21600
vitamin K supplementation | 21600
slight bleeding control | 21600
rFVIIa scheduled dosing | 21600
factor VII level correction | 21600
PT/INR correction | 21600
hemoglobin stabilization | 21600
weaned off rFVIIa | 21600
acquired factor VII deficiency diagnosis | 21600
hepatic amyloidosis | 21600
AL amyloidosis-kappa subtype | 21600
serum protein electrophoresis (no M-spike) | 21600
urine protein electrophoresis (no M-spike) | 21600
elevated serum free light chain ratio (5.65) | 21600
bone marrow biopsy declined | 21600
bortezomib treatment | 21600
dexamethasone treatment | 21600
cyclophosphamide treatment | 21600
4 cycles completed | 21600
progressive liver dysfunction | 21600
cardiac amyloidosis | 21600
cardiac MRI (amyloid infiltration) | 21600
echocardiogram (LV diastolic dysfunction) | 21600
elevated pro BNP (2,012) | 21600
normal ALT | 21600
normal AST | 21600
elevated INR (3.9) | 21600
elevated PTT (43) | 21600
creatinine (1.3) | 21600
esophageal variceal bleeding | 21600
variceal banding | 21600
severe ascites | 21600
spontaneous bacterial peritonitis | 21600
hepatic encephalopathy | 21600
bone marrow transplant evaluation | 21600
liver transplant evaluation | 21600
not a candidate (advanced disease) | 21600
GI bleeding episodes | 21600
rFVIIa administration (GI bleeding) | 21600
worsening coagulopathy | 21600
elevated PTT | 21600
colchicine treatment | 21600
prednisone treatment | 21600
completed 1 cycle | 21600
no improvement | 21600
uncontrolled upper GI bleeding | 21600
death | 21600
