23 years old | 0
female | 0
learning disability | -0
meningitis | -0
generalized abdominal pain | -48
admitted to hospital | 0
clinicobiological presentation of generalized peritonitis | 0
abdominal ultrasonography | 0
infiltration of the periappendicular fat | 0
intraperitoneal effusion | 0
septic shock | 0
median laparotomy | 0
perforation of a voluminous tumoral mass of the ceacum | 0
tumor fixed posteriorly | 0
tumor invades adjacent structures | 0
palpation of the liver | 0
palpation of the right annex | 0
no secondary lesions | 0
no nodules of carcinomatosis | 0
right mesocolon strewn with adenomegaly | 0
tumor adhered posteriorly to the second duodenum | 0
right hemicolectomy R2 | 0
ileostomy | 0
septic shock | 0
transfer to university hospital | 0
12 days stay in Intensive Care Unit | 12
pathological examination | 12
diagnosis of right colon schwannoma | 12
thoracoabdominopelvic CT scan | 48
tumoral residue at right iliac fossa | 48
no secondary site | 48
multidisciplinary meeting | 96
decision to make a complementary resection | 96
complementary resection not feasible | 96
tumoral residue invading right annex | 96
tumoral residue invading right iliac vessels | 96
tumoral residue invading right ureter | 96
restoring digestive continuity | 96
follow-up at outpatient clinic | 96
CT scanning control 2 years postoperatively | 730
tissue mass involving the small bowel | 730
mesenteric recurrence | 730
stability of the old tumoral residue | 730
exploratory laparotomy | 730
voluminous mass invading the root of the mesentery | 730
multiple parietal nodules | 730
surgical biopsies | 730
neurofibrmatous nature | 730
no adjuvant treatment | 730
multidisciplinary meeting | 730
no indication of radiotherapy or chemotherapy | 730
4 years follow-up | 1460
no complications | 1460
need for right nephrostomy | 1460
ureter compression by primary tumoral residue | 1460