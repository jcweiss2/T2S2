diabetes mellitus | 0
obesity | 0
consumed a bottle of rice wine thrice a week | 0
colonoscopy | 0
endoscopic mucosal resection | 0
preventive hemoclips applied | 0
discharged from the endoscopy room | 0
right abdominal pain | 24
tenderness | 24
rebound tenderness | 24
severe infection | 24
white blood cell count 21,460/mm3 | 24
C-reactive protein level 17.8 mg/dL | 24
blood urea nitrogen level 28 mg/dL | 24
creatinine 2.13 mg/dL | 24
lactic acid 2.4 mmol/L | 24
total bilirubin 1.7 mg/dL | 24
abdominopelvic computed tomography | 24
multiple air bubbles in the right lateral abdominal muscles | 24
broad-spectrum antibiotic therapy | 24
emergency exploratory laparotomy | 44
laparoscopic right hemicolectomy | 44
multiple-organ failure | 44
metabolic acidosis | 44
diagnosis of NF of the abdominal wall muscle | 48
urgent surgical debridement and drainage | 48
surgical debridement | 48
renal replacement therapy | 48
intensive care unit | 48
imipenem-resistant Acinetobacter baumannii | 72
extended spectrum beta-lactamase negative Escherichia coli | 72
septic shock | 840
multiple-organ failure | 840
death | 840