39 years old | 0
male | 0
Hispanic | 0
admitted to the hospital | 0
flu-like symptoms | -192
headache | -192
fatigue | -192
myalgia | -192
cough | -192
chills | -192
fever | 0
heart rate 133 beats/min | 0
blood pressure 118/76 mmHg | 0
respiratory rate 20 breaths/min | 0
oxygen saturation 94% | 0
diminished vesicular breath sounds | 0
oxygen saturation 89% | 3
oxygen supplementation via nasal cannula | 3
white blood cell count 7.8 K/uL | 0
venous blood gas pH 7.37 | 0
PaCO2 44 mmHg | 0
ferritin 635 ng/ml | 0
lactate dehydrogenase (LDH) 395 U/L | 0
multifocal infiltrates | 0
SARS-CoV-2 RNA positive | 0
intravenous fluids | 0
azithromycin | 0
ceftriaxone | 0
respiratory distress | 48
high flow nasal cannula oxygen | 48
intubation | 48
lung protective ventilation | 48
neuromuscular blockade | 48
sedation | 48
severe ARDS | 48
convalescent plasma | 48
methylprednisolone | 48
enoxaparin | 48
worsening ARDS | 144
refractory hypoxia | 144
VV-ECMO | 168
delirium | 168
Enterococcus faecalis bacteremia | 168
non-occlusive deep vein thrombosis | 168
tracheostomy | 864
decannulated | 1008
mechanical ventilation via pressure support ventilation | 1008
tracheostomy collar | 1016
SARS-CoV2 negative | 720
speech-language assessment | 720
oral diet | 720
CT chest | 720
aggressive daily rehabilitation treatment | 720
physical therapy (PT) | 720
occupational therapy (OT) | 720
ambulate independently | 1008
perform all activities of daily living (ADLs) independently | 1008
discharged home without oxygen supplementation | 1512
follow-up CT chest | 1532
complete resolution of the bilateral multifocal opacities | 1532
SARS-CoV-2 test negative | 1532
returned to baseline | 1532
no respiratory symptoms or complications | 1532