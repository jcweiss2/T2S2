40 years old | 0
Asian | 0
man | 0
parotid cancer | -87600
brain metastasis | -87600
lung metastasis | -87600
liver metastasis | -87600
bone metastasis | -87600
radiation | -87600
chemotherapy | -87600
palliative whole brain radiation (XRT) | -87600
urinary retention | -3
ascending paralysis to waist | -3
MRI | -3
large spinal tumor | -3
emergent XRT to spine | 0
rapid upper body weakness | 0
respiratory distress | 0
neuro-oncology team discussed prognosis | 0
offered palliative supportive measures | 0
offered intubation | 0
patient cognitively intact | 0
electively intubated | 0
without sedation | 0
anticipation of wife's arrival | 0
wife arrived | 24
neuro-oncology team updated wife | 24
grave prognosis | 24
patient stated "I want to die today" | 24
team restated wishes | 24
patient replied "take tube out, die today" | 24
wife requested privacy | 24
discussed withdrawal of life support | 48
patient mouthed "changed mind, want to live" | 48
feeding tube | 72
tracheotomy | 72
postoperative course | 72
pneumonia | 72
hypotension | 72
sepsis | 72
intensive care | 72
patient stated "I want to die" | 456
team advocated honoring wishes | 456
wife believed confusion | 456
patient cognitively intact | 456
patient said "take tube away, let me die" | 504
family meeting | 504
palliative care specialist involved | 504
wife disagreed to extubation | 504
wife unavailable | 504
patient condition deteriorated | 576
confused | 576
agitated | 576
wife requested meeting | 576
withdrawal of life support | 576
transferred to private room | 576
died peacefully | 578
extubation | 578
surrounded by wife, family, friends, neuro-oncology team | 578
