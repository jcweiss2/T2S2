79 years old | 0
female | 0
admitted to the hospital | 0
acute limb ischemia | -2
hypertension | -8760
atrial fibrillation | -8760
non-dialysis-dependent chronic renal failure | -8760
operated on for acute aortic embolic occlusion | -8760
bilateral femoral catheter embolectomy | -8760
started oral anticoagulation | -8760
pedal pulses | -8760
no posterior tibial pulses | -8760
irregular medication use | 0
international normalized ratio of prothrombin time | 0
arrhythmic pulse | 0
hypertensive | 0
normal femoral, popliteal and pedal pulses on right leg | 0
weak femoral pulse on left leg | 0
no distal pulses on left leg | 0
pain | 0
motor deficit | 0
grade IIb limb ischemia | 0
referred for surgery | 0
diminished creatinine clearance | 0
general anesthesia | 0
femoral access | 0
common, superficial and deep femoral arteries dissected and clamped | 0
arteriotomy | 0
embolectomy catheter used | 0
thrombi retrieved | 0
catheter progressed more than 60cm on superficial artery | 0
no significant back bleeding | 0
decision to perform angiography | 0
CO2 chosen as substitute for iodine contrast | 0
homemade water seal CO2 delivery system used | 0
injection performed through KMP 4Fr catheter | 0
patent popliteal artery | 0
patent fibular artery | 0
occlusion on mid-third of anterior tibial artery | 0
new embolectomy performed | 0
catheter progressed to foot | 0
more thrombi retrieved | 0
control angiography showed complete resolution of anterior tibial artery occlusion | 0
arteriorraphy performed | 0
pulses present on limb | 0
ischemia signs resolved | 0
no compartment syndrome signs | 0
remained in ICU | 0
no nephrotoxic agents used | 0
diuresis stimulated by furosemide | 0
developed urinary tract infection | 216
deteriorating renal function | 216
uremia | 216
dialysis started | 432
developed pneumonia | 864
septic shock | 864
required vasoactive drugs | 864
discharged to hospice care facility | 864
chronic dialysis | 864