50 years old | 0
male | 0
admitted to the hospital | 0
chronic pancreatitis | -720
epigastric abdominal pain | -48
generalized weakness | -48
chronic abdominal pain | -720
acetaminophen/oxycodone | -720
pancreatic enzyme replacement therapy | -720
blood pressure 100/92 mm Hg | 0
heart rate of 94 bpm | 0
respiratory rate of 16 breaths/min | 0
O2 saturation of 97% on room air | 0
epigastric tenderness | 0
diffuse calcifications | -720
hyperglycemic | 0
blood glucose of 703 mg/dL | 0
serum bicarbonate of 16 mmol/L | 0
ketones in the urine | 0
acetone in the blood | 0
anion gap corrected for albumin was 27 | 0
DKA | 0
NPO | 0
IV lactated Ringer’s solution with potassium | 0
IV insulin drip | 0
cardiac enzymes sent | 0
lipase sent | 0
septic workup sent | 0
cardiac enzymes within normal limits | 2
lipase elevated to 156 | 2
septic workup negative | 2
blood glucose monitored every hour | 0
electrolytes and albumin monitored every 4 h | 0
IV hydration continued | 0
potassium and dextrose adjustments | 0
anion gap closed | 24
transitioned to long-acting insulin detemir 10 Units SQ QHS | 24
diabetic diet | 26
insulin sliding scale | 24
discharged | 48
insulin aspart 3 Units TID with meals | 48
insulin detemir 10 Units QHS | 48
insulin detemir 6 Units QAM | 48
autoimmune workup for diabetes sent | 24
autoimmune workup negative | 48
ketorolac for abdominal pain | 48
follow up with primary care physician | 48
HbA1c values normal | -720
HbA1c 16% | 24