74 years old | 0
male | 0
type 2 diabetes mellitus | 0
admitted to the hospital | 0
vague abdominal and lower back pain | -168
leukocytosis | -3
white blood cell count of 25 × 10^9/L | -3
left shift | -3
recently traveled to Mexico | -672
dyspepsia | -672
upper gastrointestinal discomfort | -672
sore throat | -336
oral antibiotics | -336
magnetic resonance imaging | -3
aortic aneurysm | -3
computed tomography scan | -3
contained infrarenal aortic aneurysm rupture | -3
vancomycin | -1
piperacillin-tazobactam | -1
blood culturing | -1
autogenous NAIS reconstruction | 2
hemodynamic stability | 0
good health | 0
durable repair | 0
deep vein imaging | 0
ultrasound | 0
operating room preparation | 0
abdomen exploration | 2
right femoral vein harvested | 2
extensive retroperitoneal infection | 2
circumferential dissection | 2
infrarenal aortic clamp | 2
aorta and periaortic tissue debrided | 2
femoral vein graft sewn | 2
omentum flap created | 2
thigh wound irrigated | 2
thigh wound closed | 2
biphasic Doppler signals | 2
abdominal washout | 48
debridement | 48
extubated | 48
intensive care unit | 48
lower extremities elevated | 48
compressive bandage | 48
thigh-high compression stockings | 48
admission blood cultures | 0
intraoperative blood cultures | 2
group A streptococcus | 0
repeat blood cultures | 72
transthoracic echocardiography | 72
valvular vegetations | 72
antibiotic therapy narrowed | 72
ceftriaxone | 72
imaging studies | 336
minimal stranding | 336
omentum around aortic reconstruction | 336
prolonged ileus | 408
discharged home | 408
thigh-high stockings | 408
aspirin | 408
intravenous antibiotics | 408
follow-up with infectious disease department | 720
oral amoxicillin | 720
follow-up with vascular surgery department | 720
afebrile | 720
well-healed abdominal and right femoral incisions | 720
intact neurovascular examination | 720
stable imaging findings | 720
amoxicillin discontinued | 720
follow-up ultrasound examination | 1440
patent abdominal aorta and iliac arteries | 1440
abdominal aortic diameter | 1440
repeat CT angiography | 2520
normal graft | 2520
no aneurysm | 2520
no dissection | 2520
no stenosis | 2520
scheduled to follow-up annually | 2520
duplex ultrasound | 2520
ankle brachial index measurements | 2520