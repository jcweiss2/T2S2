59 years old | 0
Vietnamese woman | 0
presented to the emergency department following motor vehicle accident | 0
syncopal episode | 0
recent gastrointestinal illness | -48
no preceding pre-syncope | 0
no palpitations | 0
no chest pain | 0
no dyspnoea | 0
no urinary incontinence | 0
no tongue biting | 0
vomiting | -48
abdominal pain | -48
no fevers | 0
no diarrhoea | 0
received first COVID-19 vaccine | -336
heart rate 114 beats per min | 0
oxygen saturation 98% | 0
respiratory rate 16 | 0
blood pressure 120/77 | 0
afebrile | 0
alert | 0
oriented | 0
euvolaemic | 0
no murmurs on examination | 0
past medical history of thalassaemia | 0
no cardiovascular risk factors | 0
no prior history of seizures | 0
no significant family history | 0
initial ECG normal sinus rhythm | 0
fixed ST elevation anteriorly | 0
low QRS voltages | 0
cardiac troponin I 24,000 | 0
c-reactive protein 10 | 0
erythrocyte sedimentation rate 12 | 0
chest x-ray unremarkable | 0
calcified granuloma in right apex | 0
first TTE LVEF 30% | 0
normal left ventricle size | 0
moderate-severe global systolic dysfunction | 0
mild concentric increase in wall thickness | 0
severely reduced tissue Doppler velocities | 0
normal right ventricle size | 0
normal right ventricle function | 0
mild-mod aortic regurgitation | 0
moderate pericardial effusion | 0
deteriorated overnight with symptomatic hypotension | 24
bradycardia 30 beats per minute | 24
ECG high grade atrioventricular block | 24
left bundle branch block | 24
commenced on isoprenaline infusion | 24
transferred to coronary care unit | 24
expedited permanent pacemaker insertion | 24
persistently hypotensive | 48
systolic blood pressure 60 mmHg | 48
oliguric | 48
commenced on dopamine infusion | 48
conscious | 48
symptomatic episodes of brief accelerated idioventricular rhythm | 48
transferred to intensive care unit | 48
TTE LVEF 10% | 96
severe LV dysfunction | 96
global hypokinesis | 96
severely impaired RV systolic function | 96
dilated inferior vena cava | 96
endomyocardial biopsy performed | 96
florid infiltrate of lymphocytes | 96
histiocytes | 96
fewer plasma cells | 96
scattered eosinophils | 96
marked oedema | 96
cardiomyocyte necrosis | 96
occasional poorly formed granulomas | 96
loose aggregates of epithelioid histiocytes | 96
multinucleated macrophages with foamy appearing cytoplasm | 96
features consistent with giant cell myocarditis | 96
no coronary angiogram performed | 96
minimal risk factors for coronary artery disease | 96
atypical presentation for ACS | 96
global hypokinesis of LV | 96
increased LV wall thickness | 96
markedly reduced tissue Doppler velocities | 96
clinical instability | 96
commenced on methylprednisone | 96
commenced on cyclosporin | 96
developed worsening lactic acidosis | 96
intubated | 96
transferred to cardiac transplant centre | 120
biventricular assist device inserted | 120
haemorrhage | 120
coagulopathy requiring massive transfusion | 120
thoracic washout | 120
recovery of biventricular function | 120
progressive multiorgan failure | 168
hepatic encephalopathy | 168
anuric renal failure requiring dialysis | 168
distal ischaemia of all limbs | 168
digital gangrene | 168
presumed bowel ischaemia | 168
immune thrombocytopaenia | 168
treated with intravenous immunoglobulin | 168
plasma exchange | 168
polymicrobial sepsis | 168
Pseudomonas aeruginosa bacteraemia | 168
Candidaemia | 168
treated with meropenem | 168
vancomycin | 168
caspofungin | 168
LV assist device explanted | 432
redo-sternotomy | 432
tissue aortic valve replacement | 432
RV assist device explanted | 600
cerebral infarction | 600
unresponsive off sedation | 600
family meeting | 648
decision to palliate | 648
passed away | 648
