52 years old | 0
male | 0
body mass index of 23.6 kg/m2 | 0
no comorbidities | 0
began bariatric history | - 2002
began bariatric surgery | - 2002
weight 216 kg | - 2002
BMI 57.4 kg/m2 | - 2002
modified Scopinaro procedure | - 2002
weight reganance | - 2017
incisional hernia | - 2017
bariatric revisional surgery | - 2017
hernia repair | - 2017
weight 170 kg | - 2017
BMI 45.1 | - 2017
gastric pouch leak | - 2017
intra-abdominal collections | - 2017
sepsis | - 2017
conserved management | - 2017
open abdomen | - 2017
negative wound pressure therapy | - 2017
parenteral nutrition | - 2017
intravenous antibiotics | - 2017
epithelized gastrocutaneous fistula | - 2017
controlled but persistent drainage | - 2017
upper endoscopy | - 2017
fistulous orifice | - 2017
extraluminal extravasation | - 2017
recurrent left subphrenic abscess | - 2017
multiple attempts at fistula closure | - 2017
argon plasma coagulation | - 2017
internal and external drainages | - 2017
clipping | - 2017
fibrin sealants | - 2017
e-vac therapy | - 2017
stenting | - 2017
discouraged with multiple failed repair attempts | - 2017
referred for further evaluation | - 2017
multidisciplinary team discussion | - 2017
decision to proceed with an innovative endoscopic technique | - 2017
placement of a CSDO across the fistula orifice | - 2017
Occlutech muscular VSD occluder | - 2017
deployment of the CSDO | - 2017
immediate closure | - 2017
restricted oral intake | 24
liquid diet | 10
regular diet | 12
pigtail drain positioned at his left subphrenic abscess | 24
recurrence of the abscess | 24
partial dislodgment of the 8-mm mVSD CSDO | 24
sepsis | 24
computed tomography | 24
fluoroscopy | 24
recurrence of the abscess | 24
second attempt with an oversized disc | 24
Occlutech Figulla Flex II UNI 24-mm | 24
sealing the fistulous orifice | 24
former device positioned between the two discs of the new one | 24
6-month clinical and imaging follow-up | 6
upper endoscopy | 6
contrast-enhanced CT scan | 6
device engrafted | 6
significant reduction of the chronic abscess | 6
no signs of fistula recurrence | 6
pigtail was maintained in the subphrenic space | 6
occasionally drained debris from the chronic abscess | 6
removed after the follow-up imaging | 6
no drainage was observed | 6