73 years old | 0
male | 0
admitted to the hospital | 0
epigastric pain | -6
nausea | -6
hematemesis | -2
smoker | 0
pacemaker | 0
arteriovenous block | 0
pale skin | 0
blood pressure 155/70 mm Hg | 0
heart rate 85 beats/min | 0
capillary oxygen saturation of 92% | 0
diffusively tender abdomen | 0
distended abdomen | 0
no clear rigidity | 0
hemoglobin 90 mg/dL | 0
white blood count 16×10^9/L | 0
C-reactive protein 122 mg/L | 0
abdominal radiography | 0
soft tissue shadow with lamellar gas | 0
CT scan | 0
thickened stomach wall | 0
gas in intramural venous branches | 0
gas in intrahepatic portal vein branches | 0
gastroscopy | 0
stomach necrosis | 0
urgent surgery | 0
ischemic stomach body | 0
necrotic areas | 0
partial gastrectomy | 0
Roux en esophago-jejunal anastomosis | 0
postoperative course uneventful | 120
discharged | 168
free of symptoms | 8760
unremarkable gastroscopy findings | 8760
pathohistological analysis | 0
ischemic transmural necrosis | 0
edematous and inflamed smaller curvature | 0
no sign of ulcer | 0
no sign of tumor | 0
no sign of mucosal laceration | 0
polymicrobial infection | 0
Klebsiella pneumoniae | 0
Pseudomonas aeruginosa | 0
Bacteroides fragilis | 0