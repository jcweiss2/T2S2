28 years old | 0
male | 0
attended a health center | -24
fatigue | -24
anosmia | -24
dyspnea | -24
SpO2 levels were 55% | -24
nasal cannula oxygen therapy | -24
SpO2 levels improved to 75% | -24
hospitalized | 0
evaluated at an emergency department | 0
chest radiography | 0
bilateral lung infiltrates | 0
RT-PCR swab tested positive for SARS-CoV-2 infection | 0
admitted in a COVID-19 infirmary unit | 0
non-invasive ventilation support | 0
intubation | 12
invasive mechanical ventilation | 12
ventral decubitus positioning | 12
Escherichia coli detected on sputum culture | 48
methicillin-sensitive Staphylococcus aureus detected on sputum culture | 48
superinfection | 48
amoxicillin prescribed | 48
blood culture revealed methicillin-resistant Staphylococcus aureus | 48
methicillin-resistant Staphylococcus aureus dismissed | 48
steady clinical improvement | 72
extubated | 120
discharged | 168
retrosternal thoracalgia | 168
thoracalgia irradiating to the left upper limb | 168
abduction and external rotation limited due to pain | 168
soft tissue swelling of the shoulder and arm | 168
fever | 168
increased levels of C-reactive protein | 168
admitted for further investigation and treatment planning | 168
gentamicin prescribed | 168
gentamicin administered | 168
thoracic CT with intravenous contrast administration | 216
scapulohumeral synovitis | 216
intra-muscular collections | 216
glenohumeral joint fluid | 216
bilateral shoulder magnetic resonance imaging (MRI) with intravenous contrast administration | 240
infraspinatus fossa collections | 240
subscapular fossa collections | 240
capsular thickening | 240
increased signal intensity post-gadolinium administration | 240
septic arthritis | 240
rotator cuff collections | 240
myonecrosis | 240
aspiration of the infraspinatus fossa collection | 252
seropurulent fluid sent for analysis | 252
drainage catheter left on the left infraspinatus collection | 252
drainage catheter removed | 264
physical rehabilitation exercises | 264
improvement of left shoulder range of motion | 288
transferred to another hospital | 288
indication to continue physical therapy and rehabilitation exercises | 288