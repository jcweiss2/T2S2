57 years old | 0 | 0 
male | 0 | 0 
lepromatous leprosy | -720 | -720 
skin biopsy | -720 | -720 
treatment with rifampicin/clofazimine/dapsone | -720 | 0 
admitted to the hospital | 0 | 0 
abdominal distension | 0 | 0 
constipation | 0 | 0 
vomiting | 0 | 0 
10-kg weight loss | -720 | 0 
peripheral lymphadenopathy | 0 | 0 
distended abdomen | 0 | 0 
positive shifting dullness | 0 | 0 
computed tomography scan of abdomen | 0 | 0 
mural thickening of terminal ileum | 0 | 0 
enlarged mesenteric lymph nodes | 0 | 0 
mesenteric fat stranding | 0 | 0 
intra-abdominal free fluid | 0 | 0 
abdominal paracentesis | 0 | 0 
atypically large lymphocytes | 0 | 0 
flow cytometry | 0 | 0 
abnormal CD4/CD8 double-negative T-cell population | 0 | 0 
cervical lymph node biopsy | 0 | 0 
high-grade peripheral T-cell lymphoma | 0 | 0 
bone marrow examination | 0 | 0 
no involvement of T-cell NHL | 0 | 0 
stage IV lymphoma | 0 | 0 
dexamethasone | 0 | 0 
tumor-lysis syndrome precautions | 0 | 0 
deteriorated clinically | 24 | 24 
transfer to medical ICU | 24 | 24 
severe sepsis | 24 | 24 
antibiotics | 24 | 168 
antifungals | 24 | 168 
ICU care | 24 | 168 
recovered | 168 | 168 
transferred to national cancer center | 168 | 168 
EPOCH chemotherapy protocol | 168 | 1008 
CNS prophylaxis | 168 | 1008 
intrathecal methotrexate | 168 | 1008 
complete metabolic remission | 672 | 672 
febrile neutropenia episodes | 336 | 1008 
recurrent bacteremia | 336 | 1008 
generalized weakness | 336 | 336 
no sensory changes | 336 | 336 
no clear fatigability | 336 | 336 
decreased power in proximal and distal muscles | 336 | 336 
normal distal latencies | 336 | 336 
normal compound muscle action potential | 336 | 336 
normal conduction velocities | 336 | 336 
normal F waves | 336 | 336 
normal sensory nerve studies | 336 | 336 
needle electromyogram | 336 | 336 
poor recruitment effects | 336 | 336 
repetitive nerve stimulation | 336 | 336 
significant incremental response | 336 | 336 
presynaptic neuromuscular junction disorder | 336 | 336 
LEMS | 336 | 336 
intravenous immunoglobulins | 336 | 408 
improvement of motor function | 408 | 408 
ambulate | 408 | 408 
consolidation by autologous bone marrow transplant | 1008 | 1008 
recurrent bacteremia and sepsis | 1008 | 1008 
multiorgan failure | 1008 | 1008 
passed away | 1512 | 1512 
remission status | 1008 | 1512