18 years old| 0
male | 0
admitted to the hospital | 0
fever | -72
rash | -72
acne |  -672
minocycline |  -672
increased WBC count | 0
eosinophilia| 0
systemic involvement| 0
diffuse erythematous or maculopapular eruption| 0
pruritis | 0
DRESS syndrome | 0
fever persisted | 0
rash persisted | 0
discharged | 24
Separate conjunctive phrases into its component events and assign them the same timestamp (for example, the separation of 'fever and rash' into 2 events: 'fever' and 'rash')  If the event has duration, assign the event time as the start of the time interval. Attempt to use the text span without modifications except 'history of' where applicable. Include all patient events, even if they appear in the discussion; do not omit any events; include termination/discontinuation events; include the pertinent negative findings, like 'no shortness of breath' and 'denies chest pain'.  Show the events and timestamps in rows, each row has two columns: one column for the event, the other column for the timestamp.  The time is a numeric value in hour unit. The two columns are separated by a pipe '|' as a bar-separated file. Skip the title of the table. Reply with the table only. Create a table from the following case:
<|eot_id|><|start_header_id|>user<|end_header_id|>
<|eot_id|><|start_header_id|>assistant<|end_header_id|>
30 years old | 0
paralysis of both legs | -336
skin getting darker (lower limbs) | -336
pain (scrotum and penis) | -336
darkening of the scrotum and penis | -336
waist strained when playing a kite | -345
weakness | -345
loss of urge to urinate | -345
loss of urge to defecate | -345
bedwetting | -336
no haematuria | 0
no cloudy urine |EOL
7. waist strained when playing kite | -337
8. weakness | -336 (1 hour after incident)
9. loss of urge to urinate | -336
10. loss of urge to defecate | -336
