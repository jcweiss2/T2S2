30 years old | 0
    female | 0
    severe pain in abdomen | -192
    fever | -192
    giddiness | -192
    full-term normal vaginal delivery | -192
    admitted to a private nursing home | -192
    gaping of episiotomy wound | -192
    resuturing | -192
    evaluated for fever | -192
    platelet count of 50,000/cumm | -192
    worsening fever | -168
    breathlessness | -168
    hypotensive | -168
    conservatively managed | -168
    shifted to our hospital | -168
    admitted to our hospital | 0
    severely tachypneic | 0
    severe hypotension | 0
    inotropic supports | 0
    intubated | 0
    mechanically ventilated | 0
    platelet count of 40,000/cumm | 0
    deranged liver function tests | 0
    creatinine of 4.1 mg/dl | 0
    coagulopathy | 0
    international normalized ratio of 4.3 | 0
    chest X-ray bilateral infiltrates | 0
    arterial blood gas PaO2/FiO2 <100 | 0
    severe ARDS | 0
    ultrasonography abdomen normal | 0
    ultrasonography pelvis normal | 0
    two-dimensional echocardiography normal | 0
    provisional diagnosis acute febrile illness | 0
    severe sepsis | 0
    septic shock | 0
    evaluation for etiology | 0
    PCR leptospira negative | 0
    dengue IgM negative | 0
    malaria smear negative | 0
    IgM antibodies hantavirus positive | 0
    falling platelet count | 240
    coagulopathy needing blood component transfusion | 240
    severe ARDS needing lung protective ventilation | 240
    renal dysfunction | 240
    renal replacement therapy | 240
    septic shock needing broad-spectrum antibiotics | 240
    inotropic support | 240
    progressively worsening chest X-ray | 240
    alveolar hemorrhage | 240
    worsening lung function | 240
    hemodynamic support | 240
    broad-spectrum antibiotics | 240
    ribavirin started | 240
    worsening lung function | 240
    expired | 240
    multiorgan dysfunction | 240
    
    
    