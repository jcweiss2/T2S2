65 years old | 0
female | 0
diabetes mellitus | 0
bilateral cataracts | 0
uveitis | -8760
palpitations | 0
dizziness | 0
sinoatrial block | 0
right bundle branch block | 0
pacemaker implantation | 0
dual-chamber pacemaker implantation | 0
progressive dyspnoea | 144
minimal activity | 144
diuretics | 144
angiotensin receptor antagonists | 144
abnormal liver function | 144
elevated level of brain natriuretic peptide | 144
heart failure with preserved ejection fraction | 144
leg oedema | 744
complete atrioventricular block | 744
atrial-paced and ventricular-paced rhythm | 744
device interrogation | 744
worsening heart failure | 816
hospitalization | 816
junctional escape rhythm | 816
complete atrioventricular block with atrial and ventricular pacing failure | 816
biventricular systolic dysfunction | 816
giant right ventricular thrombus formation | 816
pacemaker re-programming | 816
unsuccessful | 816
cardiac arrest | 840
temporary pacing electrode | 840
inserted into the coronary sinus | 840
transferred to hospital | 864
urgent thrombectomy | 888
endomyocardial biopsy | 888
cardiac sarcoidosis | 888
infiltrative inflammatory cells | 888
epithelioid cell granulomas | 888
multinucleated giant cells | 888
steroid pulse therapy | 888
corticosteroids | 888
maintenance therapy | 888
improved left ventricular ejection fraction | 888
intravenous catecholamine support | 888
withdrawn | 888
discharged | 888
guideline-directed medical therapy | 888
heart failure with reduced ejection fraction | 888
bisoprolol | 888
enalapril | 888
spironolactone | 888
empagliflozin | 888
anti-coagulation therapy | 888
warfarin | 888
prednisolone | 888
positron emission tomography | 9360
no uptake of 18F-fluorodeoxyglucose | 9360
in the myocardium | 9360
sustained ventricular tachycardia | 10416
pacemaker upgrading | 10416
implantable cardioverter defibrillator | 10416
recurrent sustained ventricular tachycardia | 10944
refractory ventricular electrical storms | 10944
mechanical ventilation | 10944
deep sedation | 10944
intravenous administration | 10944
amiodarone | 10944
lidocaine | 10944
severe biventricular pump failure | 10944
fever | 10944
arterial hypotension | 10944
leukocytosis | 10944
bacteraemia | 10944
methicillin-resistant Staphylococcus epidermidis | 10944
Candida albicans | 10944
sepsis | 10944
death | 11136
multiple organ failure | 11136
severe pump failure | 11136
sepsis | 11136
autopsy | 11136
diffuse fibrotic tissues | 11136
both ventricles | 11136
myocardium | 11136
right ventricle | 11136
substantially replaced | 11136
fibrotic tissues | 11136
without inflammatory cell infiltration | 11136
significant fibrotic changes | 11136
anatomical sinus node | 11136
right atrium | 11136