79 years old | 0
    white | 0
    man | 0
    laparoscopic converted to open cholecystectomy | -504
    gangrenous perforated gallbladder | -504
    retrograde fundus-down approach | -504
    inability to obtain the critical view | -504
    tubular structure (thought to be a duct of Luschka) | -504
    ligated tubular structure | -504
    cystic artery ligated | -504
    cystic duct ligated | -504
    single drain placed | -504
    procedure completed | -504
    persistent high-output bilious drainage | -504
    discharged on postoperative Day 6 | -504
    drain in place | -504
    returned to outside facility | -216
    jaundice | -216
    weakness | -216
    fatigue | -216
    pain | -216
    CT scan of abdomen | -216
    nuclear cholescintigraphy scan | -216
    confirmed biliary leak | -216
    free intra-abdominal fluid | -216
    biliary peritonitis | -216
    transferred to critical care unit | -216
    placed on broad spectrum antibiotics | -216
    treated for atrial fibrillation with rapid ventricular response | -216
    bilirubin level of 17 mg/dl | -216
    profound protein-calorie malnutrition | -216
    albumin of 1.9 gm/dl | -216
    percutaneous cholangiogram performed | -216
    hilar ligation of hepatic duct | -216
    inability to pass wire or catheter distally | -216
    right posterior percutaneous cholangiogram catheter placed | -216
    right anterior percutaneous cholangiogram catheter placed | -216
    definitive biliary diversion | -216
    managed with high calorie high protein enteral nutrition | -216
    nasogastric Dobhoff tube | -216
    tolerated appropriate oral intake | -168
    scheduled for follow-up in 2 weeks | -168
    improved substantially | 0
    repeat CT scan | 0
    appropriate drainage of all abdominal fluid collections | 0
    bilirubin improved to 1.2 mg/dl | 0
    albumin of 3.1 gm/dl | 0
    prealbumin of 17.3 gm/dl | 0
    scheduled for definitive biliary reconstruction | 0
    during operation | 0
    porta dissected | 0
    common hepatic artery identified and preserved | 0
    proper hepatic artery identified and preserved | 0
    unable to palpate percutaneous biliary catheters | 0
    high placement above the hilum | 0
    multiple clips | 0
    transected CBD distally | 0
    removed numerous clips | 0
    noted bile drainage | 0
    unable to identify cholangiogram catheter | 0
    identified second tubular structure | 0
    transected second tubular structure | 0
    identified second extrahepatic bile duct | 0
    anterior percutaneous catheter identified proximally | 0
    on-table cholangiogram with fluoroscopy | 0
    two separate extrahepatic biliary systems | 0
    draining right lobe | 0
    draining left lobe | 0
    both distal ducts ligated | 0
    prevent spillage | 0
    Roux limb of jejunum created | 0
    anastomosed retrocolic | 0
    two separate hepatic ducts at hilum | 0
    drain placed | 0
    no evidence of bile leakage | 0
    discharged on postoperative Day 6 | 144
    normal hepatic function | 144
    normal bilirubin | 144
    no further complications | 144
    follow-up cholangiogram | 144
    normal intrahepatic ducts | 144
    no evidence of stricture | 144
    no evidence of leak | 144
    successful repair | 144
    cholangiogram catheters removed | 144
    discharged from clinic | 144