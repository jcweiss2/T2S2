54 years old | 0
male | 0
admitted to the hospital | 0
discomfort in the hepatic region | -672
diagnosed with cirrhosis, hypersplenism and portal hypertension | -672
multiple nodules at S4 and S5 in the liver | -672
hepatocellular carcinoma | -672
interventional surgery | -672
multiple early stage lung tumors | -672
treated with thrombopoietin | -24
treated with cryoprecipitate | -24
white blood cell count, 6.07×10^9/L | 0
hemoglobin, 124 g/L | 0
platelet count, 297×10^9/L | 0
total bilirubin, 29.3 µmol/L | 0
direct bilirubin, 11.8 µmol/L | 0
total serum protein, 59.5 g/L | 0
albumin, 32.7 g/L | 0
prothrombin time, 15.40 s | 0
partial thromboplastin activation time, 33.90 s | 0
carcinoembryonic antigen (CEA), 4.89 ng/mL | 0
carbohydrate antigen 199 (CA19-9), 269.10 U/mL | 0
carbohydrate antigen 724 (CA72-4), 7.19 U/mL | 0
cytokeratin 19 fragment (CYFRA21-1), 6.30 ng/mL | 0
hepatitis B virus DNA <5.00E+02 IU/mL | 0
Child-Pugh classification grade B | 0
Child-Pugh score of 8 points | 0
lung cancer | 0
clinical T1 N0 M0 stage IA | 0
left superior segmentectomy | 0
right superior wedge resection | 0
adenocarcinomas | 0
invasive adenocarcinoma on the left | 0
well-differentiated adenocarcinoma on the right | 0
negative margins | 0
no evidence of metastasis in the lymph nodes | 0
left thoracic duct effused 1,200 mL sanguineous drainage | 6
increased heart rate | 6
hypotension | 6
plasma transfused | 6
red blood cells transfused | 6
platelets transfused | 6
cryoprecipitate transfused | 6
atrial fibrillation | 24
dyspnea | 24
acute respiratory distress syndrome (ARDS) | 24
diffused alveolar hemorrhage (DAH) | 24
stale blood clots in the phlegm | 24
white blood cell count, 13.2×10^9/L | 48
hemoglobin, 66 g/L | 48
platelet count, 123×10^9/L | 48
prothrombin time, 15.80 s | 48
partial thromboplastin activation time, 35.40 s | 48
fibrinogen, 1.45 g/L | 48
total bilirubin, 33.7 µmol/L | 48
direct bilirubin, 15.3 µmol/L | 48
total serum protein, 50.1 g/L | 48
albumin, 33.3 g/L | 48
patchy infiltrates scattered throughout both lungs | 96
noninvasive ventilator-assisted ventilation | 96
oxygenation improved | 96
partial pressure of oxygen improved | 96
sanguineous drainage diminished | 168
Klebsiella pneumoniae | 240
Candida albicans | 240
meropenem administered | 240
voriconazole administered | 240
septicemia resolved | 288
voriconazole per os | 288
discharged from the hospital | 384
no evidence of recurrent disease | 744