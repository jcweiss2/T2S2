20 years old | 0
male | 0
Caucasian | 0
admitted to the hospital | 0
septic shock | 0
febrile | 0
tachycardia | 0
tachypnea | 0
hypotensive | 0
norepinephrine | 0
neutropenia | 0
thrombocytopenia | 0
hypokalemia | 0
recto-cecal abscess | -504
appendectomy | -504
febrile neutropenia | -504
meropenem | -504
vancomycin | -504
micafungin | -504
amikacin | -360
discontinued amikacin | -360
right arm cellulitis | -288
abscess | -288
ESBL and CRE Escherichia coli | -288
colistin | -288
loading dose of colistin | -288
maintenance dose of colistin | -288
meropenem | -288
vancomycin | -288
amphotericin B | -288
tigecycline | -168
severe reaction | -168
hypotension | -168
shortness of breath | -168
hypoxia | -168
tachycardia | -168
tachypnea | -168
flushed face | -168
leukocytosis | -168
acute kidney injury | -168
adrenaline | -168
chlorpheniramine | -168
hydrocortisone | -168
resolved leukocytosis | -144
resolved renal function | -144
discontinued norepinephrine | -144
second severe reaction | -120
hypotensive | -120
shortness of breath | -120
hypoxia | -120
flushed face | -120
generalized erythema | -120
leukocytosis | -120
acute kidney injury | -120
increased total bilirubin level | -120
discontinued colistin | -120
meropenem | -120
tigacycline | -120
amikacin | -120
resolved norepinephrine | -96
resolved laboratory results | -96
transferred to the floor | -48
piperacillin/tazobactam | -48
tigecycline | -48
amikacin | -48
ventricular fibrillation | 0
died | 0