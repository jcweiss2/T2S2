56 years old | 0
male | 0
alcohol abuse | 0
40 pack-year smoking history | 0
scrotal pain | -96
myalgia | -96
inability to walk | -96
fulminant necrosis of the scrotum | 0
necrosis of the dorsum and heels of both feet | 0
necrosis of the left middle finger | 0
intravenous benzylpenicillin | 0
intravenous flucloxacillin | 0
transfer to the regional center | 0
diagnosis of scrotal FG with concurrent multifocal NF | 0
intravenous clindamycin | 0
intravenous meropenem | 0
intravenous vancomycin | 0
surgical exploration and debridement | 0
scrotal debridement | 0
bilateral orchiectomy | 0
debridement of necrotic tissue from both feet and left middle finger | 0
admission to the intensive care unit (ICU) | 0
intravenous vasopressor support (noradrenaline) | 0
pathological analysis of scrotal tissue | 0
polymicrobial growth including Streptococcus intermedius, Escherichia coli, Klebsiella oxytoca, and Staphylococcus aureus | 0
histological examination of limb tissue | 0
transfer to a metropolitan tertiary institution | 24
further 6 days in ICU | 24
noradrenaline vasopressor support | 24
scrotal debridement | 48
left medial thigh exploration | 48
insertion of bilateral middle ear ventilation tubes | 48
scrotal wound reexploration and closure | 96
further debridement of limb wounds | 96
further debridement and received split skin grafts from the left thigh to bilateral heel wounds | 192
discharged from the metropolitan center | 720
discharged to a regional rehabilitation facility | 720
oral ciprofloxacin | 720
oral amoxicillin/clavulanate | 720
lifelong testosterone replacement therapy | 720
discharged home | 1200
full recovery | 1200
return to fruit picking | 2160