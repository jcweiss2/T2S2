47 years old| 0
    man | 0
    diabetes mellitus | 0
    presented to the emergency department | 0
    abrupt-onset severe headache | 0
    right-sided blindness | 0
    headache at occiput | -24
    right-sided blindness | 0
    COVID-19 infection | -480
    RT-PCR test | -480
    pulmonary symptoms | -480
    intensive care unit admission | -480
    no COVID-19 vaccine | -480
    drowsy | 0
    oriented to person | 0
    oriented to place | 0
    oriented to time | 0
    blood pressure 170/100 mmHg | 0
    dysarthric speech | 0
    right homonymous hemianopia | 0
    alexia without agraphia | 0
    no petechiae | 0
    no purpura | 0
    brain computed tomography | 0
    intraparenchymal hemorrhage | 0
    edema | 0
    left occipital lobe | 0
    string sign | 0
    left transverse sinus | 0
    diagnosis of hemorrhagic venous infarction | 0
    transverse sinus thrombosis | 0
    D-dimer level 1030 | 0
    platelet count 20,000 | 0
    platelet count 150,000 | -480
    peripheral blood smear | 0
    giant platelets | 0
    no schistocytes | 0
    COVID-19 RT-PCR | 0
    HCV negative | 0
    HBV negative | 0
    HIV negative | 0
    received 10 units of platelets | 0
    dexamethasone 8 mg three times daily | 0
    platelet count 49,000 | 0
    bone marrow aspiration | 0
    bone marrow biopsy | 0
    hypolobulated megakaryocytes | 0
    IVIG 20 g for 5 days | 0
    thrombocytopenia responded | 0
    platelet count 115,000 | 0
    diagnosis of ITP | 0
    discharged | 192
    prednisolone 25 mg twice daily | 192
    platelet count 140,000 | 672
    neurological symptoms improved | 672
    homonymous hemianopia improved | 672
    difficulties in reading | 672
    cerebral venous sinus thrombosis | 0
    immune thrombocytopenic purpura | 0
    SARS-CoV-2 infection | -480
    systemic inflammation | 0
    cytokine storm | 0
    direct immune-mediated post-infection mechanism | 0
    virus-induced angiitis | 0
    hemophagocytic lymphohistiocytosis ruled out | 0
    thrombotic thrombocytopenic purpura ruled out | 0
    sepsis ruled out | 0
    heparin-induced thrombocytopenia ruled out | 0
    drug-induced thrombocytopenia ruled out | 0
    COVID-19 vaccine mechanism considered | 0
    immune-mediated thrombocytopenia | 0
    anti-platelet 4-factor antibody considered | 0
