33 years old| 0
male | 0
renal transplant recipient | 0
parent-to-child kidney transplantation | -4320
end-stage renal disease | -4320
methylprednisolone | -4320
tacrolimus | -4320
mycophenolate mofetil | -4320
severe upper abdominal pain | -72
upper abdominal pain radiating towards back | -72
admitted to local hospital | -72
abdominal computed tomography | -72
ultrasonography | -72
analgesic treatment | -72
aspartate aminotransferase increased | -72
alanine aminotransferase increased | -72
referred to hospital | 0
nausea | 0
upper abdominal pain | 0
acute abdominal pain | 0
liver damage | 0
flurbiprofen tapes | 0
intravenous magnesium isoglycyrrhizinate | 0
intravenous cefoperazone sodium | 0
sulbactam sodium | 0
septic shock | 0
multiple organ dysfunction syndrome | 0
liver dysfunction | 0
acute kidney injury | 0
transferred to intensive care unit | 48
end-stage renal failure | -25920
lethargic | 0
heart rate 136 beats/min | 0
respiratory rate 23 breaths/min | 0
blood pressure 83/42 mmHg | 0
body temperature 36.8 °C | 0
abdominal tenderness | 0
high ALT | 0
high AST | 0
high alkaline phosphatase | 0
high gamma-glutamyltransferase | 0
high C-reactive protein | 0
high procalcitonin | 0
high creatinine | 0
prolonged activated partial thromboplastin time | 0
prolonged thrombin time | 0
low fibrinogen | 0
negative hepatitis A virus serology | 0
negative hepatitis B virus serology | 0
negative hepatitis C virus serology | 0
negative human immunodeficiency virus serology | 0
negative treponema pallidum serology | 0
hepatitis B surface antibodies positive | 0
hepatitis B core antibodies positive | 0
absent IgM toxoplasma antibodies | 0
absent IgM rubella virus antibodies | 0
absent IgM cytomegalovirus antibodies | 0
absent IgM herpes simplex virus 2 antibodies | 0
negative blood culture | 0
negative Epstein-Barr virus PCR | 0
normal pancreas | 0
normal spleen | 0
normal gallbladder | 0
normal common bile duct | 0
no ascites | 0
no abnormal fluid collection | 0
no focal liver lesions | 0
no intestinal obstruction | 0
no intestinal perforation | 0
no mesenteric artery thrombosis | 0
normal chest X-ray | 0
normal electrocardiogram | 0
next-generation sequencing | 0
real-time PCR | 0
IgG assays | 0
VZV IgG-negative | 0
NGS VZV positive | 0
real-time PCR VZV positive | 0
visceral disseminated VZV infection | 0
antiviral therapy | 0
intravenous acyclovir | 0
intravenous meropenem | 0
linezolid | 0
caspofungin | 0
noradrenaline | 0
terlipressin | 0
intravenous sodium bicarbonate | 0
acute liver failure | 0
disseminated intravascular coagulation | 0
acute respiratory failure | 0
acute renal injury | 0
death | 16
