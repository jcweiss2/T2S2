29 years old | 0
    female | 0
    born at 38 weeks gestation | 0
    cesarean section | 0
    failed induction | 0
    referral to tertiary neonatal ICU | 20
    suspected duodenal atresia | 20
    weight 2400 g | 0
    length 55 cm | 0
    head circumference 35 cm | 0
    stable condition | 0
    normal vital signs | 0
    afebrile | 0
    heart rate 130/minute | 0
    respiratory rate 55/minute | 0
    oxygen saturation 95-96% | 0
    normal blood investigations | 0
    normal platelets | 0
    left upper limb deformity | 0
    radial flexion | 0
    partial syndactyly | 0
    complete radial aplasia | 0
    abnormal wrist flexion | 0
    normal skeletal survey | 0
    soft abdomen | 0
    passing stool | 0
    nil per os | 0
    persistent dilated stomach | 0
    residual greenish gastric aspirate | 0
    suspicion of duodenal web | 0
    laparotomy | 48
    annular pancreas | 48
    grossly dilated stomach | 48
    grossly dilated duodenum | 48
    normal liver echogenicity | 0
    patent hepatic veins | 0
    normal gallbladder | 0
    normal kidney size | 0
    preserved cortical medullary differentiation | 0
    no ascites | 0
    spleen not visualized | 0
    repeated spleen not visualized | 0
    Howell-Jolly bodies | 0
    suspicion of asplenia syndrome | 0
    normal liver location | 0
    spleen not visualized on scan | 0
    levocardia | 0
    complex congenital heart disease | 0
    single atrium | 0
    large pyramidal appendages | 0
    single ventricle | 0
    right ventricle morphology | 0
    good ventricular function | 0
    single AV valve | 0
    dextro-transposition of great arteries | 0
    moderate pulmonary stenosis | 0
    small PDA | 0
    normal head ultrasound | 0
    choroid plexus cyst | 0
    persistent late-onset staphylococcus sepsis | 504
    prolonged antibiotic treatment | 504
    improved condition | 0
    full feeding | 0
    extubated to nCPAP | 0
    oxygen requirement 30% | 0
    prophylactic antibiotics | 0
    anti-heart failure medications | 0
    follow-up with cardiology | 0
    follow-up with orthopedics | 0
    follow-up with plastic surgery | 0
    accepted for higher-level care | 0
    diagnosed asplenia syndrome | 0
    right isomerism | 0
    congenital complex heart disease | 0
    annular pancreas | 0
    left upper limb radial aplasia | 0
    partial syndactyly | 0
    Howell-Jolly bodies confirmation | 0
    immune-compromised | 0
    increased sepsis risk | 0
    normal intestinal rotation | 0
    unavailability of corrective surgery | 0
    discharged for higher-level care | 0
