53 years old | 0
female | 0
Caucasian | 0
admitted to the Emergency Department | 0
dyspnoea | 0
chest tightness | 0
dizziness | 0
palpitations | 0
nausea | 0
vomiting | 0
oral glucose tolerance test | -2
hypoglycaemia | -2
impaired fasting glucose | -672
borderline haemoglobin A1c | -672
hypertension | -672
dyslipidaemia | -672
secondary hyperparathyroidism | -672
simvastatin | -672
calcium carbonate/cholecalciferol | -672
metoprolol | -672
losartan | -672
pale skin | 0
cool extremities | 0
weak radial pulses | 0
prolonged capillary refilling time | 0
respiratory rate 40 breaths/min | 0
oxygen saturation 80% | 0
heart rate 114 b.p.m. | 0
blood pressure 111/75 mmHg | 0
bilateral inspiratory crackles | 0
hypoxaemia | 0
metabolic acidosis | 0
hyperglycaemia | 0
elevated cardiac troponin T | 0
leucocytosis | 0
acute kidney injury | 0
sinus tachycardia | 0
hypokinesia in the mid-inferior and apical segments | 0
left ventricular ejection fraction 15% | 0
pulmonary oedema | 0
interstitial oedema | 0
cardiogenic shock | 0
norepinephrine | 12
levosimendan | 12
insulin therapy | 12
antibiotic therapy | 12
fever | 12
lactate increased | 12
urinary output decreased | 12
heart rate 122 b.p.m. | 12
systolic blood pressure 85 mmHg | 12
cardiac index 2.1 L/min/m2 | 12
mean pulmonary artery pressure 23 mmHg | 12
improved cardiac index | 24
improved left ventricular ejection fraction | 24
weaned from norepinephrine | 24
discharged home | 168
readmitted | 408
elevated metanephrine | 408
elevated normetanephrine | 408
elevated plasma methoxytyramine | 408
elevated chromogranin A | 408
pharmacological adrenergic blockade | 408
computer tomography | 408
left adrenal phaeochromocytoma | 408
left adrenalectomy | 1440
discharged home | 1536
follow-up visit | 2556
scheduled for follow-up computed tomography and lab testing | 3060