38 years old | 0
male | 0
chondrosarcoma | -504
mild compressive atelectasis | 0
wide local excision | 0
anterior chest wall defect | 0
missing ribs | 0
exposed cardiopulmonary structures | 0
rib cage reconstruction with polypropylene mesh | 0
soft tissue reconstruction with free anterolateral thigh flap | 0
nipple areola complex harvested as free graft | 0
endotracheal tube | 0
noradrenaline 0.05 µg/kg/min | 0
intraoperative hemodynamic instability | 0
vasopressin added | 48
spontaneous breathing trials unsuccessful | 0
weaning from ventilator support unsuccessful | 0
pneumothorax detected | 24
chest tube inserted | 24
normal left ventricular ejection fraction | 0
antibiotics escalated | 48
blood culture negative | 48
afebrile | 48
vacuum dressing applied | 120
polyurethane sponge and film at −125 mm Hg | 120
reduced PEEP requirement | 120
better tolerance of SBT | 120
better tolerance of PSV | 120
extubated | 192
transitioned to high-flow nasal cannula | 192
shifted out of ICU | 240
healthy flap | 240
healthy suture line | 240
healthy NAC graft | 240
discharged with NPWT | 264
satisfactory lung expansion | 264
NPWT stopped | 360
minimal residual paradoxical breathing | 360
no discomfort in breathing | 360
denied SIRS | 0
denied septic shock | 0
denied cardiogenic shock | 0
no obvious infection source | 0
blood cultures negative | 0
afebrile | 0
shock persisted | 0
no tracheostomy needed | 0
no vascular complications in free flap | 0
