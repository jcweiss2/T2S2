66 years old|0
woman|0
hospitalized to the emergency room|0
fever|0
hypotension|0
tachycardia|0
elevated leukocytes|0
elevated CRP|0
acute renal failure|0
elevated creatinine|0
decreased glomerular filtration rate (GFR)|0
leukocyturia|0
proteinuria|0
bacteria in urine|0
horseshoe kidney|0
second-degree urinary retention|0
urosepsis|0
transferred to intensive care unit|0
stent insertion|0
restricted renal function|0
computed tomography (CT) of chest|0
computed tomography (CT) of abdomen|0
computed tomography (CT) of pelvis|0
10.5 × 10 × 11 cm inhomogeneous mass|0
cystic parts adjacent to right ovary|0
contact to right ureter|0
contact to iliac vessels|0
contact to bladder|0
suspicion of infiltration of sacrum|0
gastroscopy|0
colonoscopy|0
diverticulosis|0
18F-FDG-PET|0
no metastases|0
sarcoma suspected|0
neoadjuvant radiotherapy|-168
tumor operation|-168
iliac vascular resection|-168
partial ureteral resection|-168
NET G2|-168
Ki67 10%|-168
CT scan|-168
two liver metastases|-168
refused further treatment|-168
MRI|-168
multiple liver lesions|-168
liver biopsy|-168
metastases of well-differentiated NET G2|-168
Ki67 15%|-168
68Ga-DOTATATE PET|-168
intense somatostatin receptor expression in liver lesions|-168
additional focus close to pancreas|-168
endosonographic ultrasound|-168
pathologic lymph node adjacent to head of pancreas|-168
no tumor of pancreas|-168
cancer of unknown primary NET G2|-168
slight renal impairment|-168
treated with two cycles of 177Lu-DOTATATE|-168
lanreotide every 4 weeks|-168
disease stabilization|-168
progression after PRRT|0
received everolimus|0
disease progression after 2 months|24
liver biopsy|24
NET G3|24
Ki67 34%|24
treated with capecitabine plus temozolomide|24
12 cycles|24
progression|24
cycle of PRRT|24
stabilization of disease|24
progression|168
treated with oxaliplatin and capecitabine|168
significant dose reduction|168
fatigue|168
diarrhea|168
chemotherapy discontinued|168
molecular testing|240
BRCA1 Mutation R691fs*10|240
tumor mutational burden zero|240
microsatellite stability|240
germline analysis confirmed BRCA mutation|240
started Olaparib 200 mg twice daily|240
stable liver metastases|240
upper abdominal pain|240
BRCA1 mutation|240
advanced disease|240
limited treatment options|240
individual medical treatment|240
cycle of PRRT with 225Ac-DOTATATE|240
Olaparib 100 mg twice daily|240
renal insufficiency (GFR 40 mL/min/1.73 qm)|240
treatment well tolerated|240
no relevant toxicity|240
no haematotoxicity|240
no further impairment of renal function|240
abdominal complaints disappeared|240
Olaparib restarted 200 mg twice daily|240
restaging with 68Ga-DOTATATE PET/MRI|240
decrease in liver metastases|240
stable large liver metastasis in left lobe|240
progression of smaller hepatic metastases in right lobe|240
additional TAT in combination with olaparib planned|240
