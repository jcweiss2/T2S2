37 years old | 0
    female | 0
    admitted with body mass index of 67 kg/m² | 0
    back pain | 0
    gastroesophageal reflux disease | 0
    obstructive sleep apnea | 0
    hyperlipidemia |E0
    hypertension | 0
    Da Vinci-assisted laparoscopic one-stage single-anastomosis DS procedure | 0
    terminal ileum identified | 0
    duodeno+ileal anastomosis created | 0
    sleeve gastrectomy done | 0
    staple line oversewn | 0
    duodenum transected 3 cm from pylorus | 0
    duodenal stump oversewn with running absorbable suture | 0
    two-layer hand sewn anastomosis between duodenum and ileum | 0
    anastomosis tested with methylene blue and air | 0
    drain placed in left upper quadrant | 0
    stomach removed | 0
    upper gastrointestinal study (UGI) on postoperative day 2 | -48
    bariatric phase 1 diet started | -48
    diet tolerated well | -48
    discharged on postoperative day 3 | -72
    persistent nausea | -264
    fatigue | -264
    severe abdominal pain | -264
    tachycardic | -264
    anemia | -264
    leukocytosis | -264
    significant distension | -264
    guarding | -264
    UGI negative | -264
    computed tomography of abdomen showing free fluid | -264
    taken to operating room for diagnostic laparoscopy | -264
    hemoperitoneum evacuated | -264
    active bleeding source not identified | -264
    gastroileostomy anastomosis inspected | -264
    no leakage seen with methylene blue test | -264
    attempt to explore duodenal stump unsuccessful | -264
    three large 19F Blake drains placed | -264
    transfused with 2 units PRBCs intra-operatively | -264
    kept intubated | -264
    transferred to ICU | -264
    hypotensive | -288
    unresponsive to fluids | -288
    abdominal drain increased sanguinous output | -288
    frank bile in second drain | -288
    elevated bilirubin | -288
    elevated amylase | -288
    tachycardic | -288
    taken back to OR for exploratory laparotomy | -288
    laparotomy through right subcostal incision | -288
    hemoperitoneum encountered | -288
    packing temporized gastroduodenal artery | -288
    gastroduodenal artery over-sewn | -288
    duodenal stump found with total blowout | -288
    staple line completely undone | -288
    Malecot tube placed in duodenum | -288
    purse-string suture applied | -288
    abdomen closed | -288
    drains placed | -288
    blood loss 2500 cc | -288
    received 5 units PRBCs | -288
    received 4 units fresh frozen plasma | -288
    transferred to ICU | -288
    hemorrhagic fluid collections on CT scan | -288
    atelectasis | -288
    acute thrombosis left internal jugular | -288
    acute thrombosis subclavian veins | -288
    placed on therapeutic Lovenox | -288
    placed on octreotide | -288
    intravenous piperacillin/taxobactam started | -288
    changed to cefazolin | -288
    discharged on postoperative day 17 | -408
    home health care for dressing changes | -408
    total parenteral nutrition | -408
    <|eot_id|>

  37 years old | 0
female | 0
admitted with body mass index of 67 kg/m² | 0
back pain | 0
gastroesophageal reflux disease | 0
obstructive sleep apnea | 0
hyperlipidemia | 0
hypertension | 0
Da Vinci-assisted laparoscopic one-stage single-anastomosis DS procedure | 0
terminal ileum identified | 0
duodeno-ileal anastomosis created | 0
sleeve gastrectomy done | 0
staple line oversewn | 0
duodenum transected 3 cm from pylorus | 0
duodenal stump oversewn with running absorbable suture | 0
two-layer hand sewn anastomosis between duodenum and ileum | 0
anastomosis tested with methylene blue and air | 0
drain placed in left upper quadrant | 0
stomach removed | 0
upper gastrointestinal study (UGI) on postoperative day 2 | -48
bariatric phase 1 diet started | -48
diet tolerated well | -48
discharged on postoperative day 3 | -72
persistent nausea | -264
fatigue | -264
severe abdominal pain | -264
tachycardic | -264
anemia | -264
leukocytosis | -264
significant distension | -264
guarding | -264
UGI negative | -264
computed tomography of abdomen showing free fluid | -264
taken to operating room for diagnostic laparoscopy | -264
hemoperitoneum evacuated | -264
active bleeding source not identified | -264
gastroileostomy anastomosis inspected | -264
no leakage seen with methylene blue test | -264
attempt to explore duodenal stump unsuccessful | -264
three large 19F Blake drains placed | -264
transfused with 2 units PRBCs intra-operatively | -264
kept intubated | -264
transferred to ICU | -264
hypotensive | -288
unresponsive to fluids | -288
abdominal drain increased sanguinous output | -288
frank bile in second drain | -288
elevated bilirubin | -288
elevated amylase | -288
tachycardic | -288
taken back to OR for exploratory laparotomy | -288
laparotomy through right subcostal incision | -288
hemoperitoneum encountered | -288
packing temporized gastroduodenal artery | -288
gastroduodenal artery over-sewn | -288
duodenal stump found with total blowout | -288
staple line completely undone | -288
Malecot tube placed in duodenum | -288
purse-string suture applied | -288
abdomen closed | -288
drains placed | -288
blood loss 2500 cc | -288
received 5 units PRBCs | -288
received 4 units fresh frozen plasma | -288
transferred to ICU | -288
hemorrhagic fluid collections on CT scan | -288
atelectasis | -288
acute thrombosis left internal jugular | -288
acute thrombosis subclavian veins | -288
placed on therapeutic Lovenox | -288
placed on octreotide | -288
intravenous piperacillin/taxobactam started | -288
changed to cefazolin | -288
discharged on postoperative day 17 | -408
home health care for dressing changes | -408
total parenteral nutrition | -408