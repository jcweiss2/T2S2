53 years old | 0
female | 0
blurred vision | -672
retinal ischemia | -672
cotton wool spots | -672
macular edema | -672
hypertensive retinopathy | -672
monoclonal protein | -672
immunoglobulin G (IgG) kappa type | -672
negative hypercoagulable panel | -672
normal blood cell counts | -672
elevated erythrocyte sedimentation rate | -672
elevated lactate dehydrogenase | -672
slightly elevated creatinine | -672
total immunoglobulin G | -672
abnormal free light chains (FLC) ratio | -672
high free kappa | -672
no monoclonal protein in 24-hour urine collection | -672
no significant proteinuria | -672
skeletal survey showed no lytic lesions | -672
bone marrow aspiration and biopsy showed 10%–15% plasma cells | -672
smoldering myeloma | -672
plasma cell directed therapy | -672
triple therapy with bortezomib, lenalidomide, and dexamethasone | -168
acute renal failure | -168
rise in Creatinine from 1.4 to 6.9 mg/dL | -168
urinalysis showed 1+ protein | -168
greater than five red blood cells per high power field | -168
no casts | -168
serum albumin was 3.1 g/dL | -168
hepatitis serologies were negative | -168
renal ultrasound showed normal-sized kidneys | -168
no evidence of obstruction | -168
renal biopsy | -168
endothelial swelling | -168
intimal edema | -168
concentric fibroplasia | -168
entrapped red blood cells | -168
complete or near-complete luminal obliteration | -168
no definite thrombi | -168
no fibrinoid necrosis | -168
Congo Red stain for amyloid was negative | -168
immunofluorescence showed no light chain restriction | -168
electron microscopy confirmed the absence of amyloid fibrils | -168
evidence of endothelial damage and ischemia | -168
acute tubular injury | -168
no crystals | -168
no abnormal lysosomes | -168
diagnosis of acute thrombotic microangiopathy | -168
Bortezomib was discontinued | -168
no recovery of renal function | -168
progressive decline of vision | -168
no response to intravitreal anti-VEGF | -168
partial response to steroids | -168
recurrent pericardial effusions | -2160
congestive heart failure | -2160
ejection fraction of 25% | -2160
severe left ventricular systolic dysfunction | -2160
moderate pulmonary hypertension | -2160
pulmonary hypertension detected at an echocardiogram | -2160
normal ejection fraction | -2160
primary pulmonary hypertension | -2160
cardiac arrest | -2160
resuscitated | -2160
broad antibiotic therapy | -2160
no clear infection source | -2160
echocardiogram showed moderate pericardial effusion | -2160
enlarged right atrium and right ventricle | -2160
tricuspid regurgitation | -2160
no evidence of tamponade | -2160
pulmonary artery systolic pressure (PASP) was very high | -2160
left ventricular ejection fraction was estimated at 60%–65% | -2160
pericardiocentesis | -2160
325 mL of serous fluid were drained | -2160
cytopathology and fluid cultures were negative | -2160
hematology-oncology was consulted | -2160
serum protein electrophoresis showed a 0.66 g/dL monoclonal band | -2160
IgG was 1226 mg/dL | -2160
serum kappa FLC was 340.8 mg/L | -2160
kappa/lambda FLC ratio of 16.15 | -2160
skeletal survey showed no lytic lesions | -2160
abdominal fat pad biopsy was negative for amyloid | -2160
rheumatology was consulted | -2160
low C3 levels | -2160
normal C4 | -2160
Complement Factor I was normal | -2160
Factor H (B1H) levels were normal | -2160
ADAMTS13 activity was 17% | -2160
ADAMTS13 inhibitor screen was negative | -2160
antiphospholipid antibody panel was negative | -2160
plasma VEGF and anti-myelin associated glycoprotein antibodies were ordered | -2160
multiple episodes of lactic acidosis | -2160
repeated intubations | -2160
severe right heart failure | -2160
treprostinil | -2160
cardiac arrest refractory to resuscitative efforts | -2160
partial autopsy | -2160
ulcer with fat layer exposure on the dorsal aspect of the left foot | -2160
bilateral serous pleural effusions | -2160
pericardial sac contained 200 mL of serous fluid | -2160
heart weighted 440 g | -2160
concentric left ventricular hypertrophy | -2160
right ventricle was dilated | -2160
lungs were congested | -2160
spleen weighted 100 g | -2160
multiple subcapsular wedge-shaped infarcts | -2160
no enlarged lymph nodes | -2160
kidneys were bilaterally atrophic | -2160
liver weighted 1330 g | -2160
nutmeg appearance | -2160
severe renal interstitial fibrosis | -2160
concentric fibrointimal thickening | -2160
endothelial damage and ischemia | -2160
tubules showed intracytoplasmic vacuoles | -2160
loss of microvilli | -2160
no crystals | -2160
no abnormal lysosomes | -2160
myocyte hypertrophy | -2160
minimal fibrosis | -2160
no evidence of amyloid deposition | -2160
centrolobular congestion and necrosis | -2160
right-sided heart failure | -2160
prominent cardiomegaly | -2160
right ventricular hypertrophy | -2160
severe pulmonary microvascular obliterative changes | -2160
death | 0