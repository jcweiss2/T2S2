24 years old | 0
primigravida | 0
37 weeks of gestation | 0
admitted to the hospital | 0
high grade fever | -72
decreased urine output | -72
yellowish discolouration | -72
altered sensorium | -72
disoriented | 0
febrile | 0
icteric | 0
sub-conjunctival haemorrhages | 0
fine basal crepitations | 0
receiving intravenous artesunate | -72
receiving ceftriaxone | -72
receiving doxycycline | -72
anaemia | 0
jaundice | 0
deranged liver function | 0
coagulopathy | 0
thrombocytopenia | 0
increased total leucocyte count | 0
elevated blood urea nitrogen | 0
elevated serum creatinine | 0
singleton pregnancy | 0
adequate liquor | 0
umbilical artery systolic-diastolic ratio of 2:1 | 0
mild hepato-splenomegaly | 0
non-reassuring fetal heart rate | 1
aspiration prophylaxis | 1
high-risk consent | 1
rapid sequence intubation | 1
cricoid pressure | 1
thiopental | 1
succinylcholine | 1
right internal jugular vein cannulation | 1
left radial artery cannulation | 1
anaesthesia maintained with isoflurane | 1
anaesthesia maintained with N2O-O2 mixture | 1
anaesthesia maintained with atracurium | 1
fentanyl | 2
oxytocin infusion | 2
caesarean delivery | 2
hypotension | 2
packed red blood cells transfusion | 2
fresh frozen plasma transfusion | 2
platelets transfusion | 2
noradrenaline infusion | 2
mild acidosis | 2
normal electrolytes | 2
normal serum glucose | 2
intensive care unit | 2
post-operative analgesia | 2
ultrasound guided bilateral transverse abdominis plane block | 2
pulmonary haemorrhage | 48
blood products transfusion | 48
bed side fibre-optic bronchoscopy | 48
erythematous mucosa | 48
blood clots | 48
active oozing | 48
diffuse bleeding | 48
broncho alveolar lavage | 48
Factor VIIa administration | 48
bleeding cessation | 60
reduction of inspired oxygen fraction | 60
bilateral non-homogeneous opacities | 48
acute kidney injury | 48
severe hyperbilirubinemia | 48
haemolytic uremic syndrome | 48
plasmapheresis | 72
dialysis | 72
diffuse cerebral oedema | 72
cerebroprotective measures | 72
stress ulcer prevention | 72
deep vein thrombosis prophylaxis | 72
glycemic control | 72
reducing fever | 96
improving consciousness | 96
inotropic support tapered | 96
improving urine output | 96
improving liver function test | 96
improving coagulation parameters | 96
improving Pao2/Fio2 ratio | 96
extubation | 144
discharged from the hospital | 168