70 years old | 0
    male | 0
    hypertension | 0
    chronic obstructive pulmonary disease | 0
    referred due to erythroderma | -17520
    intense pruritus | -17520
    refractory to topical corticosteroid therapy | -17520
    refractory to oral corticosteroid therapy | -17520
    shiny, bright red erythroderma | 0
    slightly indurated to palpation | 0
    bilateral axillary lymph nodes palpable | 0
    bilateral inguinal lymph nodes palpable | 0
    basophilia of 14.1% | 0
    slightly elevated LDH (253 IU/l) | 0
    skin biopsy revealed parakeratosis | 0
    dense lymphocytic infiltrate in the papillary dermis | 0
    epidermotropism | 0
    immunohistochemical analysis positive for CD2 | 0
    immunohistochemical analysis positive for CD3 |6
    immunohistochemical analysis positive for CD4 |0
    immunohistochemical analysis positive for CD5 |0
    immunohistochemical analysis negative for CD7 |0
    immunohistochemical analysis negative for CD8 |0
    numerous enlarged lymph nodes in cervical regions |0
    numerous enlarged lymph nodes in axillary regions |0
    numerous enlarged lymph nodes in inguinal regions |0
    Sézary cell count of 1031/mm3 |0
    paracortical infiltration due to Sézary syndrome |0
    Sézary syndrome diagnosis |0
    treatment with PUVA therapy |0
    treatment with interferon alpha |0
    treatment with bexarotene |0
    treatment with extracorporeal photopheresis |0
    disease progression with enlarged lymph nodes |0
    pruritus became uncontrollable |0
    LUC 56.8% |0
    basophilia 26% |0
    treatment initiation with alemtuzumab |0
    alemtuzumab 30mg subcutaneously three times a week |0
    received cotrimoxazole |0
    received famciclovir |0
    received valganciclovir |0
    marked improvement with 80% erythroderma clearance |2160
    pruritus cessation |2160
    Sézary cell count decrease to 0 |2160
    treatment withdrawal due to severe neutropenia |2880
    leukocytes 0.3 × 103/µl |2880
    neutrophils 0.12 × 103/µl |2880
    grade IV heart failure |2880
    acute exacerbation of underlying disease with bronchospasm |2880
    intensive care unit admission |2880
    recovery with supportive treatment |2880
    G-CSF therapy |2880
    no signs of clinical disease activity |11088
    no signs of haematological disease activity |11088
    