55 years old | 0  
    female | 0  
    admitted to the hospital | 0  
    fever | -24  
    cough | -24  
    progressive lower limb edema | -24  
    abdominal distention | -24  
    type 2 diabetes mellitus | 0  
    oral metformin | 0  
    oral amlodipine | 0  
    non-smoker | 0  
    no alcohol consumption | 0  
    no history of drug abuse | 0  
    mild peripheral blood leukocytosis | 0  
    thrombocytopenia | 0  
    hypoalbuminemia | 0  
    hyperbilirubinemia | 0  
    normal creatinine | 0  
    chest X-ray right-sided pleural effusion | 0  
    empirical antibiotics | 0  
    increased diuretics dosage | 0  
    ascitic fluid drained | 0  
    pleural fluid drained | 0  
    urine culture positive for Streptococcus agalactiae | 0  
    clinical improvement | 0  
    repeated chest X-ray reduction in right hydrothorax | 0  
    discharged | 168  
    oral ciprofloxacin | 168  
    oral lasix | 168  
    multivitamins | 168  
    admitted for elective liver transplant | 672  
    total hepatectomy | 672  
    transplantation with full right lobe graft | 672  
    three biliary anastomoses | 672  
    arterial anastomosis repeated twice | 672  
    transfusion of 12 units packed red blood cells | 672  
    transferred to ICU | 672  
    extubated | 696  
    re-intubated due to ARDS | 744  
    immunosuppressive therapy | 0  
    oral tacrolimus | 0  
    oral mycophenolate mofetil | 0  
    oral prednisolone | 0  
    anastomotic biliary stricture | 0  
    bile leak | 0  
    percutaneous transhepatic cholangiography | 0  
    percutaneous transhepatic biliary drainage | 0  
    internal-external biliary catheter | 0  
    pigtail catheter | 0  
    drains kept in place | 0  
    pigtail catheter removed | 504  
    internal-external PTBD catheter left in place | 504  
    right upper quadrant abdominal pain | 504  
    no fever | 504  
    no vomiting | 504  
    no change in peripheral blood leukocyte count | 504  
    no change in bilirubin | 504  
    no change in ALT | 504  
    no change in alkaline phosphatase | 504  
    increased CRP | 504  
    ultrasound right-sided sub-diaphragmatic collection | 504  
    septic screen | 504  
    IV meropenem | 504  
    PTBD catheter culture positive for E. meningoseptica | 504  
    IV meropenem changed to IV ciprofloxacin | 504  
    IV metronidazole | 504  
    repeat PTBD catheter fluid culture | 528  
    repeat culture positive for E. meningoseptica | 552  
    clinical improvement | 504  
    abdominal pain resolved | 504  
    antibiotics continued for two weeks | 504  
    asymptomatic | 672  
    normal leukocyte count | 672  
    CRP drop | 672  
    repeat fluid cultures negative | 672  
    no complications from antibiotic treatment | 672  

