67 years old | 0
female | 0
caucasian | 0
renal transplantation | 0
chronic renal failure | -672
unconfirmed chronic glomerulonephritis | -672
basiliximab | 0
tacrolimus | 0
mycophenolate mofetil | 0
prednisolone | 0
late onset of graft function | 0
haemodialysis dependent | 0
severe combined acute cellular rejection | 168
antibody mediated C4d positive rejection | 168
rabbit antithymocyte globulin | 168
plasmapheresis | 168
intravenous immunoglobulins | 168
recovery of graft function | 336
elevation of amylase | 0
elevation of lipase | 0
ultrasound examination | 0
solitary stone in gall bladder | 0
conservative therapy | 0
reduction of mycophenolate mofetil | 0
progressive sharp pain | 2160
abdominal region | 2160
temperatures exceeding 39 C | 2160
shivering | 2160
admission to surgery clinic | 2160
tacrolimus | 2160
mycophenolate mofetil | 2160
prednisolone | 2160
increased level of serum amylase | 2160
increased level of lipase | 2160
leukocytes | 2160
CRP | 2160
procalcitonin | 2160
acute contrast-enhanced CT scan | 2160
acute pancreatitis | 2160
pancreatic abscess | 2160
subphrenic abscess collections | 2160
fluid between loops of small intestine | 2160
surgical treatment | 2160
transverse laparotomy | 2160
drainage of abscess | 2160
sample collection for cultivation | 2160
severance of ligamentum gastrocolicum | 2160
opening of bursa omentalis | 2160
drainage of abscess | 2160
irrigation of abdominal cavity | 2160
discontinuation of tacrolimus | 2160
discontinuation of mycophenolate mofetil | 2160
administration of corticoids | 2160
cultivation of abscesses | 2160
Escherichia coli | 2160
meropenem | 2160
metronidazole | 2160
progressive increase in azotemia | 2160
manifestations of graft failure | 2160
CVVHD | 2160
extubation | 2160
support of vasopressors | 2160
spontaneous diuresis | 2160
follow-up CECT scan | 2160
reduction of inflammatory parameters | 2160
stabilisation of laboratory values | 2160
renewal of immunosuppressive therapy | 2160
reduction of corticoids | 2160
full sustenance | 3024
surgical wound locally bandaged | 3024
VAC system | 3024
transfer to nephrological department | 3024
discharge for home care | 3024
diagnostic rebiopsy of graft | 4320
no signs of rejection | 4320
immunosuppressive medication | 4320
tacrolimus | 4320
prednisolone | 4320
good graft function | 4320