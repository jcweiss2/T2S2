26 years old | 0
female | 0
sickle cell trait | 0
presented to the emergency department | 0
altered mental status | 0
recovered from a viral illness | -336
presented to the emergency department | -168
shortness of breath | -168
diffuse pain | -168
became acutely unresponsive | 0
30-s pulseless electrical activity arrest | 0
return of spontaneous circulation | 0
transferred to a higher acuity facility | 0
admitted to the intensive care unit | 0
multisystem organ failure | 0
acute respiratory distress syndrome | 0
acute renal failure | 0
bone marrow failure | 0
hemoglobin 5.7 g/dL | 0
platelets 57 K/μL | 0
leukocytes 27.33 K/μL | 0
neutrophil-predominant | 0
MRI of the brain | 24
diffuse scattered areas of restricted diffusion | 24
transcranial Doppler | 168
increased velocity of the left middle cerebral artery | 168
increased pulsatility indices diffusely | 168
echocardiography | 0
global hypokinesis | 0
left ventricular ejection fraction of 40% | 0
concern for sickle cell crisis | 0
thrombotic thrombocytopenic purpura | 0
schistocytes seen on peripheral blood smear | 0
started on broad-spectrum antimicrobials | 0
plasma exchange | 0
methylprednisolone | 0
hemoglobin electrophoresis | 120
confirmed HbSC disease | 120
ADAMSTS activity >10% | 120
peripheral blood smear | 120
schistocytes | 120
neutrophil-containing morulae | 120
bone marrow biopsy | 120
normocellular marrow | 120
trophozoites in multiple RBCs | 120
started on clindamycin | 120
started on atovaquone | 120
started on doxycycline | 120
anaplasmosis-induced sickle cell crisis | 120
Babesia coinfection | 120
PCR for anaplasmosis negative | 120
PCR for babesiosis negative | 120
treatment for babesiosis stopped | 120
continued for anaplasmosis | 120
neurologic examination | 144
eyes open spontaneously | 144
decerebrate posturing | 144
not following commands | 144
eculizumab treatment | 264
worsening renal function | 264
suspected atypical hemolytic uremic syndrome | 264
continued for 3 weeks | 264
transferred out of intensive care | 744
care gradually deescalated | 744
mental status not improved | 1176
discharged | 1176
tracheostomy | 1176
percutaneous endoscopic gastrostomy | 1176
