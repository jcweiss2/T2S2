64 years old | 0
male | 0
admitted to the hospital | 0
acute pancreatitis | 0
Imrie/Glassgow Score = 6 | 0
biliary pathology | 0
CT scan of the abdomen | 0
extensive edematous changes | 0
hepatoportal venous gas (HPVG) | 0
concern regarding one segment of small bowel | 0
CT mesenteric angiogram | 2
poorly enhancing segment of small bowel | 2
venous thrombosis | 2
reduction in the volume of HPVG | 2
emergency laparotomy | 2
resection of a nonviable ischemic segment of small bowel | 2
omental saponification | 2
prolonged intensive care admission | 2
multiorgan dysfunction | 2
acute kidney injury | 2
adult respiratory distress syndrome | 2
discharged to the ward | 45
readmitted to the intensive care unit | 48
overwhelming sepsis | 48
repeat imaging | 48
large peripancreatic necrotic collections | 48
interventional radiology drainages | 48
antimicrobials | 48
antifungal | 48
inotropic support | 48
deteriorated | 48
died | 62
diagnosis of acute pancreatitis | -24
underlying biliary pathology | -24
initial computed tomography (CT) scan | 0 
extensive edematous changes involving the entire pancreas | 0 
significant volume of HPVG | 0 
concern regarding one segment of small bowel | 0 
CT mesenteric angiogram | 2 
poorly enhancing segment of small bowel | 2 
concerning for venous thrombosis | 2 
significant reduction in the volume of HPVG | 2 
decision to proceed for emergency laparotomy | 2 
emergency laparotomy | 2 
resection of a nonviable ischemic segment of small bowel | 2 
omental saponification | 2 
prolonged intensive care admission | 2 
management of multiorgan dysfunction | 2 
acute kidney injury | 2 
adult respiratory distress syndrome | 2 
discharged to the ward | 45 
readmitted to the intensive care unit | 48 
overwhelming sepsis | 48 
repeat imaging | 48 
large peripancreatic necrotic collections | 48 
interventional radiology drainages | 48 
escalation in both antimicrobials | 48 
antifungal | 48 
inotropic support | 48 
deteriorated | 48 
died | 62