55 years old | 0
male | 0
alcohol abuse | 0
leukopenia | 0
shortness of breath | -48
cough | -48
fever | -48
chills | -48
confusion | -48
altered mental status | -48
unconscious | 0
no witnessed seizure | 0
no trauma | 0
last seen conscious | -12
intubated | 0
assist-control mechanical ventilation | 0
sinus tachycardia | 0
hypotension | 0
vasopressors | 0
right-sided decreased air entry | 0
diffuse crackles | 0
white blood cells 0.8 × 10^9/L | 0
absolute neutrophil count 360 mm^3 | 0
hemoglobin 8.1 g/L | 0
platelets 109,000 | 0
creatinine 3.5 mg/dl | 0
potassium 4.5 meq/L | 0
right lower lobe consolidation | 0
right pleural effusion suggested | 0
no pleural effusion | 0
bronchial secretions culture grows gram-positive diplococci | 0
Streptococcus pneumoniae | 0
ALPS syndrome | 0
admitted to intensive care unit | 0
vancomycin | 0
piperacillin/tazobactam | 0
discharged | 72
