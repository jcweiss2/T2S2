35 years old | 0
female | 0
gave birth to healthy twins | -24
in vitro fertilization | -280
facial nerve paresis | -672
severe headache | 24
generalized tonic–clonic seizures | 24
loss of consciousness | 24
arterial blood pressure 195/110 mmHg | 24
heart rate 120 beats/min | 24
eclampsia | 24
intravenous infusion of magnesium sulphate | 24
ebrantil | 24
20% manitol | 24
diazepam | 24
bilateral vision loss | 48
proteinuria 2+ | 48
cortical blindness | 48
mild right-sided facial nerve paresis | 48
hypodensity of the posterior white matter | 48
vasogenic edema | 48
T2- and fluid-attenuated inversion recovery-weighted images | 48
hyperintense signals in the white matter | 48
predominantly in the parietal and occipital regions | 48
junctions of vascular watershed zones of the brain | 48
antihypertensive therapy | 48
enalapril maleate | 72
methyldopa | 72
human albumin | 72
significant bilateral improvement of the visual function | 120
best-corrected visual acuity 1.0 | 120
bilateral peripheral relative scotoma | 120
depressed sensitivity of the paracentral left visual field | 120
right-sided partial facial nerve paresis | 120
significant regression of the edema | 168
discrete residual changes over the posterior horns of the side ventricles | 168
discharged | 216