60 years old | 0
menopausal | 0
postmenopausal metrorrhagia | 0
postmenopausal bleeding | 0
endovaginal ultrasound | 0
intracavitary image of 15 mm | 0
polyp | 0
hysteroscopic surgery | 0
polyp resection | 0
endometrial biopsy | 0
abdominal pelvic pain | 48
tachycardic | 48
febrile | 48
hypotensive | 48
saturation of 90% | 48
diffuse abdominal sensibility | 48
computed tomography (CT) scan | 48
desaturation | 48
fall of pressure to 90/50 mmHg | 48
admitted to the recovery room | 48
biological sample | 48
C-reactive protein 360 | 48
blood gases | 48
lactate 4 | 48
intubated | 48
Glasgow coma scale 12 | 48
desaturation at 80% | 48
intra-uterine collection | 48
hydroaeric level | 48
increased uterus size | 48
gynecological examination | 48
aspiration of the collection | 48
fetid blood | 48
bacteriological samples | 48
blood cultures | 48
antibiotic therapy | 48
imipinem | 48
amikacine | 48
vasoactive drug | 48
noradrenaline | 48
septic shock | 51
death | 51
sensitive Escherichia coli | 51
hypertensive | 0
amlodipine | 0
no perforation | 48
no pelvic peritonitis | 48
