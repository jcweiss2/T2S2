19 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
army officer | 0 | 0 | Factual
fever | -120 | 0 | Factual
arthralgia | -120 | 0 | Factual
myalgia | -120 | 0 | Factual
headache | -120 | 0 | Factual
productive cough | -120 | 0 | Factual
yellowish sputum | -120 | 0 | Factual
chest heaviness | -120 | 0 | Factual
dyspnea | -120 | 0 | Factual
diarrhea | -120 | 0 | Factual
reduced oral intake | -120 | 0 | Factual
no history of travelling | 0 | 0 | Factual
no recent jungle activities | 0 | 0 | Factual
no past medical illness | 0 | 0 | Factual
no previous hospitalization | 0 | 0 | Factual
no medical treatment for current condition | 0 | 0 | Factual
conscious | 0 | 0 | Factual
dehydrated | 0 | 0 | Factual
cold peripheries | 0 | 0 | Factual
febrile | 0 | 0 | Factual
temperature of 38.5°C | 0 | 0 | Factual
hypotensive | 0 | 0 | Factual
blood pressure of 81/53 mmHg | 0 | 0 | Factual
tachycardic | 0 | 0 | Factual
heart rate of 146 beats per minute | 0 | 0 | Factual
tachypnoeic | 0 | 0 | Factual
respiratory rate of 30 breaths per minute | 0 | 0 | Factual
oxygen saturation of 75-80% | 0 | 0 | Factual
coarse crepitation over both lower lung zones | 0 | 0 | Factual
tenderness at epigastric region | 0 | 0 | Factual
palpable liver | 0 | 0 | Factual
no cervical lymph nodes | 0 | 0 | Factual
no inguinal lymph nodes | 0 | 0 | Factual
no axillary lymph nodes | 0 | 0 | Factual
haemoglobin of 11.3 g/dL | 0 | 0 | Factual
low white blood cell count | 0 | 0 | Factual
neutrophil predominance | 0 | 0 | Factual
platelet count of 80 × 10^6/L | 0 | 0 | Factual
C-reactive protein of 28.28 mg/dL | 0 | 0 | Factual
acute kidney injury | 0 | 0 | Factual
serum sodium of 137 mmol/L | 0 | 0 | Factual
serum potassium of 3.7 mmol/L | 0 | 0 | Factual
serum urea of 14 mmol/L | 0 | 0 | Factual
serum creatinine of 206 μmol/L | 0 | 0 | Factual
liver function tests normal | 0 | 0 | Factual
serum albumin of 22 g/dL | 0 | 0 | Factual
creatinine kinase of 351 IU/L | 0 | 0 | Factual
arterial blood gases on room air | 0 | 0 | Factual
pH of 7.378 | 0 | 0 | Factual
pCO2 of 37 mmHg | 0 | 0 | Factual
pO2 of 52.7 mmHg | 0 | 0 | Factual
O2 saturation of 89% | 0 | 0 | Factual
HCO3 of 21.7 mmol/L | 0 | 0 | Factual
Dengue NS-1 Antigen negative | 0 | 0 | Factual
IgG and IgM antibody negative | 0 | 0 | Factual
chest radiograph showed consolidation | 0 | 0 | Factual
diagnosis of severe community acquired pneumonia | 0 | 0 | Factual
acute kidney injury | 0 | 0 | Factual
resuscitation with normal saline | 0 | 0 | Factual
non-invasive ventilation | 0 | 0 | Factual
inotropic support | 0 | 24 | Factual
intravenous ceftriaxone | 0 | 24 | Factual
intravenous azithromycin | 0 | 24 | Factual
intubation | 24 | 24 | Factual
mechanical ventilation | 24 | 72 | Factual
bronchoscopy | 24 | 24 | Factual
haemoserous and greenish secretion | 24 | 24 | Factual
repeated chest radiograph showed worsening consolidation | 24 | 24 | Factual
abscess formation | 24 | 24 | Factual
intravenous meropenem | 24 | 72 | Factual
intravenous cloxacillin | 24 | 72 | Factual
antiviral oseltamivir | 24 | 72 | Factual
continuous venous-venous haemofiltration | 24 | 72 | Factual
severe metabolic acidosis | 24 | 72 | Factual
oliguric acute kidney injury | 24 | 72 | Factual
persistent spiking of temperature | 24 | 72 | Factual
worsening of septic parameters | 24 | 72 | Factual
refractory hypotension | 24 | 72 | Factual
death | 72 | 72 | Factual
blood cultures negative | 0 | 72 | Factual
atypical bacterial and Leptospiral serologies negative | 0 | 72 | Factual
Hepatitis B/C and HIV serologies undetected | 0 | 72 | Factual
respiratory viruses screening negative | 0 | 72 | Factual
tracheal aspiration and bronchoalveolar lavage positive for MDR Acinetobacter baumannii | 0 | 72 | Factual
MDR Acinetobacter baumannii susceptible to polymyxin B | 0 | 72 | Factual
minimum inhibitory concentration of 0.5 μg/ml | 0 | 72 | Factual
MDR Acinetobacter baumannii resistant to penicillin group | 0 | 72 | Factual
MDR Acinetobacter baumannii resistant to ampicillin/sulbactam | 0 | 72 | Factual
MDR Acinetobacter baumannii resistant to third generation cephalosporins | 0 | 72 | Factual
MDR Acinetobacter baumannii resistant to fluoroquinolone | 0 | 72 | Factual
MDR Acinetobacter baumannii resistant to carbapenem group | 0 | 72 | Factual
PCR for carbapenemases genes NDM, OXA-23, OXA 24 or OXA-58 not performed | 0 | 72 | Factual