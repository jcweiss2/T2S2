55 years old | 0
male | 0
admitted to the intensive care unit | 0
motorcycle accident | -1
sternal lesions | 0
humeral lesions | 0
D4 vertebral fractures | 0
D9 vertebral fractures | 0
hypertensive pneumothorax | 0
Glasgow Coma Score of 14/15 | 0
intracapsular spleen haematoma | 0
multiple fractures of the pelvis | 0
empirical therapy with ceftazidime and gentamicin | 120
fever | 144
septic shock | 144
severe leucocytosis | 144
low platelet count | 144
vasoactive amines | 144
mechanical ventilation | 144
monolateral purulent pleural suffusion | 144
thoracic drainage | 144
blood samples taken for culture | 144
growth of pleomorphic Gram-positive microorganisms | 226
identification by 16S rRNA PCR amplification and sequencing | 226
identification of C. hongkongensis | 226
antimicrobial susceptibility testing | 226
discontinuation of empirical treatment with vancomycin and meropenem | 336
recovery from sepsis | 336