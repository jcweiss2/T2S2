54 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
pre-syncope | -0.1 | 0 | Factual
syncope | -0.1 | 0 | Factual
left-sided chest tightness | -0.1 | 0 | Factual
generalized fatigue | -336 | 0 | Factual
weight loss | -336 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
weight of 41 kg | 0 | 0 | Factual
blood pressure of 96/60 mm Hg | 0 | 0 | Factual
unremarkable cardiac examination | 0 | 0 | Factual
unremarkable respiratory examination | 0 | 0 | Factual
diffuse erythematous rash | 0 | 0 | Factual
normal sinus rhythm | 0 | 0 | Factual
raised troponin concentration | 0 | 0 | Factual
eosinophil count of 7.6 × 10^9/l | 0 | 0 | Factual
referred to cardiology | 0 | 0 | Factual
myocarditis | 0 | 0 | Possible
cardiac magnetic resonance imaging | 24 | 24 | Factual
coronary angiography | 24 | 24 | Factual
no coronary artery disease | 24 | 24 | Factual
skin biopsy | 48 | 48 | Factual
cardiac biopsy | 48 | 48 | Possible
edoxaban | 72 | 720 | Factual
prednisolone | 72 | 720 | Factual
follow-up in the rheumatology clinic | 336 | 336 | Factual
missed appointment | 720 | 720 | Factual
neck swelling | 1440 | 1440 | Factual
urgently admitted to hospital | 1440 | 1440 | Factual
eosinophil count of 19.7 × 10^9 cells/l | 1440 | 1440 | Factual
increase dose of prednisolone | 1440 | 1440 | Factual
computed tomography of neck | 1440 | 1440 | Factual
lymphadenopathy | 1440 | 1440 | Factual
T-cell lymphoma | 1440 | 1440 | Factual
cyclophosphamide therapy | 1440 | 2016 | Factual
sepsis | 1680 | 1680 | Factual
cholecystitis | 1680 | 1680 | Factual
new onset of seizures | 1680 | 1680 | Factual
reduction in consciousness | 1680 | 1680 | Factual
Glasgow Coma Scale of 9/15 | 1680 | 1680 | Factual
head CT | 1680 | 1680 | Factual
multiple bilateral acute infarctions | 1680 | 1680 | Factual
transferred to intensive care unit | 1680 | 1680 | Factual
hepatitis B | -8760 | 0 | Factual
asthma | -8760 | 0 | Factual
intravenous drug use | -8760 | 0 | Factual
excessive use of alcohol | -8760 | 0 | Factual
ischemic stroke | 1680 | 1680 | Possible
reduced GCS score | 1680 | 1680 | Factual
intracranial bleeding | 1680 | 1680 | Possible
malignancy | 1440 | 1440 | Factual
intracerebral infection | 1680 | 1680 | Possible
CMR | 24 | 24 | Factual
subendocardial late gadolinium enhancement | 24 | 24 | Factual
mild LV systolic impairment | 24 | 24 | Factual
eczematous changes | 48 | 48 | Factual
bone marrow biopsy | 48 | 48 | Factual
no increase in eosinophils | 48 | 48 | Factual
axillary lymph node biopsy | 1440 | 1440 | Factual
T-cell lymphoma | 1440 | 1440 | Factual
embolic brain event | 1680 | 1680 | Factual
intracardiac thrombus | 1680 | 1680 | Possible
apical tear | 1680 | 1680 | Factual
intramural myocardial tear | 1680 | 1680 | Factual
small apical cavity | 1680 | 1680 | Factual
mobile structures attached to dissected myocardium | 1680 | 1680 | Factual
diastolic flow in the apical cavity | 1680 | 1680 | Factual
systolic flow out of the apical cavity | 1680 | 1680 | Factual
corticosteroids | 72 | 720 | Factual
anticoagulation | 72 | 720 | Factual
palliation | 2016 | 2016 | Factual
deterioration | 2016 | 2016 | Factual
poor prognosis | 2016 | 2016 | Factual