67 years old | 0
male | 0
Caucasian | 0
admitted to the hospital | 0
coronary artery disease | -2160
type II diabetes | -2160
hypertension | -2160
peripheral vascular disease | -2160
normal renal function | 0
septic arthritis of the right knee | 0
coronary artery bypass | -672
Staphylococcus aureus infection | -672
septicemias | -168
disseminated Staphylococcus aureus infections | -168
mechanical ventilation | -168
ARDS | -168
five surgical revisions | -168
haemodynamically unstable | -264
vasopressors | -264
broad-spectrum antibiotics | -264
renal function deterioration | -360
oliguric acute renal failure | -360
sepsis | -360
nephrotoxic medication | -360
COX-2 inhibitor | -360
gentamycin | -360
ACEI | -360
continuous venovenous haemofiltration | -432
uraemia | -432
metabolic acidosis | -432
encephalopathy | -432
serum creatinine stabilization | -480
anuric ARF | -576
hydration | -576
diuretics | -576
10% pentastarch | -528
intermittent haemodialysis | -624
renal ultrasound | -624
normal sized kidneys | -624
no hydronephrosis | -624
urinary sediment | -624
dirty brown casts | -624
no eosinophilia | -624
fractional excretion of sodium | -624
renal radionuclide study | -624
bilateral hypoperfusion | -624
renal blood flow | -624
renal biopsy | -624
severe hydropic changes | -624
cytoplasm of tubular cells | -624
discharged from hospital | 4320
chronic haemodialysis | 4320