57 years old | 0 | 0 
female | 0 | 0 
menopausal | 0 | 0 
admitted to the gynecological emergency unit | 0 | 0 
left lower quadrant abdominal pain | -1008 | 0 
pelvic heaviness | -1008 | 0 
urinary frequency | -1008 | 0 
past history of 5 miscarriages | -1008 | 0 
tubal ligation | -1008 | 0 
active smoker | 0 | 0 
no medication | 0 | 0 
large and painful mass | 0 | 0 
pelvic MRI | 0 | 0 
mass measuring 18 × 17 × 12 cm | 0 | 0 
serum tumor markers were negative | 0 | 0 
surgical pelvic exploration | 672 | 672 
total hysterectomy with adnexectomy | 672 | 672 
removal of the mass | 672 | 672 
definitive histological diagnosis was leiomyosarcoma | 672 | 672 
isolated fever | 48 | 48 
laboratory evaluation | 48 | 48 
major inflammatory syndrome | 48 | 48 
contrast-enhanced computed tomography scan | 48 | 48 
abscess | 48 | 48 
blood pressure dropped | 48 | 48 
vasopressor therapy | 48 | 48 
emergency revision surgery | 48 | 48 
peritoneal cavity exploration | 48 | 48 
moderately abundant non-purulent serosanginous peritoneal fluid | 48 | 48 
adhesions to the Douglas pouch | 48 | 48 
peritonitis | 48 | 48 
antibacterial treatment with piperacillin/tazobactam and gentamicin | 48 | 48 
extubated | 72 | 72 
hemodynamic support with noradrenaline | 72 | 72 
transferred to the intensive care unit | 72 | 72 
noradrenaline requirement decreased | 96 | 96 
discontinuation of noradrenaline | 96 | 96 
decrease in inflammatory markers | 96 | 96 
microbiological analysis of the peritoneal fluid identified Gardnerella vaginalis | 96 | 96 
gentamicin was discontinued | 96 | 96 
metronidazole was added | 96 | 96 
Atopobium vaginae was identified | 120 | 120 
antibacterial susceptibility testing of Garderella vaginalis | 120 | 120 
antibacterial susceptibility testing of Atopobium vaginae | 120 | 120 
discharged from the intensive care unit | 120 | 120 
antibacterial therapy was stopped | 168 | 168 
final diagnosis was an early postoperative peritonitis-induced septic shock | 168 | 168 
Gardnerella vaginalis and Atopobium vaginae | 168 | 168 
vaginal incision in the abdominal cavity | 672 | 672 
bacterial dissemination | 672 | 672 
peritonitis | 48 | 48 
septic shock | 48 | 48 
asymptomatic carrier | 0 | 0 
vaginal flora | 0 | 0 
male urethral flora | 0 | 0 
bacterial vaginosis | 0 | 0 
secnidazole or metronidazole | 0 | 0 
antimicrobial resistance pattern testing | 120 | 120 
broad-spectrum antibacterial therapy | 48 | 48 
piperacillin/tazobactam | 48 | 48 
Gardnerella vaginalis was resistant to metronidazole | 120 | 120 
Atopobium vaginae was sensitive to metronidazole | 120 | 120 
post-caesarean septic shock | 0 | 0 
Peptostreptococcus | 0 | 0 
bacteremia after vaginal myomectomy | 0 | 0 
vertebral osteomyelitis | 0 | 0 
prostatic adenoma | 0 | 0 
tubo-ovarian abscess | 0 | 0 
endocarditis of the tricuspid valve | 0 | 0 
immunodepression | 0 | 0 
type 1 diabetes | 0 | 0 
chronic alcoholism | 0 | 0 
genital area | 0 | 0 
post-operative infection | 48 | 168 
differential diagnosis | 0 | 0