62 years old | 0
male | 0
admitted to the hospital | 0
arterial hypertension | 0
dilated heart disease of ischemic origin | 0
severe left ventricular dysfunction | 0
chronic hepatitis B infection | 0
left colostomy carrier | 0
complicated acute diverticulitis | - time unknown, assume -720 
bilateral SARS-CoV-2 pneumonia | -504
onset of symptoms | -504
Pulmonary CT | 0
severe bilateral SARS-CoV-2 lung infection | 0
high-flow oxygen therapy | 0
dexamethasone | 0
ceftriaxone | 0
piperacillin-tazobactam | 0
intubation | 0
mechanical ventilation | 0
prone position sessions | 0
severe acute respiratory distress syndrome (ARDS) | 0
PaO2/FiO2 <100mmHg | 0
APACHE II: 11 points | 0
SOFA score: 9 points | 0
nosocomial pneumonia | 264
empirical therapy | 264
meropenem | 264
linezolid | 264
P. aeruginosa (AmpC profile) | 264
tracheobronchial aspirate | 264
meropenem MIC 1 mg/L | 264
antibiotic treatment adjusted | 264
meropenem | 264
new episode of nosocomial pneumonia | 1296
secondary bacteremia | 1296
Carbapenem-resistant P. aeruginosa | 1296
meropenem MIC > 16 mg/L | 1296
initial empirical treatment | 1296
meropenem | 1296
colistin | 1296
ceftazidime-avibactam | 1296
tracheobronchitis | 1872
extensively drug-resistant P. aeruginosa | 1872
ceftazidime-avibactam resistance | 1872
ceftalozane-tazobactam | 1872
inhaled colistin | 1872
prolonged mechanical ventilation | 0
tracheostomy | 0
multiple weaning attempts | 0
Aspergillus fumigatus | - time unknown, assume 1000
Enterococcus faecium bacteremia | - time unknown, assume 1000
febrile episodes | - time unknown, assume 1000
multiple antibiotics | - time unknown, assume 1000
discharged from ICU | 2000 
transferred to a rehabilitation healthcare center | 2000