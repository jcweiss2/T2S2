78 years old | 0
female | 0
myasthenia gravis | -672
hypertension | -672
chronic kidney disease | -672
obesity | -672
proctosigmoidectomy | -240
L3-L4 laminectomy | -240
foraminotomy | -240
implantation of a percutaneous spinal cord stimulator | -168
admitted to the intensive care unit | -120
myasthenic crisis | -120
dysphagia | -120
ptosis | -120
dysarthria | -120
intubated | -120
plasma exchange | -120
prednisone | -120
pyridostigmine | -120
discharged home | -90
neurology follow up appointment | -60
mycophenolate | -60
prednisone dosage decreased | -60
admitted to the hospital | 0
right shoulder pain | 0
fever | -72
chills | -72
sweats | -72
left-hand cellulitis | -30
contrasted computerized tomography of left upper extremity | -30
soft tissue ulceration | -30
cellulitis | -30
intramuscular abscess | -30
ceftaroline | -30
doxycycline | -30
trimethoprim-sulfamethoxazole | -30
Nocardia farcinica | -30
discharged home | -30
right shoulder pain worsened | -168
persistent right shoulder pain | -168
intermittent right shoulder pain | -504
temperature | 0
heart rate | 0
respiratory rate | 0
blood pressure | 0
oxygen saturation | 0
examination of right shoulder | 0
pain with passive range of motion | 0
limited active range of motion | 0
no overlying erythema | 0
no warmth | 0
no swelling | 0
white blood cell count | 0
absolute neutrophil count | 0
c-reactive protein | 0
erythrocyte sedimentation rate | 0
comprehensive metabolic panel | 0
contrasted CT of right shoulder | 0
multi loculated collections | 0
subacromial bursa | 0
glenohumeral joint effusion | 0
bedside arthrocentesis | 24
fluid analysis | 24
white blood cell count | 24
neutrophilic | 24
lymphocytic | 24
monocytic | 24
no crystals | 24
gram stain | 24
N. farcinica | 24
operative debridement | 72
glenohumeral joint | 72
foul smelling purulent material | 72
abscesses | 72
periscapular fluid | 72
N. farcinica | 72
meropenem | 120
TMP-SMX | 120
leukocytosis | 240
CRP | 240
ESR | 240
repeat contrasted CT | 240
decreased fluid collections | 240
noncontrasted CT of chest | 240
bibasilar effusions | 240
bibasilar infiltrates | 240
scattered nodularity | 240
no abscesses | 240
noncontrasted CT of head | 240
no intracranial abscesses | 240
dual antimicrobial therapy | 240
intravenous meropenem | 240
oral high dose TMP-SMX | 240
carbapenem resistance | 720
thrombocytopenia | 720
amoxicillin-clavulanate | 720
altered mentation | 720
failure to thrive | 720
hospice care | 720