40 years old | 0
    female | 0
    lower abdominal pain | -168
    nonbilious vomiting | -168
    loose stools | -168
    occasional breathlessness | -168
    decreased urine output | -168
    fever | -72
    dry tongue | 0
    no pedal edema | 0
    no generalized lymphadenopathy | 0
    pulse rate 130/min | 0
    blood pressure 96/80 mmHg | 0
    oxygen saturation 90% | 0
    respiratory rate 34/min | 0
    body temperature 98.4°F | 0
    tenderness in right iliac fossa | 0
    no palpable mass | 0
    audible bowel sounds | 0
    hemoglobin 98 g/L | 0
    high total leukocyte count 32.98 × 109/L | 0
    platelet count 263.4 × 109/L | 0
    urea 42.83 mmol/L | 0
    creatinine 159.12 mmol/L | 0
    electrolyte tests within normal limits | 0
    total bilirubin 12.65 mmol/L | 0
    direct bilirubin 6.15 mmol/L | 0
    alanine aminotransferase 8.2 mkat/L | 0
    aspartate aminotransferase 50.9 mkat/L | 0
    alkaline phosphatase 247.6 U/L | 0
    gamma-glutamyl transferase 25.2 U/L | 0
    total protein 57 g/L | 0
    albumin 30.8 g/L | 0
    hepatitis C virus positive | 0
    bilateral moderate pleural effusion | 0
    no abnormality on echocardiography | 0
    admitted to surgical department | 0
    intravenous normal saline | 0
    pain management | 0
    supplemental oxygen | 0
    empirical intravenous antibiotic therapy | 0
    ceftriaxone 1 g every 12 h | 0
    metronidazole 500 mg every 8 h | 0
    ultrasound-guided thoracic paracentesis | 0
    purulent aspirate | 0
    pleural fluid gram staining | 0
    AFB staining | 0
    culture and antibiotic sensitivity | 0
    biochemical analysis | 0
    pleural fluid lactate dehydrogenase 68,900 U/L | 0
    serum procalcitonin elevated | 0
    abdominal ultrasound scan detected intrabdominal collection | 0
    bilateral pyothorax | 0
    intra-abdominal collection | 0
    contrast-enhanced CT scan of torso | 2
    bilateral pleural effusion | 2
    ground-glass centrilobular nodules | 2
    acute appendicitis with rupture at tip | 2
    adjacent collection | 2
    communication between peritoneal and pleural cavities | 2
    COVID-19 pneumonia differential | 0
    hollow viscus perforation with acute respiratory distress syndrome differential | 0
    disseminated tuberculosis differential | 0
    non-Hodgkin lymphoma with chylothorax differential | 0
    RT-PCR negative | 0
    erect chest X-ray bilateral pleural effusion | 0
    no free air under diaphragm | 0
    pleural fluid infective nature | 0
    adenosine deaminase 223.5 U/L | 0
    pleural fluid triglycerides normal | 0
    ultrasound scan pleural effusion | 0
    intra-abdominal collection | 0
    disseminated tuberculosis differential | 0
    appendicular perforation differential | 0
    bilateral intercostal tube drainage | 0
    exploratory laparotomy with appendectomy | 0
    retroperitoneal collection 100 ml | 0
    gangrenous appendix | 0
    small and large bowel unremarkable | 0
    no mesenteric lymphadenopathy | 0
    healthy adnexa | 0
    hypotension during surgery | 0
    noradrenaline infusion started | 0
    not extubated | 0
    postoperative ICU admission | 0
    ventilatory support | 0
    noradrenaline support adjusted | 0
    vasopressin infusion started | 0
    urine output maintained | 0
    urea 6.7 mmol/L | 0
    creatinine 97 mmol/L | 0
    tracheostomy on postoperative day 7 | 168
    total parenteral nutrition started | 168
    ionotropic support tapered | 0
    bilateral ICD removal | 0
    chest radiograph lung expansion | 0
    Klebsiella pneumoniae in intraoperative collection | 0
    K. pneumoniae in pleural fluid | 0
    antibiotics adjusted | 0
    blood culture no organism | 0
    pleural fluid AFB negative | 0
    nucleic acid amplification test negative for tuberculosis | 0
    transmural necrosis of appendix | 0
    acute inflammatory infiltrates | 0
    bacterial colonies | 0
    right ICD removal postoperative day 9 | 216
    left ICD removal postoperative day 11 | 264
    TPN through central line | 168
    Ryle’s tube feeding | 168
    oral feeds postoperative day 17 | 408
    ventilator weaning | 432
    shifted out of ICU postoperative day 18 | 432
    suture removal postoperative day 14 | 336
    high-dependency unit monitoring | 432
    discharged postoperative day 21 | 504
    no fresh complaints follow-up | 720
    daily activities without effort | 720
    