66 years old | 0
man | 0
polycystic kidney disease | 0
polycystic liver disease | 0
kidney dialysis for ten years' duration | 0
admitted to the emergency department | 0
acute abdominal pain | 0
left flank pain | -168
fever | -168
vomiting | -168
severe diffuse pain | -48
obstipation | -48
physical examination | 0
temperature of 38.5°C | 0
enlarged left kidney | 0
painful left kidney | 0
diffuse tenderness | 0
purulent urine | 0
white blood count of 10300/mm3 | 0
serum creatinine concentration of 624 μmol/ml | 0
urine culture isolated Escherichia coli | 0
X-ray abdominal exam showed small bowel dilation | 0
enhanced CT scan revealed multiple hepatic cysts | 0
bilaterally enlarged polycystic kidneys | 0
communication between heterogeneous cyst in left kidney and pericolic space | 0
soft tissue thickening in the left mesocolon | 0
increased amount of peritoneal fluid | 0
diagnosis of peritonitis | 0
laparotomy exploration | 0
generalized peritonitis | 0
150 ml purulent collection from ruptured cyst of giant polycystic left kidney | 0
peritoneal lavage | 0
drainage after debridement | 0
bacteriol analysis of the collection isolated Escherichia coli | 0
did not improve with intensive medical support | 72
parenteral antibiotic | 72
died | 72
septic shock | 72
hemodynamic instability | 72
