56 years old | 0
    woman | 0
    admitted with diagnosis of deep neck infection | 0
    neck swelling | -144
    tenderness | -144
    hypertension | -52560
    preoperative airway evaluation | 0
    Mallampatti class IV | 0
    mouth opening of less than three finger widths | 0
    right side retropharyngeal abscess | 0
    extending to the anterior and posterior cervical space | 0
    carotid space | 0
    not premedicated | 0
    blood pressure 140/83 mmHg | 0
    heart rate 110 beats/min | 0
    saturation of percutaneous oxygen (SpO2) 97% | 0
    arterial blood gas analysis | 0
    mild respiratory alkalosis due to tachypnea | 0
    respiration rate of 25 breaths/min | 0
    pH 7.50 | 0
    partial pressure of CO2 34.1 mmHg | 0
    partial pressure of O2 124.6 mmHg | 0
    O2 saturation 99% | 0
    oxygen saturation maintained above 97% throughout the procedure | 0
    preoxygenation administered via facial mask with 100% oxygen | 0
    potentially difficult intubation anticipated | 0
    indirect videolaryngoscope prepared | 0
    endotracheal tubes (ETTs) of various diameters prepared | 0
    lidocaine spray applied | 0
    indirect videolaryngoscopic airway examination performed | 0
    10% lidocaine spray administered via oral cavity | 0
    gargling | 0
    epiglottis visible | 0
    glottis not visible (Cormack and Lehane grade 3) | 0
    intubation using indirect videolaryngoscope performed under general anesthesia | 0
    sugammadex 400 mg prepared | 0
    general anesthesia induced via propofol 120 mg | 0
    rocuronium 60 mg | 0
    mask ventilation feasible | 0
    tidal volume of 300 mL achieved | 0
    peak airway pressure approximately 20 cmH2O | 0
    intubation initially attempted with 7.0 mm ID ETT | 0
    tube changed to 6.5 mm ID ETT | 0
    successfully intubated | 0
    anesthesia maintained with 1.7 volume % sevoflurane | 0
    remifentanil | 0
    2 L/min of air | 0
    2 L/min of O2 | 0
    pressure-controlled ventilation mode used | 0
    end-tidal CO2 maintained at 28–30 mmHg | 0
    pulse oximetry 100% | 0
    incision and retropharyngeal abscess drainage via transcervical approach | 0
    surgeon decided to delay wound closure | 0
    transferred directly to ICU | 0
    breathing maintained via mechanical ventilator | 0
    risk of airway obstruction after extubation | 0
    saturation well controlled at above 95% via pressure-controlled ventilation | 0
    tidal volume 450 mL | 0
    respiration rate 12 breaths/min | 0
    PEEP 5 cmH2O | 0
    FiO2 0.4 | 0
    next day in ICU | 24
    recommenced spontaneous breathing | 24
    successfully extubated | 24
    surgeon decided to perform wound closure and packing gauze removal the following day | 48
    monitored anesthesia care planned | 48
    not premedicated | 48
    noninvasive blood pressure monitoring | 48
    electrocardiography | 48
    pulse oximetry | 48
    end-tidal CO2 measurement via nasal cannula with 100% O2 at 3 L/min | 48
    sedation established via continuous infusion of dexmedetomidine at 6 µg/kg/hr | 48
    SpO2 decreased to 95% | 48
    changed to reservoir mask with 100% O2 administered at 6 L/min | 48
    SpO2 dropped to 94% | 48
    decision to use high-flow nasal cannula | 48
    high-flow nasal cannula set to 30 L/min of humidified oxygen flow | 48
    SpO2 maintained at 100% | 48
    loading dose of dexmedetomidine 6 µg/kg/hr for 10 min | 48
    dose reduced to 0.6 µg/kg/hr | 48
    prior to incision, 50 µg of fentanyl administered | 48
    after approximately 20 min | 48
    fentanyl 50 µg administered | 48
    midazolam 1 mg administered | 48
    dexmedetomidine increased to 0.7–1.0 µg/kg/hr | 48
    patient complained of ongoing discomfort | 48
    vital signs stable | 48
    no signs of bradycardia | 48
    no discomfort reported during subsequent operations | 48
    OAA/S score of 2 maintained | 48
    in recovery room, 100% O2 at 3 L/min supplied via nasal cannula | 48
    O2 saturation maintained at 96–100% | 48
    transported to general hospital room | 48
    discharged on 12th postoperative day | 288
    
    56 years old | 0
    woman | 0
    admitted with diagnosis of deep neck infection | 0
    neck swelling | -144
    tenderness | -144
    hypertension | -52560
    preoperative airway evaluation | 0
    Mallampatti class IV |: 0
    mouth opening of less than three finger widths | 0
    right side retropharyngeal abscess | 0
    extending to the anterior and posterior cervical space | 0
    carotid space | 0
    not premedicated | 0
    blood pressure 140/83 mmHg | 0
    heart rate 110 beats/min | 0
    saturation of percutaneous oxygen (SpO2) 97% | 0
    arterial blood gas analysis | 0
    mild respiratory alkalosis due to tachypnea | 0
    respiration rate of 25 breaths/min | 0
    pH 7.50 | 0
    partial pressure of CO2 34.1 mmHg | 0
    partial pressure of O2 124.6 mmHg | 0
    O2 saturation 99% | 0
    oxygen saturation maintained above 97% throughout the procedure | 0
    preoxygenation administered via facial mask with 100% oxygen | 0
    potentially difficult intubation anticipated | 0
    indirect videolaryngoscope prepared | 0
    endotracheal tubes (ETTs) of various diameters prepared | 0
    lidocaine spray applied | 0
    indirect videolaryngoscopic airway examination performed | 0
    10% lidocaine spray administered via oral cavity | 0
    gargling | 0
    epiglottis visible | 0
    glottis not visible (Cormack and Lehane grade 3) | 0
    intubation using indirect videolaryngoscope performed under general anesthesia | 0
    sugammadex 400 mg prepared | 0
    general anesthesia induced via propofol 120 mg | 0
    rocuronium 60 mg | 0
    mask ventilation feasible | 0
    tidal volume of 300 mL achieved | 0
    peak airway pressure approximately 20 cmH2O | 0
    intubation initially attempted with 7.0 mm ID ETT | 0
    tube changed to 6.5 mm ID ETT | 0
    successfully intubated | 0
    anesthesia maintained with 1.7 volume % sevoflurane | 0
    remifentanil | 0
    2 L/min of air | 0
    2 L/min of O2 | 0
    pressure-controlled ventilation mode used | 0
    end-tidal CO2 maintained at 28–30 mmHg | 0
    pulse oximetry 100% | 0
    incision and retropharyngeal abscess drainage via transcervical approach | 0
    surgeon decided to delay wound closure | 0
    transferred directly to ICU | 0
    breathing maintained via mechanical ventilator | 0
    risk of airway obstruction after extubation | 0
    saturation well controlled at above 95% via pressure-controlled ventilation | 0
    tidal volume 450 mL | 0
    respiration rate 12 breaths/min | 0
    PEEP 5 cmH2O | 0
    FiO2 0.4 | 0
    next day in ICU | 24
    recommenced spontaneous breathing | 24
    successfully extubated | 24
    surgeon decided to perform wound closure and packing gauze removal the following day | 48
    monitored anesthesia care planned | 48
    not premedicated | 48
    noninvasive blood pressure monitoring | 48
    electrocardiography | 48
    pulse oximetry | 48
    end-tidal CO2 measurement via nasal cannula with 100% O2 at 3 L/min | 48
    sedation established via continuous infusion of dexmedetomidine at 6 µg/kg/hr | 48
    SpO2 decreased to 95% | 48
    changed to reservoir mask with 100% O2 administered at 6 L/min | 48
    SpO2 dropped to 94% | 48
    decision to use high-flow nasal cannula | 48
    high-flow nasal cannula set to 30 L/min of humidified oxygen flow | 48
    SpO2 maintained at 100% | 48
    loading dose of dexmedetomidine 6 µg/kg/hr for 10 min | 48
    dose reduced to 0.6 µg/kg/hr | 48
    prior to incision, 50 µg of fentanyl administered | 48
    after approximately 20 min | 48
    fentanyl 50 µg administered | 48
    midazolam 1 mg administered | 48
    dexmedetomidine increased to 0.7–1.0 µg/kg/hr | 48
    patient complained of ongoing discomfort | 48
    vital signs stable | 48
    no signs of bradycardia | 48
    no discomfort reported during subsequent operations | 48
    OAA/S score of 2 maintained | 48
    in recovery room, 100% O2 at 3 L/min supplied via nasal cannula | 48
    O2 saturation maintained at 96–100% | 48
    transported to general hospital room | 48
    discharged on 12th postoperative day | 288
    