84 years old man | 0
    admitted to the hospital's emergency department | 0
    edema of the right leg | -168
    week-long fever | -168
    no current or past history of cardiovascular disease | 0
    no current or past history of any specific diseases | 0
    fully conscious | 0
    pulse rate 70 beats/min | 0
    blood pressure 120/80 mm Hg | 0
    temperature 37.5°C | 0
    pulsatile mass in the abdomen | 0
    white blood cells 4.6 × 103/μL | 0
    hemoglobin 11 g/dL | 0
    C-reactive protein 3.6 mg/dL | 0
    high D-dimer (62 μg/mL) | 0
    high creatinine (2.5 mg/dL) | 0
    high soluble interleukin 2 (IL-2) receptor (10,300 U/mL) | 0
    contrast-enhanced CT showed infrarenal AAA (61 mm in diameter) | 0
    contrast-enhanced CT showed bilateral common iliac artery aneurysms (left 32 mm; right 29 mm) | 0
    contrast-enhanced CT showed periaortic soft tissue density in the retroperitoneal lesion suggestive of hematoma or tumor | 0
    periaortic lesion situated centrally on the right side of the AAA | 0
    periaortic lesion extended from the level of the right renal artery to the region of the right groin | 0
    periaortic lesion compressed the inferior vena cava | 0
    periaortic lesion compressed the right urinary tract | 0
    deep venous thrombosis | 0
    hydronephrosis | 0
    vitamin K antagonist therapy started | 0
    suprarenal inferior vena cava filter placement not performed | 0
    lower leg swelling gradually decreased | 0
    plain MRI scans showed hyperintense signal at the periaortic lesion on diffusion-weighted image compatible with malignant lymphoma | 0
    hemodynamically stable | 0
    no typical symptoms of AAA rupture | 0
    open biopsy in the right groin on the fourth day after admission | 96
    diagnosis of diffuse large B-cell lymphoma | 96
    sepsis due to urinary tract infection developed | 96
    mechanical ventilation required | 96
    endotoxin adsorption therapy by polymyxin B:immobilized fiber column hemoperfusion | 96
    recovered from sepsis | 216
    recovered from respiratory failure | 216
    preliminary informed consent for AAA and malignant lymphoma treatment provided | 216
    asymptomatic | 0
    almost normal renal function | 0
    no therapeutic intervention for unilateral hydronephrosis | 0
    no therapeutic intervention for right urinary tract compression | 0
    too frail for open surgery after intensive care treatment | 0
    EVAR chosen | 0
    right internal iliac artery embolized on day 14 after admission | 336
    endovascular repair with Excluder device on day 18 after admission | 432
    left internal iliac artery embolization | 432
    completion angiography showed no endoleak | 432
    no postoperative aortic events | 432
    chemotherapy for malignant lymphoma not performed | 432
    discharged on postoperative day 49 | 1176
    follow-up CT scans obtained 2 weeks after operation showed no change in aneurysm size | 1176
    follow-up CT scans obtained 2 weeks after operation showed no change in lymphoma size | 1176
    no aortic events in 19 months after operation | 1176
    able to spend most time at home with family | 1176