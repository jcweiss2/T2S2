73 years old | 0
female | 0
admitted to the hospital | 0
hypertension | -672
melena | -24
blood pressure of 110/70 mmHg | 0
heart rate of 108 beats/min | 0
body temperature of 36.8 °C | 0
respiratory rate of 18 breaths/min | 0
no pain complaint | 0
no abdominal mass | 0
red blood cell of 2.51 × 1012/L | 0
hemoglobin of 8 g/dL | 0
white blood cell count of 21.75 G/L | 0
prothrombin of 80% | 0
urea of 14 mmol/L | 0
creatinine of 127 µmol/L | 0
infrarenal abdominal aortic aneurysm (AAA) | 0
esophagogastroduodenoscopy (EGD) | 2
small curvilinear ulcer | 2
red scars | 2
atrophic gastritis | 2
colonoscopy | 2
no bleeding point | 2
moderate upper gastrointestinal (GI) bleeding | 0
gastric ulcer | 0
resuscitated with intravenous fluid administration | 0
red blood cells transfusion | 0
platelets transfusion | 0
proton pump inhibitor infusion | 0
fasting | 0
hemodynamics remained temporarily stable | 24
no more hematochezia | 24
upper abdominal pain | 72
dizziness | 72
hypotension | 72
systolic pressure dropped rapidly to approximately 60 mmHg | 72
heart rate of 120 beats/min | 72
SpO2 of 90% | 72
gastric drainage with much bright red blood | 72
transferred to the Intensive Care Unit | 72
coma | 72
second endoscopy | 72
aggressive attempts at resuscitation | 72
normal saline | 72
packed red blood cell | 72
fresh plasma | 72
vasopressor | 72
tracheal intubation | 72
stomach filled with blood clots | 72
abdominal computed tomography (CT) scan | 72
infrarenal fusiform AAA | 72
ruptured and leaked into the second part of the duodenum | 72
aortoduodenal fistula | 72
urgent endovascular aortic repair (EVAR) | 72
placement of 3 stent graft components | 74
plugging the ruptured aneurysm with histoacryl | 74
no more presence of contrast leak into the gastrointestinal tract | 74
died | 84
multiple organ failures | 84
reversible hypovolemic shock | 84