55 years old | 0
female | 0
height 151cm | 0
weight 61kg | 0
returned from the Philippines | -168
fever | -168
cough | -168
lethargy | -168
myalgia | -168
mild asthma | 0
sleep apnoea | 0
Type 2 diabetes mellitus | 0
oral hypoglycaemics | 0
non-smoker | 0
admitted to hospital | 0
SARS CoV-2 PCR positive | 0
CT chest scan | 0
patchy bilateral air-space infiltrates | 0
ground glass density | 0
transferred to ICU | 96
intubation | 96
lung-protective ventilation | 96
septic shock | 96
multi-organ dysfunction | 96
referred for ECMO | 120
oxygenation deteriorated | 120
metabolic derangements | 120
PEEP 20 cm of H2O | 120
P/F ratio 62 | 120
echocardiography | 120
normal left ventricular systolic function | 120
mild right ventricular systolic dysfunction | 120
mild RV dilatation | 120
mild to moderate tricuspid regurgitation | 120
RESP score 1 | 120
predicted survival 57% | 120
commence VV ECMO | 240
cannulation | 240
femoral-femoral approach | 240
21F return cannula | 240
23F drainage cannula | 240
ventilation reduced | 240
tidal volume 2ml/kg | 240
PEEP 10 cmH2O | 240
respiratory rate 10 bpm | 240
thrombus in right atrium | 240
improvement in haemodynamic | 240
RV function | 240
inability to mechanically ventilate | 336
complete loss of tidal volumes | 336
ECMO dependent | 336
HRCT | 480
minimal amount of potentially recruitable lung | 480
extensive consolidation and collapse of lungs | 480
prone ventilation | 648
airway bleeding | 552
complete proximal airway occlusion | 552
anticoagulated with heparin | 552
coagulation profile | 552
mild heparinization | 552
Activated Partial Thromboplastin Time | 552
airway bleeding treated | 552
nebulised tranexamic acid | 552
cessation of heparin | 552
bronchoscopic removal of thrombus | 552
fibrous tissue strands | 552
cryotherapy | 552
direct injection of tranexamic acid | 552
epinephrine | 552
cytology of bronchial tissue | 552
bronchial cells | 552
lung isolation | 552
bronchial blocker | 552
double-lumen endotracheal tube | 552
repeat bronchoscopy | 624
ongoing bleeding | 624
sloughing of bronchial mucosa | 624
Argon plasma coagulation | 624
fibrin debris | 624
main stem bronchi | 624
prone ventilation continued | 648
improvement in aeration of lung fields | 648
ECMO circuit change out | 888
elevated D-dimer | 888
haemolysis | 888
oxygenator change out | 936
hypercalcaemia | 768
high calcium levels | 768
parathyroid hormone levels | 768
serum phosphate | 768
1,25-dihydroxy vitamin D | 768
thyroid hormone levels | 768
pamidronate disodium | 792
calcitonin | 792
normalisation of calcium levels | 1080
trials of weaning ECMO | 960
decreased ECMO gas flow | 960
stable gas exchange | 960
decannulation | 1224
removal of ECMO cannulas | 1224
open repair of femoral veins | 1224
surgical tracheostomy | 1320
weaned off ventilator support | 1320
phonate via insufflation of oxygen | 1320
awake | 1440
obeying commands | 1440
actively participating in rehabilitation | 1440
interacting with family | 1440