75 years old | 0
male | 0
admitted to the hospital | 0
fever | -168
chills | -168
dizziness | -168
remission after fever | -168
headache | -168
abdominal pain | -168
diarrhea | -168
sputum | -168
nasal congestion | -168
runny nose | -168
hypertension | -672
physical examination | 0
temperature 39.0 °C | 0
heart rate 98 bpm | 0
respiratory rate 20 breaths per minute | 0
blood pressure 139/75 mmHg | 0
oxygen saturation in room air 98% | 0
clear breath sounds in both lungs | 0
uniform heart rhythm | 0
negative neurological tests | 0
white blood cell count 7.1 × 10^9/L | 0
neutrophils 58.6% | 0
monocytes 24.4% | 0
hemoglobin 83 g/L | 0
C-reactive protein (CRP) 111.20 mg/L | 0
cell factor interleukin (IL)-6: 279.22 pg/mL | 0
cell factor IL-10 3653.30 pg/mL | 0
plasma procalcitonin 0.19 ng/mL | 0
blood amyloid A 509.5 mg/L | 0
erythrocyte sedimentation rate 71 mm/L | 0
lactate dehydrogenase 694 U/L | 0
creatine kinase 19 U/L | 0
albumin 27 g/L | 0
K+ 2.99 mmol/L | 0
Na+ 135.1 mmol/L | 0
Cl- 98.5 mmol/L | 0
calcium 1.87 mmol/L | 0
phosphorus 0.65 mmol/L | 0
normal creatinine level | 0
anti-nuclear antibody, titer 1:100 | 0
anti-SSA- | 0
anti-SCL70 | 0
TORCH test (Toxoplasma, rubella, cytomegalo, and herpes viruses) normal | 0
Plasmodium test normal | 0
fungal D-glucan test normal | 0
coronavirus disease 2019 normal | 0
hematologic fever IgM antibody normal | 0
Widder test normal | 0
Weil Felix reaction normal | 0
bilateral blood culture test results suggested the occurrence of "L. monocytogenes" | 0
cerebrospinal fluid nucleated cell count 420 × 10^6/L | 0
cerebrospinal fluid lymphocyte 75% | 0
cerebrospinal fluid lactate dehydrogenase 472 U/L | 0
cerebrospinal fluid total protein 261.3 mg/dL | 0
cerebrospinal fluid glucose 1.51 mmol/L | 0
cerebrospinal fluid chloride content (Cl-) 111.0 mmol/l | 0
cerebrospinal fluid adenosine deaminase 16 U/L | 0
cerebrospinal fluid cryptococcal smear and cryptococcal capsular antigen test negative | 0
cerebrospinal fluid culture negative | 0
cerebrospinal fluid metagenomic test results indicated the presence of "G+ bacteria, L. monocytogenes" | 0
chest computed tomography (CT) results of the patient revealed a small amount of effusion in the pleural cavities on both the sides | 0
nodules were distinctly visible in the pleura and under the pleura | 0
cranial computed tomography no obvious abnormalities | 0
chest CT of the patient’s after two weeks treatment displayed multiple nodules in both lungs | 24
scattered patchy shadows in both the lungs | 24
possible infection | 24
small amount of pleural effusion in both lungs | 24
cranial MR plain scan + water suppression + diffusion-weighted diffusion weighted imaging showed abnormal signals scattered in the sub-frontal cortex, midbrain, and posterior horns of both the sides of the ventricle | 24
lacunar foci were found to be scattered under the frontal cortex on both the sides | 24
transparent interstitial space was formed | 24
sepsis | 0
lung infection | 0
respiratory failure | 0
electrolyte imbalance: hyponatremia, hypokalemia | 0
autoimmune disease | 0
Listeria monocytic meningoencephalitis | 0
levofloxacin 0.5 g qd intravenously | 72
body temperature did not drop significantly | 72
highest body temperature was still observed to be above 39.0 °C | 72
blood culture indicated the presence of a penicillin-resistant "Staphylococcus capital subspecies" | 72
Vancomycin injection 500000 U q6h | 96
intravenous infusion for anti-infection treatment | 96
body temperature reached the normal levels | 96
Vancomycin was used for 6 d | 168
body temperature was maintained at the normal level for more than 3 d | 168
discharged from the hospital | 168
high fever again | 168
maximum body temperature of 39.7 °C | 168
chills | 168
cough | 168
sputum | 168
thick and difficult to cough up | 168
no discomfort noted such as chest pain | 168
no limb twitching | 168
pupils were sluggish in the light reflection | 168
appeared confused | 168
mentally soft | 168
could only communicate briefly | 168
muscle strength test could not cooperate | 168
voluntary activities were seen | 168
diarrhea | 168
hospitalized in the emergency intensive care unit (ICU) | 168
high-frequency oxygen inhalation | 168
anti-infective and anti-inflammatory treatment of piperacillin and tazobactam 4.5 g q8h intravenously | 168
40 mg methylprednisolone injection | 168
repeated fever | 168
body temperature was above 38.3 °C | 168
considering that atypical bacterial infections were not covered | 168
intravenous infusion of levofloxacin 0.5 g qd as an anti-infective treatment | 168
body temperature returned to normal | 168
consciousness became clear | 168
CRP dropped to 76.4 mmol/L | 168
transferred to the general ward of the Department of Respiratory Medicine for further treatment | 168
atrial fibrillation occurred suddenly | 168
unresponsiveness | 168
slurred speech | 168
shortness of breath under nasal cannula oxygen inhalation | 168
slow light reflexes | 168
stiff neck | 168
increased muscle tone | 168
wet rales in both lungs | 168
critically severe | 168
repeated fever with the body temperature fluctuating around 38.7 °C | 168
sudden blood pressure drops | 168
signs of septic shock | 168
active rehydration | 168
norepinephrine micropump was used to maintain blood pressure | 168
antibiotics were adjusted to 1 million units of vancomycin injection q12h combined with meropenem injection 1.0 g q8h | 168
bacterial encephalitis | 168
meropenem injection 1.0 g q8h | 168
trachea was observed to be intubated | 168
breathing was assisted by a ventilator | 168
condition continued to deteriorate rapidly | 168
symptoms of repeated high fever, septic shock, and multiple organ failure | 168
gradual decrease in consciousness | 168
active fluid resuscitation | 168
administered norepinephrine injection to maintain the blood pressure | 168
tracheal intubation combined with ventilator-assisted ventilation | 168
condition did not improve significantly | 168
family decided to discontinue the further treatment | 168