81 years old | 0
    male | 0
    multiple comorbidities | 0
    presented with large left pleural effusion | 0
    fever | -504
    progressive dyspnea | -504
    dry cough | -504
    left pleuritic chest pain | -504
    chronic lymphocytic leukemia | 0
    treated with Fludarabine | 0
    treated with Cyclophosphamide | 0
    treated with Rituximab | 0
    type 2 diabetes mellitus | 0
    hypertension | 0
    hyperlipidemia | 0
    chronic kidney failure | 0
    eGFR of 28 mL/min/1.73 m2 | 0
    no smoking | 0
    no alcohol abuse | 0
    fever (38.1°C) | 0
    tachycardia (105 bpm) | 0
    peripheral percutaneous oxygen saturation 100% | 0
    tachypnea | 0
    normal blood pressure | 0
    abolished left vesicular murmur | 0
    adenopathy not observed | 0
    hepatomegaly not observed | 0
    splenomegaly not observed | 0
    cardiovascular examination normal | 0
    neurologic examination normal | 0
    neutrophilia (18.7 g/L) | 0
    elevated CRP (297 mg/L) | 0
    stable lymphocytosis (242 g/L) | 0
    anemia (7.8 g/L) |; 0
    chest X-ray showed large left pleural effusion | 0
    computed tomography confirmed multiloculated left pleural effusion | 0
    first bedside pleural puncture showed citrine exudate | 0
    pleural protein 37 g/L | 0
    pleural fluid protein to serum ratio 0.61 | 0
    intravenous cefotaxime | 0
    persistence of fever | 0
    persistence of neutrophilia | 0
    severe hypoxemia | 0
    bacteriological standard culture negative | 0
    blood cultures negative | 0
    auramine stained sputum smears negative | 0
    mycobacterial cultures negative | 0
    surgical thoracentesis | 240
    evacuation of 2 liters purulent liquid | 240
    pleura thick and nodular | 240
    white pseudo-membranes | 240
    metronidazole added to cefotaxime | 240
    cytobacteriological examination negative | 240
    lymphocyte phenotyping ruled out B-cell lymphoma | 240
    multiple organ failure | 264
    intensive care unit admission | 264
    septic shock | 264
    multiple organ failure | 264
    mechanical ventilation | 264
    vasopressor infusion | 264
    renal replacement therapy | 264
    death | 288
    Gram-negative bacilli isolated from pleural culture | 288
    L. pneumophila serogroup 1 identified | 288
    urinary antigen confirmed L. pneumophila serogroup 1 | 288
    fatal pleural empyema | 288
    Legionella pneumophila resistant to all antibiotics | 288
