64 years old | 0
male | 0
Caucasian | 0
admitted to the hospital | 0
diagnosis of Fournier's gangrene | 0
septic shock | 0
hypertension | -672
mild chronic renal insufficiency | -672
diabetes mellitus type 2 | -672
oral hypoglycaemic agents | -672
progressive respiratory deterioration | -24
hemodynamic instability | -24
intensive care unit | 0
multidisciplinary approach | 0
intensivist | 0
endocrinologist | 0
urologist | 0
reconstructive surgeon | 0
hemodynamic stabilization | 0
broad-spectrum antibiotic therapy | 0
first surgical debridement | 0
temporary diverting colostomy | 0
second radical debridement | 48
suprapubic cystostomy | 48
negative pressure wound therapy | 48
polyurethane foams | 48
stapled into the wound | 48
continuous negative pressure | 48
125 mmHg | 48
daily hyperbaric oxygen therapy | 48
2.4 atmospheres absolute | 48
90 min | 48
blood culture results | 72
methicillin-resistant Staphylococcus epidermidis | 72
wound cultures | 72
Proteus mirabilis | 72
Enterococcus faecalis | 72
no signs of deep wound infection | 168
NPWT dressing changed | 168
reapplied | 168
healthy granulation tissue | 504
no sign of infection | 504
skin and soft-tissue defects | 504
primary delayed closure | 504
scrotal advancement flaps | 504
Integra dermal regeneration template | 504
temporary cover | 504
full-thickness skin defects | 504
perineum | 504
right ischial region | 504
posterior part of the scrotum | 504
NPWT re-applied | 504
dermal regenerative template | 504
bolster dressing | 504
complete contact | 504
wound bed | 504
NPWT dressing changed | 504
dermal regenerative template inspected | 504
no complications | 504
outer silicone layer removed | 720
neodermis | 720
split-thickness skin graft | 720
right inner thigh | 720
NPWT | 720
bolster dressing | 720
complete healing | 1104
discharged from the hospital | 1104
no major complications | 1104
fully recovered | 2196
satisfying functional and aesthetic result | 2196