39 years old | 0
male | 0
nursing home employee | 0
non-smoker | 0
denies use of alcohol | 0
denies use of illicit drugs | 0
admitted to the hospital | 0
skin flare-up | -168
tenderness in the right upper limb | -168
visible scratches on the proximal right upper arm | -168
sore throat | -96
fever | -96
temperature 37.7 °C | 0
heart rate 133 bpm | 0
blood pressure 72/56 mmHg | 0
30 breaths/min | 0
oxygen saturation 99% | 0
erythema of the right upper arm | 0
swelling of the right upper arm | 0
pain in the right upper arm | 0
no paralysis of the right hand | 0
no contracture of the right hand | 0
white blood cell count 2.85×10^3/μL | 0
neutrophils 95.7% | 0
hemoglobin 12.2 g/dL | 0
platelet 9.3×10^4/μL | 0
C-reactive protein 45.36 mg/dL | 0
total protein 4.9 g/dL | 0
albumin 2.2 g/dL | 0
aspartate aminotransferase 210 U/L | 0
alanine aminotransferase 156 U/L | 0
total bilirubin 1.7 mg/dL | 0
creatine kinase 709 U/L | 0
blood urea nitrogen 61 mg/dL | 0
creatinine 4.9 mg/dL | 0
sodium 129 mEq/L | 0
potassium 3.8 mEq/L | 0
chloride 89 mEq/L | 0
glucose 108 mg/dL | 0
presepsin 2146 pg/mL | 0
prothrombin time-International normalized ratio 1.32 | 0
fibrinogen 760.0 mg/dL | 0
antithrombin 3 52.7% | 0
CT scan | 0
change in CT value in the triceps brachii muscle | 0
change in CT value in the latissimus dorsi muscle | 0
LRINEC score 9 | 0
shock | 0
tachypneic state | 0
noradrenaline infusion | 0
vasopressin infusion | 0
broad-spectrum antimicrobial agents | 0
trachea intubated | 0
ventilatory assistance | 0
emergency surgery | 0
incision in the dorsal side of the triceps brachii | 0
extensive excision of the fascia | 0
contamination with pus | 0
Streptococcus pyogenes in blood cultures | 96
Streptococcus pyogenes in intraoperative drainage cultures | 96
flare of the right precordia exacerbated | 96
incision from the precordia to the medial elbow | 96
debridement of contaminated tissues | 96
nerves and vessels marked with vessel tapes | 96
fasciotomy | 120
fasciotomy | 144
transfer from intensive care unit to ward | 168
ampicillin administration | 216
clindamycin administration | 216
wounds cleaned daily | 216
wounds remained open | 216
Klebsiella aerogenes in wound cultures | 360
cefepime administration | 360
thorough debridement | 456
nerves and vessels identified by vessel tapes | 456
wound closed with full-thickness skin graft | 1080
discharged | 1944
cefepime administration until hospitalization day 36 | 864
minocycline administration | 1296
no symptoms of nerve injuries | 8760
active shoulder range of motion | 8760
active elbow range of motion | 8760
active forearm range of motion | 8760
hypertrophic scar contracture at the right axilla | 8760