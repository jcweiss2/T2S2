53 years old | 0
male | 0
admitted to the hospital | 0
diarrhea | -504
hematochezia | -504
weight loss | -504
abdominal pain | -504
petechial rash | -14
nausea | -14
vomiting | -14
dyspnea | -14
rash | -14
colonoscopy | -336
biopsies | -336
edematous mucosa | -336
friable mucosa | -336
acute inflammation | -336
chronic inflammation | -336
Crohn disease | -336
discharged from hospital | -336
worsening symptoms | -14
admitted to emergency department | 0
hypotension | 0
tachycardia | 0
anemia | 0
low calcium | 0
elevated BUN | 0
low albumin | 0
high stool lactoferrin | 0
high pro-BNP | 0
folate deficiency | 0
thiamine deficiency | 0
proteinuria | 0
hyaline casts | 0
coarse granular casts | 0
pericardial effusion | 0
pleural effusions | 0
moderate wall thickening of small bowel loops | 0
moderate wall thickening of colon | 0
enterocolitis | 0
fat pad biopsy | 24
amyloidosis | 24
Congo red staining | 24
apple green birefringence | 24
esophagogastroduodenoscopy | 24
colonoscopy | 24
biopsies | 24
petechial lesions | 24
friable mucosa | 24
elevated immunoglobulin G | 24
low immunoglobulin A | 24
elevated kappa | 24
low lambda | 24
kappa/lambda ratio | 24
M-spike | 24
IgG kappa monoclonal gammopathy | 24
elevated 24-h urine protein | 24
bone marrow biopsy | 48
kappa-restricted plasma cell neoplasm | 48
duplication of chromosome 1q | 48
gain of chromosomes 5, 9, 15 | 48
early rouleaux formation | 48
IV fluid resuscitation | 0
midodrine | 24
blood product transfusions | 24
electrolyte supplementation | 24
folate supplementation | 24
thiamine supplementation | 24
discharged from hospital | 168
worsening shortness of breath | 168
nausea | 168
vomiting | 168
diarrhea | 168
fatigue | 168
hypotension | 168
bacteremia | 168
septic shock | 168
cyclophosphamide | 168
bortezomib | 168
dexamethasone | 168
stabilized | 168
discharged from hospital | 336
outpatient follow-up | 336
new onset diarrhea | -504
intermittent hematochezia | -504
denies dyspnea | -504
denies weight loss | -504
denies fatigue | -504
denies rash | -504
vital signs stable | -504
elevated total protein | -504
referred for colonoscopy | -504
colonoscopy not completed | -504