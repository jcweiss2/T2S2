54 years old | 0
female | 0
admitted to emergency department | 0
urinary symptoms | -72
nausea | -72
diffuse abdominal pain | -72
type 2 diabetes mellitus | -78840
basal insulin 20 IU per day | -78840
home-based capillary blood glucose monitoring | -78840
denied follow-up appointments | -78840
denied prior hospitalizations | -78840
recurrent UTI | -2928
empirical antibiotics | -2928
fatigue | -72
increased urinary frequency | -72
urgency | -72
acute urinary retention | -72
Foley catheter placement | -72
diuresis | -72
non-specific management | -72
fever 39 °C | -48
vomiting | -48
blood pressure 58/36 mmHg | 0
pulse 77 bpm | 0
respiration rate 26 bpm | 0
body temperature 36 °C | 0
oxygen saturation 92% | 0
capillary blood glucose 337 mg/dL | 0
altered mental status | 0
Glasgow Coma Scale 12 | 0
capillary refill 3 s | 0
normal lung examination | 0
abdomen without peritoneal irritation | 0
vesical globus | 0
bilateral costovertebral angle tenderness | 0
Foley catheter placement | 0
hematuria | 0
IV fluids resuscitation | 0
vasopressor agents | 0
third-generation cephalosporins | 0
leukocytes 35.7 ×10³/uL | 0
neutrophils 33.4 ×10³/uL | 0
hemoglobin 11.7 g/dl | 0
platelets 138 ×10³/uL | 0
fibrinogen 981 mg/dL | 0
creatinine 4.3 mg/dL | 0
glucose 334 mg/dL | 0
urea 132 mg/dL | 0
corrected sodium 136 mEq/L | 0
potassium 5 mEq/L | 0
chloride 94 mEq/L | 0
serum osmolality 282 mOsm/L | 0
venous pH 7.31 | 0
venous PCO2 25 mmHg | 0
venous PO2 37 mmHg | 0
HCO3 12.37 mmol/L | 0
base excess -13.7 mmol/L | 0
leukocyte esterase positive | 0
nitrite test negative | 0
500 leukocytes per HPF | 0
ketones present | 0
urine culture positive for ESBL E. coli | 0
meropenem-sensitive | 0
levofloxacin-resistant | 0
non-contrast abdominal CT scan | 0
kidneys loss of anatomy | 0
gas in perirenal space | 0
gas extending through ureters and bladder | 0
pneumoperitoneum | 0
septic shock | 0
grade IV emphysematous pyelonephritis | 0
mild diabetic ketoacidosis | 0
stage 3 acute kidney injury | 0
wide spectrum carbapenem antibiotics | 0
fluid resuscitation | 0
IV insulin | 0
bilateral nephrectomy | 192
appendix removal | 192
necrosis >90% | 192
parenchymal abscesses | 192
renal vein and arteries septic thrombi | 192
acute appendicitis | 192
ICU admission | 192
CVVH renal replacement therapy | 192
death | 264
