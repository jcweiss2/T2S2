47 years old | 0
woman | 0
self-reported 11-year history of diabetes mellitus | -96288
nausea | -48
vomiting | -48
decreased oral intake | -48
back pain radiating to the neck | -48
throbbing headache | -24
levothyroxine | -336
subcutaneous long-acting insulin (glargine) | -336
topiramate | -336
canagliflozin | -336
initiated 2 weeks earlier | -336
post-thyroidectomy Graves' disease | -96288
cholecystectomy for multiple cholelithiasis | -96288
depression | -96288
fibromyalgia | -96288
hyperlipidemia | -96288
history of spinal fusion surgery | -96288
appeared volume depleted | 0
temperature 98.9°F | 0
blood pressure 118/76 mmHg | 0
regular heart rate of 91 bpm | 0
BMI 27.45 kg/m² | 0
dry mucosal membranes | 0
absence of axillary sweat | 0
mild epigastric tenderness | 0
glucose 152 mg/dL | 0
sodium 138 mEq/L | 0
potassium 4.4 mEq/L | 0
chloride 105 mEq/L | 0
total carbon dioxide 16 mEq/L | 0
anion gap 17 | 0
serum blood urea nitrogen 16 mg/dL | 0
creatinine 0.76 mg/dL | 0
arterial blood gas revealed mixed acid-base disorder | 0
anion gap metabolic acidosis | 0
non-anion gap metabolic acidosis | 0
primary respiratory acidosis | 0
pH 7.18 | 0
PCO2 47.6 mmHg | 0
bicarbonate 17 mEq/L | 0
urinalysis pH 5 | 0
2+ ketones | 0
3+ glucose | 0
unremarkable thyroid function tests | 0
unremarkable liver function tests | 0
serum lactic acid level 1 mEq/L | 0
nondiagnostic urine drug screen | 0
nondiagnostic serum drug screen | 0
withholding insulin | 0
discontinuing canagliflozin | 0
initiating intravenous volume expansion with 5 L 0.9% saline | 0
unremarkable cultures | 0
unremarkable spine MRI | 0
unremarkable lumbar puncture | 0
poor oral intake | 0
nausea partially responded to ondansetron | 0
vomiting partially responded to ondansetron | 0
serum glucose <200 mg/dL | 0
insulin not administered | 0
serum bicarbonate fell to 10 mEq/L | 0
transferred to medical intensive care unit | 0
presumed acidemia | 0
repeat arterial blood gas performed 12 hours after admission | 12
pH 7.05 | 12
PCO2 26.9 mmHg | 12
bicarbonate fell to 7 mEq/L | 12
total serum carbon dioxide content 5 mEq/L | 12
blood glucose 107 mg/dL | 12
progressive acidosis | 12
isotonic bicarbonate (150 mEq/L) in 5% dextrose initiated | 12
rate 150 mL/hour | 12
ingested soft diet | 12
blood glucose increased to 200-300 mg/dL | 12
presumptive diagnosis of atypical DKA | 12
IV infusion regular insulin 2 units/hour initiated | 12
serum bicarbonate normalized | 24
anion gap normalized | 24
regular diet resumed | 24
nausea resolved | 24
vomiting resolved | 24
abdominal discomfort resolved | 24
previously managed for type 2 diabetes | -96288
undetectable C-peptide level | 24
latent autoimmune diabetes in adults (LADA) | 24
euglycemic DKA caused by SGLT2 inhibitor | 24
optimal management of euglycemic DKA | 24
SGLT2 inhibitor-associated side effects | 24
FDA black box warning | 24
canagliflozin discontinued | 0
insulin withheld for 24 hours | -24
low insulin levels | -24
increased ketogenesis | -24
dramatic drop in systemic pH | -24
SGLT2 inhibitor-mediated glycosuria | -24
volume depletion-mediated fall in glomerular filtration rate | -24
continued ketoacidosis | -24
dramatic fall in serum bicarbonate | -24
calculated total base deficit 524 mEq | 24
exogenous bicarbonate delivered 300 mEq | 24
catabolism of circulating ketoacids | 24
improved acid-base status | 24
ketoacid production fell | 24
dextrose administration | 12
insulin administration | 12
progressive acidemia | 12
euglycemia | 12
sepsis excluded | 0
lactic acidosis excluded | 0
non-anion gap component explored | 0
topiramate-induced renal tubular acidosis considered | 0
prolonged excretion of ketoacids | 0
absence of other causes | 0
marked anion gap acidosis | 0
sporadic reports of SGLT2 inhibitor-associated DKA | 0
euglycemic DKA in type 2 diabetes | 0
onset of diabetes at age 37 | -96288
undetectable C-peptide consistent with LADA | 24
increased risk of ketoacidosis in type 1 diabetes | 24
FDA concern about SGLT2 inhibitors in type 1 diabetes | 24
effects of SGLT2 inhibitors on pancreatic islet cells | 24
delayed recognition | 24
life-threatening complications | 24
clinical pearls | 24
duality of interest | 24
