60 years old | 0
woman | 0
admitted to the emergency unit | 0
pain | -48
paresthesia | -48
coolness of the right lower leg and foot | -48
cesarean section | -48
no previous thromboembolic events | -48
cold toes | 0
capillary filling lasting more than 5 seconds | 0
absent distal pulses in both legs | 0
computed tomography angiography | 0
floating thrombus in the abdominal aorta | 0
minimal marginal flow | 0
iliac arteries with marginal atherosclerotic plaques | 0
thromboembolism of the entire right deep femoral artery | 0
thromboembolism of the left deep femoral artery | 0
sustained flow in superficial femoral arteries | 0
occluded third segment of the right popliteal artery | 0
thromboembolus spreading to the posterior tibial artery | 0
marginal recanalization | 0
surgical thromboembolectomy | 0
LMWH | 0
proton pump inhibitor | 0
analgesic therapy | 0
cefuroxime | 0
transfusions of deplasmatized red blood cells | 0
no fever | 0
no respiratory symptoms | 0
no typical COVID-19-associated symptoms | 0
positive PCR test for SARS-CoV-2 | 0
transferred to COVID-19 center | 0
amoxicillin | 24
clavulanic acid | 24
intravenous PPI | 24
subcutaneous LMWH | 24
asymptomatic SARS-CoV-2 infection | 24
recovery from surgical intervention | 24
homozygous MTHFR C677T gene mutation | 24
discharged | 336
rivaroxaban | 336
PPI | 336
admitted to intensive care unit due to acute liver injury | 2976
nausea | -672
jaundice | -24
denied hepatotoxic substances except rivaroxaban | 2976
no portal vein thrombosis | 2976
no Budd-Chiari Syndrome | 2976
no viral hepatitis | 2976
no autoimmune diseases | 2976
no metabolic diseases of the liver and biliary tract | 2976
MSCT of thorax, abdomen, and pelvis | 2976
post-COVID'19 changes in lungs | 2976
ground glass | 2976
perilobular fibrosis | 2976
normal liver hemodynamic parameters | 2976
no cirrhosis | 2976
fulminant liver failure | 2976
acute hepatocellular injury | 2976
DILI | 2976
negative COVID-19 test | 2976
grade 3 hepatic encephalopathy | 2976
transfer to National Transplant Center | 2976
rapidly progressive liver failure | 2976
hepatic coma | 2976
respiratory insufficiency | 2976
mechanical ventilation | 2976
intensive care measures | 2976
liver allocation | 2976
tonic-clonic seizures | 2976
diffuse brain edema | 2976
no brain hemorrhage | 2976
no brain ischemia | 2976
no neurological response | 2976
general condition deteriorated | 2976
death | 2976
no autopsy | 2976
