25 years old|0
female|0
pregnant|0
pre-existing heart disease|0
complete atrioventricular canal repair at 2 years of age|0
mitral regurgitation|0
left ventricular ejection fraction of 33%|0
mechanical mitral prosthesis implantation at 19 years of age|0
cardiac resynchronization therapy at 19 years of age|0
New York Heart Association Class III|0
unplanned pregnancy at 14th week of gestation|0
carvedilol 25 mg/day|0
furosemide 40 mg/day|0
warfarin with INR levels between 3.0 and 3.5|0
worsening heart failure until 30th week of gestation|0
hospitalized|0
non-invasive positive pressure ventilation|0
low-dose intravenous furosemide|0
morphine|0
carvedilol adjusted to 75 mg/day|0
improved clinical condition|0
sore throat|168
cough|168
SARS-CoV-2 positive test|168
temperature 36°C|168
blood pressure 115/75 mmHg|168
heart rate 85 b.p.m.|168
oxygen saturation 97%|168
decreased respiratory sounds in lung bases|168
systolic murmur along left sternal border|168
fever|192
myalgia|192
hypotension|192
referred to COVID-19 ICU|192
piperacillin and tazobactam|192
therapeutic unfractionated heparin|192
amiodarone|192
norepinephrine|192
dobutamine|192
acute foetal distress|192
emergency caesarean delivery at 32nd week of gestation|192
mechanical ventilation|192
multiple organ failure|192
septic shock|192
increased inflammatory biomarkers|192
increased prothrombotic biomarkers|192
worsening lung tomographic scan|192
sedation with midazolam|192
sedation with fentanyl|192
neuromuscular blockers with cisatracurium|192
lung-protective ventilation in volume control mode|192
PaO2/FiO2 167|192
FiO2 45%|192
positive end-expiratory pressure 8|192
PaO2/FiO2 240|192
furosemide|192
methylprednisolone|192
meropenem|192
fluconazole|192
polymyxin B|192
amikacin|192
daptomycin|192
clinical improvement|792
sustained haemodynamic parameters|792
sustained respiratory parameters|792
extubated|792
PaO2/FiO2 240|792
oxygen saturation 94% with 2 L/min nasal catheter|792
non-invasive ventilation with positive pressure|792
conscious|792
good clinical condition|792
acute respiratory failure|888
low cardiac output|888
major gastrointestinal bleeding|888
major airway bleeding|888
death|888
COVID-19 confirmed by necropsy|888
diffuse alveolar damage|888
viral cytopathic effects|888
small pulmonary thrombi in pulmonary capillaries|888
acute tubular necrosis|888
cerebral oedema|888
placental villous maturation appropriate for gestational age|888
increased syncytial knots|888
mild fibrin depositions|888
acute placental infarcts involving ~20% of villous tissue|888
no chronic histiocytic inter villositis|888
no deciduous acute inflammation|888
