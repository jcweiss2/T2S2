36 years old | 0
male | 0
chronic smoker | 0
alcoholic | 0
presented to the emergency ward | 0
blunt abdominal trauma | 0
resuscitation with fluids | 0
norepinephrine infusion | 0
exploratory laparotomy | 0
postoperative | 0
did not accept feeds orally | 0
did not accept feeds through nasogastric tube | 0
called for central venous access | 0
parenteral nutritional support | 0
no apparent external neck swelling | 0
no neurological deficit | 0
deranged coagulation study | 0
international normalized ratio 1.8 | 0
right IJV cannulation attempted | 0
aspirated blood during pilot puncture | 0
aspirated white purulent material | 0
abandoned IJV cannulation | 0
right subclavian vein cannulation attempted | 0
developed cough | 0
developed stridor | 0
developed increasing breathlessness | 0
intubated | 0
urgent chest X-ray | 0
chest X-ray ruled out pneumothorax | 0
transferred to Intensive Care Unit | 0
mechanical ventilation | 0
right subclavian CVC inserted | 0
aspirated material sent for acid-fast bacilli detection | 0
acid-fast bacilli positive | 0
Mycobacterium tuberculosis colonies cultured | 0
erythrocyte sedimentation rate 60 mm | 0
HIV ELISA positive | 0
CD4 count 180/μl | 0
miliary tuberculosis on chest X-ray | 0
CT neck showed retropharyngeal abscess | 0
destruction of C-5 and C-6 vertebral bodies | 0
cervical brace advised | 0
medicine consultation obtained | 0
pulmonary consultation obtained | 0
category I anti-tubercular therapy started | 0
cotrimoxazole prophylaxis | 0
antiretroviral drugs started | 168
tracheostomy performed | 0
