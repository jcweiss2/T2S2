65 years old | 0
male | 0
mixed race | 0
farmer | 0
admitted to the hospital | 0
cough | -72
greenish expectoration | -72
chest pain | -72
asthenia | -72
weight loss | -72
valvuloplasty | -2160
aortic valve replacement | -2160
Warfarin | -2160
Carvedilol | -2160
left anterior hemiblock | -2160
acute respiratory failure | 0
poor ventilatory mechanics | 0
inadequate management of secretions | 0
use of accessory muscles | 0
mixed acidosis | 0
orotracheal intubation | 0
invasive mechanical ventilation | 0
systolic blood pressure 104/54 mmHg | 0
partial oxygen saturation 80% | 0
respiratory rate 36 rpm | 0
heart rate 120 beats/min | 0
left pneumothorax | 0
thoracic drainage tube | 0
Propofol | 0
fentanyl | 0
IPPV mode | 0
tidal volume 460 ml | 0
inspiratory time 1 s | 0
flow 45 L/min | 0
positive end-expiratory pressure 5 cm of H2O | 0
respiratory rate 12-14 breaths/min | 0
fraction inspired oxygen 45% | 0
minute volume 7.3 L/min | 0
exhaled tidal volume 460 ml | 0
maximum airway pressure 29 cm of H2O | 0
plateau pressure 20 cm of H2O | 0
average pressure 10 cmH2O/L/s | 0
compliance 31.9 ml/cm of H2O | 0
arterial blood gas analysis | 0
pH 7.17 | 0
pCO2 35 mm/Hg | 0
PO2 62.8 mm/Hg | 0
HCO3 12.7 mmol/L | 0
Base excess 13.4 | 0
SO2 88.6% | 0
metabolic acidosis | 0
shock | 0
dehydration | 0
hemo-dynamic compromise | 0
tension pneumothorax | 0
central venous catheter | 0
nasogastric tube | 0
bladder catheter | 0
chest tube | 0
pneumonia | 0
tree-like infiltrate | 0
consolidations | 0
pleural effusion | 0
CT scan | 0
leukocytes 14 200 mm3 | 0
hemoglobin 8.9 g/dl | 0
hematocrit 28.9% | 0
mean corpuscular volume 77 fl/red cell | 0
mean concentration of hemoglobin 23.7 picograms/cell | 0
mean cell hemoglobin concentration 30.6 grams/deciliter | 0
red blood cell count 374 mm3 | 0
platelets 166 000 mm3 | 0
Monocytes 3.2% | 0
eosinophils 1.4% | 0
lymphocytes 3.9% | 0
neutrophils 91.3% | 0
basophils 0.2% | 0
glucose 114.3 mg/dl | 0
electrolytes | 0
sodium 141 meq/L | 0
potassium 3.2 meq/L | 0
chlorine 111 meq/L | 0
calcium 7.9 meq/L | 0
BUN 15 mg/dl | 0
creatinine 0.9 g/dl | 0
ampicillin/sulbactam | 0
clarithromycin | 0
rifampicin | 24
isoniazid | 24
pyrazinamide | 24
ethambutol | 24
bronchoscopy | 24
sharp pale palate mucosa | 24
erythematous stippling | 24
cavitary image | 24
bronchioloalveolar lavage | 24
bronchial brushing | 24
Pseudomonas aeruginosa | 28
Klebsiella pneumonia | 28
carbapenemases resistance mechanism | 28
KPC type enzyme | 28
Mycobacterium tuberculosis | 28
GeneXpert MTB/RIF System | 28
MALDI-TOF mass spectrometry | 28
Colistin | 120
nebulized amikacin | 120
new CT scan | 240
complete resolution of pneumothorax | 240
interstitial pattern | 240
left pulmonary cavern | 240
pleural effusion | 240
hemodynamic instability | 312
vasopressor | 312
inotropic support | 312
norepinephrine | 312
dobutamine | 312
atrial fibrillation | 312
rapid reverse ventricular response | 312
death | 312