23 years old | 0
female | 0
G2P1 | 0
BMI 23 | 0
admitted to the hospital | 0
labour pains | 0
fever symptoms denied | 0
shortness of breath denied | 0
cough denied | 0
sore throat denied | 0
expected delivery date | -48
afebrile | 0
temperature 37°C | 0
BP 138 mm Hg | 0
BP 89 mm Hg | 0
heart rate 103 beats/min | 0
external OS 2 cm | 0
premature rupture of membrane | 0
meconium-stained liquor | 0
fetal distress | 0
hemoglobin level 10.2gm% | 0
COVID Rapid Antigen Test positive | 0
mild cough | -168
Covishield vaccination not done | 0
emergency caesarean section | 0
healthy live born male neonate | 0
baby weighed 2.86 kg | 0
no evidence of vertical transmission | 0
RT PCR test not done | 0
baby transferred to nursery | 0
blood sent for matching | 0
1 unit of B+ blood transfused | 0
Postpartum Hemorrhage | 1
heavy vaginal bleeding | 1
atonicity of the uterus | 1
Injection carboprost | 1
tranexamic acid | 1
Inj methergine | 1
IV syntocinon | 1
per rectal misoprostol | 1
PPH persisted | 1
BP 106 mm Hg | 1
BP 64 mmHg | 1
respiratory rate 17 per min | 1
heart rate 120 beats per minute | 1
abdomen reopened | 2
uterus flabby | 2
devascularization | 2
B-lynch suture | 2
uterus partially contracted | 2
abdomen closed | 2
2 litres of blood lost | 2
3 units of B+ blood transfused | 2
oral feeding started | 16
respiratory distress | 48
O2 saturation 92% | 48
IV piperacillin/tazobactam | 48
IV metronidazole | 48
Inj pantoprazole | 48
Tab ivermectin | 48
Tab montelukast | 48
Tab cetirizine | 48
Inj ondansetron | 48
Tab zinc | 48
Tab vitamin C | 48
Capsules vitamin D | 48
Infusion paracetamol | 48
Tab paracetamol | 48
1 unit of blood transfused | 72
condition improved | 72
no tracheal intubation | 72
O2 saturation 96-98% | 72
abdominal stitches removed | 192
repeat blood report | 240
D-Dimer 9.78 mg/L | 48
C-Reactive Protein 129 mg/L | 48
WBC count 16200 /μL | 48
Haemoglobin 8.2 g/dL | 48
Interleukin 49.7 pg/mL | 48
Ferritin 224.1 ng/mL | 48
D-Dimer 3.31 mg/L | 240
C-Reactive Protein 11.6 mg/L | 240
WBC count 9300 /μL | 240
Haemoglobin 9.3 g/dL | 240
Interleukin 16.7 pg/mL | 240
Ferritin 171.6 ng/mL | 240
RT PCR negative | 336
discharged | 360