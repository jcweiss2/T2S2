45 years old | 0
man | 0
admitted to the intensive care unit | 0
fever | -1344
chills | -1344
malaise | -1344
pneumonia | -1344
prolonged fevers | -1344
Streptococcus viridans bacteremia | -1344
Mycoplasma bacteremia | -1344
intermittent fevers | -1344
30-pound weight loss | -1344
high fevers | 0
sepsis | 0
Staphylococcus capitis bacteremia | 0
freely mobile pedunculated vegetations within the thoracic aortic endograft | 0
right lower lobe consolidation | 0
collapse | 0
bilateral pleural effusions | 0
diffusely thickened native aortic wall | 0
foci of air between the graft and the native wall of the aorta | 0
open surgical explantation of the aortic endograft | 0
open surgical explantation of the left subclavian artery stent graft | 0
aortic débridement | 0
inline reconstruction with a rifampin antibiotic-soaked prefabricated Dacron graft | 0
focal abscess | 0
aortopulmonary fistula | 0
wedge resection of the left upper lobe | 0
hypothermic circulatory arrest | 0
excised infected native descending thoracic aorta | 0
Candida infection | 0
chylothorax | 0
total parenteral nutrition | 0
coil embolization | 0
Onyx glue obliteration of the thoracic duct | 0
discharged | 264
patent repair | 1440
no evidence of infection | 1440
