22 years old | 0
male | 0
Crohn's colitis | -17520
fistulectomy for complex perianal fistula | -17520
severe weight loss (25 kg during 2 years) | -17520
diarrhea | -17520
abdominal pain | -17520
recurrent perianal tenderness | -17520
mesalamine | 0
herbal medicine | 0
fistular openings | 0
subcutaneous abscess pockets | 0
severe tenderness on anus and buttock | 0
unable to maintain sitting or supine position | 0
limited social activity | 0
mild fever | 0
examination under anesthesia | 0
complicated anal fistulas | 0
perianal abscesses | 0
colonoscopy | 0
multiple and diffuse aphthous ulcerations | 0
contrast-enhanced computed tomography scan of abdomen | 0
multifocal inflammatory wall thickening | 0
thick-walled abscess pockets | 0
beaded appearance of subcutaneous small abscesses | 0
Crohn's disease activity index (CDAI) score 244 | 0
abscess drainage | 0
seton operation | 0
azathioprine (AZA) administration at 25 mg | 0
AZA dose increased to 50 mg | 336
revisit hospital | 336
high fever (39.2°C) | 336
myalgia | 336
leukocytes 180/μl | 336
segmented cells 6% | 336
hemoglobin 6.6 g/dl | 336
platelets 48,000/μl | 336
ESR 55 mm/h | 336
CRP 24.7 mg/l | 336
laboratory data within normal limits | 336
discontinuation of AZA | 336
suspected pancytopenia | 336
suspected septicemia | 336
administration of human recombinant granulocyte colony-stimulating factor | 336
broad-spectrum antibiotic therapy | 336
fever subsided | 336
cell count fully recovered | 336
Escherichia coli found on blood culture | 336
antibiotics sensitive | 336
thiopurine methyltransferase (TPMT) wild type (*1/*1) | 336
decreased frequency of bowel movements | 336
improved perianal pain | 336
improved oozing | 336
follow-up colonoscopy 3 months later | 2160
diffuse fibrotic scar | 2160
disappearance of multiple ulcerations | 2160
weight gain of 10 kg | 2160
regular follow-up | 2160
no clinical recurrence | 2160
CDAI score 114 | 2160
