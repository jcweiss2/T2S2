45 years old | 0
male | 0
South Asian | 0
farmer | 0
exposed to flood waters | -168
chest pain | 0
generalized myalgias | 0
fever | -168
flu-like symptoms | -168
resolved fever | -48
resolved flu-like symptoms | -48
nonsmoker | 0
denies alcohol use | 0
denies illicit substance use | 0
no pertinent travel history | 0
no pet history | 0
blood pressure 86/58 mm Hg | 0
heart rate 102 beats per minute | 0
pulse-oximetry 94% | 0
random blood glucose 184 mg/dL | 0
temperature 36.4 °C | 0
severely icteric | 0
S3 | 0
no murmurs | 0
decreased air entry | 0
scattered crackles bilaterally | 0
mildly distended abdomen | 0
nontender abdomen | 0
alert and oriented | 0
no neurological deficits | 0
mild pitting edema | 0
borderline cardiomegaly | 0
mild interstitial edema | 0
sinus rhythm | 0
no acute dynamic changes | 0
resuscitated with intravenous crystalloid infusion | 0
electrolytes repleted | 0
coronavirus rapid antigen test negative | 0
admitted to medical intensive care unit | 0
initiated on piperacillin-tazobactam | 0
initiated on tigecycline | 0
routine management bundle for severe sepsis | 0
excluded corticosteroid therapy | 0
respiratory failure | 24
severe hypoxemia | 24
commenced on high-flow noninvasive ventilation | 24
moderate global hypokinesis | 24
estimated ejection fraction 30-35% | 24
mild-moderate mitral regurgitation | 24
basilar bilateral air-space disease | 24
aspiration pneumonitis | 24
serologies positive for leptospirosis | 24
white cell count 19.6 | 0
hemoglobin 13.4 | 0
platelets 67 | 0
serum sodium 132 | 0
serum potassium 4.4 | 0
serum creatinine 4.3 | 0
blood urea nitrogen 81 | 0
serum calcium 9.2 | 0
serum magnesium 0.9 | 0
fasting blood sugar 84 | 0
alanine aminotransferase 73 | 0
aspartate aminotransferase 34 | 0
alkaline phosphatase 154 | 0
serum albumin 3.2 | 0
international normalized ratio 1.2 | 0
prothrombin time 14.6 | 0
activated partial thromboplastin time 34 | 0
total bilirubin 15.5 | 0
conjugated bilirubin 11.1 | 0
troponin I 1.2 | 0
creatine kinase 293 | 0
erythrocyte sedimentation rate 55 | 0
C-reactive protein 42 | 0
blood cultures negative | 0
urine culture negative | 0
human immunodeficiency virus enzyme-linked immunosorbent assay nonreactive | 0
QuantiFERON-TB GOLD negative | 0
Biofire Respiratory Panel negative | 0
COVID-19 test negative | 0
leptospirosis immunoglobulin M antibodies positive | 0
hepatitis B surface antigen negative | 0
hepatitis C IgM antibodies negative | 0
hepatitis C immunoglobulin G antibodies negative | 0
dengue IgM antibodies negative | 0
dengue IgG antibodies negative | 0
malaria thick and thin smears negative | 0
urine Legionella antigen negative | 0
atrial tachycardia | 24
atrial fibrillation | 24
ventricular tachycardia | 24
defibrillated | 24
initiated on amiodarone infusion | 24
septic shock | 48
cardiogenic shock | 48
multiorgan failure | 72
deteriorated | 72
succumbed to illness | 96
new-onset cardiomyopathy | 24
myocarditis | 24
Weil’s syndrome | 48
jaundice | 48
renal failure | 48
hepatic failure | 48
discharged | -1