43 years old | 0
female | 0
admitted to the hospital | 0
productive cough | -240
diarrhoea | -240
vomiting | -240
end-stage renal failure | -240
crescentic IgA nephropathy | -240
live related renal transplant in 1992 | -240
chronic transplant glomerulopathy | -240
tacrolimus | 0
mycophenolate mofetil | 0
sodium bicarbonate | 0
atenolol | 0
ramipril | 0
methoxy polyethylene glycol-epoetin beta (Mircera©) | 0
severe hyponatraemia | 0
serum sodium 102 mmol/L | 0
acute-on-chronic kidney injury | 0
bilateral consolidation | 0
no evidence of fluid overload | 0
septic screen negative | 0
antibiotics started | 0
transferred to intensive care unit (ICU) for CVVHD | 0
sodium concentration adjusted in dialysate fluid | 0
serum sodium correction ≤8 mmol/24 h | 0
Day 3 confusion | 72
agitated | 72
no signs of meningism | 72
intubated | 72
lumbar puncture | 72
CT brain | 72
cerebrospinal fluid unremarkable | 72
CT brain no encephalitis | 72
serum sodium 116 mmol/L | 72
condition stabilized rapidly | 72
sepsis | 72
high tacrolimus level 32 μg/L | 72
renal failure | 72
extubated | 96
regained normal cognitive function | 96
regained normal neurological function | 96
transferred to renal unit | 144
serum sodium 135 mmol/L | 144
dialysis dependent | 144
discharged | 240
no evidence of cerebral oedema | 72
no seizure activity | 72
rapid symptom resolution | 72
full neurological function | 96
