73 years old | 0
male | 0
acute on chronic COPD exacerbation | 0
Type 2 respiratory failure | 0
conventional noninvasive ventilation | 0
profound acidemia | 0
pH - 7.057 | 0
base excess - 7.5 | 0
PCO2 - 11.23 kPa | 0
PaO2 - 13.7 kPa | 0
FiO2 - 50% | 0
P: F ratio around 200 | 0
high inflammatory markers | 0
total leukocyte count (TLC) 26 × 10^9/L | 0
procalcitonin 11.2 mcg/L | 0
CRP 104 mg/L | 0
worsened renal functions | 0
oliguric | 0
appropriate antibiotics | 0
noradrenaline infusion | 0
mean arterial pressure target 70 mm Hg | 0
continuous veno8venous hemodiafiltration | 0
negative fluid balance 1.5 L | 0
hemodynamic monitoring | 0
pulse-induced contour cardiac output | 0
continued acidosis | 12
PaCO2 - 10.86 kPa | 12
failure to remove CO2 | 12
non-invasive ventilation | 12
bilateral clear chest on auscultation | 12
increased vasopressors requirements | 12
extracorporeal carbon dioxide removal (ECCO2R) instituted | 12
pump flow - 0.56 L/min | 12
sweep flow - 10 L/min | 12
sweep FiO2 - 1.0 | 12
CO2 removal 6-10 L sweep flow | 12
CO2 removal 75-100 ml/min | 12
activated partial thromboplastin time ratio 1.2-1.6 | 12
platelets monitored | 12
fibrinogen monitored | 12
Hb monitored | 12
sweep flows adjusted according to CO2 values | 12
heparin infusions avoided initially | 12
pH improved to 7.30 | 12
PaCO2 normalized to 6.5 kPa | 12
non-invasive ventilation continued | 12
bi-level positive airway pressure MODE | 12
Sats >90% | 12
pH >7.3 | 12
R/R <30 | 12
improved inflammatory markers | 12
TLC 16 × 10^9/L | 12
CRP 46 mg/L | 12
procalcitonin 0.9 mcg/L | 12
enteral nutrition continued | 12
continuous veno-venous hemodiafiltration turned off | 12
sepsis relapse | 240
acidotic | 240
worsened work of breathing | 240
sweep flows adjusted | 240
conventional ventilation not increased | 240
no increased sedation | 240
no increased paralyzing agents | 240
ECCO2R turned off after 20 days | 480
sweep flows gradually taken down | 480
minimal CO2 removal | 480
sweep flow 4 L/min | 480
CO2 removal 80 ml/min | 480
sweep flow 1 L/min | 480
CO2 removal 45 ml/min | 480
critical illness related weakness | 480
prolonged weaning | 480
rehabilitation by physiotherapy | 480
successfully decannulated | 480
discharged from ICU | 480
