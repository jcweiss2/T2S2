male | 0
infant | 0
born at 40 6/7 weeks | 0
vaginal delivery | 0
hyperemesis gravidarum | -280
prenatal labs unremarkable | -280
ultrasound unremarkable | -280
no family history of inborn errors of metabolism | 0
newborn screen collected | 24
tachypnea | 72
tachypnea resolved | 72
discharged home | 96
difficulty establishing breast feeding | 96
fever | 120
poor feeding | 120
dehydration | 120
admitted to intensive care unit | 120
rehydration | 120
sepsis evaluation | 120
newborn screen returned | 125
elevated C14:1 | 125
elevated C14:2 | 125
elevated C14 | 125
elevated C14:1/C16 | 125
VLCADD suggested | 125
cardiac evaluations normal | 125
EKG normal | 125
echocardiogram normal | 125
infectious work-up completed | 125
antibiotic medication started | 125
antiviral medication started | 125
normal glucose concentrations | 76
elevated creatine kinase | 76
rhabdomyolysis | 76
elevated BUN | 76
elevated creatinine | 76
renal dysfunction | 76
mildly elevated liver function tests | 76
aggressive hydration started | 76
10% dextrose-containing fluids started | 76
medical food low in long chain fat started | 76
MCT supplementation started | 76
CK declined | 148
creatinine improved | 148
labs improved | 148
discharged | 456
good oral intake of medical formula | 456
initial plasma acylcarnitine concentrations highly indicative of VLCADD | 125
decreased with treatment | 148
molecular DNA testing for ACADVL | 125
two mutations c.848T>C and c.751A>G | 125
c.848T>C mutation pathogenic | 125
c.751A>G mutation not previously described | 125
normal growth and development | 1024
diet treatment continued | 1024
routine plasma acylcarnitines often elevated | 1024
l-Carnitine supplementation started | 532
hospitalizations for illness | 532
poor oral intake | 532
g-tube placement | 532
no further evidence of rhabdomyolysis | 1024