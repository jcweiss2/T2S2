15 years old | 0
female | 0
admitted to the hospital | 0
tuberculosis infection | -672
positive QuantiFERON gold test | -672
iron deficiency anemia | -672
hemoglobin 97–104 g/L | -672
systemic lupus erythematosus | -672
symmetric nonerosive polyarthritis | -672
nonscarring alopecia | -672
photosensitivity | -672
Raynaud phenomenon | -672
antinuclear antibodies positive | -672
anti-Smith antibodies positive | -672
anti-ribonucleoprotein antibodies positive | -672
naproxen | -672
hydroxychloroquine | -672
corticosteroids not taken for several years | -672
started treatment with rifampin | -264
rifampin 600 mg | -264
rifampin 10 mg/kg/d | -264
tolerated rifampin well for 11 days | -253
chills | -237
myalgias | -237
chills and myalgias began a few hours after rifampin ingestion | -237
chills and myalgias resolved a few hours later | -237
stopped treatment for 3 days | -228
in-person assessment | -213
normal physical examination | -213
arthritis in 2 joints | -213
advised to resume rifampin | -213
resumed rifampin | -212
severe neck pain | -212
myalgias | -212
arthralgias | -212
shortness of breath | -212
chest pain | -212
hypotension | -212
fluid bolus | -212
febrile | -212
tachypneic | -212
tachycardic | -212
low-to-normal blood pressure | -212
no angioedema | -212
no rash | -212
no wheezing | -212
no gastrointestinal symptoms | -212
intravenous fluids | -212
empiric vancomycin | -212
empiric ceftriaxone | -212
hypotensive again | -209
diaphoretic | -209
fluid resuscitation | -209
norepinephrine infusions | -209
epinephrine infusions | -209
admitted to the intensive care unit | -209
no rash or mucous membrane involvement | -209
decreased leukocyte count | -209
low eosinophil counts | -209
hemoglobin level decreased | -207
bilirubin levels normal | -207
haptoglobin levels normal | -207
direct antiglobulin test negative | -207
blood film did not show schistocytes | -207
inflammatory markers elevated | -207
C-reactive protein level increased | -207
aspartate aminotransferase level increased | -207
complement C3 level slightly decreased | -207
complement C4 level normal | -207
creatinine kinase level normal | -207
cortisol level increased | -207
computed tomography scan of the head normal | -207
echocardiogram normal | -207
CT angiography of the neck showed localized myositis | -207
chest radiograph showed mild pulmonary edema | -207
CT imaging of the lungs showed bilateral increased septal thickening with ground glass opacities | -207
infectious work-up negative | -207
SARS-CoV-2 negative | -207
received 1 dose of rifampin in the ICU | -204
decreased blood pressure | -204
vasopressor dose increased | -204
rifampin stopped | -198
weaned off vasopressors | -183
started isoniazid for TBI | -183
completed 9 months of therapy | -183
advised to avoid rifamycin-based medications | -183
discharged | 24