65 years old | 0
female | 0
admitted to the hospital | 0
recurrent fever | -744
nausea | -168
vomiting | -168
highest body temperature 38 ℃ | -744
neutrophil count 6.96×10^9/L ↑ | 0
monocyte count 0.86×10^9/L ↑ | 0
lymphocyte percentage 14.9% ↓ | 0
red blood cell count 3.17×10^12/L ↓ | 0
hemoglobin content 87 g/L ↓ | 0
hematocrit 0.28 L/L ↓ | 0
average red blood cell hemoglobin concentration 312 g/L ↓ | 0
platelet count 363×10^9/L ↑ | 0
platelet distribution width 8.3 fl ↓ | 0
C-reactive protein (CRP) 52.01 mg/L ↑ | 0
diagnosed with secondary infectious thrombocytopenia | 0
diagnosed with gram-negative bacilli septicemia (Klebsiella pneumoniae) | 0
diagnosed with liver abscess | 0
diagnosed with bilateral lung inflammation | 0
diagnosed with type 2 diabetes | 0
diagnosed with hypertension grade 3 (extremely high risk) | 0
given vancomycin | 0
given caspofungin | 0
given dexamethasone | 0
given posaconazole oral suspension | 0
liver abscess puncture and drainage treatment | 24
inflammatory indexes decreased | 48
light perception disappeared in the left eye | 72
eyelid redness and pain | 72
purulent secretion | 72
repeated fever | 72
left-sided headache | 72
diagnosed with endogenous endophthalmitis (left) | 72
diagnosed with orbital cellulitis (left) | 72
diagnosed with rubeosis iridis (left) | 72
diagnosed with exudative retinal detachment (left) | 72
diagnosed with diabetic retinopathy (right) | 72
intravitreal injection with vancomycin and ceftazidime | 96
symptoms relieved | 120
left eyeball enucleation | 216
fever again after the operation | 216
given moxifloxacin | 216
given sulperazon | 216
temperature elevated again | 240
CT examination | 240
inflammation of both lungs | 240
pericardial effusion | 240
bilateral pleural thickening and effusion | 240
atelectasis in right inferior lobe | 240
liver cyst | 240
liver abscess | 240
right renal cyst | 240
myoma of the uterus | 240
history of hypertension | -8760
highest blood pressure 180/100 mmHg | -8760
oral valsartan | -8760
controlled blood pressure at 140/80 mmHg | -8760
no special history of other systematic diseases | 0
no history of surgery | 0
no history of blood transfusion | 0
no history of drug allergy | 0
diagnosed with sepsis | 0
diagnosed with secondary thrombocytopenia | 0
diagnosed with liver abscess | 0
diagnosed with gram-negative bacilli sepsis (Klebsiella pneumoniae) | 0
diagnosed with infection of lumbar vertebrae | 0
diagnosed with mesenteric panniculitis | 0
diagnosed with pelvic effusion | 0
diagnosed with pericardial effusion | 0
diagnosed with suppurative endophthalmitis (left) | 0
diagnosed with orbital cellulitis (left) | 0
diagnosed with retinal detachment (left) | 0
diagnosed with choroidal detachment (left) | 0
diagnosed with type 2 diabetes retinopathy (right) | 0
diagnosed with cortical senile cataract (right, immature stage) | 0
diagnosed with type 2 diabetes | 0
diagnosed with type 2 diabetes nephropathy stage I | 0
diagnosed with type 2 diabetic peripheral neuropathy | 0
diagnosed with hypertension grade 3 (extremely high risk) | 0
diagnosed with hepatic cyst | 0
diagnosed with renal cyst | 0
diagnosed with hypoproteinemia | 0
diagnosed with coronary atherosclerotic heart disease | 0
diagnosed with lacunar cerebral infarction | 0
diagnosed with moderate anemia | 0
diagnosed with risk of malnutrition | 0
convulsion with unconsciousness | 288
transferred to the respiratory intensive care unit | 288
CT examination | 288
lacunar infarction | 288
encephalomalacia | 288
bilateral pleural effusion | 288
lower lobe of the right lung insufficiently inflated | 288
intracranial infection | 288
lumbar puncture | 288
cerebrospinal fluid (CSF) analysis | 288
microbial metagenomic next-generation sequencing (mNGS) | 288
biochemistry analysis | 288
glucose <1.1 mmol/L ↓ | 288
chlorine 108 mmol/L ↓ | 288
CSF protein >3,000 mg/L ↑ | 288
mNGS results | 288
high sequence of Klebsiella pneumoniae | 288
drug-resistant gene SHV-type beta-lactamases (blaSHV) | 288
given 2 g meropenem q8h prolonged for 3 hours | 288
body temperature improved | 312
blood routine improved | 312
CRP improved | 312
CT examination | 432
pulmonary edema and pleural effusion dissipated and absorbed | 432
CSF analyses | 456
chlorine 119 mmol/L ↓ | 456
micro amount of proteins 1,107 mg/L ↑ | 456
microalbumin 816.3 mg/L ↑ | 456
immunoglobulin G 308.5 mg/L ↑ | 456
α2-macroglobulin 18.5 mg/L ↑ | 456
β2-microglobulin 2.67 mg/L ↑ | 456
discharged from the hospital | 744