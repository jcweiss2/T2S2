52 years old | 0
male | 0
admitted to the hospital | 0
complaining of colicky upper abdominal pain | -168
nausea | -168
vomiting | -168
worsened in the last 2 days | -48
pneumonia | -10080
thoracic empyema | -10080
chronic pancreatitis | -10080
acute exacerbation | -8760
hypertension | 0
stage IV chronic renal disease | 0
tobacco smoker | 0
heavy drinker | 0
denied illicit drugs use | 0
not taking any antibiotics | 0
not taking any antiemetics | 0
not taking any painkillers | 0
critically ill | 0
emaciated | 0
dehydrated | 0
tachypneic | 0
tachycardic | 0
poor peripheral perfusion | 0
blood pressure was 70/50 mmHg | 0
room air oximetry was 88% | 0
Glasgow coma scale was 15 | 0
cardiac examination was unremarkable | 0
pulmonary examination was unremarkable | 0
abdomen was distended | 0
diffusely painful | 0
rebound tenderness | 0
normal bowel sounds | 0
mild anemia | 0
leukocytosis | 0
marked left shift | 0
acute renal failure | 0
metabolic acidosis | 0
increased hepatic enzymes | 0
normal amylase | 0
normal lipase | 0
normal bilirubin | 0
normal clotting tests | 0
peritonitis | 0
exploratory laparotomy | 0
free purulent effusion | 0
edema of the intestinal loops | 0
edema of the great omentum | 0
abscess in the retro-cavity of the epiplon | 0
peritoneal lavage | 0
abscess drainage | 0
closure of the abdominal wound with a Bogotá bag | 0
referred to the intensive care unit | 0
mechanical ventilatory support | 0
vasoactive drugs | 0
hemodynamic instability | 0
died | 24
culture obtained from the abdominal cavity was positive for Escherichia coli | 24
culture obtained from the abdominal cavity was positive for Group F β-hemolytic Streptococcus | 24
culture obtained from the abdominal cavity was positive for Raoultella planticola | 24
blood culture sets were positive for Group F β-hemolytic Streptococcus | 24
blood culture sets were positive for Raoultella planticola | 24
Bacterial identification was performed using VITEK-2 compact | 24
median xipho-pubic surgical incision | 24
Bogotá bag closure of the abdomen | 24
pleural adhesion in the left hemithorax | 24
sero-hemorrhagic effusion | 24
fibrinoid material | 24
pancreas weighed 183 g | 24
distorted shape | 24
surrounded by increased fat tissue | 24
effaced lobulation | 24
mousy color | 24
intermingled by white areas of a hardened consistency | 24
purplish 3 cm pseudocyst | 24
rupture of the external wall | 24
extensive fibrosis | 24
acinar atrophy | 24
intraductal eosinophilic protein plugs | 24
chronic inflammatory infiltration | 24
fibrin | 24
peritonitis | 24
acute inflammatory infiltration | 24
venules thrombosis | 24
granulation tissue | 24
lungs atelectasis | 24
respiratory bronchiolitis | 24
tracheal squamous metaplasia | 24
myocardial hypertrophy | 24
bone marrow hypercellularity | 24
myeloid hyperplasia | 24
loss of hepatocytes centrilobular trabeculation | 24
vacuolation | 24
acute tubular necrosis | 24
acute splenitis | 24