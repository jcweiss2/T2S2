46 years old | 0
male | 0
sickle cell disease | 0
abdominal pain | -24
acute cholecystitis | -24
LC | -24
discharged home | -24
worsening abdominal pain | 0
abnormal liver function studies | 0
common bile duct transection | 0
attempted ERCP | 0
aborted ERCP | 0
transferred to hospital | 0
severe respiratory distress | 0
sickle cell crisis | 0
sinus tachycardia | 0
heart rate 156 | 0
blood pressure 173/87 | 0
pulse oximetry 92% | 0
high flow nasal cannula | 0
transferred to ICU | 0
Hematology consulted | 0
total bilirubin 15.1 mg/dl | 0
creatinine 1.1 mg/dl | 0
AST 150 U/l | 0
ALT 434 U/l | 0
Alkaline phosphatase 175 U/l | 0
White blood cells 15.3 × 10^3/cm2 | 0
hematocrit 26% | 0
hemoglobin 9.1 g/dl | 0
platelets 216 × 10^3/cm2 | 0
INR 1.5 | 0
CT angiogram | 0
multifocal pneumonia | 0
free peritoneal fluid | 0
Chest CT | 0
no pulmonary embolism | 0
repeat ERCP | 0
wide-open distal common bile duct | 0
inability to pass a wire distally | 0
Interventional radiology consulted | 0
PTC | 0
completely transected duct | 0
wire traversed into distal ductal orifice | 0
taken to operating room | 0
open surgical repair | 0
over 2 l of bilious fluid | 0
bile peritonitis | 0
portal dissection | 0
exposed PTC catheter | 0
necrosed common bile duct | 0
resected common bile duct | 0
multiple surgical clips removed | 0
cystic artery identified | 0
right and left hepatic arteries preserved | 0
PTC catheter pulled | 0
distal common bile duct orifice closed | 0
Roux-en-Y hepaticojejunostomy | 0
drain placed | 0
abdomen closed | 0
transferred to ICU | 0
extubated | 24
oxygen desaturations | 24
Hemoglobin electrophoresis | 24
elevated HgbS and C | 24
red blood cell exchange transfusion | 24
goal hemoglobin S and C <30% | 24
discharged home | 192
total bilirubin 4.1 mg/dl | 192
normal transaminases | 192
stable hematocrit 30% | 192
normal renal function | 192
seen in clinic | 672
total bilirubin 1.0 mg/dl | 672
cholangiogram | 672
no evidence of leak or stricture | 672
cholangiogram catheter removed | 672
discharged from clinic | 672