14 years old | 0
female | 0
nausea | -72
vomiting | -72
abdominal pain | -72
admitted to the local clinic | -72
diagnosis of acute viral gastroenteritis | -72
hyperglycemia | -72
ketonuria | -72
transferred to emergency unit | 0
lethargic | 0
severely dehydrated | 0
drowsy | 0
tachycardia | 0
tachypnea | 0
hypothermia | 0
normal blood pressure | 0
weight loss | -168
body mass index | 0
chest x-rays showed no specific abnormalities | 0
abdominal x-rays showed no specific abnormalities | 0
metabolic acidosis | 0
hyperglycemia | 0
ketonemia | 0
ketonuria | 0
DKA | 0
type 1 diabetes | 0
C-peptide | 0
glycosylated hemoglobin | 0
antiglutamic acid decarboxylase | 0
anti-islet cell antibodies | 0
anti-insulin antibodies | 0
fluid replacement | 0
intravenous insulin infusion | 0
hourly neurological evaluations | 0
generalized tonic seizure | 4
bradycardia | 4
cardiopulmonary arrest | 4
external cardiac massage | 4
epinephrine injection | 4
return of spontaneous circulation | 10
metabolic acidosis | 10
hypophosphatemia | 10
phosphate replacement | 10
K2HPO4 | 10
KCl | 10
brain CT scan | 10
no brain edema | 10
no intracranial pathology | 10
dexamethasone | 10
mannitol | 10
intensive care unit | 10
stuporous | 16
shallow respiration | 16
weak respiration | 16
slow respiration | 16
endotracheal intubation | 16
respiratory acidosis | 16
severe hypophosphatemia | 16
phosphate replacement increased | 16
repeat brain CT imaging | 16
no specific findings | 16
electrolyte and pH values normalized | 48
mechanical ventilation | 48
phosphate replacement increased | 48
fluid replacement | 48
potassium replacement | 48
intravenous insulin administration | 48
stable vital signs | 72
self-respiration recovered | 72
arterial blood gas levels normalized | 72
plasma phosphate increased | 72
weaning from inotropic support | 72
weaning from ventilator support | 72
transferred to general ward | 96
oral feeding | 96
multiple subcutaneous insulin injections | 96
phosphate supplementation stopped | 96
electroencephalogram | 96
no epileptiform discharges | 96
no slow waves | 96
discharged | 240
no neurologic complications | 240
no respiratory problems | 240
no further phosphate supplementation | 240