31 years old | 0\
female | 0\
non-smoking | 0\
Caucasian | 0\
no past medical history | 0\
sudden-onset severe headache | -840\
left arm numbness | -840\
SAH | -840\
grade 2 SAH | -840\
ruptured right middle cerebral artery aneurysm | -840\
percutaneous endovascular coil embolization | -816\
fever | -672\
chills | -672\
constant abdominal pain | -672\
purulent uterine discharge | -672\
sepsis | -668\
septic shock | -668\
mild disorientation | -668\
slower capillary refill | -668\
coarse rales | -668\
SOFA score 4 | -668\
invasive blood pressure 90/65 mmHg | -668\
heart rate 135/min | -668\
arterial oxygen saturation 82 % | -668\
hemoglobin 6.8 g/dL | -668\
d-dimers 4.58 μg/mL | -668\
C-reactive protein 322 mg/L | -668\
fibrinogen concentration 6.4 mL | -668\
E. coli | -668\
pulmonary nodules | -668\
enlarged uterus | -668\
complete loss of zonal anatomy | -668\
splenic metastatic lesion | -668\
β-hCG 232,085 mUI/mL | -668\
suction evacuation and curettage | -664\
choriocarcinoma | -664\
FIGO score 12 | -664\
high risk GTN | -664\
multiagent chemotherapy | -660\
low-dose etoposide | -660\
cisplatin | -660\
EMA/CO regimen | -653\
grade 3 neutropenia | -647\
G-SCF | -647\
dose reduction of etoposide | -647\
dose reduction of actinomycin D | -647\
grade 2 alopecia | -647\
grade 2 nausea | -647\
dexamethasone | -647\
ondansetron | -647\
EP/EMA regimen | -640\
grade 2 fatigue | -640\
male condoms | -640\
β-hCG normalization | -610\
disease-free for 21 months | 504