38 years old | 0
male | 0
referred with 6 month history of warm, swollen, and painful right knee | -4320
warm right knee | -4320
swollen right knee | -4320
painful right knee | -4320
initial redness of right knee | -4320
redness resolved spontaneously | -4320
first symptoms occurred 10 weeks after car accident | -2400
car accident resulting in craniocerebral trauma | -2400
coma | -2400
intracranial hypertension | -2400
required temporary ventricular drainage | -2400
during ICU stay developed sepsis with Klebsiella Pneumoniae | -2400
sepsis with Pseudomonas Aeruginosa | -2400
period of multi-organ failure | -2400
swelling of right knee noticed at start of rehabilitation | -2400
no evidence of infection in synovial fluid | -2400
no knee trauma reported during car accident | -2400
no knee trauma during hospital stay | -2400
referred for further diagnosis | -4320
clinical examination at presentation revealed warm, swollen, painful right knee | 0
no redness at presentation | 0
no other joints involved | 0
normal body temperature | 0
normal remainder of clinical examination | 0
arthrocentesis of the knee showed WBC 57000 | 0
neutrophils 90% | 0
cultures negative | 0
mycobacterial culture negative | 0
no crystals in fluid | 0
elevated CRP 43 mg/L | 0
elevated blood WBC 11500/mm³ | 0
rheumatoid factor negative | 0
anti-CCP antibodies negative | 0
anti-nuclear factor negative | 0
Borellia antibodies negative | 0
Chlamydia Trachomatis PCR negative | 0
Neisseria Gonorrhoeae PCR negative | 0
MRI showed no major cartilage problems | 0
MRI showed no meniscal lesions | 0
MRI showed no ligamental lesions | 0
MRI showed bony infarctions in femur and tibia | 0
needle arthroscopy performed | 0
hyperemic synovium | 0
hypertrophic synovium | 0
synovium covered with white film | 0
synovial biopsies obtained | 0
inflammation in synovial tissue | 0
high amount of neutrophils in synovial tissue | 0
direct cultures of synovial tissue showed Staphylococcus Warneri | 0
Staphylococcus Warneri resistant to penicillin | 0
PCR for Borrelia negative | 0
PCR for mycobacteria genus negative | 0
PCR for mycobacterium complex negative | 0
treatment with Levofloxacin initiated for 6 weeks | 0
clinical evolution showed improvement | 432
persisting swelling of knee after 6 weeks | 432
repeated needle arthroscopy | 432
synovial biopsies showed decreased inflammatory infiltrate | 432
synovial fluid WBC 3810 | 432
synovial fluid neutrophils 38% | 432
CRP 66.2 at first arthroscopy | 0
CRP 26.2 after 6 weeks | 432
discharged | 432
staphylococcus warneri infection | 0
septic arthritis due to staphylococcus warneri | 0
indolent septic arthritis | 0
negative cultures of articular fluid | 0
delay in diagnosis | 0
cultures of synovial tissue obtained | 0
diagnosis established by synovial tissue culture | 0
no prosthetic device present | 0
possible entry of S. Warneri through catheter during ICU admission | -2400
low virulence of S. Warneri | 0
slow growth of S. Warneri | 0
negative blood cultures for S. Warneri | 0
culture of vegetation tags in prosthetic valve endocarditis | 0
