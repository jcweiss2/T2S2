55 years old | 0
perimenopausal female | 0
non-insulin dependent diabetes | 0
admitted to the hospital | 0
midline lower abdominal pain | -96
dysuria | -96
lower back pain | -96
nausea | -96
vomiting | -96
vaginal bleeding | -96
amenorrhea | -216
afebrile | 0
normotensive | 0
non-tachycardic | 0
lower abdominal tenderness | 0
uterus palpable at the level of the umbilicus | 0
normal external female genitalia | 0
enlarged uterus | 0
cervix displacing anteriorly | 0
no cervical motion tenderness | 0
cervix not visualized | 0
wet prep negative | 0
endometrial biopsy | 0
leukocytosis | 0
urinalysis with nitrites | 0
urinalysis with leukocytes | 0
urinalysis with blood | 0
transvaginal ultrasound | 0
uterine masses consistent with leiomyomata | 0
thickened endometrium | 0
echogenic endometrium | 0
lobulated areas of tissue | 0
ovaries not visualized | 0
differential diagnosis | 0
acute cystitis | 0
leiomyomata | 0
degenerating fibroids | 0
underlying malignancy | 0
pain improved with acetaminophen and ibuprofen | 0
treated for acute cystitis | 0
discharged home | 0
re-presented to the emergency room | 96
worsening suprapubic pain | 96
fevers | 96
chills | 96
nausea | 96
vomiting | 96
ongoing vaginal bleeding | 96
no malodorous discharge | 96
lower abdominal and suprapubic tenderness | 96
hypotensive | 96
leukocytosis | 96
elevated lactate | 96
CT of the abdomen and pelvis | 96
fibroid uterus | 96
pelvic free fluid | 96
expanded endometrial cavity | 96
hyperdensity within the mass | 96
sepsis due to urinary source | 96
evaluation for gynecologic source | 96
evaluation for gastrointestinal source | 96
crystalloid for fluid resuscitation | 96
norepinephrine for blood pressure support | 96
broad spectrum antibiotics | 96
admitted to the Medical Intensive Care Unit | 96
leukocytosis improved | 96
lactate improved | 96
persistently hypotensive | 96
mildly tachycardic | 96
afebrile | 96
serial physical and laboratory exams | 96
antibiotics continued | 96
clinical condition deteriorated | 105
worsening leukocytosis | 105
lactic acidosis | 105
increasing pressor support | 105
antibiotics broadened | 105
urine output | 105
distinct lower abdominal guarding | 105
decision to proceed to operating room | 105
exploratory laparotomy | 105
source control | 105
intrauterine source | 105
consented for exploratory laparotomy | 105
total abdominal hysterectomy | 105
bilateral salpingo-oophorectomy | 105
pressor support | 105
intraoperative findings | 105
enlarged uterus | 105
necrotic intrauterine mass | 105
foul-smelling intrauterine mass | 105
gross inspection | 105
no obvious myometrial invasion | 105
total abdominal hysterectomy | 105
bilateral salpingo-oophorectomy | 105
estimated blood loss | 105
abdomen and pelvis irrigated | 105
Blake drain placed | 105
fascia closed | 105
subcutaneous tissue irrigated | 105
sterile gauze packed | 105
pressor support decreased | 105
urine output increased | 105
extubated in the operating room | 105
transferred to Surgical Intensive Care Unit | 105
weaned off vasopressors | 120
blood cultures | 120
Clostridium species | 120
Bacteroides vulgatus | 120
antibiotics narrowed | 120
ampicillin-sulbactam | 120
clindamycin | 120
post-operative care | 120
transferred out of SICU | 192
meeting post-operative milestones | 192
maintained on IV antibiotics | 288
white blood cell count normalized | 288
discharged home | 288
wound-vac | 288
amoxicillin-clavulanate | 288
metronidazole | 288
surgical pathology | 288
pT1a carcinosarcoma | 288
myometrial invasion | 288
presented at multi-disciplinary tumor board | 288
adjuvant carboplatin | 288
paclitaxel | 288
vaginal brachytherapy | 288