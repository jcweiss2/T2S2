19 years old | 0
woman | 0
diagnosed with hydatidiform mole | 0
vaginal bleeding | -216
fresh blood | -216
clots | -216
vesicle-like tissue | -24
married | -35040
spontaneous full-term singleton birth | -17520
no significant complications | -17520
fourth antenatal visit | 0
midwife visits | -720
referred to obstetrician | -720
first ultrasound screening | -720
suspected molar pregnancy | -720
referred to hospital for curettage | -720
vital signs normal | 0
22- to 22-week-sized uterus | 0
speculum examination insignificant bleeding | 0
no mass infiltration | 0
anemia | 0
hemoglobin 8.1 g/dL | 0
hematocrit 23.8% | 0
leukocytes 9630/uL | 0
platelets 396000/µL | 0
β-hCG 1000×103 mIU/mL | 0
normal thyroid function | 0
triiodothyronine 1.6 mg/dL | 0
free T4 1.5 mg/dL | 0
decreased thyroid stimulating hormone | 0
chest X-ray no abnormalities | 0
ultrasound enlarged uterus | 0
uterine cavity vesicular appearance | 0
suspected molar pregnancy | 0
blood transfusion | 0
vacuum curettage | 0
hospital admission | 0
left labia minora mass | 120
mass 3×3×2 cm | 120
suspected hematoma | 120
vacuum curettage performed | 120
blood loss 3000 cc | 120
sharp curettage | 120
uterine mass removed | 120
conservative management | 120
pain in genital area | 124
conscious | 124
deteriorated vital signs | 124
shock | 124
blood pressure 90/60 mmHg | 124
pulse 130 bpm | 124
vulvar mass 6×5×4 cm | 124
perforation 0.5×0.5 cm | 124
active bleeding | 124
emergency evacuation | 124
hematoma incised | 124
blood clot evacuated | 124
vesicle-like tissue in mass | 124
fragile tissue bleeding | 124
bleeding controlled with sutures | 124
suspected stage II GTN | 124
histopathological examination | 124
chronic villi with cystic dilatation | 124
hydrophilic avascular degeneration | 124
cytotrophoblasts | 124
syncytiotrophoblasts | 124
excessive proliferation | 124
normal cell nuclei | 124
blood clot in decidua | 124
no malignant tumor cells | 124
complete mole with excessive proliferation | 124
reevaluation of histopathology | 124
partial hydatidiform mole in vagina | 124
embolism suspected | 124
partial hydatidiform mole in uterus | 124
p53 positive 20% | 124
transferred to ICU | 124
intubated | 124
oxygen saturation 80% | 124
condition never improved | 124
prolonged intubation | 124
hypoxia | 124
massive blood loss during surgery | 124
postoperative hemoglobin 2.3 g/dL | 124
hemoglobin increased to 9 g/dL | 124
bilateral pneumonia | 528
leukocytosis 18460/µL | 528
sepsis | 528
antibiotics | 528
pulmonary edema | 96
metabolic encephalopathy | 96
died due to sepsis | 528
