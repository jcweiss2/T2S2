33 years old | 0
female | 0
cesarean section | 0
term | 0
polyhydramnios | -672
nonconsanguineous marriage | 0
Zoladex implant | -1416
dysmorphic | 0
weighed 2.370 kg | 0
47 cm long | 0
microcephaly | 0
head circumference 29 cm | 0
severely deformed nose | 0
stenotic nostril | 0
cul-de-sac | 0
hypotelorism | 0
cleft palate | 0
microphthalmia | 0
micrognathia |&0
respiratory distress | 0
admitted to NICU | 0
septic workup | 0
severe respiratory distress | 4
endotracheal intubation | 4
CBC normal | 0
blood electrolytes normal | 0
blood gases normal | 0
chest X-Ray normal | 0
atrial septal defect | 0
patent ductus arteriosus | 0
kidneys normal | 0
lateral ventricle dilatation | 0
absent septum pellucidum | 0
holoprosencephaly | 0
fused cerebral hemisphere | 0
fused thalami | 0
mono-nostril | 0
lobar holoprosencephaly | 0
skeletal survey normal | 0
karyotype 46 XX | 0
feeding by orogastric tube | 72
gram-negative sepsis | 336
Pseudomonas aeruginosa | 336
DIC | 336
died | 336
