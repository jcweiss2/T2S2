22 years old | 0
    female | 0
    Malay ethnicity | 0
    presented to the haematology department | 0
    fever | -168
    left axillary swelling | -168
    no past medical history | 0
    no family history | 0
    non-smoker | 0
    does not consume alcohol | 0
    works as a bank clerk | 0
    pale | 0
    left axillary swelling of 5 x 5 cm | 0
    firm | 0
    non-tender | 0
    no discharge | 0
    no palpable lymph nodes | 0
    no organomegaly | 0
    normochromic normocytic anaemia | 0
    haemoglobin 5.5 g/dL | 0
    leucocytosis 22 x 10^9/L | 0
    thrombocytopenia 30 x 10^9/L | 0
    no coagulopathy | 0
    peripheral blood smear presence of blasts | 0
    abnormal promyelocytes | 0
    faggot cells | 0
    bone marrow aspirate presence of blasts | 0
    trephine biopsy hypercellular marrow | 0
    blast population expressing myeloperoxidase | 0
    lacking CD34 | 0
    lacking CD3 | 0
    marrow flow cytometry aberrant myeloid cells | 0
    CD117 | 0
    cMPO | 0
    CD13 | 0
    CD33 | 0
    CD38 | 0
    lacking CD34 | 0
    lacking HL-DR | 0
    PML-RAR-alpha fusion gene detected | 0
    left axillary swelling histology diffuse monomorphic infiltrates | 0
    neoplastic cells | 0
    fine nuclear chromatin | 0
    moderate rim of basophilic cytoplasm | 0
    immunohistochemistry positive for MPO | 0
    CD13 | 0
    CD33 | 0
    CD68 | 0
    CD117 | 0
    negative for CD34 | 0
    negative for HLA-DR | 0
    granulocytic sarcoma | 0
    diagnosed high-risk APML | 0
    Modified Sanz score 2017 | 0
    dexamethasone prophylaxis | 0
    differentiation syndrome prophylaxis | 0
    ATRA 45 mg/m2 daily | 0
    arsenic trioxide 0.15 mg/kg | 0
    idarubicin | 0
    culture-negative neutropenic sepsis | 14
    Type 1 respiratory failure | 14
    intubated | 14
    intensive care unit admission | 14
    no alveolar haemorrhage | 14
    diffuse nodular pulmonary infiltrations | 14
    no pulmonary embolism | 14
    serum galactomannan not detected | 14
    antimicrobial treatment | 14
    responded to antimicrobials | 14
    induction therapy | 0
    consolidation therapy | 0
    maintenance therapy | 0
    complete molecular remission | 720
    