36 years old | 0
female | 0
subarachnoid haemorrhage | -672
rupture of a right-sided middle cerebral artery aneurysm | -672
secondary vasospastic malignant infarction | -672
haemicraniectomy | -672
posthaemorrhagic cerebrospinal fluid circulatory dysfunction | -672
implantation of a ventriculoperitoneal shunt | -672
left-sided hemiparesis | -672
able to communicate on a basic level | -672
able to execute simple actions | -672
deterioration of condition | -336
unresponsive to external stimuli | -336
vegetative dysfunction | -336
vomiting | -336
extreme sweating | -336
tachypnoea | -336
tachycardia | -336
correction of suspected overdrainage of the ventriculoperitoneal shunt | -168
cranioplastic skull reconstruction | -168
unresponsive wakefulness syndrome | -168
weaning from respirator | -168
breathing spontaneously through a tracheal cannula | -168
infected decubiti | -168
upper limb phlegmon | -168
pneumothorax | -168
anaemia | -168
anovesical fistula | -168
multiple infections | -168
pneumonia | -168
urinary tract infection | -168
catheter-associated sepsis | -168
rhythmic myoclonus | -168
tremor | -168
levetiracetam | -168
valproic acid | -168
clonazepam | -168
no seizures | -168
no epileptic activity | -168
poor prognosis | -168
transfer to university hospital | 0
re-evaluation of prognosis and treatment options | 0
cranial CT | 0
MRI of the brain | 0
superficial siderosis | 0
laminar necrosis | 0
temporal, frontal and opercular atrophies | 0
widened ventricle of the right hemisphere | 0
PET with 18F-fluorodeoxyglucose | 0
normal glucose metabolism | 0
cerebral glucose metabolism | 0
focal neurological deficit | 0
global brain dysfunction | 0
tapering off oral baclofen | 0
intrathecal baclofen | 0
reduction and stop of levetiracetam, valproic acid and clonazepam | 0
lamotrigine | 0
no epileptiform activity | 0
amantadine | 0
improvement of consciousness | 16
improvement of tetraparesis | 16
improvement of myoclonus | 16
speaking valve | 16
speech apraxia | 16
retrograde amnesia | 16
full orientation | 16
ability to communicate | 16
ability to move all extremities | 16
reduced spasticity | 16
transfer to neurorehabilitation centre | 88
fully oriented patient | 88
mild cognitive deficits | 88
decanulation | 88
eating autonomously | 88
standing with help | 88
walking with difficulty | 88