32 years old|0
obese|0
male|0
Turkish|0
lymphoma with plasmablastic differentiation|0
tumor lysis syndrome|0
septic shock|0
HIV diagnosis|-672
dolutegravir/abacavir/lamivudine (DTG/ABC/3TC) administration|-672
admitted to ICU|0
nasogastric tube administration of DTG/ABC/3TC|0
meropenem administration|0
linezolid administration|0
anidulafungin administration|0
Cp-DTG measurement|96
meropenem Cp through (12.4 mg/L)|96
meropenem Cp peak (35.4 mg/L)|96
linezolid Cp through (1.7 mg/L)|96
linezolid Cp peak (11.9 mg/L)|96
anidulafungin Cp through (2.1 mg/L)|96
anidulafungin Cp peak (5.8 mg/L)|96
undetectable CpDTG including peak|96
acute inflammation from septic shock and tumor lysis syndrome|0
biomarker elevation (ferritin 123280 ng/mL)|0
biomarker elevation (C-reactive protein 24 mg/dL)|0
biomarker elevation (D-dimer 5359 mcg/mL)|0
biomarker elevation (procalcitonin 91 ng/mL)|0
hyperlactatemia (9.5 mmol/L)|0
high norepinephrine requirements (3.6 mg/hour)|0
trophic enteral feeding|0
high gastric retention episodes|0
EF intolerance leading to intestinal mucosa atrophy|0
decreased dolutegravir absorption|0
hypoalbuminemia (1.4 g/dL)|0
hyperbilirubinemia (4.5 mg/dL)|0
fever up to 40ºC|0
rifampin treatment|-72
double dose dolutegravir reduction|-72
continuous venovenous hemodialysis|96
negligible dolutegravir removal by hemodialysis|96
minimal DTG elimination by kidneys (<1%)|0
