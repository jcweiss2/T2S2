57 years old | 0
female | 0
menopausal | 0
admitted to the gynecological emergency unit | 0
left lower quadrant abdominal pain | -504
pelvic heaviness | -504
urinary frequency | -504
past history of 5 miscarriages | -0
tubal ligation | -0
active smoker | 0
no medication | 0
large and painful mass | 0
pelvic MRI | 0
mass measuring 18 × 17 × 12 cm | 0
no lymphadenopathy | 0
no ascites | 0
no peritoneal implants | 0
uterus and adnexa were normal | 0
serum tumor markers were negative | 0
surgical pelvic exploration | 168
30-centimeter mass of the left broad ligament | 168
no ascites | 168
no peritoneal carcinomatosis | 168
uterus and right adnexa were normal | 168
total hysterectomy with adnexectomy | 168
removal of the mass | 168
definitive histological diagnosis was leiomyosarcoma | 168
isolated fever | 48
laboratory evaluation | 48
major inflammatory syndrome | 48
leukocytes 15,000/μL | 48
C-reactive protein 317 mg/dL | 48
contrast-enhanced computed tomography scan | 48
bilobed air and fluid collection | 48
abscess | 48
blood pressure dropped | 48
vasopressor therapy | 48
noradrenaline | 48
emergency revision surgery | 48
peritoneal cavity exploration | 48
moderately abundant non-purulent serosanginous peritoneal fluid | 48
adhesions to the Douglas pouch | 48
peritonitis | 48
antibacterial treatment with piperacillin/tazobactam and gentamicin | 48
microbiological samples | 48
extubated | 72
hemodynamic support with noradrenaline | 72
transferred to the intensive care unit | 72
noradrenaline requirement decreased | 96
discontinuation of noradrenaline | 96
decrease in inflammatory markers | 96
microbiological analysis of the peritoneal fluid | 96
Gardnerella vaginalis | 96
gentamicin discontinued | 96
metronidazole added | 96
Atopobium vaginae | 120
antibacterial susceptibility testing | 120
Garderella vaginalis resistant to metronidazole | 120
Garderella vaginalis susceptible to penicillin G | 120
Garderella vaginalis susceptible to amoxicillin/clavulanate | 120
Garderella vaginalis susceptible to cefotaxim | 120
Garderella vaginalis susceptible to clindamicin | 120
Garderella vaginalis susceptible to vancomycin | 120
Atopobium vaginae susceptible to all tested antibacterials | 120
piperacillin/tazobactam active against both bacteria | 120
final diagnosis | 120
early postoperative peritonitis-induced septic shock | 120
caused by Gardnerella vaginalis and Atopobium vaginae | 120
discharged from the intensive care unit | 168
antibacterial therapy stopped | 168