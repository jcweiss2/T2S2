18 years old | 0
female | 0
admitted to the hospital | 0
severe headache | -24
periorbital and mid-facial swelling | -24
fever | -14
headache | -14
light pain in the right ear | -14
purulent secretion from the ear | -14
swelling and redness of the skin behind the right ear | -14
tinnitus | -14
hearing disorder | -14
diagnosed with right acute mastoiditis | -14
treated with antibiotics | -14
painkillers and anti-inflammatory drugs | -14
anorexia | -10
high fever | -10
confusion | -10
arterial hypertension | -672
ACE inhibitors | -672
marked right facial and periorbital swelling | 0
blepharoptosis | 0
chemosis | 0
proptosis | 0
visual acuity of 7/12 on her right eye | 0
intraocular pressures in both eyes were normal | 0
no relative afferent pupillary defect | 0
color vision was normal | 0
fundoscopy revealed no signs of optic disc swelling | 0
abnormal eye movements | 0
pain on right eye movement | 0
no clinical evidence of right optic nerve compression | 0
no trigeminal sensory deficit | 0
febrile | 0
conscious, but somnolent | 0
no other neurological deficits | 0
blood cultures were taken | 0
inflammatory parameters were significantly elevated | 0
white blood cells count 18×104/L | 0
erythrocyte sedimentation rate 67 mm/h | 0
C-reactive protein 250 mg/L | 0
renal and liver functions within normal limits | 0
tests for vasculitis, HIV, and diabetes were all negative | 0
prothrombin G20210A mutation (PT20210A) | 0
coagulation profile and urinalysis were both normal | 0
MRI of the brain revealed non-opacification of the right cavernous sinus | 0
received empirically high-dose intravenous Ceftriaxone | 0
anticoagulation with Enoxaparin | 0
positive for Streptococcus pneumoniae | 0
shortness of breath | 48
referred to the Intensive Care Unit (ICU) | 48
non-invasive mechanical ventilation | 48
antibiotics were changed to Amikacin and Piperacillin–Tazobactam | 48
chest X-ray revealed unilateral homogeneous opacification on right lobar lung | 48
bronchial aspirate culture confirmed hospital acquired pneumonia | 48
control contrast-enhanced magnetic resonance angiography (CE–MRA) | 96
persistence of the lacunar image in the right cavernous sinus | 96
ophthalmological symptoms improved | 96
periorbital swelling has been diminishing | 96
discharged on oral anticoagulant – Acenocoumarol | 168
follow-up CT venogram will indicate resolution of the thromboses | 168
made a full recovery | 168