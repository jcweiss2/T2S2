76 years old | 0
female | 0
shortness of breath | -1
dysphagia | -1
nausea | -1
neck discomfort | -1
morbid obesity | -6120
laparoscopic adjustable gastric band | -6120
esophageal dilation | -2040
intermittent dysphagia | -2040
removal of LAGB | -336
noncontrast computed tomography of the chest | 0
dilated esophagus | 0
right lateral diverticulum | 0
impacted food bolus | 0
endoscopy | 0
intubation | 0
partial removal of food bolus | 0
inability to wean off mechanical ventilation | 24
severe sepsis | 24
acute respiratory distress syndrome | 24
tracheostomy | 24
surgical gastrostomy tubes | 24
discharged to long-term acute care hospital | 720
achalasia | 0
outflow tract obstruction | 0
pseudoachalasia | 0
Zenker diverticulum | 0
mass lesion | 0
paraesophageal hernia | 0
bariatric procedure | 0
high esophageal lumen pressure | -6120
esophageal musculature weakness | -6120
dysphagia | -1
impactions | -1
removal of LAGB without identification of mass lesion or hernia | -336
manometry | 0
fluoroscopy | 0