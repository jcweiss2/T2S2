2 years old | 0
female | 0
admitted to the hospital | 0
painless limping | 0
walking on tiptoe | 0
premature birth | -8760
low birth weight | -8760
neonatal sepsis | -8760
parenteral antibiotics | -8760
septic arthritis | -8760
overlooked septic arthritis | -8760
no surgical drainage | -8760
no ultrasound-guided repeated aspiration | -8760
pelvic obliquity | 0
Trendelenburg-Duchenne gait | 0
limited right hip abduction | 0
internal rotation | 0
lower-extremity length discrepancy | 0
shortening of right femur | 0
viable femoral head | 0
decreased neck-shaft angle | 0
relative overgrowth of greater trochanter | 0
proximally migration | 0
shortening of femoral neck | 0
severe coxa vara | 0
femoral neck pseudoarthrosis | 0
vertical orientation of the capital physis | 0
Hilgenreiner-epiphyseal angle 75° | 0
Choi Type IIIB | 0
Johari classification Group V | 0
proximal femoral valgus osteotomy | 24
adductor tenotomy | 24
adductor soft tissue release | 24
correction of neck shaft angle | 24
lateral approach | 24
subperiosteal detachment of vastus lateralis muscle | 24
closing wedge valgus osteotomy | 24
internal fixation | 24
partial weight bearing | 24
postoperative management | 24
successful correction of Trendelenburg gait | 168
restored right lower extremity alignment | 168
corrected lower-extremity length discrepancy | 168
transfer of greater trochanter | 168
restoring normal tension to pelvitrochanteric muscles | 168
improving mechanical efficiency | 168
Hilgenreiner-epiphyseal angle 35° | 168
acetabular depth improvement | 720
consolidation of osteotomy | 1020
hardware removal | 1020
no hip pain | 1560
better hip range of motion | 1560
flexion 100° | 1560
extension 10° | 1560
abduction 40° | 1560
adduction 45° | 1560
internal rotation 30° | 1560
external rotation 45° | 1560
no difficulties with recreational activities | 1560
osteotomy healed | 1560
squatting | 1560
running | 1560
climbing stairs | 1560
walking without limp | 1560
no pain in hip | 1560
shortening reduced | 1560
x-ray of hip showed relatively well formed head | 1560
neck shaft angle 136° | 1560
union of previous pseudoarthrosis | 1560