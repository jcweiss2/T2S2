64 years old | 0
male | 0
hypertension | -672
liver cirrhosis | -672
alcohol use disorder | -672
acute mild and intermittent chest pain | -24
dizziness | -24
nausea | -24
palpitations | -24
admitted to the hospital | 0
fever | -24
elevated high sensitivity troponin | 0
normocytic anemia | 0
thrombocytopenia | 0
hypertriglyceridemia | 0
hyponatremia | 0
hypoalbuminemia | 0
elevated liver function enzymes | 0
hyperbilirubinemia | 0
non-ST-elevation myocardial infarction | 0
demand ischemia | 0
severe left ventricular hypertrophy | 0
impaired diastolic dysfunction | 0
lethargic | 24
intermittently agitated | 24
confused | 24
slightly febrile | 24
tachycardic | 24
hypotensive | 24
euvolemic | 24
scleral icterus | 24
jaundice | 24
abdomen soft and non-tender | 24
normoactive bowel sounds | 24
abdomen distended with shifting dullness | 24
worsening liver enzymes | 24
elevated ammonia level | 24
elevated lactic acid | 24
elevated procalcitonin | 24
new acute renal failure | 24
leukocytosis | 24
transferred to the Intensive Care Unit | 24
liver shock | 24
multi-factorial encephalopathy | 24
intubated | 24
started on vasopressors | 24
treated with NAC | 24
treated with rifaximin | 24
treated with lactulose | 24
treated with empiric antibiotics | 24
blood cultures returned positive for Listeria monocytogenes | 48
acute blood loss anemia | 48
possible gastrointestinal hemorrhage | 48
underwent an emergency esophagogastroduodenoscopy | 48
esophageal varices banded | 48
abdominal venous ultrasound | 48
abdominal paracentesis | 48
EEG revealed severe diffuse encephalopathy | 48
lumbar puncture | 48
cerebral spinal fluid cultures returned positive for Listeria monocytogenes | 72
treated with intravenous ampicillin | 72
treated with gentamicin | 72
gentamicin discontinued | 96
rhabdomyolysis | 96
required hemodialysis | 96
extubated | 120
transferred back to the medical floors | 120
continued to receive hemodialysis | 120
continued to receive intravenous ampicillin | 120
continued to receive lactulose | 120
minimal improvement in kidney function | 120
minimal improvement in mentation | 120
repeat ammonia level still elevated | 168
total bilirubin elevated | 168
transitioned to comfort care | 168