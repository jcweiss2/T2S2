27 years old | 0
    female | 0
    sickle cell disease (SSD) | 0
    autosplenectomy | 0
    Crigler-Najjar syndrome | 0
    cholecystectomy | 0
    acute sickle cell pain crisis | 0
    bilateral arm pain | 0
    back pain | 0
    leg pain | 0
    new-onset dyspnea on exertion | -24
    denied chest pain | 0
    hydroxyurea | -8760
    right lower extremity ulcer | -8760
    Voxelotor | 0
    chronic complaint of fatigue | 0
    anemia | 0
    Voxelotor 1.5 g oral daily | 0
    sickle cell pain crises approximately twice yearly | 0
    hemodynamically stable | 0
    hydromorphone | 0
    intravenous fluids | 0
    normal saline | 0
    supplemental oxygen | 0
    anemia | 0
    chest X-ray (CXR) negative for cardiopulmonary infiltrates | 0
    admitted to medical floor | 0
    hydromorphone | 0
    transitioned to Oxycontin | 0
    maintenance fluids | 0
    bedside incentive spirometry | 0
    Voxelotor discontinued | 0
    significant decrease in blood counts | 24
    bicytopenia | 24
    anemia | 24
    thrombocytopenia | 24
    worsening hemolysis | 24
    hyperkalemia | 24
    worsening renal function | 24
    hypoxia | 24
    oxygen saturation 70% | 24
    oxygen supplementation with Venturi-Mask | 24
    clinical suspicion for thrombotic thrombocytopenic purpura (TTP) | 24
    LDH 2646 U/L | 24
    over 4 schistocytes/HPF | 24
    calculated PLASMIC score 4 | 24
    intermediate risk for severe ADAMTS13 deficiency | 24
    transferred to MICU | 24
    double-lumen Shiley central venous catheter (SCVC) placed | 24
    total plasma exchange therapy (TPE) | 24
    RBCs transfusion | 24
    high-dose intravenous methylprednisolone | 24
    ADAMTS13 level activity 64.9% | 24
    platelets improved | 48
    creatinine improved | 48
    LDH improved | 48
    stable after 2 days of plasma exchange | 48
    discharged home | 72
    home voxelotor restarted | 72
    lower dose | 72
    acute painful crisis | 0
    acute coronary syndrome | 0
    acute papillary necrosis | 0
    multiorgan failure | 24
    widespread vasoAocclusive crisis | 24
    thrombocytopenia | 24
    microangiopathic hemolytic anemia (MAHA) | 24
    generalized weakness | 24
    gastrointestinal upset | 24
    neurologic changes | 24
    renal dysfunction | 24
    fever | 24
    sepsis | 24
    acute elevation of renal and hepatic markers | 24
    improvement with plasma exchange | 48
    SCD with multiorgan failure | 24
    TPE-related complications | 72
    paresthesia secondary to hypocalcemia | 72
    bleeding complications | 72
    catheter-related sepsis | 72
    thrombosis | 72
    hypotension | 72
    systemic infection | 72
    fatality | 72
    acute injury to renal and hepatic circulation | 24
    improvement after plasma exchange | 48
    multi-organ failure with SS crises | 24
    vasoocclusion | 24
    organ ischemia | 24
    organ failure in 2-3 organ systems | 24
    thrombocytopenia | 24
    renal dysfunction | 24
    reversal of dysfunction | 72
    
    
    