64 years old | 0
    male | 0
    hypertension | 0
    medication non-adherence | 0
    liver cirrhosis | 0
    active alcohol use disorder | 0
    presented to the Emergency Department | 0
    acute mild and intermittent chest pain | -24
    dizziness | -24
    nausea | -24
    palpitations | -24
    pain started the morning prior to presentation | -24
    resolved spontaneously | -24
    re-emerged throughout the next day | -24
    last shot of alcohol | -72
    reported drinking 1 shot of ethanol 3 times weekly | 0
    recent increased use of acetaminophen | 0
    generalized chronic body aches | 0
    unable to quantify the amount | 0
    denied use of herbal supplements | 0
    denied use of vitamins | 0
    denied use of other over-the-counter medications | 0
    alert | 0
    oriented | 0
    examination unremarkable | 0
    hemodynamically stable | 0
    temperature of 38.7°C | 0
    heart rate of 94 beats per min | 0
    respiratory rate of 18 breaths per min | 0
    blood pressure of 113/55 mmHg | 0
    peripheral oxygen saturation of 97% | 0
    elevated high sensitivity troponin | 0
    normocytic anemia | 0
    hemoglobin 9.2 g/dL | 0
    MCV 84 fL | 0
    thrombocytopenia | 0
    hypertriglyceridemia | 0
    HDL <8 mg/dL | 0
    hyponatremia | 0
    hypoalbuminemia | 0
    elevated liver function enzymes | 0
    ALP 117 unit/L | 0
    AST 900 unit/L | 0
    ALT 169 unit/L |+0
    hyperbilirubinemia | 0
    creatinine kinase within normal limits | 0
    brain natriuretic peptide within normal limits | 0
    lipase levels within normal limits | 0
    baseline hemoglobin approximately 9 to 10 g/dL | 0
    baseline platelets 20 to 30 K/mm3 | 0
    no indication of an active bleed | 0
    electrocardiogram showed normal sinus rhythm | 0
    left axis deviation | 0
    unchanged from previous imaging | 0
    no ST- or T-wave changes | 0
    chest X-ray unremarkable | 0
    admitted to the medical floors | 0
    non-ST-elevation myocardial infarction | 0
    demand ischemia | 0
    2-dimensional echocardiogram | 0
    transesophageal echocardiogram | 0
    preserved ejection fraction | 0
    severe left ventricular hypertrophy | 0
    impaired diastolic dysfunction | 0
    no evidence of valvular defects | 0
    no evidence of infective endocarditis | 0
    scheduled for a stress test | 0
    noted to be lethargic | 24
    Critical Care Unit consulted | 24
    acute encephalopathy | 24
    intermittently agitated | 24
    confused | 24
    lethargic | 24
    slightly febrile | 24
    temperature of 39.2°C | 24
    tachycardic | 24
    blood pressure of 76/41 mmHg | 24
    euvolemic | 24
    scleral icterus | 24
    jaundice | 24
    soft abdomen | 24
    non-tender abdomen | 24
    normoactive bowel sounds | 24
    distended abdomen | 24
    shifting dullness | 24
    worsening liver enzymes | 24
    ALP 131 unit/L | 24
    AST 4698 unit/L | 24
    ALT 1143 unit/L | 24
    total bilirubin 12.7 mg/dL | 24
    ammonia level of 166 mcmol/L | 24
    lactic acid of 5.7 mmol/L | 24
    procalcitonin of 11.33 ng/mL | 24
    acetaminophen level <10 mcg/mL | 24
    salicylate level <2.5 mg/dL | 24
    new acute renal failure | 24
    BUN 22 mg/dL | 24
    creatinine 1.54 mg/dL | 24
    leukocytosis | 24
    segmented neutrophils 78% | 24
    bands 17% | 24
    transferred to the Intensive Care Unit | 24
    liver shock | 24
    multi-factorial encephalopathy | 24
    computerized tomography scan of the brain without contrast | 24
    no gross intracranial hemorrhage | 24
    no midline shift | 24
    no hydrocephalus | 24
    worsening lethargy | 24
    intubated for airway protection | 24
    started on vasopressors | 24
    norepinephrine | 24
    hemodynamic instability secondary to sepsis | 24
    treated with NAC | 24
    treated with rifaximin | 24
    treated with lactulose | 24
    empiric antibiotics | 24
    intravenous vancomycin 1000 mg daily | 24
    cefepime 500 mg daily | 24
    blood cultures returned positive for Listeria monocytogenes | 24
    not a candidate for liver transplantation | 24
    recent alcohol use | 24
    no acute or chronic viral hepatitis | 24
    evidence of previous immunity from vaccinations | 24
    no evidence of HIV | 24
    no evidence of CMV | 24
    no evidence of EBV | 24
    no evidence of HSV infections | 24
    complicated with acute blood loss anemia | 24
    possible gastrointestinal hemorrhage | 24
    requiring multiple transfusions | 24
    transfusions of platelets | 24
    transfusions of red blood cells | 24
    transfusions of fresh frozen plasma | 24
    emergency esophagogastroduodenoscopy | 24
    actively bleeding grade II esophageal varices | 24
    banded esophageal varices | 24
    abdominal venous ultrasound | 24
    no portal vein thrombosis | 24
    bidirectional flow in the right hepatic vein | 24
    intrinsic liver disease | 24
    abdominal paracentesis | 24
    no evidence of spontaneous bacterial peritonitis | 24
    EEG revealed severe diffuse encephalopathy | 24
    Listeria septicemia | 24
    worsening mentation | 24
    lumbar puncture | 24
    treated with intravenous ampicillin 2000 mg every 6 h | 24
    treated with gentamicin 80 mg daily | 24
    cerebral spinal fluid cultures returned positive for Listeria monocytogenes | 24
    worsening renal function | 24
    gentamicin discontinued | 48
    CSF contained 2290 mm3 red blood cells | 24
    CSF contained 658 mm3 white blood cells | 24
    segmented neutrophils 95% | 24
    glucose 19 mg/dL | 24
    protein 68 mg/dL | 24
    complicated by rhabdomyolysis | 24
    creatinine 6.9 mg/dL | 24
    CK 1493 unit/L | 24
    sepsis | 24
    liver shock | 24
    required hemodialysis | 24
    lactic acid normalized | 24
    procalcitonin normalized | 24
    extubated | 24
    transferred back to the medical floors | 24
    continued to receive hemodialysis 3 times weekly | 24
    minimal improvement in kidney function | 24
    continued to receive 21 full days of intravenous ampicillin | 24
    lactulose 3 times daily | 24
    minimal improvement in mentation | 24
    repeat ammonia level elevated | 24
    total bilirubin of 33.4 mg/dL | 24
    encephalopathy | 24
    hemodynamic instability | 24
    hepatic failure | 24
    renal failure | 24
    no improvement | 24
    seen by the Palliative Care Unit | 24
    transitioned to comfort care | 24
    family reported no recent consumption of deli meat | 24
    no recent consumption of cheeses | 24
    no recent consumption of smoked fishes | 24
    no recent consumption of raw chicken | 24
    no known outbreaks in the area | 24
    