87 years old | 0
man | 0
brought in by ambulance | 0
fever of 38.0°C | 0
general fatigue | 0
denied history of trauma | 0
denied history of falls | 0
endoscopic sphincterotomy for choledocholithiasis | -7920
percutaneous coronary intervention for ischemic heart disease | -70080
took warfarin potassium | 0
took aspirin | 0
took antidiabetic medications | 0
took diuretics | 0
heart rate of 115 per minute | 0
blood pressure of 92/61 mmHg | 0
respiratory rate of 13 per minute | 0
body temperature of 36.2°C | 0
Glasgow coma scale E4 | 0
Glasgow coma scale V4 | 0
Glasgow coma scale M4 | 0
height 164 cm | 0
body weight 70 kg | 0
body mass index 26.0 kg/m2 | 0
moderate abdominal pain | 0
tenderness in the epigastrium | 0
hemoglobin 9.6 g/dL | 0
white blood cell count 23170/µL | 0
platelet count 13.6 × 10^4/µL | 0
total bilirubin 1.0 mg/dL | 0
alanine transaminase 843 IU/L | 0
aspartate aminotransferase 339 IU/L | 0
lactate dehydrogenase 1278 U/L | 0
alkaline phosphatase 947 U/L | 0
blood urea nitrogen 40.5 mg/dL | 0
creatinine 3.06 mg/dL | 0
prothrombin time 18.3 seconds | 0
prothrombin time % 44% | 0
international normalized ratio 1.6 | 0
activated partial thromboplastin time 38.4 seconds | 0
procalcitonin 251 ng/mL | 0
C-reactive protein 17.4 mg/dL | 0
lactate 33 mg/dL | 0
brain natriuretic peptide 1206 ng/mL | 0
α-Fetoprotein 0.7 ng/mL | 0
sepsis | 0
anemia | 0
liver dysfunction | 0
renal dysfunction | 0
heart failure | 0
coagulopathy | 0
swelling not detected | 0
wall thickening of the gallbladder not detected | 0
subcapsular high density area of the liver | 0
subcapsular hemorrhage | 0
small amount of free fluid around the spleen | 0
initial diagnosis of sepsis due to cholangitis | 0
initial diagnosis of sepsis due to liver damage | 0
admitted to intensive care unit | 0
treated with intravenous antibiotics | 0
meropenem hydrate | 0
endoscopic retrograde cholangiography performed | 0
no stone in the bile duct | 0
endoscopic nasobiliary drainage performed | 0
treated with noradrenaline | 0
treated with dobutamine hydrochloride | 0
blood culture positive for klebsiella oxytoca | 24
meropenem hydrate administered | 24
hemoglobin 7.5 g/dL | 72
white blood cell count 19030/µL | 72
C-reactive protein 30.1 mg/dL | 72
procalcitonin 279.6 ng/mL | 72
blood urea nitrogen 50.1 mg/dL | 72
creatinine 2.57 mg/dL | 72
anemia progressed | 72
required 2 units of blood transfusion | 72
renal damage slightly improved | 72
infection not controlled | 72
inflammatory markers remained high | 72
contrast-enhanced abdominal CT performed | 72
intrahepatic low density areas | 72
subcapsular low density areas | 72
gallbladder wall defect | 72
small amount of free fluid around the liver | 72
small amount of free fluid around the spleen | 72
hemorrhagic fluid obtained through paracentesis | 72
transhepatic perforation of acute cholecystitis suspected | 72
emergency interventional radiology | 72
percutaneous transhepatic gallbladder drainage attempted | 72
high echogenic debris in the gallbladder | 72
drainage tube inserted into the gallbladder | 72
90 mL red-yellow pus aspirated | 72
orifice of fistula | 72
contrast medium drained into intrahepatic secondary abscess | 72
contrast medium drained into intraperitoneal cavity | 72
percutaneous abscess drainage attempted | 72
150 mL hemorrhagic fluid aspirated | 72
abdominal angiography attempted | 72
no extravasation | 72
no hepatic artery aneurysm | 72
no cystic artery aneurysm | 72
transhepatic gallbladder perforation confirmed | 72
hemoperitoneum confirmed | 72
sepsis confirmed | 72
PTGBD and percutaneous abscess drainage performed | 72
general condition improved | 72
emergency laparotomy avoided | 72
culture of red-yellow pus positive for enterococcus avium | 72
culture of red-yellow pus positive for enterococcus gallinarum | 72
culture of red-yellow pus positive for klebsiella oxytoca | 72
culture of intrahepatic abscess positive for enterococcus gallinarum | 72
repeat blood culture negative | 120
antibiotics changed to sulbactam sodium/ampicillin sodium | 168
sulbactam sodium/ampicillin sodium administered | 168
contrast-enhanced CT showed reduction in intrahepatic abscess | 408
contrast-enhanced CT showed reduction in subcapsular hematoma | 408
cholangiography via PTGBD tube revealed recanalization of cystic duct | 408
orifice of fistula not detected | 408
no stone in the gallbladder | 408
no stone in the bile duct | 408
discharged | 792
