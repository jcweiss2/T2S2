14 years old | 0
male | 0
brought to the emergency department | 0
near-drowning incident | -?
loss of consciousness | -?
brief bystander CPR performed | -?
hemodynamically stable | 0
fully conscious | 0
complained of abdominal pain | 0
diffuse abrasions on torso | 0
abdomen soft | 0
no peritoneal signs | 0
chest x-ray performed | 0
pneumoperitoneum | 0
CT scan revealed pneumomediastinum | 0
intraabdominal free fluid | 0
concern for hollow viscus perforation | 0
taken emergently to operating room | 0
laparotomy performed | 0
gross contamination with food debris | 0
total GE junction disruption | 0
hemodynamically labile | 0
damage control procedure performed | 0
distal esophagus stapled closed | 0
proximal stomach stapled closed | 0
four drains placed | 0
mediastinal drain placed | 0
gastrostomy tube placed | 0
no surgical proximal esophageal diversion | 0
large bore nasogastric tube placed | 0
intraabdominal drains placed | 0
fascia closed | 0
transferred to ICU | 0
ICU stay complicated by septic shock | 24
respiratory failure | 24
prolonged intubation | 24
deep venous thrombosis | 24
pulmonary embolism | 24
bilateral pleural effusions | 24
general deconditioning | 24
parenteral nutrition started | 24
extubated on postoperative day 18 | 432
fluoroscopic evaluation demonstrated esophageal leak | 432
mediastinal drain controlled leak | 432
stomach negative for leak | 432
enteral nutrition initiated via G tube | 432
discharged on day 50 | 1200
nasogastric tube retained | 1200
mediastinal drain retained | 1200
three months after initial injury | 2160
underwent Ivor-Lewis esophagectomy | 2160
gastric pull-up for anastomosis | 2160
partial left lateral decubitus position | 2160
midline abdominal incision | 2160
gastric conduit made | 2160
right thoracotomy performed | 2160
distal esophagus identified | 2160
stomach advanced into chest | 2160
end-to-end anastomosis stapler used | 2160
leak test performed | 2160
jejunostomy tube placed | 2160
extubated on postoperative day 3 | 2160
nutritionally supported with enteral feeds | 2160
esophagram on day 7 | 2160
no leak at anastomosis | 2160
immediate stomach emptying | 2160
initiated on liquid diet | 2160
discharged on day 10 | 2160
most recent clinic visit 5 months post-reconstruction | 3600
tolerates regular diet | 3600
gaining weight | 3600
recovering well | 3600
no declarations of interest | 0
written informed consent obtained | 0
ethical approval exempt | 0
authors meet authorship criteria | 0
