73 years old | 0
female | 0
hypertension | 0
syphilis | 0
type 2 diabetes mellitus | 0
altered mental status | 0
mechanical fall | -744
pruritic scalp | -744
purulent drainage from sinuses on the scalp | -744
temperature of 97.9°F | 0
heart rate of 127 bpm | 0
respiratory rate of 22 breaths/min | 0
blood pressure of 144/80 mmHg | 0
oxygen saturation of 98% | 0
oriented to person | 0
oriented to place | 0
not oriented to time | 0
face erythematous | 0
face edematous | 0
scalp erythematous | 0
scalp edematous | 0
right ear erythematous | 0
right ear edematous | 0
large fluctuant mass | 0
purulent drainage | 0
posterior auricular mass | 0
hyperglycemia | 0
anion gap metabolic acidosis | 0
serum bicarbonate of 20 | 0
ketonuria | 0
extensive multifocal scalp swelling | 0
admitted to the intensive care unit | 0
diabetic ketoacidosis | 0
cellulitis of the scalp | 0
underlying abscesses | 0
continuous infusion of insulin | 0
intravenous Vancomycin | 0
intravenous Cefepime | 0
incision and drainage of scalp lesion | 48
subgaleal abscess | 48
MRSA | 72
paranasal sinus CT | 72
transesophageal echocardiogram | 72
pulse irrigation of the wounds | 96
sharp debridement | 96
serial bedside debridements | 96
scalp wound | 96
right posterior auricular wound | 96
split-thickness skin grafts | 120
definitively closed | 120
discharged | 768
intravenous Vancomycin | 0