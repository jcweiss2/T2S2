16 years old | 0\
primigravida | 0\
admitted to the emergency room | 0\
pregnancy diagnosis of 37.6 weeks of gestation | -672\
viable intrauterine pregnancy | -672\
fetal heart rate of 143 beats per minute | -672\
fetus situated longitudinally with cephalic presentation | -672\
back to the left | -672\
cervix 6 cm dilated | -672\
70% effaced | -672\
station +1 | -672\
intact membranes | -672\
mild edema of the extremities | -672\
normal osteotendinous reflexes | -672\
obstetrical ultrasound | -672\
pregnancy of 37+0 weeks of gestation | -672\
posterior body placenta maturation grade III | -672\
amniotic fluid index of 8.7 cm | -672\
biophysical profile of 8/8 | -672\
Hadlock of 34.2% | -672\
weight of 3033 grams | -672\
continue labor monitoring | -672\
spontaneous rupture of the membranes | -5\
labor progressed | -5\
effective labor | -5\
4 contractions every 10 minutes | -5\
contractions lasted 40 to 45 seconds | -5\
no need for uterotonic agents | -5\
moved to the labor room | -1\
fully dilated | -1\
100% clearance | -1\
station of +3 | -1\
fetus in left occiput anterior position | -1\
live newborn delivered | 0\
Apgar scores of 7 and 9 | 0\
gestational age of 40 weeks | 0\
height 48 cm | 0\
weight of 2650 grams | 0\
Schultze mechanism | 0\
placenta came out with normal characteristics | 0\
grade III uterine inversion | 0\
manual reinversion maneuvers | 0\
total blood loss of 1200 mL | 0\
UA | 0\
oxytocin | 0\
carbetocin | 0\
misoprostol | 0\
persistent uterine inversion | 0\
exploratory laparotomy | 1\
general anesthesia | 1\
surgery room | 1\
reinversion | 1\
UA persisted | 1\
PPH | 1\
Hayman hemostatic suture | 1\
no response | 1\
bilateral ligation of the anterior trunk of the hypogastric artery | 1\
immediate recovery of uterine tone | 1\
cessation of PPH | 1\
uterus regained tone | 1\
postligation bleeding | 1\
50 mL of the total blood loss | 1\
transfused 2 bags of packed red blood cells | 2\
gasometry showed a hemoglobin level of 7 g | 2\
transferred to the recovery room | 2\
transferred to the medical intensive care unit | 2\
transferred to a hospital room | 24\
normal diet | 24\
ambulation | 24\
spontaneous uresis | 24\
normal peristalsis | 24\
breastfeeding | 24\
discharged | 48