73 years old | 0
male | 0
massive splenomegaly | 0
polycythaemia vera | 0
myelofibrosis | 0
mild valvular heart disease | 0
scheduled for splenectomy | 0
admitted | 0
negative real-time PCR test for CoV-2 | 0
early postoperative course uneventful | 0
splenectomy-related decrease in platelet count | 0
CoV-2 positive | 0
exposure to infected patient | 0
clinical features consistent with non-severe CoV-2 disease | 0
transferred to surgical CoV-2 unit | 0
care of multidisciplinary team | 0
surgeons | 0
infectious disease consulting service | 0
sudden worsening of general condition | 0
non-severe-to-severe CoV-2 disease | 0
appearance of dyspnoea | 0
elevation in D-dimer up to 30946 ng/mL | 0
chest CT scan | 0
multiple bilobar ground-glass opacities | 0
interstitial pneumonia | 0
massive left pleural effusion | 0
no signs of pulmonary embolism | 0
left chest tube inserted | 0
improvement of dyspnoea | 0
severe hypotension | 312
massive drop in haemoglobin levels until 55 g/L | 312
mild prolongation of prothrombin time (PT) values of 1.21 of international normalised ratio | 312
abdomen CT scan | 312
thrombosis in the remnant of the splenic vein | 312
splenomesenteric confluence | 312
large blood collection in the left hypochondrium | 312
no signs of active bleeding | 312
supported with three units of packed red blood cells | 312
unit of platelets | 312
urgent surgical exploration | 312
diffuse peritoneal bleeding spots | 312
abdominal lavage | 312
haemostatic patches positioning | 312
no parameters of multiple organ failure | 312
admitted to the intensive care unit (ICU) | 312
extubated | 312
re-posted to the surgical CoV-2 unit | 312
developed fever | 312
hypoxaemia | 312
initially treated with high-flow oxygen support | 312
required mechanical ventilation | 312
sequential organ failure assessment score 5 | 312
ICU mortality risk of 20.2% | 312
blood cultures | 312
urine cultures | 312
pleural liquid cultures | 312
microbiological isolation | 312
samples for cytomegalovirus DNA | 312
cytomegalovirus DNA negative | 312
pleural liquid sample showed Staphylococcus epidermidis | 312
Bacillus licheniformis | 312
blood cultures positive for S. hominis | 312
general conditions did not improve | 312
failed on postoperative day 22 in the ICU | 528
discharged | 528
death | 528
