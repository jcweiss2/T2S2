70 years old | 0
female | 0
Caucasian | 0
presented to emergency department | 0
worsening shortness of breath | 0
productive cough | -72
nasal congestion | -72
diarrhea | -72
vomiting | -72
hypertension | -inf
tobacco use | -inf
no significant surgical history | 0
no significant family history | 0
in distress | 0
pale appearance | 0
oxygen saturation 77% on room air | 0
blood pressure 94/53 mmHg | 0
heart rate 122 bpm | 0
temperature 36.8 °C | 0
poor air movement | 0
diminished breath sounds at the bases bilaterally | 0
no audible wheezing | 0
no crackles | 0
arterial blood gas pH 7.30 | 0
pCO2 43 mmHg | 0
pO2 48 mmHg | 0
lactic acid 4.4 mmol/L | 0
leukocyte count 25,000/mm3 | 0
bandemia 21% | 0
hemoglobin 13.2 g/dL |1
hematocrit 40.2% | 0
platelet count 199,000/mm3 | 0
chest x-ray hazy bibasilar opacities | 0
no pleural effusion | 0
no pneumothorax | 0
noninvasive bi-level ventilation | 0
oxygen saturation increased to 93% | 0
shortness of breath improved | 0
desire not to be intubated | 0
desire not to be resuscitated | 0
blood cultures obtained | 0
urine cultures obtained | 0
respiratory virus panel | 0
influenza panel | 0
urine streptococcal antigen | 0
urine legionella antigen | 0
piperacillin-tazobactam | 0
vancomycin | 0
admitted to medical intensive care unit | 0
antimicrobial changed to ceftriaxone | 0
antimicrobial changed to azithromycin | 0
blood cultures grew Pasteurella multocida | 24
organism sensitive to all antibiotics tested | 24
de-escalated to ceftriaxone monotherapy | 24
other cultures negative | 24
viral panels negative | 24
owns sixteen indoor cats | 24
denied recent scratches | 24
denied recent bites | 24
skin intact | 24
no evidence of scratches | 24
no evidence of bites | 24
no tetanus shot administered | 24
noninvasive ventilation weaned | 72
transitioned to venturi mask | 72
hemodynamics stable | 72
off vasopressor support | 72
leukocytosis improved | 72
lactic acidosis resolved | 72
bilateral pleural effusions visualized | 72
right effusion more prominent | 72
thoracentesis performed | 72
1000 mL straw-colored fluid removed | 72
transudate by Light's criteria | 72
gram stain negative | 72
culture negative | 72
remained hypoxic | 144
CT angiogram performed | 144
multifocal pneumonia right middle lobe | 144
multifocal pneumonia right lower lobe | 144
multifocal pneumonia left lower lobe | 144
moderate sized right pleural effusion | 144
no pulmonary embolism | 144
discharged home | 144
home oxygen | 144
IV ceftriaxone | 144
14 days of treatment | 144
