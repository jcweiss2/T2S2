53 years old | 0
    male | 0
    admitted to the hospital | 0
    exertional dyspnea | -168
    productive cough | -960
    extended thymectomy | -3360
    lymphoepithelioid type of thymoma | -3360
    adjuvant radiotherapy (45 Grays) | -3360
    sarcoidosis | -1440
    imaging study | -1440
    transbronchial lung biopsy | -1440
    new cavitary lesion detected on HRCT | -240
    anti-tuberculosis chemotherapeutic regimen | -240
    blood pressure 90/60 mmHg | 0
    body temperature 39.3℃ | 0
    pulse rate 152 beats per minute | 0
    respiration rate 32 breaths per minute | 0
    inspiratory crackles in both lower lung fields | 0
    chest roentgenogram haziness | 0
    disseminated nodules in both lung fields | 0
    conglomerated cavities in right upper lobe | 0
    multiple micronodular densities on chest CT | 0
    multiple cavitary nodules in right upper lobe | 0
    condition worsened compared to CT 10 days previous | 0
    new ground glass opacity (GGO) in both lower lobes | 0
    white blood cell count 3500 cells/mm3 | 0
    hemoglobin 15.2 g/dL | 0
    platelet count 253,000 cells/mm3 | 0
    erythrocyte sedimentation rate 36 mm/h | 0
    C-reactive protein 17.29 mg/dL | 0
    mildly elevated AST 81 U/L | 0
    normal renal function | 0
    HIV test negative | 0
    arterial blood gas pH 7.44 | 0
    PaCO2 34.0 mmHg | 0
    PaO2 60.5 mmHg |#%
0
    HCO3 22.8 mmol/L | 0
    SaO2 91.9% | 0
    admitted to intensive care unit | 0
    bronchoalveolar lavage (BAL) | 0
    BAL fluid cell count 119/µL | 0
    BAL cell differential 30% macrophages | 0
    BAL cell differential 60% lymphocytes | 0
    CD4/CD8 ratio 7/46 | 0
    BAL cell differential 10% neutrophils | 0
    PCR positive for Pneumocystis jirovecii | 0
    DFA positive for Pneumocystis jirovecii | 0
    culture negative for cytomegalovirus | 0
    trimethoprim/sulfamethoxazole administered | 0
    methylprednisolone administered | 0
    neutrophil dihydrorhodamine test normal | 0
    T lymphocytes (CD3) 290/µL | 0
    B lymphocytes (CD19) 0/µL | 0
    CD4 148/µL | 0
    CD8 132/µL | 0
    IgG 507 mg/dL | 0
    IgA 31 mg/dL | 0
    IgM <3 mg/dL | 0
    video-assisted thoracoscopic biopsy | 0
    diffuse thickening of alveolar wall with fibrosis | 0
    lymphocyte infiltration | 0
    acid-fast bacilli smear negative | 0
    immunohistochemical analysis negative for CMV | 0
    immunohistochemical analysis negative for HSV | 0
    immunohistochemical analysis negative for adenovirus | 0
    Good's syndrome diagnosis | 0
    supportive ventilatory care | 0
    antibiotic treatment for acute respiratory distress syndrome | 0
    hypogammaglobulinemia persisted | 0
    regular IVIG infusions | 0
    pneumonia not improved | 0
    diarrhea not improved | 0
    infection worsened | 0
    Candida albicans in pleural fluid culture | 0
    Candida albicans in catheter tip culture | 0
    septic shock | 2160
    multi-organ failure | 2160
    death | 2160