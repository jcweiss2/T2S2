35 years old | 0
Hispanic | 0
female | 0
admitted to the hospital | 0
chronic pancreatitis | -672
alcoholic liver disease | -672
alcohol abuse | -672
10/10 diffuse abdominal pain | -72
abdominal pain radiating to the thorax | -72
previous admission | -168
acute chronic pancreatitis | -168
pancreatic pseudocyst | -168
necrosis | -168
current smoker | 0
16-pack year history | 0
consuming 1 to 2 glasses of alcohol daily | -720
abstinent from alcohol ingestion | -720
denied any history of illicit drug use | 0
blood pressure 91/55 | 0
pulse 114 bpm | 0
respiratory rate 18 | 0
T 98.1°F | 0
99% saturation on room air | 0
abdomen was markedly distended | 0
diffusely tender to palpation | 0
positive fluid wave | 0
voluntary guarding | 0
leukocytosis | 0
white blood cell 16.9 | 0
hemoglobin 10.3 | 0
sodium 130 | 0
lipase 149 | 0
liver function tests within normal limits | 0
repeat computed tomographic abdomen and pelvis with contrast | 0
significant increase in ascites | 0
multiple pancreatic cysts | 0
10 mm fluid density lesion | 0
enlarged peripancreatic fluid | 0
paracentesis | 0
2 L of ascitic fluid removed | 0
WBC 8423 | 0
RBC 1570 | 0
PMN 82% | 0
protein 3.2 | 0
amylase 5507 | 0
lactate dehydrogenase 478 | 0
serum-ascites albumin gradient 0.1 | 0
endoscopic retrograde cholangiopancreatography | 0
5 Fr by 9 cm plastic stent placed | 0
transferred to the intensive care unit | 24
acute respiratory distress syndrome | 24
arterial blood gas | 24
pH 7.36 | 24
PCO2 30 | 24
PO2 50 | 24
HCO3 18.8 | 24
100% FiO2 | 24
non-rebreathing mask | 24
vasopressor support | 24
mean arterial pressure 65 | 24
septic shock | 48
leukocytosis | 48
ceftriaxone 2000 mg | 48
spontaneous bacterial peritonitis treatment | 48
IV meropenem | 48
serial CT scans | 72
post ERCP imaging | 72
intubated | 72
acute respiratory failure | 72
tracheostomy | 96
percutaneous endoscopic gastrostomy feeding tube | 96
3 additional paracentesis procedures | 120
4 L removed | 120
3 L removed | 144
2 L removed | 168
Jackson-Pratt drains | 168
interval CT of the abdomen | 168
increase in size of the pancreatic pseudocyst | 168
loculated mesenteric collections | 168
serosal implants | 168
surgical consultation | 168
hyperdense material | 168
hemorrhagic pancreatitis | 168
interventional radiology | 192
drained the pseudocysts | 192
1.6 L of dark purulent fluid | 192
hemoglobin stabilized | 192
8.5 g/dL | 192
CT abdomen scans | 216
resolving pseudocyst collections | 216
pancreatic edema | 216
bilateral pleural effusions | 216
thoracentesis | 216
600 mL of fluid removed | 216
transudative pattern | 216
WBC 664/mm3 | 216
RBC 1580/mm3 | 216
PMN 62% | 216
glucose 81 mg/dL | 216
protein 2.2 g/dL | 216
LDH 232 µ/L | 216
Pseudomonas aeruginosa health care–associated pneumonia | 240
IV meropenem | 240
Clostridium difficile–associated diarrhea | 240
oral vancomycin | 240
IV metronidazole | 240
weaned off the ventilator | 1224
transitioned to a trach collar | 1224
second ERCP | 1248
common bile duct stent removal | 1248
PEG tube removal | 1248
discharged to a subacute rehabilitation facility | 2448
1.5 LPM supplemental oxygen | 2448
nasal cannula | 2448