60 years old | 0
male | 0
hypothyroidism | -720
alcohol abuse | -720
admitted to an outside hospital | -720
found unresponsive | -720
subacute, rapidly progressive cognitive decline | -720
sepsis | -720
aspiration pneumonia | -720
accidental opioid overdose | -720
accidental benzodiazepine overdose | -720
acute respiratory failure | -720
intubation | -720
ICU admission | -720
rehabilitation | -720
discharged home | -720
mental status not back to baseline | -720
behavioral changes | -24
re-admitted to outside hospital | 0
progressive neuropsychiatric decline | 0
decreased awareness | 0
decreased engagement with surroundings | 0
near akinetic mutism | 0
elevated protein at 86 mg/dL | 0
T2-weighted image hyperintensities in bilateral basal ganglia | 0
increased T2-weighted image signal of white matter in bilateral cerebral hemispheres | 0
intermittent left-sided frontotemporal slowing | 0
sharp waves | 0
diffuse slowing | 24
trial of lacosamide | 0
3-day course of IVMP 1 gr/day | 0
transferred to Tampa General Hospital | 24
awake and alert | 24
non-verbal | 24
unable to follow commands | 24
unable to mimic commands | 24
required assistance with activities of daily living | 24
meaningful movements limited | 24
no focal weakness | 24
no asymmetric weakness | 24
serum laboratory testing unrevealing | 24
mildly elevated CRP | 24
mildly elevated ESR | 24
repeat lumbar puncture | 24
OP 22 cmH2O | 24
mildly elevated protein 70 mg/dL | 24
MRI white matter changes | 24
continuous video EEG | 24
slow background | 24
intermittent generalized and rhythmic slow | 24
no epileptogenic activity | 24
CT chest, abdomen, pelvis negative | 24
steroid responsive encephalopathy with thyroiditis considered | 24
5-day course of IVMP 1 gr/day | 24
no clinical improvement | 24
administration of non-prescription opioids | -720
administration of non-prescription benzodiazepines | -720
injectable anabolic steroids | -720
testosterone enanthate | -720
dianabol | -720
application of insecticides | -720
application of rodent-repellents | -720
treated with IVIG 2 gm total | 48
brain biopsy performed | 72
spongiform changes | 72
reactive gliosis | 72
absence of inflammation | 72
discharged to rehabilitation facility | 96
slowly significant clinical improvement | 144
alert and attentive | 8760
non-dysarthric speech | 8760
normal speech content | 8760
following commands | 8760
mild expressive aphasia | 8760
fully ambulatory | 8760
MMSE score 23/30 | 8760
moderately extensive chronic deep white matter changes | 8760
genetic evaluation negative | 8760
continued clinical improvement | 8760
toxin-induced leukoencephalopathy | 72
non-FDA approved anabolic steroids | -720
opioids | -720
benzodiazepines | -720
insecticides | -720
rodent-repellents | -720
elevated protein (CSF) | 0
normal CSF glucose | 0
normal CSF encephalitis panel | 0
normal CSF VDRL | 0
normal CSF cytology | 0
normal CSF West Nile virus | 0
normal CSF 14-3-3 | 0
normal CT head | 0
normal MRI brain | 0
normal MRA head and neck | 0
normal cerebral angiogram | 0
negative autoimmune panel | 24
negative paraneoplastic panel | 24
negative protein 14-3-3 | 24
negative infectious workup | 24
negative metabolic panel | 24
negative heavy metal panel | 24
negative genetic evaluation | 8760
