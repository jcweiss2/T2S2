61 years old | 0
male | 0
admitted to the hospital | 0
hypertension | -672
squamous cell carcinoma of the skin | -672
cyst removal | -672
fever | -72
confusion | -72
rash | -72
TMP-SMX | -336
surgery | -336
excision | -336
wound infected | -336
squamous cell skin lesions removal | -336
altered mental status | 0
sinus tachycardia | 0
mild tenderness in the right upper quadrant | 0
healing excisions | 0
sutured wound | 0
diffuse petechiae | 0
maculopapular rash | 0
no mucosal/oral involvement | 0
no bullae or pustules | 0
no gross motor or sensory deficits | 0
white blood cell count of 5.1 × 10 ³/uL | 0
no eosinophils or monocytes | 0
platelet count of 13 × 10 ³/uL | 0
sodium of 122 mmol/L | 0
creatinine of 2.77 mg/dL | 0
blood urea nitrogen of 50 mg/dL | 0
Aspartate aminotransferase of 238 units/L | 0
Alanine aminotransferase of 79 units/L | 0
Prothrombin time of 12.4 s | 0
International normalized ratio of 1.1 | 0
Partial thromboplastin time of 65 s | 0
sepsis | 0
lactic acid of 1.8 mmol/L | 0
fluid resuscitation | 0
blood cultures drawn | 0
vancomycin | 0
piperacillin/tazobactam | 0
platelet transfusion | 0
transferred to ICU | 0
plasmapheresis | 0
Infectious Disease consultation | 0
Nephrology consultation | 0
Hematology/Oncology consultation | 0
peripheral smear | 0
no schistocytes | 0
elevated fibrinogen | 0
elevated D-dimer | 0
ADAMTS13 activity of 34.9 % | 0
G6PD value within normal limits | 0
renal studies | 0
2+ hemoglobin | 0
trace RBC's | 0
FeNA of 2.79 mEq/L | 0
intrinsic renal injury | 0
TMP-SMX discontinued | 0
mentation returned to baseline | 72
maculopapular rash disappeared | 72
lab values corrected | 96
transferred out of ICU | 96
discharged | 120