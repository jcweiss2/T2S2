28 years old | 0
male | 0
admitted to the hospital | 0
iron deficiency anemia | -672
intermittent diarrhea | -672
rectal bleeding | -672
cirrhotic appearance of the liver | -672
splenomegaly | -672
gastric varices | -672
elective esophagogastroduodenoscopy (EGD) | 0
lesions consistent with gastric varices | 0
glue injection | 0
exsanguinating hemorrhage | 0
admission to the intensive care unit | 0
resuscitation | 0
hemodynamic stability | 0
loose stools | -8760
occasional blood | -8760
heavy drinking | -8760
iatrogenic upper gastrointestinal hemorrhage | 0
variceal bleeding | 0
portal hypertension | 0
cirrhosis of uncertain etiology | 0
repeated EGD | 24
general anesthesia | 24
Sengstaken-Blakemore tube | 24
CT angiogram | 24
no active bleeding | 24
provisional diagnosis of portal hypertension | 24
cirrhosis | 24
rescue transjugular intrahepatic portosystemic shunt (TIPS) | 48
removal of the Sengstaken-Blakemore tube | 72
episodes of melena | 96
further admission to the intensive care unit | 96
third EGD | 120
oozing gastric varices | 120
multiple bandings | 120
glue injections | 120
further attacks of melena | 144
TIPS patency | 144
Doppler ultrasonography | 144
CT angiography | 144
inconclusive TIPS patency | 144
cirrhosis of the liver with uncertain etiology | 168
high United Kingdom Model for End-Stage Liver Disease score | 168
transfer to the regional liver transplantation unit | 168
TIPS venogram | 192
migration of glue | 192
inferior vena cava (IVC) | 192
right atrium (RA) | 192
pulmonary embolization | 192
repeat CT scan | 216
good patency of the TIPS | 216
distribution of glue cast | 216
mobile glue cast in the RA | 216
embolized pieces in branches of the pulmonary arteries | 216
transthoracic echocardiography | 240
mobile echogenic, standlike structures within the RA | 240
normal biventricular size and function | 240
cardiology team consultation | 264
potential retrieval options | 264
anticoagulation with therapeutic low-molecular-weight heparin | 264
liver failure | 288
cardiopulmonary bypass machine | 288
open heart removal | 288
comprehensive work-ups | 312
magnetic resonance cholangiopancreatography | 312
sigmoidoscopy | 312
final diagnosis of cirrhosis of the liver due to primary sclerosing cholangitis | 312
overlapping ulcerative colitis | 312
migration of glue used to treat gastric varices | 312
multidisciplinary discussion | 336
consensus on glue retrieval options | 336
IR approach | 336
standby rescue cardiothoracic team | 336
fluoroscopy by the IR team | 360
no visible radiopaque glue cast | 360
echocardiogram | 360
presence of an echogenic glue cast | 360
lipiodol dissolved | 360
radiolucent Histoacryl glue remained in the RA | 360
IR option no longer feasible | 360
multidisciplinary meeting | 384
direct atrial extraction by the cardiothoracic team | 384
liver transplantation surgery | 384
cardiopulmonary bypass machine support | 384
waiting list for liver transplantation | 408
glue cast removal by direct extraction | 408
liver transplantation surgery | 408