9 years old | 0
neutered male | 0
domestic shorthair cat | 0
presented to tertiary referral hospital | 0
acute hemodynamic decompensation | 0
weakness | -72
suspected lower urinary tract disease | -72
no history of trauma | 0
indoor only | 0
severe cardiovascular collapse | -72
obtunded | 0
prolonged capillary refill time | 0
bradycardia (70 beats/min) | 0
hypothermia (35°C) | 0
weak femoral pulses | 0
low blood pressure (undetectable via Doppler) | 0
initial resuscitation (lactated Ringer's solution bolus) | 0
fluid rate for dehydration replacement | 0
ultrasound: free abdominal fluid | 0
no pleural/pericardial effusion | 0
no B-lines in thorax | 0
ECG: atrial standstill with idioventricular escape rhythms | 0
severe metabolic acidosis | 0
hyperkalemia | 0
presumptive diagnosis of uroabdomen | 0
calcium gluconate administration | 0
sodium bicarbonate administration | 0
abdominocentesis: serosanguinous fluid | 0
[Creatinine]abdominal-fluid/[Creatinine]serum = 6.09 | 0
[K+]abdominal-fluid/[K+]plasma = 2.28 | 0
intracellular bacteria (cocci) in abdominal fluid | 0
ceftazidime administration | 0
percutaneous central venous line placement | 0
urinary catheter placement | 0
difficulty in urinary catheter passage | 0
concern for urethral obstruction | 0
lactated Ringer's solution bolus | 0
cardiovascular response monitoring | 0
systolic blood pressure increased to 110 mmHg | 0
heart rate increased to 180 beats/min | 0
capillary refill time <2 seconds | 0
ECG: sinus rhythm | 0
external heat support | 0
temperature normalization | 0
tramadol administration | 0
peritoneal dialysis initiation | 0
peritoneal dialysis solution (lactated Ringer's with dextrose and heparin) | 0
dialysate volume exchange | 0
increased dialysate volume over 12 hours | 0
improved blood gas analysis at 8 hours | 8
brighter and more responsive | 8
fluid retention: dialysate OUT > dialysate IN | 0
diagnostic abdominal ultrasound at 18 hours | 18
large volume of gravity-dependent sediment in bladder | 18
suspected bladder rupture | 18
fever | 18
clindamycin administration | 18
stable condition | 36
azotemia improvement | 36
glucose and lactate improvement | 36
peritoneal dialysis catheter removal | 36
retrograde contrast cystography: bladder rupture | 36
exploratory laparotomy | 36
surgical correction of bladder rupture | 36
bladder biopsy for culture | 36
postoperative ultrasound: bilateral pleural effusion | 36
echocardiogram: no cardiac disease or fluid overload | 36
negative fluid balance (240 ml) | 36
clinical euvolemia | 36
thoracocentesis | 36
pleural fluid analysis: transudate | 36
[Creatinine]pleural/[Creatinine]plasma = 2.38 | 36
diagnosis of urothorax | 36
uneventful recovery | 36
no respiratory distress | 36
pleural effusion resolution | 36
Klebsiella pneumoniae and Mannheimia haemolytica culture | 36
Micrococcus and Staphylococcus species culture | 36
enrofloxacin administration | 36
discharged after 4 days | 96
follow-up ultrasound: no abdominal or pleural fluid | 168
