11 years old | 0 | 0 
female | 0 | 0 
admitted to the hospital | 0 | 0 
fever | -72 | 0 
vomiting | -72 | 0 
generalized abdominal pain | -72 | 0 
rash on palms and trunk | 0 | 0 
severe drowsiness | 0 | 0 
lethargy | 0 | 0 
no conjunctivitis | 0 | 0 
no lymphadenopathy | 0 | 0 
respiratory rate 25/min | 0 | 0 
oxygen saturation 93% | 0 | 0 
harsh breathing with crackles | 0 | 0 
tachycardia | 0 | 0 
hypotension | 0 | 0 
abdomen tender to palpation | 0 | 0 
right lower quadrant tenderness | 0 | 0 
white blood cell count 13.5 × 10^3/μL | 0 | 0 
red blood cell count 3.5–5.8 × 10^6/mm^3 | 0 | 0 
erythrocyte sedimentation rate 82 mm/h | 0 | 0 
C-reactive protein 298.5 mg/L | 0 | 0 
procalcitonin 18.45 mcg/L | 0 | 0 
abdominal ultrasound showing enlarged appendix | 0 | 0 
emergency laparotomy appendectomy | 0 | 24 
postoperative course toxic | 24 | 48 
hemodynamic implications | 24 | 48 
tachycardia | 24 | 48 
hypotension | 24 | 48 
fractional shortening | 24 | 48 
oxygen therapy | 24 | 72 
bronchopneumonia | 24 | 72 
ceftriaxone and amikacin treatment | 24 | 72 
imipenem treatment | 48 | 72 
positive history of contact with COVID-19 | 0 | 0 
positive serology of SARS-CoV-2 | 24 | 24 
ferritin elevated | 24 | 24 
IL6 elevated | 24 | 24 
high-sensitivity troponin elevated | 24 | 24 
D-dimer elevated | 24 | 24 
enoxaparin treatment | 24 | 72 
IV immunoglobulin treatment | 48 | 72 
aspirin treatment | 48 | 168 
red blood cell transfusion | 48 | 48 
systemic corticosteroids treatment | 72 | 168 
dobutamine treatment | 72 | 120 
vasoactive drugs discontinued | 120 | 120 
afebrile | 96 | 168 
clinical symptoms improved | 96 | 168 
arterial pressure stable | 96 | 168 
no pathogenic agents detected | 96 | 168 
histopathological examination showing catarrhal appendicitis | 168 | 168 
D-dimer downward trend | 168 | 168 
troponemia resolved | 168 | 168 
inflammatory parameters normal | 168 | 168 
LV function improved | 168 | 168 
discharged | 168 | 168 
follow-up outpatient visit | 336 | 336 
blood tests normalized | 336 | 336 
COV-2 IgG elevated | 336 | 336 
abdominal and cardiac ultrasounds normal | 336 | 336 
follow-up outpatient visits planned | 336 | 720