33-week gestation | 0
    preterm | 0
    male | 0
    delivered through precipitous vaginal delivery | 0
    respiratory distress | 0
    intubated | 0
    mechanically ventilated | 0
    surfactant | 0
    caffeine | 0
    apnea of prematurity | 0
    ampicillin | 0
    amikacin | 0
    concern of neonatal sepsis | 0
    hypotensive | -72
    normal saline boluses | -72
    dobutamine drip | -72
    increased concern for sepsis | -72
    cefepime | -72
    negative blood cultures | 72
    clinical condition improved | 72
    antibiotics discontinued | 72
    routine cranial ultrasound normal | 72
    echocardiogram normal | 72
    cranial circumference 31 cm | 72
    normal neurological examination | 72
    abdominal distention | 144
    pain on examination | 144
    necrotizing enterocolitis suspected | 144
    vancomycin | 144
    meropenem | 144
    pneumatosis intestinalis not observed | 144
    portal venous gas not observed | 144
    negative blood cultures | 144
    2 weeks antimicrobial treatment | 144
    clinical improvement | 144
    enteral feedings started | 144
    cranial circumference increased to 34 cm | 432
    bulging anterior fontanelle | 432
    alert | 432
    active | 432
    normal neurological examination | 432
    cefepime initiated | 432
    hypernatremia | 432
    enteral sterile water drip | 432
    ventricular puncture | 432
    CSF collected | 432
    no leukocytes in CSF | 432
    CSF glucose decreased | 432
    CSF protein elevated | 432
    cranial ultrasound hydrocephalus | 432
    no intraventricular hemorrhage | 432
    no mass seen | 432
    MRI hydrocephalus | 432
    right frontoparietal cerebral arteriovenous malformation | 432
    MR angiography confirmed mycotic aneurysm | 432
    Candida lusitaniae isolated | 504
    methicillin-resistant Staphylococcus epidermidis | 504
    vancomycin | 504
    amphotericin B | 504
    neurosurgery consulted | 504
    severe apnea | 504
    hypotonia | 504
    lethargy | 504
    resuscitation failed | 504
    aneurysm rupture suspected | 504
    death | 504
    