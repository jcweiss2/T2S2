61 years old | 0
male | 0
dyspnea | -120
fever | -120
COVID-19 | 0
hospitalized | 0
bilateral lung infiltrates | 0
severe dyspnea | 0
hydroxychloroquine | 0
azithromycin | 0
favipiravir | 0
clinical deterioration | 144
ICU admission | 144
tachypnea | 144
high oxygen demand | 144
moderate respiratory distress | 144
oxyhemoglobin saturation 91% | 144
CRS | 144
severe lymphopenia 100/mm3 | 144
hyperferritinemia 1271 ng/mL | 144
prone positioning | 144
high-flow oxygen support | 144
first dose tocilizumab 400 mg IV | 144
acute hypoxemic respiratory failure | 168
second dose tocilizumab | 168
intubation | 168
worsening hypoxemia | 168
accessory muscle use | 168
paradoxical abdominal respiration | 168
central venous catheter placement | 168
mechanical ventilation | 168
extubation | 264
ICU discharge | 264
right shoulder pain | 288
chest pain | 288
pain radiating to right arm | 288
pain exacerbated by sneezing | 288
pain exacerbated by coughing | 288
pain exacerbated by deep breathing | 288
pain exacerbated by movements | 288
afebrile | 288
normal bilateral upper extremity strength | 288
normal glenohumeral range of motion | 288
painful active right shoulder movements | 288
painful passive right shoulder movements | 288
right parasternal redness | 288
right parasternal warmth | 288
right parasternal swelling | 288
costochondral joint pain | 288
referred pain distribution | 288
unremarkable chest radiograph | 288
elevated CRP 15 mg/L | 288
normal leukocyte count | 288
moderate lymphopenia 1000/mm3 | 288
bilateral diffuse ground glass opacities | 288
crazy-paving pattern | 288
consolidation | 288
subcutaneous swelling second and third right costal cartilage | 288
right glenohumeral joint degeneration | 288
Tietze syndrome diagnosis | 288
paracetamol 1g/day for 3 days | 288
progressive pain increase | 288
pain spread to neck | 288
diclofenac 50 mg q.i.d. | 288
tramadol 50 mg q.i.d. | 288
IV methylprednisolone 40 mg for 3 days | 288
sternoclavicular joint swelling | 288
sternoclavicular joint redness | 288
sternoclavicular joint tenderness | 288
MRI chest and right shoulder | 288
fluid collection right sternoclavicular joint | 288
chest cavity abscess | 288
chest wall abscess | 288
inflammatory changes post-contrast MRI | 288
central avascular area in abscess | 288
CT-guided aspiration | 288
purulent liquid 10 mL | 288
Gram stain PMNs without bacteria | 288
acid-fast stain negative | 288
MSSA culture | 288
beta-lactam allergy | 288
IV linezolid for 2 weeks | 288
clindamycin 300 mg t.i.d. | 288
decreased abscess diameter at follow-up | 576
decreased abscess content at follow-up | 576
