33 years old | 0
    woman | 0
    abnormal uterine bleeding | -4320
    endometrial ablation | -4320
    dysuria | -4320
    grayish vaginal discharge | -4320
    malodorous vaginal discharge | -4320
    white blood cell count 16 × 103 cells/mm³ | 0
    hematocrit 39% | 0
    levofloxacin prescribed | 0
    hospitalized | 72
    multiple syncopal events | 72
    blood pressure 74/24 mmHg | 0
    afebrile | 0
    no rash | 0
    cool extremities | 0
    obesity | 0
    benign abdominal exam | 0
    no cervical motion tenderness | 0
    no cervical discharge | 0
    no pelvic abnormality | 0
    negative urine β-human chorionic gonadotropin | 0
    white blood cell count 60 × 103 cells/mm³ | 0
    hematocrit 42% | 0
    platelets 38 × 103 cells/mm³ | 0
    lactate 6.5 mmol/L | 0
    CT scan abdomen and pelvis showing ascites | 0
    pelvic ultrasound unremarkable | 0
    empiric antibiotic therapy with vancomycin | 0
    empiric antibiotic therapy with cefepime | 0
    empiric antibiotic therapy with metronidazole | 0
    transferred to intensive care unit | 0
    white blood cell count 113 × 103 cells/mm³ | 12
    hematocrit 58% | 12
    received 12 liters IV normal saline | 12
    lactate 13.5 mmol/L | 12
    tobramycin added | 12
    clindamycin added | 12
    doxycycline added | 12
    vasopressor support | 0
    required massive IV fluid resuscitation | 24
    received 26 liters IV fluid in first 24 hours | 24
    received 51 liters IV fluid by 72 hours | 72
    disseminated intravascular coagulation (DIC) | 72
    received 46 units blood product | 72
    pericardial effusion | 0
    cardiac tamponade | 0
    pericardial drain placement | 0
    removal of 1500 mL transudative fluid | 0
    bilateral pleural effusions | 0
    bilateral chest tube placement | 0
    4 liters per day transudative fluid output | 0
    exploratory laparotomy | 0
    negative for intra-abdominal infection | 0
    negative for viscous perforation | 0
    massive ascites | 0
    hyperemic uterus | 0
    no vaginal Staphylococcus aureus | 0
    no vaginal yeast | 0
    negative cervical gonorrhea | 0
    negative cervical chlamydia | 0
    marked neutrophilia | 0
    no hematologic malignancy | 0
    negative bone marrow biopsy for malignancy | 0
    negative HIV-1 antibody | 0
    negative blood cultures | 0
    negative urine cultures | 0
    negative pleural fluid cultures | 0
    negative pericardial fluid cultures | 0
    negative peritoneal fluid cultures | 0
    negative sputum cultures | 0
    profound anasarca | 0
    unable to perform repeat pelvic exam | 0
    unable to perform ophthalmologic exam | 0
    clinical picture consistent with toxin-mediated process | 0
    suspected Clostridium sordellii | 0
    plasmapheresis started on hospital day 3 | 72
    improvement in hemodynamics | 72
    fluid removal with venovenous hemofiltration | 72
    edema improved | 96
    pupils fixed and dilated | 96
    CT head scan showing diffuse cerebral edema | 96
    CT head scan showing tonsillar herniation | 96
    family meeting convened | 96
    life support withdrawn | 96
    death | 96
    autopsy showing diffuse edema | 96
    autopsy showing DIC in all organs | 96
    diffuse endometrial necrosis | 96
    Gram-positive rods in endometrial tissue | 96
    Clostridium species confirmed | 96
    negative C sordellii PCR | 96
    positive Clostridium bifermentans PCR | 96
    negative postmortem endometrial cultures | 96