59 years old | 0 | 0 
female | 0 | 0 
blood type O | 0 | 0 
Rh positive | 0 | 0 
liver cancer | -672 | 0 
transarterial embolization | -336 | -336 
sorafenib | -304 | -168 
dizziness | -168 | -168 
skin ulcers | -168 | -168 
radiation therapy | -14 | -14 
Piggyback LT | 0 | 0 
hepatitis B | 0 | 0 
entecavir | 0 | 0 
HBV serology test | 0 | 0 
HBsAg | 0 | 0 
anti-HBs | 0 | 0 
HBeAg | 0 | 0 
anti-HBe | 0 | 0 
anti-HBc | 0 | 0 
human immunodeficiency virus | 0 | 0 
hepatitis A | 0 | 0 
hepatitis C | 0 | 0 
donor | 0 | 0 
21 years old | 0 | 0 
male | 0 | 0 
blood type O | 0 | 0 
Rh positive | 0 | 0 
HLA class-I | 0 | 0 
HLA class-II | 0 | 0 
A11 | 0 | 0 
A30 | 0 | 0 
B13 | 0 | 0 
DR11 | 0 | 0 
DR15 | 0 | 0 
DQ6 | 0 | 0 
DQ7 | 0 | 0 
A2 | 0 | 0 
B13 | 0 | 0 
B46 | 0 | 0 
DR14 | 0 | 0 
DR15 | 0 | 0 
DQ5 | 0 | 0 
DQ6 | 0 | 0 
blood products | 0 | 0 
irradiated | 0 | 0 
filtered | 0 | 0 
transfusion | 0 | 0 
transplantation process | 0 | 0 
acute renal failure | 0 | 24 
hematoma | 0 | 24 
hepatitis B immunoglobulin | 24 | 24 
immunosuppressive drugs | 24 | 0 
steroids | 24 | 0 
tacrolimus | 24 | 0 
hemodialysis | 24 | 168 
fresh frozen plasma | 24 | 168 
leukocyte-depleted red blood cells | 24 | 168 
active bleeding | 24 | 168 
renal function | 168 | 0 
pathological analyses | 168 | 168 
HCC | 168 | 168 
massive tumor necrosis | 168 | 168 
liver function | 240 | 0 
AST | 240 | 0 
ALT | 240 | 0 
GGT | 240 | 0 
ALP | 240 | 0 
fever | 240 | 408 
PCT | 240 | 312 
rash | 408 | 504 
obscure red spots | 408 | 408 
itching | 408 | 408 
Nikolsky sign | 408 | 408 
tacrolimus | 408 | 408 
sirolimus | 408 | 408 
mycophenolate mofetil | 408 | 408 
sputum culture | 408 | 408 
Acinetobacter baumannii | 408 | 408 
MRSA | 408 | 408 
erythematous macules | 456 | 456 
papules | 456 | 456 
limbs | 456 | 456 
palms | 456 | 456 
neck | 456 | 456 
face | 456 | 456 
oral examination | 456 | 456 
white ulcers | 456 | 456 
buccal mucosa | 456 | 456 
lips | 456 | 456 
bone marrow suppression | 456 | 456 
WBC | 456 | 456 
PLT | 456 | 456 
HGB | 456 | 456 
intensive care unit | 456 | 456 
dermatologist | 456 | 456 
gamma globulin | 456 | 456 
skin biopsy | 456 | 456 
FISH | 456 | 456 
peripheral blood | 456 | 456 
abdominal incision | 504 | 504 
sutured | 504 | 504 
bone marrow aspiration | 576 | 576 
bone marrow pathology | 576 | 576 
granulocytes | 576 | 576 
red blood cells | 576 | 576 
megakaryocytes | 576 | 576 
macrophages | 576 | 576 
neutrophils | 576 | 576 
platelets | 576 | 576 
bone marrow cell | 576 | 576 
megakaryocyte | 576 | 576 
platelet | 576 | 576 
FISH analysis | 600 | 600 
donor lymphocytes | 600 | 600 
skin biopsy | 600 | 600 
epidermal dyskeratosis | 600 | 600 
basic vacuolization | 600 | 600 
lymphocytic infiltrates | 600 | 600 
GVHD | 600 | 600 
differential diagnoses | 600 | 600 
bacterial | 600 | 600 
fungal | 600 | 600 
viral | 600 | 600 
drug reactions | 600 | 600 
toxic epidermal necrolysis | 600 | 600 
hemophagocytic syndrome | 600 | 600 
blood culture | 600 | 600 
virus | 600 | 600 
serological tests | 600 | 600 
MDT | 600 | 600 
steroids | 600 | 600 
tacrolimus | 600 | 600 
G-CSF | 600 | 600 
meropenem | 600 | 600 
voriconazole | 600 | 600 
rash | 600 | 720 
general condition | 600 | 720 
ferritin | 720 | 720 
esophageal | 720 | 720 
oral ulcers | 720 | 720 
temperature | 840 | 840 
hallucinations | 840 | 840 
skin | 840 | 840 
bone marrow | 840 | 840 
mucosal epithelium | 840 | 840 
immunodeficiency | 840 | 840 
infections | 840 | 840 
MRSA | 840 | 840 
Acinetobacter baumannii | 840 | 840 
Enterococcus faecalis | 840 | 840 
septic shock | 1008 | 1008 
MODS | 1008 | 1008 
death | 1008 | 1008