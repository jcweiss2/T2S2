47 years old | 0
female | 0
admitted to the hospital | 0
skin ecchymosis | 0
vaginal bleeding | 0
white blood cell count of 7.91×10^9/l | 0
hemoglobin level of 84 g/l | 0
platelet count of 14×10^9/l | 0
prothrombin time 16.9 s | 0
activated partial thromboplastin time 40.7 s | 0
fibrinogen level 1.66 g/l | 0
d-dimer level 20 μg/mL | 0
bone marrow smear hypercellularity | 0
96.5% abnormal promyelocytic granulocytes | 0
Auer bodies | 0
strongly positive peroxidase staining | 0
immunophenotype positivity for myeloperoxidase | 0
CD13 positivity | 0
CD33 positivity | 0
HLA-DR positivity | 0
CD56 positivity | 0
initial diagnosis of APL | 0
treatment with ATRA | 0
treatment with ATO | 0
chest tightness | 336
dyspnea | 336
systemic edema | 336
pleural effusion | 336
differentiation syndrome | 336
chest computed tomography scan | 336
color Doppler ultrasound | 336
white blood cell count 9.4×10^9/l | 336
hemoglobin level 59 g/l | 336
platelet count 38×10^9/l | 336
prothrombin time 18.3 s | 336
fibrinogen level 0.91 g/l | 336
d-dimer level 20 μg/mL | 336
karyotype 45, X, –X, del(9)(q13q22), t(11;12)(p15;q13) | 336
PML–RARA fusion transcript negative | 336
IDH2 mutation 37.68% | 336
TET2 mutation 49.72% | 336
ASXL1 mutation 100% | 336
TP53 mutation 54.75% | 336
WT1-exon7 mutation 100% | 336
WT1-exon9 mutation 43.77% | 336
discontinuation of ATRA | 336
discontinuation of ATO | 336
diuretic detumescence | 336
ventilator-assisted respiratory therapy | 336
second bone marrow smear 95.5% abnormal promyelocytic granulocytes | 336
occasional Auer body | 336
positive peroxidase staining 100% | 336
no remission | 336
complete resistance to ATRA | 336
complete resistance to ATO | 336
switched to IA regimen | 336
idarubicin | 336
cytarabine | 336
severe pulmonary infection | 336
antibiotics for 2 weeks | 336
infection controlled | 336
low WBC count | 336
low platelet count | 336
third bone marrow smear 10.5% blasts | 336
HIAG chemotherapy regimen | 336
homoharringtonine | 336
GCSF | 336
complete remission | 336
consolidation therapy with HIAG regimen | 1464
severe pulmonary infection | 1464
septic shock | 1464
metabolic acidosis | 1464
heart failure | 1464
intensive care unit admission | 1464
recovered after 1 month | 1464
refusal of allo-HSCT | 1464
two cycles of half-dose CAG regimen | 1872
aclarubicin hydrochloride | 1872
cytarabine | 1872
GCSF | 1872
two cycles of HA regimen | 1872
homoharringtonine | 1872
minimal residual disease negative | 1872
leukemia-free at 24-month follow-up | 4320
