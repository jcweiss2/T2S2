82 years old | 0
male | 0
hypertension | 0
tobacco consumption | 0
alcohol consumption | 0
axillary lymph node growth | -8760
cervical lymph node growth | -8760
biopsy | -8760
metastatic MCC diagnosis | -8760
staging PET 68-Ga DOTANOC | -8760
supradiaphragmatic lymph node metastases | -8760
pembrolizumab treatment start | -8760
objective clinical response | -8760
acute anorexia | -8760
mental confusion | -8760
emergency department referral | -8760
obnubilated | -8760
dehydrated | -8760
hyperglycemia (1,350 mg/dL) | -8760
acute kidney injury grade 3 | -8760
hyponatremia | -8760
hypercalcemia | -8760
hyperphosphatemia | -8760
ketonuria (20 mg/dL) | -8760
respiratory arrest | -8760
bradycardia | -8760
hypotension | -8760
orotracheal intubation | -8760
mechanic ventilation | -8760
aminergic support | -8760
mixed metabolic acidemia | -8760
ICU admission | -8760
progressive clinical stability | -8760
increased amylase | -8760
increased lipase | -8760
low C peptide (0.4 ng/mL) | -8760
no anti-GAD antibodies | -8760
no anti-TPO antibodies | -8760
no anti-Tg antibodies | -8760
normal pituitary function | -8760
normal thyroid function | -8760
diabetic ketoacidosis diagnosis | -8760
inaugural insulinopenic type 1 diabetes | -8760
possible pancreatitis | -8760
intensive insulin therapy | -8760
support therapy | -8760
oncology ward transfer | -8760
clinical condition improvement | -8760
corticosteroid therapy | -8760
insulin therapy | -8760
immunotherapy discontinuation | -8760
basal bolus insulin therapy (30 U/day) | -8760
dysarthria | 0
ataxia | 0
oncology ward admission | 0
chest-abdomen-pelvis computed tomography | 0
partial response | 0
axillary lymph node metastasis persistence | 0
brain MRI | 0
neural-axis MRI | 0
electromyography | 0
mild axonal sensorimotor polyneuropathy | 0
ANA positive (≥1/640) | 0
other autoimmune markers negative | 0
vitamin assays negative | 0
viral serologies negative | 0
lumbar puncture | 0
slight proteinorachia (54 mg/dL) | 0
absent pleocytosis | 0
intrathecal antibody synthesis | 0
mirror banding profile (pattern 4) | 0
cytology negative | 0
immunofluorescence assay | 0
fine granular IgG staining | 0
immunoblot negative | 0
recombinant cells negative | 0
methylprednisolone pulse therapy | 0
worsening dysarthria | 24
worsening ataxia | 24
dysphagia | 24
readmission | 24
methylprednisolone cycle | 24
intravenous immunoglobulin | 24
no clinical response | 24
nasogastric tube placement | 24
gastric mucosa infiltration | 24
MCC progression | 24
palliative care | 24
death | 720
