8 years old | 0
female | 0
spayed | 0
domestic shorthair cat | 0
admitted to the hospital | 0
lethargy | -23
pain | -23
elevated body temperature | 0
hypotensive | 0
tachypneic | 0
puncture wounds | 0
mild hyperglycemia | 0
normal white blood cell count | 0
normal packed cell volume | 0
normal total protein | 0
negative for retroviral disease | 0
mild diffuse bronchointerstitial pulmonary pattern | 0
normal abdomen | 0
normal skeletal structures | 0
soft tissue swelling | 0
gas noted dorsal to the lumbar spine | 0
cellulitis | 0
intravenous crystalloid fluid boluses | 0
lactated Ringer’s solution | 0
buprenorphine | 0
hospitalization declined | 0
discharged home | 0
oral transmucosal buprenorphine | 0
oral amoxicillin/clavulanic acid | 0
re-presented to the hospital | 23
obtunded | 23
hypoglycemic | 23
septic suppurative inflammation | 23
subcutaneous fluid pocket | 23
aerobic culture | 23
abdominal ultrasound | 23
normal venous blood gas | 23
admitted to the intensive care unit | 23
ampicillin–sulbactam | 23
enrofloxacin | 23
metronidazole | 23
vitamin C | 23
maropitant citrate | 23
famotidine | 23
fentanyl constant rate infusion | 23
dextrose | 23
LRS with 5% dextrose and 40 meq/l potassium chloride | 23
sedated with fentanyl and midazolam | 23
wound debrided and lavaged | 23
wet-to-dry tie over bandage | 23
double-lumen catheter | 23
indwelling urinary catheter | 23
attempt to place an arterial catheter | 23
norepinephrine CRI | 23
dopamine CRI | 23
vasopressin CRI | 23
hydrocortisone CRI | 23
more responsive | 48
able to lift its head | 48
dextrose supplementation discontinued | 48
wet-to-dry bandage replaced | 48
IV enrofloxacin, ampicillin–sulbactam, metronidazole, maropitant, hydrocortisone CRI and vitamin C continued | 48
norepinephrine, dopamine and vasopressin CRIs continued | 48
dopamine dose decreased | 48
norepinephrine dose decreased | 48
vasopressin dose unchanged | 48
able to maintain sternal recumbency | 72
ate a small amount of food | 72
motor function and pain sensation present | 72
unable to stand or walk | 72
less painful | 72
fentanyl CRI decreased | 72
wet-to-dry bandage changed | 72
norepinephrine and vasopressin doses decreased | 72
CRIs eventually discontinued | 72
MAP stayed between 70 and 80 mmHg | 72
anesthetized | 120
7 mm Jackson-Pratt drain placed | 120
wound closed | 120
briefly hypotensive | 120
treated with dopamine | 120
hypotension resolved | 120
dopamine discontinued | 120
recheck PCV | 120
anemia suspected | 120
blood type performed | 120
given one unit of compatible feline packed red blood cells | 120
started eating readily | 120
transitioned to oral amoxicillin/clavulanic acid, enrofloxacin and OTM buprenorphine | 120
culture of the wound reported | 120
oral enrofloxacin discontinued | 120
paws on the right thoracic and right pelvic limbs became swollen | 144
edematous and cold to the touch | 144
right cephalic IV catheter and right dorsal pedal arterial catheters removed | 144
vascular access via the central venous catheter maintained | 144
paws continued to be cold to the touch, painful and became discolored | 168
skin on the paw pads started to slough | 168
line of demarcation dividing affected tissue and normal healthy skin noted | 168
strong pedal pulses detected | 168
clopidogrel started | 168
normotensive | 168
continued wound care | 168
daily wet-to-dry bandage changes | 168
hydrotherapy | 168
discharged | 264
soft padded bandages in place | 264
paws fully healed | 336
ambulatory with mild residual pelvic limb weakness | 336