60 years old | 0
male | 0
nonsmoker | 0
admitted to the hospital | 0
facial edema | -480
neck edema | -480
right upper limb edema | -480
mass on right chest | -480
computed tomography scan | 0
retroperitoneal lymphadenopathy | 0
pericardial effusion | 0
metastases in mediastinum | 0
bilateral adrenal gland metastases | 0
right thoracic wall nodule | 0
multiple bone metastases | 0
fecal examination for occult blood | 0
biopsy of right thoracic wall nodule | 0
low differentiated lung adenocarcinoma | 0
pemetrexed and nedaplatin for chemotherapy | 0
acute abdominal pain | 168
acute peritonitis | 168
abdominal CT scan | 168
free air in peritoneal cavity | 168
massive ascites | 168
emergency surgery | 168
dirty ascites | 168
hyperemia and edema in small intestinal wall | 168
pus adhesion in omentum and small intestine surface | 168
grey nodules in mesentery | 168
perforations of jejunum | 168
intestinal resection | 168
end-to-end anastomosis | 168
pathological diagnosis of metastatic lung adenocarcinoma | 168
immunohistochemical analysis | 168
tumor cells positive for CK7 and TTF-1 | 168
septic shock | 360
death | 360