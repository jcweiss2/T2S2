74 years old | 0 | 0 
male | 0 | 0 
hypertension | 0 | 0 
insulin-dependent diabetes mellitus type 2 | 0 | 0 
diabetic retinopathy | 0 | 0 
weight loss | -168 | 0 
iron deficiency anemia | -168 | 0 
tumor in the colon ascendens | -168 | 0 
liver metastases | -168 | 0 
right hemicolectomy | 0 | 0 
low-grade pT3cN0 adenocarcinoma | 0 | 0 
absence of metastases in 24 excised lymph nodes | 0 | 0 
lymphovascular growth | 0 | 0 
no vascular or perineural growth | 0 | 0 
activated BRAF mutation in exon 15 (V600E) | 0 | 0 
loss of expression of MLH1 and PMS2 | 0 | 0 
mismatch repair-deficient (MMR-D)/microsatellite-instable (MSI) tumor | 0 | 0 
initiated therapy with pembrolizumab | 0 | 0 
symptoms of a cold | -168 | 7 
leukocytosis | -168 | 7 
slight increase in C-reactive protein | -168 | 7 
dry coughing | 7 | 22 
no fever | 7 | 22 
increase in AST and ALT | 7 | 22 
ICI-induced hepatitis grade 2 | 7 | 22 
initiated prednisolone therapy | 22 | 22 
decrease in C-reactive protein and AST | 22 | 29 
increase in white blood cells and neutrophils | 22 | 29 
dyspnea | 22 | 29 
elevation of troponin T | 22 | 29 
septal hypokinesia | 22 | 29 
no dynamic change over time in troponin T | 22 | 29 
somnolence | 29 | 29 
difficulty walking | 29 | 29 
dysarthria | 29 | 30 
hoarseness | 29 | 30 
pain in neck and right leg | 29 | 30 
difficulty raising right leg | 29 | 30 
increased dose of prednisolone | 30 | 30 
no signs of stroke | 30 | 30 
increased creatine kinase and myoglobin levels | 30 | 30 
ICI-induced myositis | 30 | 30 
gradual decrease in creatinine levels | 30 | 30 
antibodies against acetylcholine receptor and titin | 30 | 30 
albumin in cerebrospinal fluid | 30 | 30 
unable to sit up | 30 | 34 
severe dysarthria and dysphagia | 30 | 34 
absent reflexes | 30 | 34 
intubated | 34 | 34 
given methylprednisolone | 34 | 37 
given intravenous immunoglobulins | 34 | 37 
given infliximab | 37 | 37 
better muscle strength in hands | 37 | 38 
carbon dioxide retention | 38 | 39 
noninvasive ventilation | 38 | 39 
sinus bradycardia | 38 | 39 
death | 39 | 39 
significant stenosis of the right coronary artery | 39 | 39 
no fibrosis or signs of recent myocardial infarction | 39 | 39 
softened tongue | 39 | 39 
no surgical complication after hemicolectomy | 39 | 39 
metastasis in the right liver lobe | 39 | 39 
pronounced inflammatory infiltration of lymphocytes | 39 | 39 
fibrosis in the intercostal musculature, diaphragm, cervical musculature and tongue | 39 | 39 
hepatocellular cancer (HCC) | 39 | 39 
fibrosis stage 2–3 according to Batts and Ludwig | 39 | 39 
respiratory insufficiency due to polymyositis | 39 | 39