67 years old | 0
    African-American man | 0
    achy, non-radiating pain in his chest | -72
    acute left foot pain | -72
    fatigue | -72
    malaise | -72
    chest pain aggravated by deep breathing | 0
    chest pain aggravated by coughing | 0
    chest pain aggravated by sitting up | 0
    chest pain aggravated by moving | 0
    denied nausea | 0
    denied vomiting | 0
    denied sweating | 0
    End Stage Renal Disease (ESRD) | -157248
    hemodialysis via right femoral catheter | -26208
    non-ischemic heart failure with reduced ejection fraction | 0
    pericardial effusion | 0
    low-grade follicular cell lymphoma | 0
    non-compliant with outpatient chemotherapy | -17472
    stroke | 0
    deep vein thrombosis (DVT) | 0
    pulmonary embolism (PE) | 0
    paroxysmal atrial fibrillation | 0
    chronic obstructive pulmonary disease (COPD) | 0
    hepatitis C infection | 0
    chronic anemia | 0
    medication non-adherence | 0
    multiple dialysis catheter placements | 0
    AV fistula creation | 0
    atrial flutter ablation | 0
    hernia repair | 0
    nuclear stress test | -8760
    ejection fraction of 27% | -8760
    elevated troponin of 0.965 | 0
    troponin decreased to 0.674 | 72
    White Blood Cell (WBC) count of 9.0 × 103/mL | 0
    71.3% neutrophils | 0
    ECG no changes compared to previous studies | 0
    nuclear stress test showed LV ejection fraction of 17% | 72
    moderate size perfusion defect in the inferior wall | 72
    mild to moderate severity perfusion defect in the inferior wall | 72
    reversible apical inferior wall ischemic changes | 72
    two episodes of low-grade fever | 48
    maximum temperature of 38.1 °C | 48
    blood cultures drawn from peripheral veins | 48
    growth of gram-positive rods (diphtheroid) | 48
    transthoracic echocardiogram | 48
    mobile echo-density measuring 2.9 cm | 48
    vegetation on mitral valve chordae | 48
    severe mitral annular calcification | 48
    moderate mitral regurgitation | 48
    mild mitral stenosis | 48
    mildly thickened aortic valve leaflets | 48
    aortic annular calcification | 48
    mild to moderate tricuspid regurgitation | 48
    repeat blood cultures | 72
    isolation of the same organism | 72
    vancomycin started during hemodialysis | 72
    femoral permcath replaced by temporary trialysis catheter | 72
    samples sent to Mayo Clinic | 72
    organism identified as Corynebacterium jeikeium | 72
    resistant to penicillin | 72
    resistant to ceftriaxone | 72
    resistant to meropenem | 72
    sensitive to vancomycin | 72
    vancomycin continued | 72
    repeated blood cultures | 120
    still positive for diphtheroid | 120
    cultures became negative | 216
    new femoral permcath inserted | 216
    discharged | 216
    Corynebacterium jeikeium endocarditis | 72
    vancomycin continued with each dialysis session for 6 weeks | 216
    fully recovered | 216
    dialysis catheter malfunction | 4032
    no out-patient repeat echocardiogram | 4032

    