59 years old | 0
female | 0
blood type O | 0
Rh positive | 0
admitted to the hospital | 0
segment-V space-occupying lesion | -365
liver cancer | -365
transarterial embolization | -365
sorafenib | -304
dizziness | -91
skin ulcers | -91
computed tomography scan | -30
radiation therapy | -14
Piggyback LT | 0
hepatitis B | 0
entecavir | 0
HBV serology test | 0
hepatitis B virus | 0
human immunodeficiency virus | 0
hepatitis A | 0
hepatitis C | 0
donor | 0
brain death | 0
car accident | 0
HLA class-I | 0
HLA class-II | 0
blood products | 0
irradiated | 0
filtered | 0
transplantation process | 0
acute renal failure | 24
hematoma | 24
hepatitis B immunoglobulin | 24
immunosuppressive drugs | 24
steroids | 24
tacrolimus | 24
hemodialysis | 48
fresh frozen plasma | 48
leukocyte-depleted red blood cells | 48
active bleeding | 48
renal function | 120
pathological analyses | 120
HCC | 120
massive tumor necrosis | 120
liver function | 240
improvement | 240
fever | 240
procalcitonin | 240
PCT | 240
rash | 312
obscure red spots | 312
chest | 312
no itching | 312
Nikolsky sign | 312
negative | 312
tacrolimus | 408
sirolimus | 408
mycophenolate mofetil | 408
immune suppression | 408
sputum culture | 408
Acinetobacter baumannii | 408
methicillin-resistant Staphylococcus aureus | 408
MRSA | 408
rash advanced | 456
erythematous macules | 456
papules | 456
limbs | 456
palms | 456
neck | 456
face | 456
oral examination | 456
white ulcers | 456
buccal mucosa | 456
lips | 456
bone marrow suppression | 456
severe | 456
WBC count | 456
platelet count | 456
hemoglobin | 456
intensive care unit | 456
dermatologist | 456
gamma globulin | 456
skin biopsy | 456
fluorescence in situ hybridization | 456
FISH | 456
peripheral blood | 456
abdominal incision | 552
split | 552
sutured | 552
bone marrow aspiration | 624
bone marrow pathology | 624
no special lesions | 624
granulocytes | 624
red blood cells | 624
megakaryocytes | 624
macrophages | 624
neutrophils | 624
platelets | 624
bone marrow cell morphology | 624
proliferating | 624
active | 624
megakaryocyte production | 624
reduced | 624
platelet levels | 624
decreased | 624
FISH analysis | 624
donor lymphocytes | 624
skin biopsy specimens | 624
epidermal dyskeratosis | 624
basic vacuolization | 624
lymphocytic infiltrates | 624
grade-1 acute lt-GVHD | 624
differential diagnoses | 624
bacterial infections | 624
fungal infections | 624
viral infections | 624
drug reactions | 624
toxic epidermal necrolysis | 624
hemophagocytic syndrome | 624
blood culture | 624
negative | 624
allergies | 624
drugs | 624
virus | 624
serological tests | 624
macrophages | 624
neutrophils | 624
platelets | 624
bone marrow biopsy | 624
collective findings | 624
clinical course | 624
consistent | 624
diagnosis | 624
lt-GVHD | 624
multidisciplinary team | 680
treatment plan | 680
steroids | 680
tacrolimus | 680
immune suppression | 680
granulocyte colony-stimulating factor | 680
G-CSF | 680
hematopoiesis | 680
meropenem | 680
voriconazole | 680
anti-infective therapy | 680
rash | 680
reduced | 680
general condition | 680
deteriorate | 680
serum ferritin | 680
increased | 680
esophageal ulcers | 680
oral ulcers | 680
worsen | 680
eating | 680
difficulty | 680
temperature | 1128
rose | 1128
hallucinations | 1128
septic shock | 1320
multiple organ dysfunction syndrome | 1320
MODS | 1320
death | 1320