60 years old | 0
man | 0
presented with scrotal pain | -0
fever (103°F) | -0
fatigue | -0
tachycardic (130 beats per minute) | -0
hypotensive (103/40 mm Hg) | -0
started on vancomycin | -0
started on Zosyn | -0
admitted under medicine service | 0
kidney function worsened | 24
switched antibiotics to meropenem | 24
creatinine level continued to rise | 24
prednisone (40 mg daily) | 0
spike fevers | 24
blood cultures negative | 24
urine cultures negative | 24
sputum cultures negative | 24
CT chest negative | 24
CT abdomen negative | 24
CT pelvis negative | 24
antibiotics stopped | 24
macular rash | -168
rash progressed to axillary area | -168
rash involved chest | -168
rash involved head | -168
rash involved neck | -168
rash involved abdomen | -168
incendiary mental status | -168
skin lesions worsened with bullae and vesicles | -168
dermatology team involved | -168
skin biopsy performed | -168
local steroid cream initiated | -168
AGEP diagnosis | -168
rash became pustular | -216
fever (109°F) | -216
transferred to ICU | -216
cooling protocol initiated | -216
pulse steroids administered | -216
fever subsided | -216
rash improvement observed | -216
decreased progression of sloughing | -216
acute kidney injury resolved | -216
steroids tapered | -216
pulse steroids completed | -216
skin biopsy | 0
urine analysis | 0
CT chest/abdomen/pelvis | 0
CBC | 0
BMP | 0
coagulation | 0
differential diagnosis (AGEP, DRESS, von Zumbusch psoriasis, Steven Johnson syndrome, leukocytoclastic vasculitis, Sneddon-Wilkinson disease, cutaneous candidiasis) | 0
PAN | -0
paroxysmal atrial fibrillation | -0
hypertension | -0
dyslipidemia | -0
non-insulin dependent diabetes mellitus | -0
prior admissions for PAN flares | -0
history of septic shock | -17520
prior failure on cyclophosphamide | -0
prednisone treatment | -0
cyclophosphamide treatment | -0
septic shock history | -17520
no calcium channel blockers | 0
negative blood cultures | 24
negative urine cultures | 24
negative sputum cultures | 24
no infection focus found | 24
pulse steroids initiated | -216
immunosuppressive management considered | -216
penicillin avoidance | -216
steroids weaned | -216
supportive care | -216
symptomatic treatment for pruritus and inflammation | -216
systemic corticosteroids used | -216
autoimmune process suspected | -216
T cell-mediated neutrophilic inflammation | -216
CD4+ T cells involvement | -216
cytotoxic CD8+ T cells involvement | -216
inflammatory cytokines and chemokines involved | -216
CXCL8 production | -216
GM-CSF production | -216
reduced neutrophil apoptosis | -216
neutrophil infiltrate on biopsy | -216
dermal edema on biopsy | -216
intra- and subcorneal spongiform | -216
superficial interstitial mid-dermal infiltrate | -216
leukocytosis with neutrophil count >7,000 cells/mm3 | 0
mild eosinophilia | 0
high fever (>38°C) | 0
non-follicular sterile pustules | 0
edematous erythema | 0
acute kidney injury | 0
neutrophilia | 0
cyclic fevers | 0
sloughing progression | -216
mental status decline | -168
bullae and vesicles | -168
axillary area involvement | -168
chest involvement | -168
head involvement | -168
neck involvement | -168
abdomen involvement | -168
ICU transfer | -216
cooling protocol | -216
pulse steroids | -216
pulse steroids completion | -216
steroid taper | -216
rash resolution | -216
kidney injury resolution | -216
fever resolution | -216
systemic manifestations improvement | -216
pruritus | 0
skin inflammation | 0
prior cyclophosphamide failure | -0
prednisone and cyclophosphamide combination | -0
autoimmune etiology considered | -216
PAN flares | -0
immunosuppressive therapy considered | -216
self-limiting AGEP | -216
favorable prognosis | -216
unresponsiveness to antibiotics | -216
negative cultures | 24
clinical suspicion of autoimmune process | -216
use of systemic steroids | -216
dramatic improvement | -216
self-resolving AGEP | -216
prednisone continuation | 0
cyclophosphamide continuation | -0
pulse steroids effectiveness | -216
AGEP as autoimmune manifestation | -216
PAN and AGEP association | -216
T cell proliferation involvement | -216
neutrophilic proliferation involvement | -216
autoimmune process in PAN | -216
severe fevers | -216
ICU admission | -216
kidney involvement | 0
high grade fever | -216
neutropenia | 0
cholestasis | 0
hepatic involvement | 0
no family history of psoriasis | 0
no psoriasis | 0
tender erythematous nodules | 0
purpura | 0
livedo reticularis | 0
ulcers | 0
bullous eruption | 0
vesicular eruption | 0
subcorneal pustular dermatosis (Sneddon-Wilkinson disease) differential | 0
leukocytoclastic vasculitis differential | 0
cutaneous candidiasis differential | 0
DRESS syndrome differential | 0
Steven Johnson syndrome differential | 0
von Zumbusch psoriasis differential | 0
intra- and subcorneal spongiform on biopsy | -216
prior septic shock | -17520
prior PAN flares | -0
prior prednisone use | -0
septic shock 2 years prior | -17520
no identifiable infection source | -17520
no insulin dependent diabetes | 0
biopsy proven PAN | -0
scrotal pain | -0
tachycardic | -0
hypotensive | -0
rash progression | -168
skin lesions worsening | -168
dermatology consultation | -168
AGEP diagnosis confirmed | -168
local steroid cream | -168
rash pustular | -216
high fever (109°F) | -216
cooling | -216
rash improvement | -216
sloughing decreased | -216
kidney injury resolved | -216
CT imaging | 0
coagulation studies | 0
differential diagnoses | 0
no infection focus | 24
immunosuppressive consideration | -216
pruritus treatment | -216
inflammation treatment | -216
autoimmune etiology | -216
PAN association | -216
T cell involvement | -216
neutrophilic proliferation | -216
kidney function recovery | -216
cholestasis excluded | 0
hepatic involvement excluded | 0
psoriasis excluded | 0
skin lesions differentials | 0
biopsy findings | -216
negative candidiasis | 0
unresponsive to antibiotics | -216
prior immunosuppressive failure | -0
autoimmune process management | -216
clinical suspicion high | -216
systemic manifestations | -216
mental status change | -168
AGEP confirmed | -168
improvement observed | -216
self-limiting course | -216
favorable outcome | -216
