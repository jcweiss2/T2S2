45 years old | 0
female | 0
presented to ED | 0
fevers | -168
headache | -168
arthralgias | -168
nausea | -168
fatigue | -168
neck pain | -168
tachycardic | -168
afebrile | -168
no rash | -168
viral illness | -168
discharged from ED | -48
worsening confusion | -48
combativeness | -48
dyspnea | -48
ataxia | -48
multiple recent bug bites | -168
pet dogs not up to date on flea and tick medication | -168
tachycardic | -48
hypotensive | -48
toxic appearance | -48
maculopapular rash | -48
no bites or ticks | -48
low blood pressure | -48
fluid resuscitation | -48
MRI of brain | -48
lumbar puncture | -48
WBC 16/HPF | -48
protein 49 mg/dL | -48
glucose 51 mg/dL | -48
albumin 32.91 mg/dL | -48
RBC 4/HPF | -48
vancomycin | -48
meropenem | -48
acyclovir | -48
doxycycline | -48
fever | -24
admitted to ICU | -24
leukocytosis | -24
lactate 2.1 mmol/L | -24
decreased kidney function | -24
thrombocytopenia | -24
anemia | -24
abnormal liver function | -24
pro time 16.5 sec | -24
prothrombin time 37.4 sec | -24
INR 1.3 | -24
d-dimer 11.28 ug/mL | -24
fibrinogen 268 mg/dL | -24
albumin 2.3 g/dL | -24
intubation | 0
acute hypoxic respiratory failure | 0
chest CT | 0
bilateral pleural effusions | 0
pulmonary alveolar and interstitial edema | 0
atelectasis | 0
echocardiogram | 0
ejection fraction 49% | 0
mildly reduced left ventricular systolic function | 0
mild global hypokinesis | 0
R. typhi IgM 1:1024 | 0
R. Rickettsii IgM 1:1024 | 0
IgG 1:128 | 0
echovirus Ab 1:80 | 0
antibiotics de-escalated | 24
doxycycline | 24
fever resolved | 48
extubated | 48
transferred from ICU to floor | 48
discharged home | 168
doxycycline | 168
resolution of symptoms | 336
no need to repeat titers | 336