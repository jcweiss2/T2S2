73 years old | 0
    female | 0
    hypertension | 0
    syphilis | 0
    type 2 diabetes mellitus | 0
    acute altered mental status | 0
    mechanical fall | -720
    pruritic scalp | -720
    purulent drainage from sinuses on the scalp behind right ear | -720
    temperature 97.9°F | 0
    heart rate 127 bpm | 0
    respiratory rate 22 breaths/min | 0
    blood pressure 144/80 mmHg | 0
    oxygen saturation 98% on room air | 0
    oriented to person | 0
    oriented to place | 0
    not oriented to time | 0
    erythematous face | 0
    erythematous scalp | 0
    erythematous right ear | 0
    edematous face | 0
    edematous scalp | 0
    edematous right ear | 0
    large fluctuant mass over occipital scalp | 0
    large fluctuant mass over parietal scalp | 0
    purulent drainage over occipital scalp | 0
    purulent drainage over parietal scalp | 0
    posterior auricular mass | 0
    no active drainage of posterior auricular mass | 0
    hyperglycemia 700 | 0
    anion gap metabolic acidosis | 0
    serum bicarbonate 20 | 0
    ketonuria | 0
    non-contrast head CT | 0
    extensive multifocal scalp swelling | 0
    right temporal swelling | 0
    right posterior parietal swelling | 0
    left frontal swelling | 0
    no acute intracranial abnormalities | 0
    admitted to ICU | 0
    diabetic ketoacidosis | 0
    cellulitis of the scalp | 0
    concern for underlying abscesses | 0
    continuous infusion of insulin | 0
    broad-spectrum coverage | 0
    intravenous Vancomycin | 0
    intravenous Cefepime | 0
    incision and drainage of scalp lesion | 48
    10-cm subgaleal abscess | 48
    purulence evacuated | 48
    MRSA in blood cultures | 72
    continued intravenous Vancomycin | 72
    continued intravenous Cefepime | 72
    paranasal sinus CT with contrast | 72
    no sinus involvement | 72
    transesophageal echocardiogram | 72
    no endocarditis | 72
    returned to operating room on day 4 | 96
    returned to operating room on day 5 | 120
    pulse irrigation of wounds | 96
    pulse irrigation of wounds | 120
    sharp debridement | 96
    sharp debridement | 120
    plastic surgery involvement | 96
    plastic surgery involvement | 120
    serial bedside debridements | 96
    serial bedside debridements | 120
    scalp wound 20 cm length | 96
    scalp wound 10 cm width | 96
    scalp wound 2 cm depth | 96
    right posterior auricular wound 7 cm x 7 cm x 2 cm | 96
    split-thickness skin grafts from right thigh | 168
    scalp wound closure | 168
    posterior auricular wound closure | 168
    100% graft take on postoperative day 7 | 264
    discharged on day 32 | 768
    intravenous Vancomycin course completion | 768
    7-week course | 768
    no graft rejection | 264
    wound bed free of purulent drainage | 264
    WBC down trending | 264
    sepsis resolving | 264
    hyperpigmentation around graft | 768
    skin graft healed well | 768