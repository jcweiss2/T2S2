33 years old | 0
male | 0
admitted to the hospital | 0
fever | -24
altered mental status | -24
nausea | -48
vomiting | -48
diarrhea | -48
food poisoning | -48
CT of the head | -24
CT of the abdomen | -24
CT of the pelvis | -24
discharged from ER | -24
HIV diagnosed | -2190
CD4+ cell count 1782 cells/mm3 | -720
HIV-1 RNA level < 20 copies/mL | -720
antiretroviral therapy | -1095
dolutegravir/lamivine/abacavir | -1095
vaccinations against Hib | -1095
vaccinations against S. pneumoniae | -1095
vaccinations against N. meningitidis | -1095
nasopharyngitis | -240
Group A Streptococcus test | -240
negative Group A Streptococcus test | -240
supportive care | -240
secondary syphilis | -1095
secondary syphilis | -1095
temperature 39.1 °C | 0
heart rate 114 beats/min | 0
respiratory rate 32 breaths/min | 0
blood pressure 163/94 mm Hg | 0
oxygen saturation 100% | 0
weight 83 kg | 0
body mass index 24.8 | 0
Glasgow Coma Scale score 11 | 0
nuchal rigidity | 0
agitation | 0
pupils equal and reactive to light | 0
dental caries | 0
lactic acid level 14.79 mmol/L | 0
sodium 143 mmol/L | 0
potassium 3.1 mmol/L | 0
chloride 109 mmol/L | 0
CO2 12 mmol/L | 0
BUN 14 mg/dL | 0
creatinine 1.1 mg/dL | 0
glucose 74 mg/dL | 0
calcium 7.9 | 0
anion gap 26 mmol/L | 0
WBC 3.5 × 103/µL | 0
hemoglobin 12.7 g/dL | 0
platelet 95 × 103/µL | 0
INR 1.6 | 0
PT 18.9 s | 0
alkaline phosphatase 226 IU/L | 0
toxicology screen positive for marijuana | 0
ethanol level < 10 mg/dL | 0
CD4+ cell count 182 cells/mm3 | 0
CT of the head unremarkable | 0
blood cultures | 0
lumbar puncture | 0
yellow/turbid cerebrospinal fluid | 0
glucose < 10 mg/dL | 0
protein 1185 mg/dL | 0
WBC 2663/µL | 0
negative cryptococcal antigen | 0
nonreactive VDRL test | 0
Gram smear of CSF fluid | 0
gram-negative diplococci | 0
vancomycin | 0
ceftriaxone | 0
ampicillin | 0
acyclovir | 0
dexamethasone | 0
intubated | 12
increased difficulty breathing | 12
drop in blood pressure | 24
PEA arrest | 24
cardiopulmonary resuscitation | 24
return of spontaneous circulation | 24
vasopressors | 24
dilated and non-reactive pupils | 24
repeat CT of the head | 24
increased edema | 24
increased effacement of basil cisterns | 24
mild increase in temporal horns | 24
unresponsive | 24
EEG complete suppression | 24
expired | 48
NTHi biotype I | 48
autopsy report | 48
cause of death | 48
sepsis | 48
meningitis | 48
NTHi | 48