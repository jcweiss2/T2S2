26 years old | 0
female | 0
nulliparous | 0
severe hypogastric pain | -24
no response to analgesics | -24
uterine myomatosis | -168
prescribed with analgesics | -168
abnormal uterine bleeding | -168
abdominal pain | -168
depressible and tender abdomen | 0
slight increase in volume in the hypogastrium | 0
no abnormal laboratory findings | 0
reverse transcription PCR for severe acute respiratory syndrome coronavirus 2 | 0
negative result | 0
mass located in the posterior wall of the uterus | 0
T1- and T2-weighted hyperintense component | 0
T1-weighted hyperintense halo | 0
materials with high T1-weighted fat-saturation signal | 0
content with high T2-weighted fat-saturation signal | 0
diffusion-weighted images | 0
apparent diffusion coefficient map | 0
low apparent diffusion coefficient value | 0
leiomyoma with red degeneration | 0
pyomyoma | 0
laparoscopic myomectomy | 0
intraoperative large myoma | 0
peripherally hypovascularized | 0
friable tissue in its center | 0
sepsis symptoms | 12
hypotension | 12
tachycardia | 12
fever | 12
respiratory distress | 12
drowsiness | 12
admitted to the intensive care unit | 12
oxygen therapy | 12
fluid resuscitation | 12
empiric antibiotic therapy | 12
anemia | 12
leukocytosis with bandemia | 12
high C-reactive protein levels | 12
procalcitonin | 12
pCO2 | 12
HCO3 | 12
BEb | 12
lactate | 12
histopathologic report | 12
uterine leiomyoma with coagulative and liquefactive necrosis | 12
tissue culture | 12
gram-negative cocci bacteria | 12
antibiotic treatment adjusted | 12
normalization of inflammatory markers | 12
clinical improvement | 12
discharged | 72