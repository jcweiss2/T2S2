65 years old | 0
male | 0
visited general surgery outpatient clinic | 0
presumptive cholangiocarcinoma | 0
previously healthy | 0
unremarkable medical history | 0
preoperative evaluations | 0
complete blood cell counts (CBCs) | 0
chemistry | 0
C-reactive protein (CRP) elevated | 0
total bilirubin | 0
direct bilirubin | 0
MELD score | 0
vital signs within normal limits | 0
axillary body temperature 36.7°C | 0
preoperative chest radiography | 0
transthoracic echocardiography | 0
imaging studies indicated tumor | 0
enlarged lymph node | 0
probable metastasis | 0
bilateral invasion of bile duct | 0
unresectable tumor | 0
planned LDLT | 0
donor hepatectomy | 0
intraoperative frozen biopsy | 0
anesthesia induced | 0
endotracheal intubation | 0
BIS monitoring | 0
arterial cannulation | 0
warming blanket applied | 0
fluid warming system prepared | 0
body temperature monitored | 0
body temperature 36.7°C | 0
retractor placed | 0
inhalant anesthetic changed | 0
anesthesia maintained | 0
sevoflurane gas eliminated | 0
lymph node excised | 0
common bile duct clamped | 0
frozen biopsy specimens negative | 0
LDLT continued | 0
nasogastric tube placed | 0
AVA catheter inserted | 0
pulmonary artery catheter inserted | 0
body temperature 36.9°C | 0
CBT measured | 0
initial CBT 37.6°C | 0
fluid warming system turned off | 0
warming blanket cooling mode | 0
room temperature adjusted | 0
laparoscopic approach | 0
converted to open hepatectomy | 0
CBT rose to 39.5°C | 0
vital signs within normal range | 0
reactive tachycardia | 0
no blood products administered | 0
no medicine except anesthetics | 0
no signs of malignant hyperthermia | 0
ETCO2 within normal range | 0
arterial blood gas analysis normal | 0
no allergic reactions | 0
device error ruled out | 0
preoperative CBCs normal | 0
vital signs normal | 0
chest radiographs normal | 0
thyroid function tests normal | 0
BIS monitored | 0
common bile duct clamping related | 0
bile drained | 0
CBT declined | 0
total duration clamping 5 hours | 0
anhepatic phase began | 0
CBT 37.5°C | 0
CBT decreased to 36.9°C | 0
warming blanket turned on | 0
fluid warming system turned on | 0
CBT maintained | 0
anesthesia time 14 hours | 0
crystalloid administered | 0
colloid administered | 0
albumin administered | 0
cell saver blood administered | 0
urine output | 0
transferred to ICU | 0
tympanic temperature 37.6°C | 0
WBC count increased | 0
CRP stable | 0
total bilirubin increased | 0
direct bilirubin increased | 0
chest radiographs no change | 0
cultures negative | 0
transferred to general ward | 120
fifth postoperative day | 120
no complications | 120
hyperthermia | 0
fever | 0
tachycardia | 0
hypothermia | 0
mild reactive tachycardia | 0
hyperthermia during LDLT | 0
bile congestion | 0
inflammatory response | 0
postoperative labs | 0
postoperative imaging | 0
postoperative monitoring | 0
intraoperative complications | 0
postoperative care | 0
recovery | 0
discharge | 120
