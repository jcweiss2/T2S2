69 years old | 0 | 0 
male | 0 | 0 
admitted to the hospital | 0 | 0 
Child–Pugh class C cirrhosis | 0 | 0 
slipping on wet grass and falling on his left side | -1 | -1 
Glasgow coma score 15/15 | 0 | 0 
vital signs within normal limits | 0 | 0 
pulse rate 78/min | 0 | 0 
RR 13/min | 0 | 0 
BP 113/54 mm Hg | 0 | 0 
SpO2-100% in air | 0 | 0 
left hip tenderness | 0 | 0 
no ecchymosis to the abdomen, flank or thigh | 0 | 0 
radiograph of his pelvis revealed an undisplaced fracture of his left acetabulum | 0 | 0 
liver dysfunction | 0 | 0 
pH 7.271 | 0 | 0 
base excess minus 7.3 | 0 | 0 
PT 18.2 | 0 | 0 
INR-1.5 | 0 | 0 
APTT ratio 1.42 | 0 | 0 
platelets 73 | 0 | 0 
bilirubin 63 mmol/l | 0 | 0 
Hb 124 g/l | 0 | 0 
18 g intravenous cannula inserted | 0 | 0 
warmed Hartmanns one litre infusion commenced | 0 | 0 
referred to the Orthopaedic on call team | 1 | 1 
initial delay due to pressure in the Emergency department | 0 | 1 
blood pressure dropped to 75/51 mm Hg | 2 | 2 
tachycardic | 2 | 2 
serum lactate 9 mmol/l | 2 | 2 
FAST examination revealed intraabdominal fluid | 2 | 2 
treated for sepsis in the Emergency department | 2 | 4 
intensive care, orthopaedic and general registrar attended the patient | 4 | 4 
pH 7.227 | 4 | 4 
base excess of −17.9 | 4 | 4 
serum lactate of 16.3 mmol/l | 4 | 4 
Hb 75 g/l | 4 | 4 
arterial blood pressure 90/60 mm Hg | 4 | 4 
pulse rate 90/min | 4 | 4 
left lower abdominal quadrant and upper thigh swollen with ecchymosis | 4 | 4 
diagnosis of haemorrhagic shock | 4 | 4 
massive transfusion pathway activated | 4 | 4 
four units of Blood transfused | 4 | 6 
four units of FFP transfused | 4 | 6 
two adult therapeutic doses of platelets transfused | 4 | 6 
10 units of cryoprecipitate transfused | 4 | 6 
noradrenaline infusion to maintain MAP > 65 mm Hg | 4 | 24 
pelvic binder in place | 4 | 24 
CT scan | 6 | 8 
CT abdomen confirmed the fracture of the left acetabulum | 8 | 8 
significant haematoma on left pelvic sidewall adjacent to the fracture | 8 | 8 
8 mm enhancing nodule suggestive of an internal iliac artery pseudoaneurysm | 8 | 8 
ill-defined blush of contrast within the haematoma | 8 | 8 
extra-peritoneal haematoma inseparable from the bladder | 8 | 8 
cirrhotic liver | 8 | 8 
6.7 cm infra-renal aortic aneurysm | 8 | 8 
transferred to the intensive care unit | 8 | 8 
invasive cardiovascular monitoring | 8 | 120 
CT Angiogram | 48 | 50 
no arterial bleed | 50 | 50 
prophylactic embolization | 50 | 50 
gelfoam embolization of anterior and posterior division segmental branches of the left internal iliac artery | 50 | 52 
10 lb skeletal traction applied | 52 | 52 
discharged to the orthopaedic ward | 120 | 120 
uncontrollable bleeding from his pin site | 120 | 120 
skeletal traction removed | 120 | 120 
continuous pressure applied to the wound | 120 | 120 
died on 30 January 2017 | 1224 | 1224 
end stage liver failure | 1200 | 1224 
hepatic encephalopathy | 1200 | 1224