32-week pregnant female | 0  
    decreased fetal movement | -168 (four weeks prior to admission)  
    fetal ultrasound | 0  
    normal cardiac activity | 0  
    fetal ascites | 0  
    edematous bowel loops | 0  
    antenatal scan showing ascites | 0  
    torch testing | 0  
    small bowel obstruction considered | 0  
    emergency cesarean section | 0  
    abdominal distention at birth | 0  
    mass felt on right umbilicus | 0  
    stabilization in neonatal ICU | 0  
    upper gastrointestinal contrast study | 24  
    normal C-loop of duodenum | 24  
    malrotation ruled out | 24  
    altered nasogastric aspirates | 24  
    serial X-ray | 24  
    absence of dye flow beyond proximal jejunal loops | 24  
    hemoglobin 6 gm% | 24  
    bowel gangrene suspected | 24  
    volvulus suspected | 24  
    emergency laparotomy at 6 hours of life | 6  
    volvulus | 6  
    gangrene of 45 cm distal ileum | 6  
    mesenteric defect | 6  
    proximal healthy 75 cm small intestine | 6  
    resection of gangrenous segment | 6  
    ileostomy | 6  
    preserved ileocecal junction | 6  
    elective stoma closure after 75 days | 1800 (75 days * 24 hours/day)  
    uneventful hospital course | 1800  
    child now 5 years old | 1800  
    no disease sequelae | 1800  
    
