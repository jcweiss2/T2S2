29 years old | 0
male | 0
admitted to intensive care unit | 0
persistent fever | -336
swelling of right knee joint | -240
pain of right knee joint | -240
fever with chills | -336
drenched in the rain | -336
took 999® cold particles | -336
drop in body temperature | -336
shortness of breath | -240
fatigue after physical activity | -240
oliguria | 0
frothy urine | 0
foul-smelling urine | 0
hypothermia 37°C | 0
heart rate 100 beats/min | 0
respiratory rate 20 breaths/min | 0
blood pressure 138/80 mmHg | 0
laboratory tests indicative of infection | 0
ultrasound color doppler showing cavity effusion | 0
synthial thickening in right knee joint | 0
thoracic CT showing pneumonia | 0
hepatic cyst in S7 segment |# 一、题目
