59 years old | 0
male | 0
admitted to the hospital | 0
decreased general well-being | 0
somnolent | 0
cachexia | 0
arterial hypotension | 0
heart rate of 90 bpm | 0
respiratory frequency of 25 per minute | 0
urinary incontinence | 0
severe necrosis of the scrotum and perineum | 0
necrosis had spontaneously perforated | 0
smell suggesting moist gangrene | 0
inflammatory syndrome | 0
hemoglobin 6.7 | 0
leukocytes 9.8 | 0
fibrinogen 8.7 | 0
C-reactive protein 327 | 0
procalcitonin 7.24 | 0
partial thromboplastin time 42.3 | 0
Bacteroides pyogenes colonization | 0
Staphylococcus haemolyticus colonization | 0
Escherichia coli colonization | 0
Clostridium innocuum colonization | 0
Enterococcus faecium colonization | 0
Enterococcus faecalis colonization | 0
Candida albicans colonization | 0
non-albicans Candida colonization | 0
injury of the right lumbar plexus | 0
diagnosis of FG | 0
calcified chronic pancreatitis | -120
pancreatic pseudocyst | -120
stent applied | -120
stent dislocated | -120
sigmoidoscopy | 24
colostomy | 24
sigmoidal anus praeter | 24
debridement of the scrotum and peritoneum | 24
surgical necrosis removal | 48
repeated debridement | 48
antimicrobiotic protection | 48
transferred from intensive care unit to urologic ward | 72
debridement | 72
suprapubic catheter change | 72
subcutaneous testicle relocation | 72
released from hospital | 168
plastic surgery | 168
skin transplantation | 168
right testicle repositioned | 168
vacuum therapy | 168
rejection and necrosis of transplanted skin | 192
necrotic areas removed | 192
vacuum therapy continued | 192
released from hospital | 216
ileus induced by adhesion pathology | 240
laparotomy | 240
adhesiolysis | 240
released from hospital | 264
control examination | 744
operated areas showed no indications of inflammation | 744
edges were smooth and easily movable | 744
wounds were dry and well covered | 744
testicles were slightly smaller | 744
scrotal skin was slightly raised | 744
preputium was tight | 744
balanitis developed | 744
arbitrary anal sphincter contractions were not possible | 744
recommended to attend another stationary intervention | 744
vacuum patch therapy | 744
digital cleaning of the ampulla recti | 744
check up on the micturition features | 744
balanitis therapy | 744
circumcision | 744