72 years old | 0
female | 0
treated diabetes | -8760
hypertension | -8760
hyperlipidemia | -8760
candidiasis | -720
HIV-1 | -720
CD4+ T-lymphocyte count 32 cells/μL | -720
VL 16,600 copies/mL | -720
abacavir (ABC) | -696
lamivudine (3TC) | -696
raltegravir (RAL) | -696
continuous ART | -696
CD4 cell count 265 cells/μL | -24
VL below the lower limit of detection | -24
abdominal pain | 0
vomiting | 0
decreased level of consciousness | 0
tachycardia | 0
labored polypnea | 0
Glasgow Coma Scale score 13 | 0
metabolic acidosis | 0
hyperlactacidemia | 0
intestinal ischemia | 0
ART suspended | 0
emergency laparotomy | 0
NOMI | 0
subtotal small bowel resection | 0
jejunostomy | 0
lactic acidosis resolved | 24
intensive care | 24
CD4 cell count 163 cells/μL | 504
VL 49,600 copies/mL | 504
HIV-1 subtype B | 504
no drug-resistant mutation | 504
R5 tropism | 504
single-dose administration of ARVs | 600
darunavir (DRV) | 600
ritonavir (RTV) | 600
lopinavir (LPV) | 600
etravirine (ETR) | 600
maraviroc (MVC) | 600
RAL | 600
plasma ARV concentrations measured | 600
Cmax of LPV and RTV below the lower limit of detection | 602
Cmax of MVC 0.580 μg/mL | 602
Cmax of RAL 0.566 μg/mL | 602
Cmax of DRV 2.18 μg/mL | 603
Cmax of ETR 2.09 μg/mL | 603
continuous ART resumed | 600
DRV 600 mg | 600
RTV 200 mg | 600
ETR 200 mg | 600
MVC 300 mg | 600
plasma ARV concentrations measured under repeated administrations | 744
Cmin of MVC 0.45 μg/mL | 744
Cmin of DRV 1.72 μg/mL | 744
Cmin of ETR below the lower limit of detection | 744
3TC 150 mg | 744
tube feeding initiated | 768
Cmin and Cmax values determined again | 1032
Cmin of MVC above the target trough | 1032
Cmax of DRV 1.1 μg/mL | 1032
Cmin of DRV below the lower limit of detection | 1032
ETR and RTV administration discontinued | 1032
dosing intervals of ARVs changed | 1032
VL decreased to 32 copies/mL | 1696
catecholamine-resistant sepsis | 2144
catheter-related bloodstream infection | 2144
death | 2144