86 years old | 0
female | 0
admitted to the hospital | 0
anorexia | -72
vomiting | -72
appendectomy | 0
right incarcerated femoral hernia | 0
small bowel obstruction | 0
severe pain | 0
redness | 0
palpable bulge | 0
white blood cell count 17.1 × 10^9/L | 0
C-reactive protein 6.13 mg/dL | 0
incarcerated ileum perforation | 0
hemorrhage necrosis | 0
necrotic ileum resection |#ERROR
