36 weeks and 0 days gestational age | 0
    female | 0
    spontaneous vaginal delivery | 0
    birth weight 2356 g | 0
    Apgar scores 9 | 0
    Apgar scores 9 | 0
    no meconium staining | 0
    respiratory distress | 0
    resuscitation with positive pressure ventilation | 0
    admitted to neonatal intensive care unit | 0
    mechanical ventilator | 0
    sepsis work-up | 0
    blood cultures | 0
    no antibiotics administered | 0
    fever | 16
    convulsions | 16
    drowsiness | 16
    pale appearance | 16
    cold extremities | 16
    cyanosis of extremities | 16
    poor capillary refill | 16
    body temperature 38.8°C | 16
    pulse 170 beats per minute | 16
    blood pressure 60/35 mmHg | 16
    respiratory rate 80 breaths per minute | 16
    oxygen saturation 87% | 16
    normal cardiovascular examination | 16
    clear lungs on auscultation | 16
    soft abdomen | 16
    not distended abdomen | 16
    slightly increased muscle tone | 16
    no skin rash | 16
    no subcutaneous hemorrhage | 16
    disseminated intravascular coagulation | 16
    cerebrospinal fluid high cell count 8.15 × 10^9/L | 16
    cerebrospinal fluid glucose 0.06 mmol/L | 16
    gram-negative rod organisms in CSF | 16
    bilateral adrenal hemorrhage | 0
    suspected adrenal insufficiency | 0
    decreased blood pressure 50/30 mmHg | 72
    increased urine output 10 mL/kg/h | 72
    urine specific gravity 1.005 | 72
    urine osmolality 160 mOsm/kg H2O | 72
    serum sodium 155 mmol/L | 72
    serum osmolality 332 mOsm/kg H2O | 72
    serum antidiuretic hormone 1.3 pg/mL | 72
    diagnosis of early-onset neonatal meningitis | 0
    diagnosis of Waterhouse-Friderichsen syndrome | 0
    positive blood cultures for E. coli | 0
    positive CSF cultures for E. coli | 24
    antibiotics treatment | 0
    hydrocortisone 10 mg/kg/day | 0
    normal blood pressure | 24
    no vasoactive agents needed | 24
    no further steroid therapy | 72
    regression of adrenal hemorrhage | 24
    negative blood cultures after 36 hours | 36
    negative CSF cultures after 36 hours | 36
    antibiotics continued until day of life 22 | 528
    diagnosis of central diabetes insipidus | 96
    intravenous vasopressin 0.3 mU/kg/h | 96
    urine output decreased to 4 mL/kg/h | 144
    urine osmolality improved to 213 mOsm/kg H2O | 144
    vasopressin dose reduced | 144
    vasopressin discontinued after day of life 12 | 288
    cerebral MRI bilateral encephalomalacia | 240
    cerebral MRI minor bleeding | 240
    cerebral MRI splenial lesion | 240
    no brain abscess | 240
    no ventriculitis | 240
    no pituitary gland abnormality | 240
    serum thyroid-stimulating hormone normal | 840
    serum thyroid hormone normal | 840
    serum adrenocorticotropic hormone normal | 840
    early morning cortisol 1.9 µg/dL | 840
    normal corticotropin-releasing hormone stimulation test | 840
    no central adrenal insufficiency | 840
    normal auditory brainstem response testing | 840
    normal electroencephalography | 840
    discharged on day of life 45 | 1080
    no respiratory assistance | 1080
    no feeding tube | 1080
