76 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
pancreatic adenocarcinoma | -672 | 0 | Factual
metastasis to the liver | -672 | 0 | Factual
diastolic heart failure | -672 | 0 | Factual
atrial fibrillation | -672 | 0 | Factual
coronary artery disease | -672 | 0 | Factual
severe hyponatremia | 0 | 0 | Factual
sodium level of 116 mmol/L | 0 | 0 | Factual
x-ray findings consistent with pneumonia | 0 | 0 | Factual
broad-spectrum antibiotics | 0 | 24 | Factual
fluid for hyponatremia | 0 | 24 | Factual
jugular vein distention | 0 | 0 | Factual
lower extremity pitting edema | 0 | 0 | Factual
transthoracic echocardiogram (TTE) | 0 | 0 | Factual
normal left ventricular cavity size | 0 | 0 | Factual
mildly reduced systolic function | 0 | 0 | Factual
septal flattening | 0 | 0 | Factual
left atrial enlargement | 0 | 0 | Factual
suspected MV vegetation | 0 | 0 | Factual
severe mitral regurgitation | 0 | 0 | Factual
tricuspid regurgitation | 0 | 0 | Factual
elevated RV systolic pressure | 0 | 0 | Factual
type 2 and type 3 pulmonary arterial hypertension | 0 | 0 | Factual
ill-defined thickening in the TV leaflets | 0 | 0 | Factual
afebrile | 0 | 0 | Factual
leukocytosis | 0 | 0 | Factual
recent urethral instrumentation | -24 | 0 | Factual
blood cultures | 0 | 24 | Factual
infectious disease specialist consultation | 0 | 0 | Factual
transesophageal echocardiogram (TEE) | 24 | 24 | Factual
normal left ventricular size and function | 24 | 24 | Factual
normal RV size and function | 24 | 24 | Factual
hypermobile interatrial septum | 24 | 24 | Factual
no left atrial or left atrial appendage thrombus | 24 | 24 | Factual
vegetations on the MV leaflets | 24 | 24 | Factual
severe mitral regurgitation | 24 | 24 | Factual
systolic flow reversal in the pulmonary vein | 24 | 24 | Factual
vegetation on the TV leaflet | 24 | 24 | Factual
tricuspid regurgitation | 24 | 24 | Factual
RVSP 47 mm Hg | 24 | 24 | Factual
negative blood cultures | 24 | 24 | Factual
polymerase chain reaction testing negative | 24 | 24 | Factual
workup for antiphospholipid syndrome unremarkable | 24 | 24 | Factual
marantic (nonbacterial) endocarditis | 24 | 24 | Factual
discontinued apixaban | -24 | 0 | Factual
recommended low molecular weight heparin or unfractionated heparin | 24 | 24 | Factual
computed tomography imaging of the head | 24 | 24 | Factual
discontinued broad-spectrum antibiotics | 24 | 24 | Factual
started on enoxaparin | 48 | 48 | Factual
expired | 168 | 168 | Factual