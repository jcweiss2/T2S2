35 years old | 0
male | 0
admitted to the hospital | 0
back pain | -336
intermittent fever | -336
oral levofloxacin | -336
infection of unknown origin | -336
severe back pain | 0
shortness of breath | 0
fatigue | 0
several-week history of fever | -168
blood pressure 129/65 mm Hg | 0
heart rate 110 beats/min | 0
temperature 102 °F | 0
respiratory rate 35 breaths/min | 0
vegetations on the tricuspid valve | 24
necrotizing bilateral pneumonia | 48
large retropharyngeal abscess | 48
epidural abscess at T8-T9 | 48
spinal cord compression | 48
active IVDU of methamphetamine | -10080
chronic hepatitis C | -10080
type 2 diabetes mellitus | -10080
IV vancomycin | 0
IV ceftriaxone | 0
intubated on a mechanical ventilator | 96
IV nafcillin | 96
drainage of the abscesses | 192
decompressive laminectomy | 192
bacteremia | 0
cardiothoracic surgery | 384
catheter-based aspiration therapy | 384
FlowTriever system | 384
Triever24 aspiration catheter | 384
Triever20 Curve aspiration catheter | 384
intracardiac echocardiography | 384
aspiration catheter navigated | 384
vegetation removed | 384
debulking therapy | 384
tricuspid valve regurgitation improved | 384
extubated | 408
discharged home | 624
IV ampicillin and sulbactam | 624
follow-up echocardiography | 1056
tricuspid valve free of vegetation | 1056
mild tricuspid regurgitation | 1056
7-month clinic visit | 1584