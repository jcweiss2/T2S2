60 years old | 0 | 0 
female | 0 | 0 
hepatitis C-related cirrhosis | 0 | 0 
recurrent hepatic encephalopathies | 0 | 0 
chronic portal vein thrombosis | 0 | 0 
admitted to the hospital | 0 | 0 
liver transplantation | 0 | 0 
construction of an end-to-side anastomosis | 0 | 0 
end-to-end bile duct anastomosis | 0 | 0 
massive venous bleeding from local varices | 0 | 0 
iliac conduit construction | 0 | 0 
recovered well after surgery | 0 | 0 
normal liver graft function | 0 | 0 
stenosis of the bile duct anastomosis | -1680 | -1680 
biliary leakage | -1680 | -1680 
elevated liver enzymes | -1680 | -1680 
treated with a pigtail | -1680 | -1680 
FCSCEMS insertion | -840 | -840 
persisting leakage | -840 | -420 
stent extraction | -420 | -420 
hepatitis C reinfection | -420 | 0 
recurrent stenosis of the biliary anastomosis | -420 | 0 
ERCP | -420 | 0 
balloon dilatations | -420 | 0 
placements of pigtails | -420 | 0 
stent placements | -420 | 0 
biopsy-proven significant fibrosis | -1680 | -1680 
treated with pegylated interferon and ribavirin | -100 | 0 
elective ERCP | 0 | 0 
recovery of 3 plastic double-pigtails | 0 | 0 
cholangiogram | 0 | 0 
large portobiliary fistula | 0 | 0 
hemobilia | 0 | 0 
FCSEMS placement | 0 | 0 
prophylactic antibiotic treatment with ciprofloxacin | 0 | 48 
septic shock | 48 | 48 
admitted to the intensive care unit | 48 | 48 
hemodynamic support | 48 | 48 
empiric broad-spectrum antibiotic treatment | 48 | 48 
computed tomography | 48 | 48 
angiography | 48 | 48 
chronic obliteration of the iliac conduit | 48 | 48 
partial perfusion of the hepatic artery by gastroduodenal collaterals | 48 | 48 
anuric kidney failure | 48 | 48 
continuous venovenous hemofiltration | 48 | 96 
intermittent hemodialysis | 96 | 672 
recovered well | 672 | 672 
evaluation for liver re-transplantation | 672 | 672 
FCSEMS replacement | 4032 | 4032 
extraction of the lying FCSEMS | 4032 | 4032 
no evidence of persisting leakage | 4032 | 4032 
no relevant stenosis | 4032 | 4032 
follow-up | 4032 | 6312 
no evidence of recurrent stenosis or portobiliary fistula | 6312 | 6312 
no further endoscopic intervention | 6312 | 6312