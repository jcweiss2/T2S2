16 years old | 0
female | 0
lost consciousness | -20
CPR applied | -20
admitted to Emergency Department | 0
ECPR performed | 20
ECMO established | 40
heparin administered | 40
spontaneous heart rate returned | 60
transferred to ICU | 80
no history of drug or food allergy | 0
body temperature 35°C | 0
heart rate 112 bpm | 0
blood pressure 85/52 mm Hg | 0
deep coma | 0
no pupillary reflex | 0
pupil size 6 mm | 0
balanced salt administered | 0
lansoprazole administered | 0
anti-infective administered | 0
no urine output | 0
CRRT started | 120
shivering | 144
left lower extremity edema | 144
papaverine administered | 144
thermotherapy applied | 144
pupillary reflex resumed | 144
sedative and analgesic drugs stopped | 144
sedative and analgesic drugs continued | 144
left lower extremity swelling worsened | 192
blood flow to left lower extremity restricted | 192
ECMO stopped | 192
blood flow to left lower extremity resumed | 192
CRRT continued | 192
enteral nutrition started | 216
anti-infective therapy switched | 240
breathed spontaneously | 264
tracheostomy performed | 264
ventilator withdrawn | 272
diarrhea developed | 336
high fever | 336
shock | 336
sputum culture positive for Acinetobacter baumannii | 336
nasogastric feeding replaced by parenteral nutrition | 336
metronidazole administered | 336
Smecta administered | 336
tigecycline administered | 336
Bifidobacterium, Lactobacillus, Enterococcus, and Bacillus cereus administered | 336
body temperature decreased | 336
diarrhea not improved | 336
vancomycin administered | 360
metronidazole administered | 360
diarrhea not mitigated | 360
bedside colonoscopy suggested PMC | 384
anti-infectives changed | 384
treatment strategy adjusted | 384
diarrhea not ameliorated | 384
dark red diarrhea observed | 432
hematochezia worsened | 432
poisoning symptoms worsened | 432
first FMT performed | 432
diarrhea improved | 432
second FMT performed | 456
third FMT performed | 464
diarrhea further mitigated | 464
nasogastric feeding of lactose-free formula milk started | 472
diarrhea reduced | 472
fourth FMT performed | 528
diarrhea further improved | 528
tracheotomy closed | 552
coronary computed tomography angiography performed | 576
origin of right coronary artery at top of sinus | 576
rehabilitation therapy started | 600
discharged | 1056
restored self-care ability | 1056