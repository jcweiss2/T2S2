11 years old | 0
    male | 0
    sliding in the supine position | -72
    iron bar entered body from right site of anus | -72
    iron bar exited from loin | -72
    waited for an hour until fire department arrived | -72
    fire department cut iron bar into 140 cm piece | -72
    taken to nearest state hospital | -72
    transferred to emergency service of our hospital | -72
    met by team in emergency service | 0
    informed by 112 emergency services operator | 0
    slightly hypothermic | 0
    intermediate overall condition | 0
    no active hemorrhaging | 0
    normal abdomen | 0
    difficulty in breathing | 0
    chest x-ray examination | 0
    abdominal x-ray examination | 0
    performed under supervision of Pediatric Surgery | 0
    performed under supervision of Orthopedics | 0
    performed under supervision of Brain Surgery | 0
    performed under supervision of Anesthesiology | 0
    performed under supervision of Radiology | 0
    patient's pain increased | 0
    breathing difficulty increased | 0
    successfully intubated on stretcher | 0
    computed tomography (CT) performed | 0
    no abdominal injury detected in CT | 0
    no chest injury detected in CT | 0
    considering possibility of rectosigmoid injury | 0
    considering possibility of retroperitoneal injury | 0
    laparotomy performed to remove iron bar | 0
    tetanus vaccination performed | 0
    antibiotic treatment started | 0
    ampicillin/sulbactam | 0
    amikacin | 0
    ornidazole | 0
    patient carefully placed in supine position | 0
    abdominal region opened | 0
    hematoma 5–6 cm in diameter at sigmoid colon mesentery | 0
    abdominal skin closed | 0
    placed in face-down position | 0
    main goal to shorten iron bar to avoid more injuries | 0
    appropriate tools not available at hospital | 0
    fire department urgently called | 0
    fire department reported three types of bar cutters | 0
    scissor-type cutter would cause more injuries | 0
    spiral cutter cannot cut such bar | 0
    spiral-type cutter that can cut iron by transmitting heat | 0
    cutter used | 0
    cold water continuously poured to prevent burning | 0
    shortened iron bar pulled out in controlled manner | 0
    iron bar removed | 0
    oxygen and nitrous oxide container tubes present | 0
    high heat and pressure almost caused explosion | 0
    light exudate containing bone pieces came from wound | 0
    Orthopedics stated no intervention required | 0
    Brain Surgery stated no intervention required | 0
    wound washed and cleaned | 0
    lumbar exit hole closed with suture | 0
    long Penrose drain placed into entry hole | 0
    patient placed in supine position | 0
    abdominal cavity examined once more | 0
    cavity closed | 0
    patient remained in intensive care unit for two days | 48
    discharged with full recovery on 11th day | 264
    control lumbar spinal MRI | 264
    subcutaneous degenerative changes at L4-L5 levels | 264
    degenerative changes in nerve roots at S2–S5 levels | 264
    electromyography findings normal | 264
    no problems while walking | 264
    no problems defecating | 264
    no problems urinating | 264
    no problems after 14th postoperative month | 4032
    
    
    