28 years old | 0
    woman | 0
    transported emergently to the hospital | 0
    fever | -72
    abdominal pain | -72
    confusion | 0
    blood pressure of 80/50 mm Hg | 0
    heart rate of 120 beats/min | 0
    respiratory rate of 32 breaths/min | 0
    body temperature of 38.3 °C | 0
    abdominal tenderness | 0
    rebound tenderness | 0
    abdominal rigidity | 0
    cervical motion tenderness | 0
    small amounts of cervical bleeding | 0
    grayish-white cervical fluids | 0
    foul-smelling cervical fluids | 0
    arterial blood gas pH of 7.35 | 0
    HCO3 level of 15.5 mmol/L | 0
    lactate level of 6.9 mmol/L | 0
    white blood cell count of 0.9 × 10^9/L | 0
    C-reactive protein level of 33.98 mg/dL | 0
    contrast-enhanced computed tomography (CT) | 0
    HPVG | 0
    pneumatosis intestinalis | 0
    mesenteric emphysema | 0
    free air | 0
    ascites | 0
    small intestinal wall thickening | 0
    emergency laparotomy | 0
    concerns of intestinal ischemia | 0
    concerns of gastrointestinal perforation | 0
    opaque ascites | 0
    no perforation | 0
    no necrosis | 0
    inflammatory redness of uterus | 0
    inflammatory redness of fallopian tubes | 0
    edema of uterus | 0
    edema of fallopian tubes | 0
    right fallopian tube adhered | 0
    abdominal cavity washed with physiological saline | 0
    abdomen closed | 0
    gram staining of opaque ascites | 0
    large number of neutrophils | 0
    gram-negative cocci | 0
    short rods | 0
    diagnosed with septic shock | 0
    pelvic peritonitis | 0
    treated in ICU | 0
    administered minocycline 200 mg/day | 0
    administered ceftriaxone 2 g/day | 0
    administered metronidazole 1500 mg/day | 0
    negative Neisseria gonorrhoeae in ascites | 0
    negative Chlamydia trachomatis in ascites | 0
    negative Neisseria gonorrhoeae in vaginal fluid | 0
    negative Chlamydia trachomatis in vaginal fluid | 0
    negative Neisseria gonorrhoeae in urine | 0
    negative Chlamydia trachomatis in urine | 0
    negative Neisseria gonorrhoeae in pharynx | 0
    negative Chlamydia trachomatis in pharynx | 0
    negative HIV-RNA PCR | 0
    detected F. necrophorum in blood | 7*24
    detected F. necrophorum in ascites | 7*24
    detected Gardnerella vaginalis in ascites | 7*24
    detected Gardnerella vaginalis in vaginal fluid | 7*24
    detected Mobiluncus species in vaginal fluid | 7*24
    no bacteria detected in urine | 7*24
    no bacteria detected in pharynx | 7*24
    no bacteria detected in stool | 7*24
    CT revealed resolution of HPVG | 8*24
    CT revealed resolution of pneumatosis intestinalis | 8*24
    patient left ICU | 12*24
    untreated bacterial vaginosis (BV) prior to admission | -3*168
    postcoital bleeding | -3*168
    dyspareunia | -3*168
    cloudy vaginal fluid | -3*168
    odorous vaginal fluid | -3*168
    multiple sexual partners | 0
    receptive oral sex | 0
    no intrauterine device | 0
    no condom use | 0
    no upper respiratory symptoms | 0
    no antibiotics used | 0
    no signs of pharyngeal tonsillitis | 0
    pharyngeal swab culture test negative | 0
    no thrombophlebitis | 0
    no pulmonary nodules | 0
    Lemierre's syndrome ruled out | 0
    no abnormalities in gingiva | 0
    no abnormalities in urinary tract | 0
    circulatory failure | 0
    suspected fatal intestinal necrosis | 0
    coexistence of HPVG and PI | 0
    inflammation of uterus | 0
    inflammation of fallopian tubes | 0
    adhesion of fallopian tubes | 0
    opaque ascites observed | 0
    gas-producing bacterium F. necrophorum detected | 7*24
    HPVG and PI disappeared | 8*24
    patient never used intrauterine devices | 0
    method of transfer from partner's oral cavity | 0
    F. necrophorum not grown in vaginal fluid culture | 0
    growth of Gardnerella vaginalis in vaginal fluid | 7*24
    growth of Gardnerella vaginalis in ascites | 7*24
    signs of BV 3 weeks prior | -3*168
    Gram stain findings polymorphic | 0
    negative Gram stain for other Fusobacterium species | 0
    no declarations of interest | 0