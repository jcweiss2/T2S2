18 years old | 0
male | 0
non-smoking | 0
hypertension | 0
chronic cough | -168
dyspnea | -168
50-pound weight loss | -168
nausea | -168
vomiting | -168
cachexic | -168
scleral icterus | -168
jaundice | -168
mucous membranes dry | -168
normal bowel sounds | -168
no pain | -168
no distension | -168
no organomegaly | -168
decreased breath sounds | -168
tachycardic | -168
hypotensive | -168
hyponatremia | -168
elevated alkaline phosphatase | -168
elevated total bilirubin | -168
elevated aspartate aminotransferase | -168
elevated alanine aminotransferase | -168
innumerable pulmonary parenchymal nodules | -168
large mass in the lingula | -168
large mass in the left lower lobe | -168
pleural effusion | -168
abdominal ultrasonography | -168
severely dilated common bile duct | -168
moderately distended gall bladder | -168
computed tomography | -168
large heterogeneous mass in the pancreatic head | -168
grossly dilated common bile duct | -168
enlarged retroperitoneal lymph nodes | -168
biopsy of lung mass | -168
biopsy of pancreatic head | -168
cell clusters with high nuclear pleomorphism | -168
prominent nuclei | -168
TTF-1 positive | -168
CK-7 positive | -168
p63 negative | -168
metastases to the brain | -168
radiation therapy | -168
adjunctive chemotherapy | -168
widespread tumor burden | -168
obstructive jaundice | -168
jaundice persisted | -168
severe pneumonia | -168
sepsis | -168
death | 72