45 years old | 0
male | 0
admitted to the hospital | 0
cardiac transplantation | 0
ischaemic cardiomyopathy | 0
atrial fibrillation | 0
atrial flutter | 0
hypertension | 0
dyslipidaemia | 0
depression | 0
mild rejection | 336
tacrolimus | 336
mycophenolate mofetil | 336
prednisolone | 336
first-degree heart block | 840
second-degree heart block | 840
isoprenaline | 840
methylprednisolone | 840
increased prednisolone dose | 840
postoperative ICU course | -720
recurrent sepsis | -720
dialysis-dependent acute kidney injury | -720
haemopericardium | -720
peripheral limb ischaemia | -720
below-knee amputation | -720
severe upper abdominal pain | 960
weaning from mechanical ventilation | 960
reduced haemoglobin | 960
elevated white cell count | 960
reduced platelets | 960
elevated bilirubin | 960
elevated gamma-GT | 960
elevated alkaline phosphatase | 960
raised transaminases | 960
hyperdense haemobilia | 960
haemoperitoneum | 960
gallbladder wall defect | 960
contiguous haematoma | 960
emergency laparoscopic cholecystectomy | 960
abdominal washout | 960
necrotic gallbladder | 960
perforated gallbladder | 960
moderate-volume haemoperitoneum | 960
bradycardic | 960
loss of cardiac output | 960
successful resuscitation | 960
chest compressions | 960
epinephrine infusion | 960
no collection | 216
no biliary obstruction | 216
protracted recovery | 216
cardiac arrest | 216
AICD insertion | 216
fungal infective endocarditis | 216
post-transplant lymphoproliferative disorder | 216
pulmonary embolism | 216
discharged from ICU | 1800
inpatient rehabilitation | 1800
readmission to ICU | 1800
sepsis | 1800
hypotension | 1800
resolved AKI | 1800
returned home | 5760
physical rehabilitation | 5760
ongoing antirejection regimen | 5760
everolimus | 5760
tacrolimus | 5760
prednisolone | 5760
ongoing physiotherapy | 5760
occupational therapy | 5760
lower limb prostheses consideration | 5760
no long-term sequelae | 5760
acalculous cholecystitis | 5760
ACC | 5760
gallbladder perforation | 5760
Niemeier type 1 perforation | 5760
surgical vagotomy | 5760
gallbladder dysmotility | 5760
stasis | 5760
gallbladder ischaemia | 5760
ischaemic cardiomyopathy | 5760
steroid administration | 5760
prolonged ICU stay | 5760
sepsis | 5760
AKI | 5760
peripheral limb ischaemia | 5760
below-knee amputation | 5760
masked ACC signs | 5760
hepatic enzyme derangement | 5760
cholestatic disease | 5760
polypharmacy | 5760
non-contrast CT | 5760
synchronous haemobilia | 5760
haemoperitoneum | 5760
coagulopathy | 5760
vascular rupture | 5760
targeted ultrasound | 5760
gallbladder wall defect confirmation | 5760
haematoma traversal | 5760
inconclusive clinical picture | 5760
emergency cholecystectomy | 5760
0. Admission to hospital (day 40 post-transplant) | 0
Medical history: atrial fibrillation, atrial flutter, hypertension, dyslipidaemia, depression | 0
Ischaemic cardiomyopathy (reason for transplant) | 0
Day 14: mild rejection | (14-40)*24 = -624 hours
Treatment with tacrolimus, mycophenolate mofetil, prednisolone | -624
Day 35: first-degree heart block, second-degree heart block | (35-40)*24 = -120 hours
Treatment with isoprenaline, methylprednisolone, increased prednisolone dose | -120
Recurrent sepsis, dialysis-dependent AKI, haemopericardium, peripheral limb ischaemia | timestamp corresponding to day 30: (30+40)*24? Wait, no. Wait, day 30 post-transplant is 30 days after transplant, and the main admission is at day 40. So relative to day 40, day 30 is 10 days before, so -10*24 = -240 hours.
Below-knee amputation at day 30 | -240
Severe upper abdominal pain | 0
Weaning from mechanical ventilation | 0
Investigations: reduced hemoglobin, elevated WBC, reduced platelets, elevated bilirubin, gamma-GT, alkaline phosphatase, transaminases | 0
CT findings: hyperdense haemobilia, haemoperitoneum, gallbladder wall defect | 0
Ultrasound findings: contiguous haematoma, defect in gallbladder fundus | 0
Treatment: emergency laparoscopic cholecystectomy, abdominal washout | 0 (within hours)
Surgery findings: necrotic gallbladder, perforated, haemoperitoneum | 0
Outcome during surgery: bradycardic, loss of cardiac output, resuscitation, chest compressions, epinephrine infusion | 0
Follow-up after 9 days: no collection, no biliary obstruction | +216 hours
Protracted recovery complications: cardiac arrest, AICD insertion, fungal endocarditis, lymphoproliferative disorder, pulmonary embolism | after surgery, but timing unclear. Since these occur after the follow-up, perhaps timestamp +216, but the case states "ensued" after surgery, so maybe same day? Unclear, so approximate.
Readmission to ICU for sepsis, hypotension | timestamp +840
Resolved AKI | timestamp +840
Ongoing treatments: everolimus, tacrolimus, prednisolone | 5760
Physiotherapy, occupational therapy, prostheses consideration | 5760
No long-term sequelae | 5760
mild rejection | -624 (day 14)
tacrolimus | -624
mycophenolate mofetil | -624
prednisolone | -624
first-degree heart block | -120 (day 35)
second-degree heart block | -120
isoprenaline | -120
methylprednisolone | -120
increased prednisolone dose | -120
recurrent sepsis | -240 (day 30)
dialysis-dependent AKI | -240
haemopericardium | -240
peripheral limb ischaemia | -240
below-knee amputation | -240
severe upper abdominal pain | 0
weaning from mechanical ventilation | 0
reduced haemoglobin | 0
elevated white cell count | 0
reduced platelets | 0
elevated bilirubin | 0
elevated gamma-GT | 0
elevated alkaline phosphatase | 0
raised transaminases | 0
hyperdense haemobilia | 0
haemoperitoneum | 0
gallbladder wall defect | 0
contiguous haematoma | 0
emergency laparoscopic cholecystectomy | 0
abdominal washout | 0
necrotic gallbladder | 0
perforated gallbladder | 0
moderate-volume haemoperitoneum | 0
bradycardic | 0
loss of cardiac output | 0
successful resuscitation | 0
chest compressions | 0
epinephrine infusion | 0
discharged from ICU | 1800 (75 days post-transplant: 75-40=35 days=840 hours. Wait, 75 days post-transplant minus 40 days would be 35 days, which is 35*24=840 hours. So discharged from ICU at +840 hours)
