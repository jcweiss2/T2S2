21 years old | 0
male | 0
body mass index 28.2 | 0
91.1kg | 0
admitted to the intensive care unit | 0
acute hypoxic/hypercapnic respiratory failure | 0
acute kidney injury | 0
septic shock | 0
heroin use | -72
diagnosed with methicillin-susceptible Staphylococcus aureus pneumonia | 0
intubated | 12
propofol for induction | 12
creatinine increased to 1.8 mg/dl | 24
urine sediment evaluation | 24
bright pink pellet | 24
amorphous crystals | 24
urine acidified | 24
urine alkalized | 24
polychromatic birefringence rhomboid uric acid crystallization | 24
amorphous urate crystals | 24
given i.v. fluids | 24
serum creatinine returned to baseline | 48
extubated | 72
discharged | 96
pink urine syndrome | 24
low urine pH | 24
urate excretion | 24
insulin resistance | -72
hypertriglyceridemia | -72
type 2 diabetes mellitus | -72
metabolic syndrome | -72
oxidative stress | -72
heme oxygenase-1 pathway | -72
propofol administration | 12
antidiuretic hormone release | 12
urate excretion increased | 24
urine osmolality increased | 24
urine output reduced | 24
urate clearance | 24
renal tubular function | 24
acute prerenal AKI | 0
GFR | 0
tubular function | 0
urate physiology | -72
uric acid crystallization | 24
nephrolithiasis | -72
urine pH | 24
ammoniagenesis | -72
renal tubular sodium-hydrogen exchanger | -72
insulin stimulates | -72
PI3K-SGK1 | -72
ammonia production | -72
urine sediment | 24
urine color | 24
urine pH | 24
urate concentration | 24
urine temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink pigment | 24
uricine | 24
urohematoporphyrin | 24
uroporphyrin | 24
coproporphyrin | 24
urohematin | 24
urocyanin | 24
indirubin | 24
indigotin | 24
uroerythrin | 24
purpurin | 24
skatol red | 24
nephrorosein | 24
urorosein | 24
uricine | 24
bilirubin metabolism | -72
heme oxygenase-1 | -72
oxidative stress | -72
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
propofol | 12
antioxidant activity | 12
anti-inflammatory activity | 12
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24
urate excretion | 24
urine color | 24
urate concentration | 24
urine pH | 24
temperature | 24
urate solubility | 24
uric acid precipitation | 24
pink urine syndrome | 24
insulin resistance | -72
propofol administration | 12
chronic hyperuricemia | -72
urate clearance | 24
acidic urine | 24
GFR | 24
chronic oxidative stress | -72
heme oxygenase-1 pathway | -72
Nrf2 | 12
heme oxygenase-1 | 12
bilirubin | 24
carbon monoxide | 24
ferritin | 24
free iron | 24
urinary uricine | 24