four-month-old | 0
mulatto | 0
male | 0
admitted to the hospital | 0
lesions miliaria rubra-like | -720
on the neck | -720
on the folds of the upper limbs | -720
on the folds of the lower limbs | -720
referred to a pediatrician | -720
prescribed a powder formulation with bismuth subgallate and zinc oxide | -720
prescribed a cream with ketoconazole, betamethasone dipropionate and neomycin sulfate | -720
applied for one month throughout the body | -720
no improvement in the condition | -672
prescribed prednisolone | -672
potassium permanganate in topical solution | -672
prescribed a single-dose ampoule of betamethasone, intramuscularly | -672
lesions spread to the trunk | -672
lesions spread to the face | -672
lesions spread to the scalp | -672
lesions became crusty | -672
referred to the dermatology clinic | -672
diagnosis of "severe seborrheic dermatitis" | -672
mother followed throughout pregnancy | -1300
mother presented all negative serological tests | -1300
mother denied any type of intercurrence | -1300
mother needed topical treatment for scabies during pregnancy | -1300
child born healthy | -1300
multiple erythematous papules | 0
crusted and erythematous lesions disseminated in the body | 0
mainly affecting the trunk | 0
mainly affecting the scalp | 0
nail dystrophy | 0
fissures in the abdomen | 0
hypoactive | 0
tachycardic | 0
febrile | 0
cushingoid facies | 0
anasarca | 0
main diagnostic hypothesis was crusted or Norwegian scabies | 0
associated with secondary infection and sepsis | 0
mother complained of important pruritus | 0
grandparents complained of important pruritus | 0
mother presented erythematous and hyperchromic papules | 0
grandparents presented erythematous and hyperchromic papules | 0
dermoscopy several parasites | 0
skin biopsy | 0
laboratory tests requested | 0
infant hospitalized in a pediatric hospital | 0
histopathology revealed tunnels in the horny layer with the presence of the parasite | 24
laboratory tests revealed significant leukocytosis | 24
laboratory tests revealed left shift | 24
laboratory tests revealed thrombocytopenia | 24
laboratory tests revealed increased levels of inflammatory markers | 24
intravenous antibiotic therapy | 24
topical application of permethrin lotion 1% once daily | 24
contact isolation | 24
family members treated with oral ivermectin | 24
family members treated with topical permethrin lotion 5% | 24
patient presented improvement of cutaneous lesions | 240
condition evolved with septic shock | 240
treatment instituted in the intensive care unit | 240
cardiac arrest | 240
death | 240