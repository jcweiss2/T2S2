29 years old | 0
female | 0
admitted to the hospital | 0
self-inflicted gunshot injury | -1008
abdominal injury | -1008
epigastrium wound | -1008
left hypochondrium wound | -1008
left lumbar area wound | -1008
laparotomy | -1008
perforation in the antrum of the stomach | -1008
multiple small bowel perforations | -1008
primary surgical repair | -1008
bilateral lateral retroperitoneal hematomas | -1008
transferred to ICU | -1008
pulmonary embolism | -504
disseminated intravascular coagulation | -504
managed with blood products | -504
recovered | -168
discharged home | -168
left iliac fossa pain | -336
watery stool | -336
reduced hemoglobin level | -336
raised serum C-reactive protein | -336
abdominal CT scan | -336
left-sided retroperitoneal collection | -336
contrast extravasation | -336
urinoma formation | -336
colonic fistula | -336
referred to trauma center | -336
cystoscopy | -336
retrograde pyelogram | -336
complete transection of the left upper ureter | -336
left percutaneous nephrostomy | -336
left-sided pigtail drain | -336
antibiotics | -336
sepsis workup | -336
multi-drug-resistant coliform | -336
clear urine draining | -336
repeat CT scan | -168
reduction in size of left-sided urinoma | -168
peripherally enhancing collection | -168
right side of the pelvis | -168
compressing urinary bladder | -168
pigtail drain insertion | -168
minimal dark reddish fluid | -168
discharged | -168
elective surgery | 0
cystoscopy | 0
extra-luminal compression of the bladder | 0
intraoperative findings | 0
dense fibrosis | 0
left end-to-end ureteric anastomosis | 0
ureteroureterostomy | 0
double J stent | 0
colonoscopy | 0
methylene blue instillation | 0
negative fistula testing | 0
discharged from hospital | 72
outpatient department | 144
flexible cystoscopy | 144
removal of left DJS | 144