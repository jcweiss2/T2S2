46 years old | 0
female | 0
presented to the emergency department | 0
headaches | -1008
posterior neck pain | -1008
nausea | -1008
loss of appetite | -1008
blurry vision | -1008
head trauma | -1344
domestic abuse incident | -1344
no hospitalization | -1344
no surgical intervention | -1344
last menstrual cycle | -1344
normal menstrual cycles | -1344
HIV/AIDS | 0
CD4 count 124 cells/μL | 0
chronic hepatitis B infection | 0
cocaine abuse | 0
remote history of infectious endocarditis | 0
low-grade fever 100.4 °F | 0
hypotension 76/51 mm Hg | 0
normal respiratory rate 17 breaths/min | 0
tachycardic heart rate 126 beats/min | 0
oxygen saturation 96% | 0
cachectic | 0
acute distress | 0
neurologic examination no abnormalities | 0
cardiovascular examination tachycardia | 0
no significant findings on physical exam | 0
no formal visual field examination | 0
moderate hyponatremia | 0
hypochloremia | 0
elevated creatinine level | 0
acute kidney injury | 0
hypoalbuminemia | 0
anemia | 0
leukopenia | 0
negative pregnancy test | 0
computed tomography scan hypoenhancing hypodense mass in sella | 0
MRI centrally necrotic mass with thick peripheral wall enhancement | 0
no evidence of sinusitis | 0
admitted to neurologic intensive care unit | 0
intravenous fluid resuscitation | 0
empiric broad-spectrum antibiotics | 0
vancomycin | 0
cefepime | 0
metronidazole | 0
fluconazole | 0
central hypothyroidism | 0
secondary adrenal insufficiency | 0
low insulin-like growth factor-1 | 0
low prolactin level | 0
oral levothyroxine | 0
stress dose hydrocortisone 50 mg every 6 hours | 0
normal urine osmolality | 0
high urine output | 48
increased thirst | 48
decreased urine osmolality 186 mOsm/kg | 48
increased blood osmolality 315 mOsm/kg | 48
urine sodium 29 mmol/L | 48
diabetes insipidus | 48
oral desmopressin 50 μg daily | 48
normalized urine output | 48
normalized urine osmolality | 48
condition improved | 0
vital signs stabilized | 0
repeat MRI after 10 days | 240
decreased mass size | 240
thickening peripheral wall | 240
continued broad-spectrum antibiotics | 240
diagnosed with pituitary abscess | 0
negative blood cultures | 0
no lumbar puncture | 0
no surgical intervention | 0
6-week antibiotic regimen | 0
repeat MRI 11 months | 7920
pituitary destruction | 7920
persistent central hypothyroidism | 0
oral hydrocortisone | 0
no menstrual cycles | 0
secondary hypogonadism | 0
self-discontinued desmopressin | 0
no polyuria | 0
no polydipsia | 0
discontinued desmopressin | 0
normal sodium levels | 0
normal serum osmolality | 0
no fever | 0
hypotension | 0
adrenal insufficiency | 0
septic shock | 0
resolved diabetes insipidus | 0
pituitary dysfunction | 0
endocrinopathies | 0
permanent hypothyroidism | 0
permanent adrenal insufficiency | 0
