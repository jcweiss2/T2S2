40 years old | 0
male | 0
admitted to hospital | 0
chest pain | -5
back pain | -5
tearing-like pain | -5
computed tomography angiography | -5
acute type A aortic dissection | -5
hypertension | -6720
heavy smoking | -72000
persistent tearing pain | 0
renal function test | 0
creatinine | 0
imaging examinations | 0
thoracic and abdominal aorta CTA | 0
aortic false lumen formation | 0
ascending aortic and total aortic arch replacement | 0
stented elephant trunk implantation | 0
general anesthesia | 0
cardiopulmonary bypass | 0
transferred to ICU | 0
red blood cells transfusion | 0
plasma transfusion | 0
cryoprecipitate transfusion | 0
platelets transfusion | 0
lung protective ventilation | 0
fluid management | 0
airway secretion clearance | 0
severe ARDS | 0
oxygenation index | 0
prone positioning | 6
bedside chest radiography | 6
diffuse exudation | 6
oxygenation index improvement | 12
prone position ventilation | 12
drain patency assessment | 12
circulatory changes monitoring | 12
blood gas analysis | 12
intermittent short-term prone positioning | 24
oxygenation index improvement | 24
diffuse exudation reduction | 48
discharged | 96