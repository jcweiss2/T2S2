27 years old | 0
    pregnant | 0
    Japanese | 0
    female | 0
    traveled to Southeast Asia | -8760
    diarrhea without abdominal pain | -504
    abdominal pain | -168
    watery diarrhea | -168
    watery diarrhea more than 10 times per day | -168
    mucous bloody stools | -168
    admitted to emergency department | 0
    severe acute enteritis | 0
    spontaneous preterm birth | 24
    newborn died | 24
    anemia | 0
    hypoalbuminemia | 0
    sigmoidoscopy | 0
    reddish edematous mucosa | 0
    adherent mucopurulent exudate | 0
    bacterial culture negative | 0
    Clostridioides difficile toxin negative | 0
    suspected severe ulcerative colitis | 0
    high-dose intravenous corticosteroid therapy planned | 0
    deterioration of consciousness | 0
    signs of peritoneal irritation | 0
    transferred to tertiary referral hospital | 0
    Glasgow Coma Scale score E3V4M6 | 0
    temperature 37.3°C | 0
    blood pressure 150/100 mmHg | 0
    pulse rate 122 beats/min | 0
    respiratory rate 22 breaths/min | 0
    percutaneous oxygen saturation 92% | 0
    distended abdomen | 0
    peritoneal irritation | 0
    anemia (Hb 10.4 g/dL) | 0
    thrombocytopenia (136,000 platelets/mm3) | 0
    prolonged coagulation (PT-INR 1.23) | 0
    elevated inflammatory response (CRP 21.1 mg/dL) | 0
    hypoalbuminemia (serum albumin 1.2 g/dL) | 0
    computed tomography | 0
    edematous changes in colorectum | 0
    loss of haustra | 0
    large amount of residue in lumen | 0
    no megacolon | 0
    no gastrointestinal perforation | 0
    stool cultures negative | 0
    CMV antigenemia test negative | 0
    managed in ICU | 0
    sigmoidoscopy | 48
    squalid ochre-colored pseudomembrane | 48
    blood | 48
    edematous reddish-purple mucosa | 48
    no granularity | 48
    no small yellowish spots | 48
    biopsies taken | 48
    suspected parasitic infection | 48
    periodic acid-Schiff staining | 72
    E. histolytica trophozoites identified | 72
    general condition worsened | 96
    required ventilator management | 96
    diagnosed with fulminant amebic enteritis | 96
    intravenous metronidazole initiated | 96
    inflammatory markers improved | 168
    diarrhea disappeared | 168
    fever disappeared | 168
    weaned off ventilator | 168
    diarrhea recurred | 480
    fever recurred | 480
    prolonged malnutrition | 480
    stool cultures negative | 480
    colonoscopy | 480
    pseudomembrane disappeared | 480
    multiple punched-out ulcers | 480
    no trophozoites | 480
    no inclusion bodies | 480
    CMV antigenemia test positive | 480
    suspected CMV enteritis | 480
    intravenous ganciclovir | 480
    symptoms improved | 480
    laboratory data improved | 480
    abdominal distension | 1440
    colonoscopy | 1440
    Gastrografin enema | 1440
    severe stenosis rectum to transverse colon | 1440
    liquid nutritional supplements | 1440
    difficulty ingesting meals | 1440
    subtotal colectomy | 1440
    ileorectal anastomosis | 1440
    wall thickening with inflammation | 1440
    stenosis rectosigmoid junction | 1440
    active inflammation | 1440
    fibrosis | 1440
    fibrotic stenosis | 1440
    no E. histolytica trophozoites | 1440
    no intranuclear inclusion bodies | 1440
    postoperative course good | 1440
    general condition improved | 1440
    discharged | 4800
    fulminant amebic enteritis | 96
    CMV enteritis | 480
    intestinal stenosis | 1440
    <|eot_id|>
    27 years old | 0
pregnant | 0
Japanese | 0
female | 0
traveled to Southeast Asia | -8760
diarrhea without abdominal pain | -504
abdominal pain | -168
watery diarrhea | -168
watery diarrhea more than 10 times per day | -168
mucous bloody stools | -168
admitted to emergency department | 0
severe acute enteritis | 0
spontaneous preterm birth | 24
newborn died | 24
anemia | 0
hypoalbuminemia | 0
sigmoidoscopy | 0
reddish edematous mucosa | 0
adherent mucopurulent exudate | 0
bacterial culture negative | 0
Clostridioides difficile toxin negative | 0
suspected severe ulcerative colitis | 0
high-dose intravenous corticosteroid therapy planned |0
deterioration of consciousness | 0
signs of peritoneal irritation | 0
transferred to tertiary referral hospital | 0
Glasgow Coma Scale score E3V4M6 | 0
temperature 37.3°C | 0
blood pressure 150/100 mmHg | 0
pulse rate 122 beats/min | 0
respiratory rate 22 breaths/min | 0
percutaneous oxygen saturation 92% | 0
distended abdomen | 0
peritoneal irritation | 0
anemia (Hb 10.4 g/dL) | 0
thrombocytopenia (136,000 platelets/mm3) | 0
prolonged coagulation (PT-INR 1.23) | 0
elevated inflammatory response (CRP 21.1 mg/dL) | 0
hypoalbuminemia (serum albumin 1.2 g/dL) | 0
computed tomography | 0
edematous changes in colorectum | 0
loss of haustra | 0
large amount of residue in lumen | 0
no megacolon | 0
no gastrointestinal perforation | 0
stool cultures negative | 0
CMV antigenemia test negative | 0
managed in ICU | 0
sigmoidoscopy | 48
squalid ochre-colored pseudomembrane | 48
blood | 48
edematous reddish-purple mucosa | 48
no granularity | 48
no small yellowish spots | 48
biopsies taken | 48
suspected parasitic infection | 48
periodic acid-Schiff staining | 72
E. histolytica trophozoites identified | 72
general condition worsened | 96
required ventilator management | 96
diagnosed with fulminant amebic enteritis | 96
intravenous metronidazole initiated | 96
inflammatory markers improved | 168
diarrhea disappeared | 168
fever disappeared | 168
weaned off ventilator | 168
diarrhea recurred | 480
fever recurred | 480
prolonged malnutrition | 480
stool cultures negative | 480
colonoscopy | 480
pseudomembrane disappeared | 480
multiple punched-out ulcers | 480
no trophozoites | 480
no inclusion bodies | 480
CMV antigenemia test positive | 480
suspected CMV enteritis | 480
intravenous ganciclovir | 480
symptoms improved | 480
laboratory data improved | 480
abdominal distension | 1440
colonoscopy | 1440
Gastrografin enema | 1440
severe stenosis rectum to transverse colon | 1440
liquid nutritional supplements | 1440
difficulty ingesting meals | 1440
subtotal colectomy | 1440
ileorectal anastomosis | 1440
wall thickening with inflammation | 1440
stenosis rectosigmoid junction | 1440
active inflammation | 1440
fibrosis | 1440
fibrotic stenosis | 1440
no E. histolytica trophozoites | 1440
no intranuclear inclusion bodies | 1440
postoperative course good | 1440
general condition improved | 1440
discharged | 4800
fulminant amebic enteritis | 96
CMV enteritis | 480
intestinal stenosis | 1440