38 years old | 0
female | 0
returned from Bali | -336
no pre travel consultation | -336
no malaria prophylaxis | -336
close contact with people in poor water and sanitation conditions | -336
saw rats around accommodation | -336
mosquito bites | -336
contact with dogs and cats | -336
asymptomatic | -168
fever | -168
chills | -168
malaise | -168
myalgia | -168
conjunctival congestion | -168
admitted to emergency department | 0
initial blood tests | 0
chest X-Ray | 0
malaria test | 0
dengue test | 0
discharged home | 0
symptomatic treatment with acetaminophen | 0
re-evaluated in ambulatory | 48
fever persisted | 48
malaise | 48
myalgia | 48
relative neutrophilia | 48
elevated hepatic aminotransferases | 48
elevated LDH | 48
mildly increased C-reactive protein | 48
admitted to Infectious Diseases Ward | 48
blood samples collected for culture | 48
serologic screen | 48
shortness of breath | 96
respiratory rate of 32/minute | 96
SatO2 90-92% on room air | 96
hypotension | 96
headache | 96
nausea | 96
macular rash | 96
arterial blood gas examination | 96
respiratory alkalosis | 96
pO2/FiO2 ratio of 327 | 96
hyperlactacidemia | 96
chest X-ray | 96
bilateral interstitial infiltrate | 96
admitted to ICU | 96
volume expansion with IV fluids | 96
IV ceftriaxone | 96
IV doxycycline | 96
oseltamivir | 96
oxygen support | 96
improved progressively | 120
no need of invasive ventilation | 120
no need of vasopressive support | 120
oliguria reverted | 120
transient decrease in hemoglobin | 120
worsening thrombocytopenia | 120
coagulopathy | 120
recovered spontaneously | 120
afebrile | 192
discharged from ICU | 192
fully recovered | 240
discharged from hospital | 312
chest X-ray | 312
resolution of pulmonary infiltrates | 312
molecular diagnostic test | 312
positive for Rickettsia spp. subgroup Typhus | 312
serum samples sent to CEVDI | 312
immunofluorescence assay | 312
seroconversion | 312
antibodies levels | 312
IgM 1:2048 | 312
IgG 1:4096 | 312
molecular detection for rickettsial DNA | 312
nested-PCR | 312
sequence characterization | 312
BLAST analysis | 312
R. typhi | 312
gltA gene fragment | 312
99% identity with R. typhi sequences | 312