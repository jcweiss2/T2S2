7 years old | 0
female | 0
admitted to the hospital | 0
periodic fever | -144
headache | -144
abdominal pain | -144
watery diarrhea | -144
projectile vomiting | -144
severe headache | -144
lethargy | -144
conjugated pneumococcal vaccines | - time unknown
Haemophilus influenzae type b vaccines | - time unknown
no contact with contaminated foods | - time unknown
no contact with domestic animals | - time unknown
mental status intact | 0
neck stiffness | 0
Bruzinski sign positive | 0
Kernig sign positive | 0
no abnormality in motor function | 0
no abnormality in muscle strength | 0
sensation intact | 0
deep tendon reflexes hyper-reactive | 0
white blood cell counts 21,150/µL | 0
segmented neutrophils 89% | 0
lymphocytes 6.3% | 0
ESR 57 mm/hr | 0
CRP 9.52 mg/dL | 0
fasting blood sugar 169 mg/dL | 0
cerebrospinal fluid examination | 0
white blood cells 1,500/µL | 0
segmented neutrophils 30% | 0
red blood cells 250/µL | 0
sugar 25 mg/dL | 0
protein 117 mg/dL | 0
no bacteria on gram staining | 0
PCR for tuberculosis negative | 0
herpes simplex virus antibody test negative | 0
co-agglutination test negative | 0
cryptococcus antigen test negative | 0
antibiotic treatment with ceftriaxone | 0
antibiotic treatment with amikacin | 0
steroid injections | 0
continued fever | 24
severe headache | 24
vomiting | 24
altered mental status | 24
stuporous | 24
delirious | 24
vancomycin added to treatment | 24
brain MRI | 24
no brain edema | 24
diplopia | 24
fever continued | 48
headache continued | 48
pain in both legs | 48
worsening mental status | 48
repeated CSF examination | 48
repeated blood tests | 48
white blood cell count 37,860/µL | 48
segmented neutrophils 88.2% | 48
lymphocytes 5.3% | 48
ESR 50 mm/hr | 48
CRP 17.19 mg/dL | 48
fasting blood sugar 142 mg/dL | 48
CSF white blood cell count 2,000/µL | 48
CSF red blood cell count 250/µL | 48
CSF sugar 73 mg/dL | 48
CSF protein 319 mg/dL | 48
gram-positive rods on gram staining | 48
L. monocytogenes identified | 48
ampicillin added to treatment | 48
antimicrobial susceptibility test | 48
IgG 872 mg/dL | 48
IgA 208 mg/dL | 48
IgM 257 mg/dL | 48
IgE 960 IU/mL | 48
C3 113 mg/dL | 48
C4 28.2 mg/dL | 48
CH50 51.1 U/mL | 48
CD3 61.3% | 48
CD4 32.7% | 48
CD8 35.2% | 48
CD19 17% | 48
ultrasound of thymus normal | 48
confused conversation | 72
no voluntary movement | 72
pupillary reflexes slow | 72
nystagmus | 72
muscle strength decreased | 72
respiratory difficulty | 72
semicoma level | 72
transferred to intensive care unit | 72
ventilator support initiated | 72
CT of brain | 72
hydrocephalus | 72
parenchymal edema | 72
brain stem extrusion | 72
extraventricular drainage | 72
repeated extraventricular drainage | 120
repeated extraventricular drainage | 312
CSF examination | 408
white blood cell count 32/µL | 408
red blood cell count 3,100/µL | 408
sugar 99 mg/dL | 408
protein 169 mg/dL | 408
no bacteria on gram staining | 408
no bacteria on blood and CSF cultures | 408
ventriculoperitoneal shunt procedure | 528
off ventilator support | 600
responded appropriately | 600
language no longer confused | 600
stable vital signs | 744
transferred from intensive care unit | 744
brain CT | 912
communicating hydrocephalus | 912
ventriculostomy | 912
parenchymal edema | 912
discharged | 1464