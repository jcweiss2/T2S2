30 years old | 0
    gravida 1 | 0
    para 0 | 0
    admitted to a local hospital | 0
    21 weeks gestation | 0
    preterm labor | 0
    negative GBS screen | -120
    complete antenatal steroid course | -72
    betamethasone intramuscular | -72
    started on latency antibiotics | -47
    ampicillin intravenous | -47
    azithromycin oral | -47
    magnesium for neuroprotection | -48
    male neonate | 0
    23 and 4/7 weeks gestational age | 0
    delivered vaginally | 0
    prolonged rupture of membranes for 58 hours | -58
    BW 0.595 kg | 0
    initially vigorous | 0
    intubation | 0
    surfactant for respiratory distress | 0
    APGAR score 5 | 1
    APGAR score 6 | 5
    APGAR score 8 | 10
    admitted to NICU | 0
    high-frequency oscillator | 0
    caffeine intravenous | 0
    umbilical catheters inserted | 0
    evaluation for bacterial infection | 0
    empiric therapy of ampicillin | 0
    empiric therapy of gentamicin | 0
    discontinued antibiotics | 48
    nil per os | 0
    total parenteral nutrition | 0
    trialed on conventional mechanical ventilation | 22
    failed mechanical ventilation | 60
    respiratory acidosis | 60
    transferred to facility | 72
    admitted to NICU | 72
    leukocytosis | 99
    WBC 19.8K/µL | 99
    bandemia 15% | 99
    septic workup | 99
    blood culture obtained | 99
    unable to draw UVC | 99
    empiric ampicillin | 99
    empiric cefepime | 99
    abdomen discolored | 99
    abdominal radiograph | 99
    gasless abdomen | 99
    blood culture positive | 99.6
    M. morganii | 99.6
    line removed | 99.6
    full sepsis workup | 120
    repeat blood cultures | 120
    peripheral blood culture | 120
    UVC blood culture | 120
    lumbar puncture | 120
    nonsterile urine culture | 120
    broadened antibiotics | 120
    meropenem | 120
    ampicillin | 120
    CSF analysis | 120
    7 RBCs/µL | 120
    1 WBC/mm³ | 120
    206 mg/dL protein | 120
    78 mg/dL glucose | 120
    CSF culture Enterococcus faecalis | 120
    nonsterile urine culture Staphylococcus epidermis | 120
    nonsterile urine culture M. morganii | 120
    nonsterile urine culture E. faecalis | 120
    peripheral culture M. morganii | 120
    UVC culture negative | 120
    clinical improvement | 120
    clinical worsening on DOL 8 | 192
    bilious emesis | 192
    increased abdominal discoloration | 192
    never on enteral feeds | 0
    oral care with colostrum | 24
    abdominal radiograph free air | 192
    spontaneous intestinal perforation | 192
    peritoneal drain placed | 192
    intraoperative peritoneal culture M. morganii | 192
    vancomycin | 192
    fluconazole | 192
    M. morganii sensitivities | 192
    ampicillin | 192
    cefepime | 192
    14-day antibiotic course | 336
    placental maternal culture E. coli | 0
    placental maternal culture Streptococcus viridans | 0
    placental maternal culture coagulase negative Staphylococcus | 0
    placental maternal culture Enterococcus | 0
    placental maternal culture Bacillus fragilis | 0
    placental fetal culture Prevotella | 0
    improved clinically | 192
    enteral feeds advanced | 192
    full enteral feeds | 192
    dexamethasone | 720
    extubated | 720
    weaned to room temperature | 2520
    patent ductus arteriosus treated with acetaminophen | 720
    bilateral germinal matrix hemorrhages | 720
    normalized ventricles | 2520
    corrected full-term cranial ultrasound | 2520
    left periventricular cyst | 2520
    stage 2 retinopathy | 2520
    discharged home | 3024
    seen in follow-up | 3024
    feeding therapy | 3024
    infant development services | 3024
    physical therapy | 3024
    normal cognitive skills | 3024
    normal expressive language | 3024
    normal fine motor | 3024
    normal gross motor | 3024
    normal sensory processing | 3024
    mild receptive language delay | 3024
    mild social emotional delay | 3024
    normal brain MRI | 3024