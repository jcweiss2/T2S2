62 years old | 0
Saudi woman | 0
admitted to King Khalid University Hospital (KKUH) | 0
laparoscopic sigmoid resection | 0
diverticula in the sigmoid | 0
diverticula in the distal descending colon | 0
fever | 72
temperature of 38.9°C | 72
septic screening | 72
urinary tract infection | 72
antibiotics started | 72
low hemoglobin | 72
blood transfusion | 72
hypotensive | 72
blood pressure 85/52 mmHg | 72
oxygen saturation 94% | 72
pulse rate 110/min | 72
transfusion stopped | 72
hydrocortisone started | 72
transferred to surgical intensive care unit (SICU) | 72
dopamine given | 72
dopamine continued for 1 week | 72
transfusion of 1 unit packed RBCs continued | 72
transferred back to general ward | 120
follow-up WBC count 12.7 | 120
blood culture showed Escherichia coli | 120
urine culture showed Klebsiella pneumonia | 120
antibiotic changed | 120
abdominal pain | 168
abdominal distention | 168
WBC 13.8 | 168
computed tomography (CT) showed few air bubbles in abdominal cavity | 168
air bubbles in retroperitoneal | 168
air bubbles extending into mediastinum | 168
bowel air at serosal surface of gallbladder | 168
bowel air at serosal surface of omentum | 168
anastomotic leakage | 168
taken back to operating room | 168
diagnostic laparoscopy | 168
laparoscopic Hartmann's sigmoid resection performed | 168
transferred to SICU postoperatively | 168
intubated | 168
inotrope started | 168
CT scan after 10 days | 240
no drainable intra-abdominal collection | 240
discharged | 240
diverticulosis | -4320
previous admissions for diverticulitis | -4320
increased urea | -4320
increased creatinine | -4320
increased potassium | -4320
increased white blood cells (WBCs) | -4320
decreased red blood cells (RBCs) | -4320
decreased hemoglobin | -4320
decreased hematocrit | -4320
decreased bicarbonate | -4320
anastomotic leakage (AL) increases morbidity | -4320
anastomotic leakage (AL) increases mortality | -4320
diverticula in the distal descending colon |6
fever |72
temperature of 38.9°C |72
septic screening |72
urinary tract infection |72
antibiotics started |72
low hemoglobin |72
blood transfusion |72
hypotensive |72
blood pressure 85/52 mmHg |72
oxygen saturation 94% |72
pulse rate 110/min |72
transfusion stopped |72
hydrocortisone started |72
transferred to surgical intensive care unit (SICU) |72
dopamine given |72
dopamine continued for 1 week |72
transfusion of 1 unit packed RBCs continued |72
transferred back to general ward |120
follow-up WBC count 12.7 |120
blood culture showed Escherichia coli |120
urine culture showed Klebsiella pneumonia |120
antibiotic changed |120
abdominal pain |168
abdominal distention |168
WBC 13.8 |168
computed tomography (CT) showed few air bubbles in abdominal cavity |168
air bubbles in retroperitoneal |168
air bubbles extending into mediastinum |168
bowel air at serosal surface of gallbladder |168
bowel air at serosal surface of omentum |168
anastomotic leakage |168
taken back to operating room |168
diagnostic laparoscopy |168
laparoscopic Hartmann's sigmoid resection performed |168
transferred to SICU postoperatively |168
intubated |168
inotrope started |168
CT scan after 10 days |240
no drainable intra-abdominal collection |240
discharged |240
diverticulosis |-4320
previous admissions for diverticulitis |-4320
increased urea |-4320
increased creatinine |-4320
increased potassium |-4320
increased white blood cells (WBCs) |-4320
decreased red blood cells (RBCs) |-4320
decreased hemoglobin |-4320
decreased hematocrit |-4320
decreased bicarbonate |-4320
anastomotic leakage (AL) increases morbidity |-4320
anastomotic leakage (AL) increases mortality |-4320
