50 years old | 0
male | 0
Japanese | 0
admitted to the hospital | 0
fever | -336
loss of appetite | -336
watery diarrhea | -336
heavy drinker | -8760
consumed approximately 250 g of alcohol per day | -3360
increased WBC count | -336
C-reactive protein level increased | -336
total bilirubin level increased | -336
prothrombin time increased | -336
hepatomegaly | -336
splenomegaly | -336
diffuse edematous colon | -336
infectious enteritis | -336
abstained from alcohol | -336
prescribed antibiotics | -336
WBC count increased | -336
total bilirubin level increased | -336
prothrombin time decreased | -336
renal failure progressed | -336
transferred to hospital | -336
jaundice | 0
anuria | 0
ascites | 0
pretibial edema | 0
hepatic encephalopathy | 0
flapping tremor | 0
WBC count increased | 0
total bilirubin level increased | 0
aspartate aminotransferase increased | 0
alanine aminotransferase increased | 0
NH3 increased | 0
albumin decreased | 0
blood urea nitrogen increased | 0
creatinine increased | 0
C-reactive protein level increased | 0
procalcitonin increased | 0
prothrombin time increased | 0
interleukin-6 increased | 0
tumor necrosis factor-alpha increased | 0
diagnosed with severe AH | 0
Maddrey discriminant function score calculated | 0
Glasgow alcoholic hepatitis score calculated | 0
infection with multidrug resistance bacteria | 0
received plasma exchange | 0
received hemodialysis | 0
received antibiotics | 0
granulocytapheresis performed | 168
WBC count decreased | 168
total bilirubin level decreased | 168
pro-inflammatory cytokines decreased | 168
interleukin-6 decreased | 168
tumor necrosis factor-alpha decreased | 168
diarrhea improved | 336
fever improved | 336
laboratory parameters improved | 336
renal failure improved | 336
discharged from hospital | 1680