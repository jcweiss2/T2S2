35 years old | 0
female | 0
admitted to the hospital | 0
history of three episodes of generalized tonic–clonic seizures | -3
urinary incontinence | -3
altered sensorium | -3
headache | -3
unsafe abortion | -240
severe fatigue | -240
shortness of breath | -240
pedal edema | -240
husband expired | -1095
severe anemia | -240
blood transfusion | -240
transfused five units of blood | -240
no history of hypertension | 0
vital signs were normal | 0
drowsy | 0
not obeying commands | 0
withdraws limbs to painful stimuli | 0
deep tendon reflexes were sluggish | 0
withdrawal response was seen in plantar reflex | 0
no signs of meningeal irritation | 0
normal hemoglobin | 0
neutrophilic leukocytosis | 0
urinary tract infection | 0
elevated C-reactive protein | 0
normal ESR | 0
normal liver function tests | 0
normal renal function tests | 0
dimorphic anemia | 0
normal coagulation profile | 0
normal autoantibodies | 0
normal neoplastic markers | 0
increased protein level in cerebrospinal fluid | 0
normal chest radiography | 0
normal arterial blood gas analysis | 0
bilateral occipital, parietal, frontal cortex and subcortical white matter T2/Fluid-attenuated inversion recovery (FLAIR) hyperintensities | 0
bilateral temporal–occipital epileptiform discharges | 0
incomplete right bundle branch block | 0
admitted to intensive care unit | 0
managed with intravenous fluids | 0
managed with antibiotics | 0
managed with antiepileptics | 0
monitoring of blood pressure | 0
improved symptomatically | 168
normal sensorium | 168
normal leukocyte counts | 168
normal vital signs | 168
discharged | 168
follow-up after 1 week | 336
uneventful follow-up | 336