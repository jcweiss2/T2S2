37 years old | 0
female | 0
transposition of the great arteries | -0
ventricular septal defect | -0
pulmonary stenosis | -0
surgical correction | -0
atrial switch procedure | -0
Mustard operation | -0
ventricular septal defect closure | -0
valved conduit implant | -0
high-grade atrioventricular block | -168
pacemaker implant | -168
drug-resistant pneumonia | -112
i.v. antibiotics | -112
fever spikes | -56
hospitalization | -56
septic shock | 0
severe acute respiratory failure | 0
mechanical ventilation | 0
multiple mobile vegetations | 0
mitral valve leaflets | 0
intraventricular abscess | 0
systemic embolization | 0
necrosis of extremities | 0
pulmonary infarction | 0
ischemic areas in spleen | 0
ischemic areas in kidneys | 0
cerebral haemorrhage | 0
methicillin-resistant Staphylococcus aureus | 0
antibiotic therapy | 4
daptomycin | 4
infected pacemaker lead extraction | 6
temporary device implant | 6
urgent neurosurgical procedure | 8
haematoma evacuation | 8
multiorgan failure | 16
death | 20