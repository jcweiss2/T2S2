62 years old | 0
male | 0
caucasian | 0
admitted to the hospital | 0
dyspnea | 0
cough | 0
body condition loss | 0
non-small cell lung cancer | -24
high PD-L1 expression | -24
tumor mass | -24
bilateral necrotic adrenal metastases | -24
hypertension | -24
chronic obstructive pulmonary disease | -24
peripheral arterial disease | -24
exertional dyspnea | 0
productive cough | 0
decrease in right apical vesicular lung sound | 0
painless palpable mass in the right hypochondrium | 0
bronchial fibroscopy | 0
wild-type Streptococcus pneumoniae | 0
amoxicillin-clavulanic acid | 2
fever | 4
chills | 4
new fibroscopy | 4
blood culture samples | 4
leukocyte count grew | 6
anaerobic blood bottle culture positive | 4
Gram-positive coccobacilli | 4
central venous catheter | -1
chemo-immunotherapy cycle | 5
Carboplatin-Pemetrexed-Pembrolizumab | 5
granulocyte colony-stimulating factor | 5
Catabacter hongkongensis | 9
respiratory status declined | 11
oxygen flow rate | 11
hypotensive | 11
oliguria | 11
poor peripheral perfusion | 11
hyperlactatemia | 11
vascular filling | 11
piperacillin-tazobactam | 11
amikacin | 11
septic shock | 23
imipenem/cilastatin | 21
death | 27