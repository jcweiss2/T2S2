67 years old|0
    female|0
    obese|0
    plasma cell leukemia|0
    generalized tiredness|-24
    altered sensorium|-24
    treatment for malignancy for 2 years|-17520
    patent airway|0
    bilateral crackles at lung base|0
    respiratory rate 30 cycles/min|0
    Spo2 70% in room air|0
    feeble peripheral pulses|0
    un-recordable blood pressure|0
    heart rate 120 bpm|0
    responding to verbal stimulus|0
    normal finger stick glucose levels|0
    pale|0
    jugular venous distension|0
    bilateral pitting pedal edema|0
    muffled heart sounds|0
    no audible murmurs|0
    no friction rubs|0
    no focal neurologic deficits|0
    bilaterally equal pupils|0
    other physical exam findings within normal limits|0
    started on IV fluid resuscitation|0
    cautious monitoring for volume overload worsening|0
    failed to respond to fluid therapy|0
    started on vasopressor|0
    started on inotrope supports|0
    intubated in ED|0
    clinical features consistent with BECK's triad|0
    diagnosed with cardiac tamponade|0
    placed on continuous cardiac monitoring|0
    supplemental oxygen through ventilator|0
    bedside goal-directed ECHO performed|0
    diagnosed with massive pericardial effusion|0
    right ventricular collapse during diastole|0
    plethoric IVC|0
    emergency pericardiocentesis|0
    counseling and consent|0
    performed procedure with central venous catheter under sonographic guidance|0
    used PHASED ARRAY probe (2.5–5 MHz)|0
    revealed 42 mm thickness effusion inferiorly|0
    aseptic precautions|0
    marked area inferior to left xiphoid under sterile conditions|0
    local anesthetic applied|0
    trocar needle introduced angled at 30°|0
    aiming toward left shoulder|0
    pericardial sac punctured|0
    pericardial fluid aspirated|0
    noted needle tip in pericardium|0
    active aspiration performed using 3-way stopcock valve with syringe|0
    250 ml of fluid aspirated|0
    patient reassessed|0
    well perfused|0
    audible heart sounds|0
    normal JVD|0
    heart globally expanded within pericardium|0
    aspiration stopped|0
    transferred to intensive care team|0
    further management|0
    placement of pericardial drain insitu|0
    cardiac tamponade|0
    pericardial effusion|0
    pericardiocentesis|0
    right ventricular collapse|0
    plethoric inferior vena cava|0
    globally expanded heart|0
    