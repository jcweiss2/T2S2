35 years old | 0
female | 0
admitted to her local hospital | 0
fever | 0
tachycardia | 0
neutropenia | 0
tonsillitis | 0
suspected sepsis | 0
diagnosis of thyroid storm | 0
autoimmune hyperthyroidism | -8760
treated with thionamide | -8760
thionamide discontinued | -8688
signs and symptoms of hyperthyroidism | -672
free thyroxine | -672
free triiodothyronine | -672
thionamide and non-selective beta-blocker prescribed | -672
thionamide discontinued | -48
admitted to hospital | 0
treatment with beta-blocker | 0
treatment with antibiotics | 0
treatment with glucocorticoids | 0
treatment with iodine solution | 72
circulatory collapse | 96
pulseless electrical activity | 96
cardiopulmonary resuscitation | 96
return of spontaneous circulation | 96
transferred to university hospital | 96
severe biventricular cardiac failure | 96
inotropic support with dobutamine | 96
recurrent cardiac arrests | 96
established on V-A ECMO support | 96
iodine solution dosages increased | 96
levosimendan infusion started | 96
complete recovery of myocardial function | 168
V-A ECMO circuit discontinued | 168
extubated | 168
surgery with total thyroidectomy | 288
discharged | 672
no cognitive sequelae | 672
normalized cardiac function | 672
close follow-up by endocrinologist | 672
Grave’s disease | -8760
Grave’s ophthalmopathy | 96
severe lactic acidosis | 96
pulmonary embolism suspected | 96
computed tomography pulmonary angiography | 96
thrombolysis | 96
CT scan performed | 96
pulmonary embolism excluded | 96
coronary angiography | 96
normal coronary arteries | 96
intra-aortic balloon pump inserted | 96
thyroid hormone levels normalized | 168
beta-blockers discontinued | 168
levosimendan commenced | 168
myocardial function recovered | 168
total thyroidectomy performed | 288
levothyroxine substitution started | 288