38 years old | 0
male | 0
Caucasian | 0
living in Tanzania | 0
admitted to the hospital | 0
fever | -144
chills | -144
cough | -144
history of asthma | -144
treated for bronchitis | -144
left upper quadrant abdominal pain | -120
abdominal pain radiated to left shoulder | -120
severe hypotension | -120
malaria blood slide positive | -120
ultrasound showed fluid in abdomen | -120
given artesunate | -120
referred to facility | -120
sick-looking | 0
mildly pale | 0
jaundiced | 0
tachycardia | 0
normal blood pressure | 0
slightly distended abdomen | 0
mild generalized tenderness | 0
no acute peritonitis | 0
low hemoglobin | 0
normal red cell indices | 0
Mean Corpuscular Volume | 0
Mean Corpuscular Hemoglobin | 0
repeat blood slide for malaria showed parasitemia | 0
Plasmodium falciparum | 0
management for severe malaria started | 0
parenteral artemether | 0
oral doxycycline | 0
CT scan abdomen with intravenous contrast | 0
free peritoneal fluid | 0
no obvious splenic rupture | 0
no contrast extravasation | 0
monitored closely in intensive care unit | 0
repeat hemoglobin levels | 0
hemoglobin continued to fall | 16
resuscitation with two pints whole blood | 16
abdominal distension worsened | 16
abdominal pain worsened | 16
exploratory laparotomy | 16
frank blood | 16
no purulence | 16
no fecal contamination | 16
spleen enlarged | 16
splenic laceration | 16
laceration actively bleeding | 16
splenectomy | 16
postoperatively recovered | 24
discharged home | 192
atovaquone/proguanil for malaria prophylaxis | 192
asplenic state | 192