22 years old | 0
male | 0
admitted to intensive care unit (ICU) | 0
fever | -240
cough | -192
sputum production | -192
respiratory distress | -24
altered sensorium | -24
no history of hospitalization within past 1 year | -8760
altered sensorium | 0
tachycardic | 0
tachypnea | 0
hypotensive | 0
heart rate-130/min | 0
blood pressure-90/60 mm Hg | 0
hypoxemia | 0
right lower lobe consolidation | 0
haemoglobin-9.3 g% | 0
white blood cell (WBC) count-3,500/cu.mm | 0
platelets-80,000/cu.mm | 0
serum creatinine-1.8 mg/dl | 0
normal liver function test | 0
normal general blood picture | 0
intubated | 0
mechanical ventilation | 0
bronchoalveolar lavage (BAL) | 0
blood samples sent for culture and sensitivity testing | 0
provisional diagnosis of acute febrile illness | 0
pneumonia | 0
septic shock | 0
started on piperacillin-tazobactum | 0
vancomycin | 0
antimalarials | 0
tests for malaria | 0
tests for leptospirosis | 0
tests for dengue | 0
tests for typhoid | 0
all tropical infective profile tests negative | 0
PaO2/FiO2 ratios 100 | 0
ventilated as per acute respiratory distress syndrome (ARDS) net protocol | 0
prone ventilation | 0
blood cultures positive for MRSA | 0
BAL cultures positive for MRSA | 0
i.v. vancomycin added | 0
PaO2/FiO2 ratios improved (P/F > 300) | 168
extubated | 168
continuing hypoxia | 168
respiratory rate of 28-30/min | 168
computed tomography pulmonary angiogram | 96
high resolution computed tomography chest | 96
patchy consolidation with cavity in lateral basal segment of right lower lobe | 96
pulmonary angiogram normal | 96
continued on vancomycin for 3 weeks | 168
respiratory rate settled | 672
discharged after 28 days of ICU stay | 672
diffuse consolidation with air bronchograms | 96
consolidation and areas of cavitation | 96
right-sided pleural effusion | 96
no hemoptysis | 0
bronchoscopy showed no hemorrhage | 0
diffuse cavitations and necrosis | 96
MRSA resistant to penicillinase-resistant penicillins | 0
MRSA sensitive to macrolides | 0
MRSA sensitive to quinolones | 0
MRSA sensitive to linezolid | 0
MRSA sensitive to clindamycin | 0
MRSA sensitive to vancomycin | 0
leucopenia | 0
low platelet count | 0
severe hypoxemia | 0
cavitary pulmonary infiltrates | 96
no airway bleeding | 0
ARDS | 0
inotrope support | 0
artificial ventilation | 0
severe leucopenia | 0
WBC counts less than 2500/cu.mm | 0
leucopenia as ominous prognostic factor | 0
Panton-Valentine leukocidin (PVL) affinity for neutrophils leading to lysis | 0
WBC count as inverse biomarker of PVL burden | 0
no prior MRSA infection | -8760
no indwelling devices | -8760
CA-MRSA pneumonia | 0
necrotizing pneumonia | 0
multiorgan failure | 0
shock | 0
no pulmonary embolism | 96
patchy consolidation | 96
cavity in right lower lobe | 96
no Klebsiella pneumonia | 0
no Pseudomonas aeruginosa | 0
no Nocardia | 0
no Actinomyces | 0
no anaerobes | 0
community-acquired pneumonia | 0
CA-MRSA | 0
