6-day-old premature female newborn | 0
    18-year-old gravida one woman | 0
    fever | -168
    prolonged premature rupture of membranes | -168
    admitted to the hospital | 0
    betamethasone | 0
    ampicillin | 0
    gentamicin | 0
    worsening maternal respiratory distress | 0
    mechanical ventilation | 0
    failure to progress after induction | 0
    PPROM | -168
    suspected chorioamnionitis | 0
    emergency cesarean section delivery | 0
    born at 28 weeks and 1 day gestation | 0
    birth weight 1140 gm | 0
    mechanical ventilation at birth | 0
    intravenous ampicillin | 0
    intravenous gentamicin | 0
    discontinued ampicillin | 48
    discontinued gentamicin | 48
    blood cultures negative | 48
    extubated successfully | 24
    noninvasive ventilation | 24
    less active | 96
    temperature instability | 96
    bradycardia | 96
    vancomycin | 96
    cefotaxime | 96
    multiple episodes of apnea | 96
    deteriorating bradycardic spells | 96
    desaturation | 96
    hypercarbia | 96
    re-intubated | 96
    synchronized intermittent mandatory ventilation | 96
    antibiotics changed to cefepime | 96
    antibiotics changed to fluconazole | 96
    antibiotics changed to acyclovir | 96
    increasing metabolic acidosis | 120
    worsening respiratory failure | 120
    high frequency oscillating ventilation | 120
    condition continued to deteriorate | 120
    hypotensive | 120
    poor perfusion despite vasopressors | 120
    blood products | 120
    bedside echocardiogram revealed normal-appearing heart | 120
    patent ductus arteriosus | 120
    left-to-right shunt | 120
    pulmonary hypertension | 120
    small pericardial effusion | 120
    moderately decreased left ventricular function | 120
    signs of low cardiac output | 120
    sepsis | 120
    severe metabolic acidosis | 120
    disseminated intravascular coagulation | 120
    antibiotic therapy | 120
    antifungal therapy | 120
    antiviral therapy | 120
    cardiopulmonary arrest | 160
    passed away | 160
    mucocutaneous culture sampled | 96
    HSV positive | 160
    placental pathology third-trimester placenta | 0
    moderate intervillous fibrosis | 0
    no evidence of chorioamnionitis | 0
    no funisitis | 0
    autopsy normally developed premature female infant | 0
    no dysmorphic features | 0
    no congenital anomalies | 0
    body weight 1525 gm | 0
    serous fluid in right pleural cavity | 0
    serous fluid in left pleural cavity | 0
    serous fluid in pericardial sac | 0
    serosanguineous ascites | 0
    normal-sized heart | 0
    unremarkable immature myocardium | 0
    open ductus arteriosus | 0
    open foramen ovale | 0
    hemorrhagic right upper lobe | 0
    hemorrhagic middle lobe | 0
    thickened septa | 0
    saccular stage of development | 0
    disorganized large cells without cilia | 0
    viral nuclear inclusions | 0
    diffuse fibrin plugs in bronchioles | 0
    diffuse alveolar hemorrhage | 0
    bloody mucus in stomach | 0
    normal mucosa | 0
    liver weight 65 gm | 0
    red-brown parenchyma | 0
    centrilobular congestion | 0
    hemorrhage around portal areas | 0
    hemorrhage under the capsule | 0
    viral inclusions in hepatocyte nuclei | 0
    margination of chromatin | 0
    molding | 0
    HSV positive in hepatocytes | 0
    peripelvic hemorrhage | 0
    no herpetic infection in kidneys | 0
    karyorrhexis | 0
    perivascular cell fragments | 0
    unremarkable CNS | 0
    microglial nodules in midbrain | 0
    microglial nodules in thalamus | 0
    HSV isolated from postmortem lung cultures | 0
    resolving hyaline membrane disease | 0
    disseminated HSV infection of liver | 0
    disseminated HSV infection of lung | 0
    disseminated HSV infection of brain | 0
    ascites | 0
    pleural effusion | 0
    persistent ductus arteriosus | 0
    involution of thymus | 0
    medullary congestion | 0
    pelvic hemorrhage of kidneys | 0
    