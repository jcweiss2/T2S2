78 years old | 0
male | 0
admitted to the hospital | 0
dyspnea | -240
shortness of breath | -240
cough | -240
anosmia | -240
myalgia | -240
hypertension | -6720
Valsartan | -6720
tachycardia | 0
normal core temperature | 0
hypertension | 0
tachypnea | 0
low oxygen saturation | 0
reduced level of consciousness | 0
SARS-CoV-2 RNA positive | 0
elevated plasma lactate | 0
low albumin | 0
elevated C-Reactive Protein | 0
elevated high sensitivity troponin | 0
elevated creatine kinase myocardial band | 0
diffuse bilateral ground-glass opacities | 0
mild pleural effusion | 0
cardiomegaly | 0
atrial fibrillation | 0
reduced left ventricular ejection fraction | 0
high pulmonary arterial pressure | 0
mildly enlarged left ventricle | 0
moderate to severe left ventricular dysfunction | 0
mild diastolic dysfunction | 0
mild mitral valve regurgitation | 0
normal septal thickness | 0
intubation | 0
transfer to ICU | 0
low systemic vascular resistance | 0
low cardiac output | 0
low delivery of oxygen | 0
cardiogenic shock | 0
septic shock | 0
Hydroxychloroquine treatment | 0
Dexamethasone treatment | 0
Intravenous Immunoglobulin treatment | 0
Ascorbic acid treatment | 0
Melatonin treatment | 0
broad-spectrum antibiotics | 0
vasopressor treatment | 0
amiodarone treatment | 0
Midodrine treatment | 0
echocardiographic measurement on day 25 | 600
left ventricular ejection fraction 25% on day 25 | 600
pulmonary arterial pressure 38 mmHg on day 25 | 600
moderate left ventricular dysfunction on day 25 | 600
right ventricular dilation on day 25 | 600
follow-up assessment on day 35 | 840
left ventricular ejection fraction 35% on day 35 | 840
pulmonary arterial pressure 55 mmHg on day 35 | 840
mild right ventricular dilation on day 35 | 840
improved respiratory distress on day 35 | 840
follow-up assessment on day 42 | 1008
left ventricular ejection fraction 45% on day 42 | 1008
pulmonary arterial pressure 45 mmHg on day 42 | 1008
mild right ventricular dilation on day 42 | 1008
discharge from ICU | 1008
respiratory arrest | 1056
cardiopulmonary resuscitation | 1056
death | 1056