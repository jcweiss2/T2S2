14 years old | 0
male | 0
Joubert syndrome | -26208
chronic renal failure | -26208
peritoneal dialysis | -26208
vomiting | -168
intolerance to food intake | -168
hyponatremia | 0
hypopotassemia | 0
hospitalized | 0
supplementation treatment | 0
blood culture | 0
urine culture | 0
peritoneal fluid culture | 0
febrile episodes | 0
IV antibiotherapy with tazobactamDampicillin | 0
Candida spp. growth in peritoneal culture | 0
liposomal amphotericin B | 0
peritoneal dialysis catheter removal | 0
anuric | 0
volume overload | 0
intermittent hemodialysis therapy | 0
abdominal ultrasound | 0
complicated fluidDfilled cystic lesions in pancreatic loge | 0
multiple cortical cysts in kidneys |;0
abdominal CT scan | 0
large cystic lesions compressing gastrointestinal system and intraabdominal organs | 0
loculated fluid collections in peripancreatic area | 0
pediatric surgery evaluation | 0
surgery planned | 0
cyst observed on anterior abdominal wall | 0
cyst rupture | 0
aspiration of 2500 cc serohemorrhagic fluid | 0
cardiac arrest | 0
erythrocyte suspension transfusion | 0
fluid support | 0
adrenaline infusion | 0
noradrenaline infusion | 0
transfer to intensive care unit | 0
blood pressure 55D35 mmHg | 0
heart rate 90 bpm | 0
pupils bilaterally dilated with absent light reflex | 0
capillary refill time 6D7 seconds | 0
arterial blood gas pH 7.15 | 0
PaCO2 41.8 mmHg | 0
PaO2 82.8 mmHg | 0
base excess D13.2 mmolDL | 0
HCO3 14 mmolDL | 0
lactate 16 mmolDL | 0
BUN 87 mgDL | 0
creatinine 2.7 mgDL | 0
mechanical ventilation | 0
saline solution bolus doses | 0
hypotension persistence | 0
dopamine infusion | 0
dobutamine infusion | 0
adrenaline infusion increased | 0
noradrenaline infusion increased | 0
erythrocyte suspension for hemoglobin 2.8 grDL | 0
thrombocyte suspension for platelet count 22.000Dmm3 | 0
4 erythrocyte suspensions over 12 hours | 0
IV fresh frozen plasma | 0
procalcitonin 12.59 ngDLmL | 0
combined antibiotherapy with meropenem | 0
vancomycin | 0
amikacin | 0
metronidazole added | 0
IV steroid administered | 0
femoral vein catheter insertion | 0
PiCCO monitoring | 0
cardiac index 6.5 LDminute | 0
SVRI 338 dynesDsecondDcm5Dm2 | 0
GEDI 780 mLDm2 | 0
EVLWI 15 mLDkg | 0
SBP 67 mmHg | 0
DBP 32 mmHg | 0
MAP 46 mmHg | 0
pulse rate 106Dminute | 0
TP bolus 10 µgDkg | 0
family consent obtained | 0
blood pressure increase after TP | 0
SBP 94 mmHg | 0
DBP 45 mmHg | 0
MAP 60 mmHg | 0
TP infusion 1 µgDkgDminute | 0
noradrenaline dose reduced to 0.7 µgDkgDminute | 0
cardiac index decrease | 0
heart rate decrease | 0
SVRI increase | 0
GEDI increase | 0
EVLWI increase | 0
CVVH initiated | 0
1000 cc ultrafiltrate aspirated | 0
BUN 27 mgDL | 0
creatinine 1.9 mgDL | 0
GEDI decrease | 0
ELWI decrease | 0
ischemic manifestations on right big toe | 9
TP infusion discontinuation | 9
SBP 69 mmHg | 10
DBP 46 mmHg | 10
MAP 54 mmHg | 10
cardiac arrest | 13
cardiopulmonary resuscitation | 13
patient death | 13
