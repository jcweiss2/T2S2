Here is the table of events and timestamps:

29 years old | 0
male | 0
hospitalized for cardiogenic shock | -672
diagnosed with biventricular failure | -672
imaging concerning for myopericarditis and constrictive physiology | -672
peripherally inserted central catheter (PICC) line placed | -672
discharged on milrinone | -672
presented to Emergency Department with septic shock | -144
PICC line removed | -144
started on IV vancomycin and piperacillin/tazobactam | -144
transferred to intensive care unit for vasopressor support | -144
Chryseobacterium indologenes grew from his admission PICC line and peripheral blood cultures | -120
PICC line dressing became contaminated with tap water | -120
antibiotics were changed to ciprofloxacin and piperacillin/tazobactam | -120
he was weaned off vasopressor support | -96
underwent pericardiectomy | -72
completed 14 days of antibiotics | -72
discharged from the hospital off inotropes with stable vital signs and labs | -72
seen in outpatient cardiology clinic, remains in good health with no evidence of recurrent infection | 672
progressive fatigue and dyspnoea on exertion for 2–3 months | -1008
hospitalized for non-ischaemic cardiomyopathy | -1008
diagnosed with non-ischaemic cardiomyopathy | -1008
computed tomography angiography of the coronary arteries revealed cardiomegaly | -1008
echocardiogram showed biventricular failure | -1008
cardiac magnetic resonance imaging showed a left ventricular ejection fraction (EF) of 23% | -1008
diastolic septal bounce and a concentrically thickened pericardium | -1008
atrial flutter with rapid ventricular response requiring radiofrequency ablation | -1008
cardiogenic shock | -1008
stabilized on inotrope therapy | -1008
discharged on home milrinone infusion via a peripherally inserted central catheter (PICC line) | -1008
fever of 38.7°C (101.8°F) and chills for 1 day at home | -96
tachycardia with a heart rate in the 110s | -96
blood pressure of 96/57 mmHg | -96
heart that was tachycardic, but normal rhythm without any murmurs, rubs, or gallops | -96
no signs of elevated jugular venous pressure and he did not have lower extremity oedema | -96
bilateral radial and dorsalis pedis pulses were equal and 2+ bilaterally | -96
lungs were clear to auscultation bilaterally in the anterior and posterior lung fields with a normal work of breathing | -96
no redness or drainage around the PICC line | -96
Chest X-ray showed no abnormalities | -96
electrocardiogram was significant for sinus tachycardia | -96
sinus tachycardia, normal axis, RSR′ pattern in V1, QRS duration of 90 ms, and non-specific T wave flattening in the inferolateral leads | -96
removed his PICC line | -96
became febrile to 39.5°C (103.1°F) and developed severe rigours as well as hypotension with blood pressure in 70s/40s mmHg | -96
elevated lactate level of 5.5 mmol/L | -96
blood cultures were drawn both peripherally and from the PICC line | -96
started on empiric vancomycin and piperacillin/tazobactam | -96
transferred to the cardiac intensive care unit for vasopressor support | -96
Gram-negative rods which later speciated as Chryseobacterium indologenes | -96
PICC line as the most likely source of infection | -96
antibiotics were changed to ciprofloxacin and piperacillin/tazobactam | -96
he was weaned off vasopressor support | -48
underwent pericardiectomy | -24
completed 14 days of antibiotics | -24
discharged from the hospital off inotropes with stable vital signs and labs | -24
seen in outpatient cardiology clinic, remains in good health with no evidence of recurrent infection | 672