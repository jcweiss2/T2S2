55 years old | 0
female | 0
gastric adenocarcinoma | -672
abdominal metastases | -672
surgery | -672
poorly differentiated adenocarcinoma | -672
signet-ring cell carcinoma | -672
CerbB-2 2+ | -672
Ki67+ | -672
Syn− | -672
CgA− | -672
CerbB-2 gene amplification negative | -672
first-line palliative chemotherapy | -504
oxaliplatin | -504
S-1 | -504
stable disease | -336
maintenance treatment | -336
S-1 | -336
cardiac obstruction | -240
ENFTP | -240
second-line chemotherapy | -168
albumin-bounded paclitaxel | -168
oxaliplatin | -168
obstructive symptoms relieved | -84
feeding tube removed | -84
grade 4 neutropenia | -84
rh-GCSF | -84
disease progression | -56
best supportive care | -56
incomplete gastrointestinal obstruction | -56
apatinib | 0
nausea | 0
vomiting | 0
abdominal pain | 0
blood pressure rose | 0
gastrointestinal hemorrhage | 456
fecal occult blood test positive | 456
hematemesis | 456
apatinib stopped | 480
severe abdominal pain | 480
gastrointestinal perforation | 480
septic shock | 480
emergency operation | 480
purulent ascites | 480
perforated ulcer | 480
miliary nodules | 480
ileal tumor | 480
metastatic signet-ring cell carcinoma | 480
MODS | 528
death | 744