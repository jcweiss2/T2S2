84 years old | 0
male | 0
admitted to the hospital | 0
edema of the right leg | -168
fever | -168
no history of cardiovascular disease | 0
no specific diseases | 0
fully conscious | 0
pulse rate 70 beats/min | 0
blood pressure 120/80 mm Hg | 0
temperature 37.5°C | 0
pulsatile mass in the abdomen | 0
white blood cells 4.6 × 10^3/μL | 0
hemoglobin 11 g/dL | 0
C-reactive protein 3.6 mg/dL | 0
high levels of D-dimer | 0
high levels of creatinine | 0
high levels of soluble interleukin 2 receptor | 0
infrarenal AAA | 0
bilateral common iliac artery aneurysms | 0
periaortic soft tissue density | 0
deep venous thrombosis | 0
hydronephrosis | 0
vitamin K antagonist therapy | 0
suprarenal inferior vena cava filter placement not performed | 0
lower leg swelling decreased | 24
plain MRI scans | 24
hyperintense signal at the periaortic lesion | 24
compatible with malignant lymphoma | 24
open biopsy | 96
diagnosis of diffuse large B-cell lymphoma | 96
sepsis due to urinary tract infection | 96
mechanical ventilation | 96
endotoxin adsorption therapy | 96
recovered from sepsis | 216
recovered from respiratory failure | 216
preliminary informed consent | 216
no therapeutic intervention for unilateral hydronephrosis | 216
no therapeutic intervention for right urinary tract compression | 216
EVAR | 432
right internal iliac artery embolization | 336
left internal iliac artery embolization | 432
completion angiography | 432
no postoperative aortic events | 432
no chemotherapy for malignant lymphoma | 1176
discharged | 1176
follow-up CT scans | 1192
no change in the size of aneurysm | 1192
no change in the size of lymphoma | 1192