pre-syncope | -0.1
syncope | 0
left-sided chest tightness | 0
generalized fatigue | -96
weight loss | -96
diffuse erythematous rash | 0
unremarkable cardiac examination | 0
unremarkable respiratory examination | 0
normal sinus rhythm | 0
raised troponin concentration | 0
eosinophil count of 7.6 × 10^9/l | 0
myocarditis | 0
coronary angiography | 12
no evidence of coronary artery disease | 12
skin biopsy | 24
cardiac biopsy | 24
discharged | 48
edoxaban | 48
prednisolone | 48
follow-up in the rheumatology clinic | 336
missed appointment | 720
neck swelling | 720
urgently admitted to hospital | 720
rise in eosinophil count | 720
increase the dose of prednisolone | 720
lymphadenopathy | 720
T-cell lymphoma | 720
chemotherapy with cyclophosphamide | 720
sepsis | 744
cholecystitis | 744
new onset of seizures | 744
reduction in consciousness | 744
Glasgow Coma Scale of 9/15 | 744
multiple bilateral acute infarctions | 744
transfer to the intensive care unit | 744
history of hepatitis B | 0
history of asthma | 0
history of intravenous drug use | 0
history of excessive use of alcohol | 0
ischemic stroke | 744
reduced GCS score | 744
seizures | 744
intracranial bleeding | 744
malignancy | 744
intracerebral infection | 744
diffuse subendocardial late gadolinium enhancement | 720
mild LV systolic impairment | 720
eczematous changes | 720
no increase in eosinophils | 720
T-cell lymphoma | 720
infarcts involving the frontal, parietal, and left temporo-occipital regions | 744
apical tear | 768
intramural myocardial tear | 768
small apical cavity | 768
mobile structures attached to dissected myocardium | 768
diastolic flow in the apical cavity | 768
systolic flow out of the apical cavity | 768
cardiac thrombus | 768
cyclophosphamide therapy | 768
partial response | 768
reduction of the eosinophil count | 768
palliation | 840