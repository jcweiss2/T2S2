55 years old | 0
male | 0
admitted to the hospital | 0
alcohol use | -2160
necrotizing biliary pancreatitis | -2160
acute portal vein thrombus | -2160
anticoagulation with therapeutic enoxaparin | -2160
large multiloculated peripancreatic fluid collections | -2160
peripancreatic walled-off necrosis (WON) | -2160
EUS-guided cystogastrostomy procedures | -168
lumen-apposing metal stent | -168
double-pigtail catheter | -168
endoscopic necrosectomies | -84
removal of the initial lumen-apposing metal stent | -84
pigtail catheter | -84
placement of 2 double-pigtail catheters | -84
subsequent necrosectomy | -42
replacement of the double-pigtail catheters | -42
persistent WON | -24
inferoposterior extension of peripancreatic necrotic collections | -24
worsening abdominal pain | -12
fevers | -12
sepsis | 0
white blood cell count 29.6 | 0
hemoglobin 8.7 g/dL | 0
international normalized ratio 1.3 | 0
hypotensive | 120
tachycardic | 120
lactic acidosis | 120
worsening anemia | 120
hemoglobin 5.3 g/dL | 120
international normalized ratio 1.9 | 120
activated partial thromboplastin time 26 | 120
retroperitoneal hematoma | 120
intraperitoneal hemorrhage | 120
enoxaparin discontinued | 120
massive transfusion protocol | 120
administration of protamine sulfate | 120
computed tomography angiography | 144
active arterial bleeding | 144
interventional radiology angiogram | 168
L2 and L3 distal lumbar artery focal pseudoaneurysms | 168
extravasation | 168
coil embolization | 168
exploratory laparotomy | 192
evacuation of retroperitoneal and intraperitoneal hematomas | 192
electrical cautery | 192
subsequent surgeries | 240
re-exploration | 240
cholecystectomy | 240
nonobstructive ileus | 240
pleural effusion | 240
thoracentesis | 240
bacteremia | 240
hydronephrosis | 240
esophagogastroduodenoscopy | 720
dilation of the posterior cystogastrostomy | 720
necrosectomy | 720
2 double-pigtail stents | 720
discharged | 720