18 years old | 0
male | 0
admitted to the hospital | 0
fever | -192
abdominal discomfort | -192
anorexia | -192
vomiting | -192
normal before the onset of symptoms | -192
no significant past medical history | 0
no history of alcohol intake | 0
no drug abuse | 0
no blood transfusions | 0
generalized abdominal mild tenderness | 0
febrile | 0
dehydrated | 0
tachycardia | 0
toxic look | 0
low blood pressure | 0
decreased urine output | -24
thrombocytopenia | -24
leukopenia | -24
elevated transaminases | -24
hemoglobin 12 g/dL | -24
bilirubin within normal limits | -24
admitted to the ICU | 0
enteric fever | 0
malaria | 0
leptospirosis | 0
normal hemoglobin | 24
leukopenia | 24
thrombocytopenia | 24
deranged liver function tests | 24
grossly deranged kidney function tests | 24
urea 208 mg/dL | 24
creatinine 12.2 mg/dL | 24
uric acid 16.5 mg/dL | 24
started on hemodialysis | 24
negative tests for malaria | 24
negative IgM anti-HAV | 24
negative IgM anti-HEV | 24
negative HBsAg | 24
negative dengue serology | 24
proteinuria | 24
hematuria | 24
no casts | 24
normal chest X-ray | 24
normal 2D-echocardiography | 24
hepatosplenomegaly | 24
splenic infarcts | 24
bulky distal body and tail of pancreas | 24
mild ascites | 24
elevated amylase | 24
elevated lipase | 24
multiorgan involvement | 24
negative autoimmune workup | 24
ruled out rickettsia | 24
ruled out post streptococcal glomerulonephritis | 24
negative Weil–Felix | 24
negative ASO titer | 24
negative COVID-19 RT-PCR | 24
negative leptospiral serology | 24
negative urine culture | 24
myalgia | 48
leg pains | 48
elevated creatinine phosphokinase | 48
blood culture grew S. enterica serovar typhi | 96
complicated by acute hepatitis | 96
complicated by acute pancreatitis | 96
complicated by splenic infarcts | 96
complicated by acute renal failure | 96
complicated by rhabdomyolysis | 96
started on intravenous antibiotics | 96
blood transfusions | 96
hemodialysis | 96
lower gastrointestinal bleeding | 120
drop in hemoglobin | 120
fresh frozen plasma transfusions | 120
vitamin K injections | 120
afebrile | 168
no gastrointestinal bleed | 168
hemoglobin stabilized | 168
good urine output | 168
creatinine 2.4 mg/dL | 168
discharged on intravenous antibiotics | 168
follow-up | 216
kidney function within normal limits | 216
transaminases within normal limits | 216
creatinine phosphokinase within normal limits | 216