75 years old | 0
male | 0
admitted to the hospital | 0
fever | -168
chills | -168
dizziness | -168
remission after fever | -168
hypertension | 0
no headache | 0
no abdominal pain | 0
no diarrhea | 0
no sputum | 0
no nasal congestion | 0
no runny nose | 0
temperature 39 °C | 0
heart rate 98 bpm | 0
respiratory rate 20 breaths per minute | 0
blood pressure 139/75 mmHg | 0
oxygen saturation 98% | 0
clear breath sounds | 0
uniform heart rhythm | 0
negative neurological tests | 0
white blood cell count 7.1 × 109/L | 0
neutrophils 58.6% | 0
monocytes 24.4% | 0
hemoglobin 83 g/L | 0
CRP 111.20 mg/L | 0
IL-6 279.22 pg/mL↑ | 0
IL-10 3653.30 pg/mL↑ | 0
procalcitonin 0.19 ng/mL | 0
blood amyloid A 509.5 mg/L↑ | 0
erythrocyte sedimentation rate 71 mm/L | 0
lactate dehydrogenase 694 U/L↑ | 0
creatine kinase 19 U/L↓ | 0
albumin 27 g/L↓ | 0
K+ 2.99 mmol/L↓ | 0
Na+ 135.1 mmol/L↓ | 0
Cl. 98.5 mmol/L↓ | 0
calcium 1.87 mmol/L↓ | 0
phosphorus 0.65 mmol/L↓ | 0
normal creatinine | 0
anti-nuclear antibody positive | 0
anti-SSA positive | 0
anti-SCL70 positive | 0
normal TORCH test | 0
normal Plasmodium test | 0
normal fungal D-glucan test | 0
normal coronavirus disease 2019 | 0
normal hemorrhagic fever IgM antibody | 0
normal Widder test | 0
normal Weil Felix reaction | 0
bilateral blood culture positive for L. monocytogenes | 0
cerebrospinal fluid nucleated cell count 420 × 106/L | 0
cerebrospinal fluid lymphocyte 75% | 0
cerebrospinal fluid lactate dehydrogenase 472 U/L | 0
cerebrospinal fluid total protein 261.3 mg/dL | 0
cerebrospinal fluid glucose 1.51 mmol/L | 0
cerebrospinal fluid chloride 111.0 mmol/L | 0
cerebrospinal fluid adenosine deaminase 16 U/L | 0
cerebrospinal fluid cryptococcal smear negative | 0
cerebrospinal fluid cryptococcal capsular antigen test negative | 0
cerebrospinal fluid culture negative | 0
cerebrospinal fluid metagenomic test positive for L. monocytogenes | 0
CRP changes | 0
IL>6 changes | 0
IL>10 changes | 0
PCT changes | 0
chest CT small pleural effusion | 0
nodules in pleura and subpleura | 0
no cranial CT abnormalities | 0
multiple lung nodules | 0
scattered patchy shadows | 0
possible infection | 0
pleural effusion decreased | 0
cranial MR abnormal signals | 0
lacunar foci under frontal cortex | 0
transparent interstitial space | 0
sepsis | 0
lung infection | 0
respiratory failure | 0
electrolyte imbalance | 0
hyponatremia | 0
hypokalemia | 0
autoimmune disease | 0
Listeria monocytic meningoencephalitis | 0
levofloxacin administration | 0
fever persisted | 0
blood culture penicillin-resistant Staphylococcus | 0
vancomycin administration | 0
temperature normalization | 24
vancomycin stopped | 168
discharged | 168
high fever recurrence | 192
maximum temperature 39.7 °C | 192
chills | 192
cough | 192
thick sputum | 192
no chest pain | 192
no limb twitching | 192
sluggish pupillary light reflex | 192
confusion | 192
soft mentality | 192
brief communication | 192
uncooperative muscle strength test | 192
voluntary activities | 192
diarrhea | 192
ICU admission | 192
high-frequency oxygen inhalation | 192
piperacillin/tazobactam administration | 192
methylprednisolone administration | 192
repeated fever | 192
levofloxacin administration | 192
temperature normalization | 192
CRP reduction | 192
transfer to respiratory ward | 192
atrial fibrillation | 192
unresponsiveness | 192
slurred speech | 192
shortness of breath | 192
slow light reflexes | 192
stiff neck | 192
increased muscle tone | 192
wet rales | 192
critical condition | 192
blood pressure drops | 192
septic shock | 192
active rehydration | 192
norepinephrine micropump | 192
vancomycin adjustment | 192
meropenem administration | 192
ICU transfer | 192
methylprednisolone reduction | 192
methylprednisolone stopped | 192
unconsciousness | 216
tongue base fallback | 216
shortness of breath | 216
stiff neck | 216
limb tremor | 216
heart rate 40 bpm | 216
tracheal intubation | 216
ventilator-assisted breathing | 216
condition deterioration | 216
repeated high fever | 216
septic shock | 216
multiple organ failure | 216
decreased consciousness | 216
fluid resuscitation | 216
norepinephrine administration | 216
ventilator-assisted ventilation | 216
treatment discontinued | 216
