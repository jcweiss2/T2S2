84 years old | 0
female | 0
diabetes mellitus | 0
hypertension | 0
paroxysmal atrial fibrillation | 0
old cerebrovascular event (left middle cerebral artery infarction) | 0
no residual weakness | 0
ambulatory | 0
acceptable cardiorespiratory status | 0
fall | -168
admitted to the hospital | 0
left intertrochanteric femur fracture | 0
Gama nailing of the femur | 24
postoperative course uneventful | 24 to 168
right-sided hemiparesis | 168
altered mental status | 168
Glasgow coma scale (GCS) 10/15 (E4, V1, M5) | 168
NCCT of the brain suggested bilateral CSF hygroma | 168
referred to a neurosurgeon | 168
left parietal Burr hole and evacuation of CSF hygroma | 168
extubated | 168
remained in ICU for neuro observation | 168
GCS 15/15 (E4, V5, M6) | 168
persistent right-sided hemiparesis | 168
generalized tonic-clonic seizures | 174
GCS dropped to 5/15 (E1, V1, M3) | 174
immediate intubation | 174
continuous infusion of fentanyl | 174
continuous infusion of midazolam | 174
mechanical ventilation | 174
antiepileptic levetiracetam | 174
NCCT of the brain revealed near-complete evacuation of bilateral CSF hygroma | 174
development of "Mount Fuji" sign | 174
management included maintenance in flat position | 174
100% oxygen | 174
sedation | 174
brain-protective measures | 174
left frontoparietal decompressive craniectomy | 174
kept in ICU under sedation | 174
repeat NCCT of the brain showed near-complete resolution of pneumocephalus | 216
sedation stopped | 216
GCS 9/15 (E4, V1, M4) | 216
tracheotomy | 408
ventilator-associated pneumonia | 600
sepsis | 600
acute kidney injury | 600
multi-organ failure | 600
death | 600
no residual weakness |#
