64 years old | 0
male | 0
white | 0
admitted to the hospital | 0
HIV/AIDS | -13440
CD4 count <10 cells/mm3 | 0
antiretroviral therapy | -8760
Kaposi Sarcoma (KS) | -10080
radiation | -10080
pancytopenia | -10080
filgrastim | -10080
left orbital apex syndrome | -24
Aspergillus fumigatus sinusitis | -24
isavuconazonium sulfate | -24
discontinued isavuconazonium sulfate | 0
liposomal amphotericin-b | 0
voriconazole | 0
discontinued liposomal amphotericin-b | 24
voriconazole changed to posaconazole | 312
fever | 480
elevated lactate | 480
absolute neutrophil count greater than 1000 cells/mm3 | 480
blood cultures | 480
urinalysis | 480
chest x-ray | 480
increasing drainage from KS lesions | 480
broad empiric antibiotic therapy | 480
IV vancomycin | 480
IV cefepime | 480
encephalopathy | 528
rigors | 528
persistent fever | 528
hypotension | 528
tachypnea | 528
cefepime changed to piperacillin/tazobactam | 528
IV fluid bolus | 528
Wound Care Team consulted | 528
potential new infection of right thigh KS lesion | 528
increased sloughing and drainage | 528
musty odor | 528
blood culture positive for P. mendocina | 528
PICC line removed | 504
catheter tip culture | 504
repeat blood cultures | 504
antibiotic susceptibilities | 528
Etest | 528
ceftazidime | 528
levofloxacin | 528
meropenem | 528
piperacillin/tazobactam | 528
antibiotic therapy adjusted to ceftazidime | 528
total 10-day course | 912
source of infection unclear | 912
open wound | 912
blood cultures cleared | 912
infection successfully treated | 1056
discharged | 1056