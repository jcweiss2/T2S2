36+6 weeks gestation | 0  
    female | 0  
    birth weight of 3776 g | 0  
    hepatitis B carrier mother | 0  
    hepatitis B immunoglobulin received | 0  
    hepatitis B vaccine received | 0  
    grunting | 5  
    nasal flaring | 5  
    subcostal retractions | 5  
    borderline saturations in room air | 5  
    continuous positive airway pressure (CPAP) support | 5  
    respiratory distress worsened | 5  
    transferred to Neonatal Intensive Care Unit (NICU) | 5  
    intubated | 13  
    high frequency oscillatory ventilation | 13  
    nitric oxide | 13  
    hyaline membrane disease | 13  
    surfactant required | 13  
    umbilical venous catheter (UVC) inserted | 13  
    umbilical arterial catheter inserted | 13  
    malpositioning of UVC in right portal vein | 13  
    UVC readjusted | 13  
    septic work up | 24  
    intravenous penicillin | 24  
    intravenous gentamicin | 24  
    renal impairment (oliguria <1 ml/hour) | 24  
    gentamicin discontinued | 24  
    cefotaxime added | 24  
    full blood count unremarkable | 0  
    CRP 0.2 mg/L | 0  
    CRP 24 mg/L | 12  
    CRP 170 mg/L | 48  
    blood culture at birth grew SGp | 0  
    SGp sensitive to penicillin | 0  
    SGp sensitive to clindamycin | 0  
    ear swab cultures showed SGp | 0  
    ear swab cultures showed Escherichia coli | 0  
    Escherichia coli sensitive to ceftriaxone | 0  
    Escherichia coli sensitive to co-trimoxazole | 0  
    Escherichia coli sensitive to cefotaxime | 0  
    Escherichia coli resistant to ampicillin | 0  
    Escherichia coli resistant to gentamicin | 0  
    lumbar puncture deferred | 24  
    lumbar puncture performed | 96  
    CSF negative for meningitis | 96  
    CRP 48 mg/L | 96  
    fever 38.6°C | 120  
    Infectious Disease team involved | 120  
    conjugated hyperbilirubinemia | 120  
    renal function normalized | 120  
    CRP 165 mg/L | 120  
    blood culture repeated | 120  
    amikacin added | 120  
    blood culture sterile | 120  
    umbilical lines removed | 120  
    urine analysis unremarkable | 120  
    echocardiogram negative for structural heart disease | 120  
    echocardiogram negative for infective endocarditis | 120  
    liver abscess identified via ultrasound | 144  
    afebrile | 144  
    extubated | 144  
    penicillin stopped | 240  
    amikacin stopped | 240  
    cefotaxime continued | 240  
    liver abscess regression | 672  
    needle aspiration of liver abscess | 840  
    biopsy of liver abscess | 840  
    aspirate scanty | 840  
    biopsy obtained | 840  
    histopathology compatible with abscess | 840  
    Gram-stain negative | 840  
    acid-fast stain negative | 840  
    fungal stains negative | 840  
    bacterial cultures sterile | 840  
    fungal cultures sterile | 840  
    liver abscess further resolution | 888  
    parenteral antibiotics discontinued | 840  
    oral co-amoxiclav continued | 840  
    liver abscess significant resolution at 3 months | 2160  
    liver abscess 0.9x0.3x0.4 cm at 16 months | 11232  
    dystrophic calcification | 11232  
    growth assessment appropriate | 11232  
    neurodevelopmental assessment appropriate | 11232  
    Hepatitis B surface antibody 947 miu/L at 9 months | 6480  
    no maternal group B streptococcal colonization | 0  
    no prolonged rupture of membranes | 0  
    no maternal pyrexia | 0  
    maternal blood counts unremarkable | 0  
    maternal urine analysis unremarkable | 0  
    no meconium stained liquor | 0  
    no chest pain | 0  
    no shortness of breath | 0  
    no neurological symptoms | 0  
    no health care worker transmission | 0  
    no chorioamnionitis | 0  
    no CLABSI | 0  