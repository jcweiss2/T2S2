23 years old | 0
female | 0
AB+ blood group | 0
admitted to the hospital | 0
pseudotumor cerebri | -672
treated by acetazolamide | -672
C-section delivery | -72
diffuse abdominal rebound tenderness | -72
guarding | -72
laparotomy | -72
small bowel gangrene | -72
resected bowel segments | -72
stoma creation | -72
septic shock | -48
gangrene of the stoma | -48
resected remnant of the small intestine | -48
gastrodouodenostomy tube insertion | -48
transferred to the intestinal rehabilitation unit | -48
parenteral nutrition | -48
listed on the waiting list for small intestinal transplantation | -48
blood group AB+ | -48
negative flow panel reactive assay | -48
anti-human leukocyte antigen antibodies | -48
positive bacterial culture from central venous catheters | -336
pulmonary thromboembolism | -336
donor found | -192
donor's blood group O+ | -192
small intestine transplantation | 0
methylprednisolone | 0
thymoglobulin | 0
rituximab | 0
weaned from the ventilator | 6
tacrolimus | 0
mycophenolate mofetil | 0
prednisolone | 0
small bowel biopsy | 120
no rejection | 120
oral nutrition started | 120
hemoglobin level dropped | 240
hypotension | 240
tachycardia | 240
AB+ RBC transfusion | 240
hemoglobin level dropped again | 264
AB+ RBC transfusion | 264
acute jaundice | 288
total bilirubin level increased | 288
exploratory laparotomy | 288
small intestinal hernia | 288
hernia reduction | 288
Lactate dehydrogenase increased | 288
reticulocyte count increased | 288
haptoglobin level decreased | 288
indirect bilirubinemia | 288
positive Direct antiglobulin test | 336
O+ RBC transfusion | 336
intravenous immunoglobulin transfusion | 432
plasmapheresis | 432
hemolysis decreased | 432
discharged | 1032
cytomegalovirus infection | 1032
acute rejection | 1032
treated | 1032
admitted again | 1104
neck soft tissue abscess | 1104
died of sepsis | 1104