16 years old | 0
    male | 0
    admitted to the hospital | 0
    sore throat | -24
    fatigue | -24
    myalgias | -24
    fever | -24
    left forearm soreness | -24
    temperature of 39.1°C | -24
    heart rate of 143 beats per min | -24
    dry mucus membranes | -24
    mild cervical lymphadenopathy | -24
    mild erythema of the posterior pharyngeal wall | -24
    tachycardia | -24
    mild tenderness on left forearm | -24
    elevated creatinine level | -24
    blood cultures obtained | -24
    vancomycin | -24
    ceftriaxone | -24
    admitted for possible sepsis | -24
    forearm soreness evolved into swollen, tender, erythematous area | 24
    recalled sleeping in a basement where spiders were noted | 24
    developed worsening hypotension | 24
    blood pressure decreased from 109/53 to 82/39 mmHg over 12 hours | 24
    persistent tachycardia | 24
    unresponsive to fluid challenge | 24
    transfer to pediatric ICU | 24
    management of decompensated shock | 24
    ionotropic support initiated | 24
    intra-arterial access obtained | 24
    transaminitis | 48
    increased bilirubin | 48
    increased C-reactive protein | 48
    leukocytosis | 48
    coagulation profile consistent with DIC | 48
    differential diagnosis of septic shock vs loxoscelism | 48
    medical toxicology consultation | 72
    left arm became increasingly tender | 72
    developing vesicular areas | 72
    darkening, necrotic-appearing base | 72
    skin swab submitted for ELISA | 72
    ELISA positive for Loxosceles venom | 72
    became dyspneic | 72
    chest X-ray revealed mild pulmonary edema | 72
    echocardiogram showed ejection fraction of 55% | 72
    hemoglobin dropped from 12.6 to 7.9 gm/dL | 144
    increase in LDH | 144
    increase in bilirubin | 144
    increase in plasma free hemoglobin | 144
    intravascular hemolysis | 144
    transfused with packed red blood cells | 144
    methylprednisolone initiated | 144
    developed tachycardia with diffuse T-wave changes | 144
    EKG concerning for myocarditis | 144
    B-type natriuretic peptide elevated to 1309 pg/mL | 144
    troponin-I elevated to 0.29 ng/mL | 144
    creatine kinase-muscle/brain elevated to 7.6 ng/mL | 144
    cardiac MRI demonstrated myocarditis | 144
    ejection fraction of 45% | 144
    myocarditis therapy initiated with IV immunoglobulins | 144
    bumetanide administered | 144
    favorable clinical response to therapy | 144
    decreasing troponin-I | 168
    decreasing B-type natriuretic peptide | 168
    normalization of EKG | 168
    improved cardiac function on repeat echocardiogram | 168
    hemoglobin reached nadir of 5.9 gm/dL | 168
    transfusions on days 7 and 8 | 168
    plasmapheresis performed on days 8, 9, 10, and 13 | 168
    hematological laboratory results normalized | 312
    laboratory values continued improving | 312
    discharged home on day 20 | 480
    wound responded to standard outpatient wound care | 480
    follow-up outpatient echocardiogram was normal | 480
    