49 years old | 0
female | 0
admitted to the hospital | 0
nausea | -48
vomiting | -48
fever | -48
diarrhea | -48
oliguria | -24
apathy | -24
type 2 diabetes mellitus | -6720
poor appetite | -48
poor sleep | -48
weight loss | -48
coma | 0
involuntary movements | 0
temperature 37.8 °C | 0
heart rate 130 beats/min | 0
respiration 28 breaths/min | 0
blood pressure 70/50 mmHg | 0
bowel sounds 6 beats/min | 0
urine output less than 0.5 mL/kg/min | 0
white blood cells 9.4 × 10^9/L | 0
neutral granulocytes 94.5% | 0
platelet count 5.2 × 10^10/L | 0
procalcitonin 0.4 ng/mL | 0
T-cell subpopulation analysis | 0
liver damage | 0
aspartate aminotransferase 923 U/L | 0
alanine aminotransferase 410 U/L | 0
total bilirubin 27.6 µmol/L | 0
serum creatinine 380 µmol/L | 0
metabolic acidosis | 0
respiratory alkalosis | 0
blood gas pH 7.46 | 0
partial pressure of carbon dioxide 25 mmHg | 0
bicarbonate level 17.8 mmol/L | 0
base excess -5.0 mmol/L | 0
lactate level 1.2 mmol/L | 0
liver ultrasound multiple mixed-density shadows | 0
NMLA | 0
sepsis | 0
septic encephalopathy | 0
septic shock | 0
SA-AKI | 0
secondary immune deficiency | 0
APACHE II score 18 | 0
SOFA score 11 | 0
cefoperazone-sulbactam | 1
fluid resuscitation | 3
noradrenaline | 3
imipenem | 3
linezolid | 3
glutathione injection | 3
computed tomography of the liver | 48
CRRT combined with HP proposed | 72
CRRT combined with HP refused | 72
CRRT combined with HP performed | 72
CRRT mode continuous venovenous hemofiltration | 72
blood flow rate 120 mL/h | 72
HA380 membrane filter | 72
CRRT and HP treatment terminated | 168
WBC decreased | 120
PCT decreased | 120
IL-6 decreased | 120
lactate decreased | 120
renal function improved | 120
SCr levels decreased | 120
immune function improved | 120
CD8+ T-cells increased | 120
APACHE II score decreased | 120
SOFA score decreased | 120
discharged | 504
recovered | 672