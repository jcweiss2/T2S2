62 years old | 0
female | 0
admitted to the hospital | 0
shortness of breath | -168
hemoptysis | -168
intermittent yellow sclera | -720
heavy alcohol consumption | -720
tachypneic | 0
tachycardiac | 0
respiratory distress | 0
nonrebreather mask | 0
broad-spectrum antibiotic therapy | 0
transferred to PCU | 0
bilevel positive airway pressure | 0
scleral icterus | 0
dried blood on lips and chin | 0
diffuse crackles over bilateral lower lung fields | 0
bilateral lower extremity pitting edema | 0
elevated white blood cell count | 0
low hemoglobin | 0
low platelet count | 0
low albumin | 0
elevated alkaline phosphatase | 0
elevated AST | 0
elevated ALT | 0
elevated bilirubin | 0
elevated lactate | 0
elevated BNP | 0
elevated high-sensitivity troponin | 0
elevated D-Dimer | 0
elevated INR | 0
prolonged PT | 0
bilateral multifocal patchy opacities on chest x-ray | 0
extensive patchy parenchymal airspace opacities on CT chest | 0
diffusely heterogeneous enhancement and nodularity throughout the liver parenchyma on CT abdomen | 0
severe respiratory acidosis | 24
intubation | 24
IV steroids | 24
bronchoalveolar lavage | 24
erythematous airways | 24
bloody return on lavage | 24
benign respiratory epithelium with reactive changes on cytology | 24
acute inflammation on cytology | 24
macrophages on cytology | 24
red blood cells on cytology | 24
negative acid-fast stain | 24
negative cultures | 24
negative Pneumocystis jiroveci smear | 24
negative autoimmune disease workup | 48
negative infectious disease workup | 48
positive human metapneumovirus by PCR | 48
vasopressors | 96
prone position | 192
hemodialysis | 216
severe acute kidney injury | 216
acidosis | 216
disseminated intravascular coagulation | 264
scattered small bilateral subarachnoid hemorrhages on CT head | 264
cardiac arrest | 264
death | 264