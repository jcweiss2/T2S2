63 years old | 0
male | 0
admitted to the hospital | 0
generalized weakness | -168
ESRD | -6720
haemodialysis | -6720
systolic heart failure | -6720
coronary artery disease | -6720
hypertension | -6720
type II diabetes | -6720
WBC 3.1 cells*109L | 0
tachycardia 96 bpm | 0
fever 39.5°C | 0
blood pressure 160/90 mmHg | 0
respiratory rate 18 | 0
oxygen saturation 96% | 0
haemoglobin 86 g/L | 0
platelets 112 cells*109L | 0
haematocrit 0.26 fraction | 0
INR 1.5 | 0
APTT 36.3 s | 0
AST 59 | 0
ALT 33 | 0
total bilirubin 10.26 μmol/L | 0
splenomegaly | 0
vancomycin | 0
cefepime | 0
metronidazole | 0
serology for hepatitis negative | 0
serology for human immunodeficiency virus negative | 0
serology for cytomegalovirus negative | 0
serology for heparin-induced-thrombocytopenia antibody negative | 0
serology for herpes simplex virus negative | 0
serology for heterophile antibody test negative | 0
serology for parvovirus B19 negative | 0
serology for legionella negative | 0
serology for mycoplasma negative | 0
coagulopathy | 24
peak INR level 2.7 | 24
peak APTT 48 s | 24
transaminitis | 24
AST 1034 Units/L | 24
ALT 217 Units/L | 24
total bilirubin 22.23 μmol/L | 24
TB-QuantiFERON indeterminate | 0
autoimmune workup negative | 0
EBV DNA polymerase chain reaction positive | 0
ferritin > 33.7 nmol/L | 0
soluble CD25 14 158 units/ml | 0
triglycerides > 2.89 mmol/L | 0
fever > 38.5°C | 0
elevated CD25 | 0
high ferritin | 0
elevated TG | 0
cytopenia | 0
dexamethasone | 168
etoposide | 168
bone marrow biopsy | 168
epithelial granulomas | 168
histiocytes containing phagocytized nucleated cells | 168
histiocytes with phagocytized erythrocytes | 168
acid-fast bacilli negative | 168
RIPE therapy | 336
miliary pattern TB | 336
chest CT | 336
pulmonary nodules | 336
anti-tuberculosis treatment | 336
WBC counts decline | 504
cell counts increase | 504
patient expired | 504
mycobacterium TB complex growth | 504