21 years old | 0
female | 0
admitted to the hospital | 0
state of shock | 0
respiratory distress | 0
vague abdominal discomfort | 0
abdominal distension | 0
fever | -336
cough | -336
breathing difficulty | -336
loose stools | -336
abdominal sepsis | 0
peritonism | 0
normal bowel sounds | 0
intubated | 0
mechanical ventilation | 0
ionotropic support | 0
coronavirus disease intensive care unit | 0
negative IgM/IgG rapid test | 0
COVID-19 real-time polymerase chain reaction test | 0
positive COVID-19 real-time polymerase chain reaction test | 0
haemoglobin: 7.2 g/dl | 0
total leucocyte count: 16 × 109/L | 0
platelet count: 99 × 109/L | 0
ultrasound abdomen | 0
large well defined thick-walled collection | 0
percutaneous pigtail drainage | 0
purulent output | 0
chest X-ray | 0
bilateral lower lobe atelectasis | 0
prominent bronchovascular markings | 0
contrast-enhanced computed tomography scan of thorax | 0
bilateral basal atelectasis | 0
ground-glass opacities | 0
CO-RADS score of 4 | 0
contrast enhanced computed tomography of the abdomen | 0
sealed off perforation | 0
localised large pelvic collection | 0
exploratory laparotomy | 24
faecopurulent peritoneal collection | 24
dense interbowel adhesions | 24
greater omentum smeared to the clumped bowel loops | 24
adhesiolysis | 24
five perforations in the distal ileum | 24
jejunal perforation | 24
primary repair | 24
loop ileostomy | 24
nasojejunal tube | 24
repeat second COVID-19 real time sample test | 120
negative COVID-19 real time sample test | 120
stomal viability | 120
pinprick test | 120
fresh blood | 120
lubricated transparent tube | 120
pink mucosa | 120
nasojejunal tube feeding | 48
histopathological examination | 120
granulomatous inflammation | 120
acid-fast bacilli | 120
Ziehl-Neelsen staining | 120
GenXpert-Mtb/Rif | 120
Mycobacterium tuberculosis | 120
anti-tubercular regime | 120
low output enterocutaneous fistula | 168
conservative management | 168
sepsis subsided | 336
oral feeds | 336
nasojejunal tube removed | 336
discharged | 720