92 years old | 0
female | 0
admitted to the hospital | 0
fever | -48
myalgia | -48
anorexia | -48
general weakness | -48
hypertension | -672
insect bite | -48
leukopenia | 0
thrombocytopenia | 0
elevated liver enzymes | 0
aspartate aminotransferase | 0
alanine aminotransferase | 0
ceftriaxone | 0
SFTSV detected | 0
SFTSV viral load | 0
conservatively treated | 0
stable | 0
sudden-onset pneumonia | 96
respiratory failure | 96
chest X-ray | 96
high-resolution computed tomography | 96
bronchiolitis | 96
bronchial wall thickening | 96
cefepime | 96
vancomycin | 96
voriconazole | 96
Aspergillus galactomannan antigen | 96
mechanical ventilation | 120
intensive care unit | 120
septic shock | 120
multifocal consolidations | 120
intravenous immunoglobulin | 144
died | 264
respiratory failure | 264
refractory hypotension | 264
metabolic acidosis | 264