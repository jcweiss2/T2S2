35 years old | 0
male | 0
admitted to cardiology unit | 0
unremitting fever | -360
chest pain | -360
abdominal pain | -360
palpitation | -360
stable vitals | 0
critical general conditions | 0
unspecific ECG abnormalities | 0
endocarditis | 0
aortic valve leaflets involved | 0
mitral valve leaflets involved | 0
optimal medical therapy initiated | 0
high risk for cardiac surgery | 0
multiorgan failure | 0
pulmonic failure | 0
kidney failure | 0
metabolic failure | 0
septic condition | 0
daily echocardiographic examination | 0
cardiorespiratory arrest | 120
high-quality chest compressions | 120
advanced cardiac life support | 120
ROSC | 136
echocardiographic check | 136
right atrial thrombus formation | 136
endovenous heparin administration | 136
continued chest compressions | 136
thrombus disappearance | 140
moved to intensive care department | 140
poor prognosis | 140 
cardiac thrombus formation | 136 
mechanical circulatory support | -120 
left ventricular thrombus formation | -120 
ventricular fibrillation | -120 
blood clots dissolution | -120 
blood clots dissemination | -120 
optimized chest compressions | 0
prompt defibrillation | 0
effective feedback of chest compressions | 0
chest conformation | 0
underlying cardiac disease | 0
rescuer approach | 0
Virchow's triad | 0
forward blood flow ceasing | 120
thrombolytic agents | 0
heparin therapy | 136
primary right heart thrombus | -120
serial echocardiographic examinations | 0
blood sludge | 136
septic syndrome | 0
hypercoagulability | 0
infectious agents | 0
coagulation cascade activation | 0
platelet aggregation | 0
pro-thrombotic responses | 0
acidosis | 0
tissue hypoperfusion | 0
liver transplantation | -120
heparin treatment | -120
intravenous heparin | 136
prothrombotic conditions | 0
spontaneous echo contrast | 136
cardiac POCUS | 0
ultrasound-implemented CPR algorithm | 0
time loss | 0
fast-track examinations | 0
ROSC prediction | 0
unshockable rhythm | 0
fast cardiac ultrasound protocol | 0
skilled operators | 0
rhythm check | 0
four-chamber apical view | 0
subcostal view | 0
ventricular function assessment | 0
potential complications assessment | 0
cardiac ultrasound | 0
routine use during CPR | 0
early causative screening | 0
cardiac function information | 0
potential complications information | 0 
patient consent | 0 
financial support | 0 
conflicts of interest | 0