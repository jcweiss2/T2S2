25 years old | 0
male | 0
admitted to the hospital | 0
high-grade fever | -144
diffuse abdominal pain | -48
hematemesis | -48
anemia | 0
thrombocytopenia | 0
hyperbilirubinemia | 0
raised transaminases | 0
normal coagulation profile | 0
normal renal function | 0
dengue NS1 antigen positive | 0
malaria antigen negative | 0
malaria smear negative | 0
dense bilateral lower lobe consolidation | 0
acute respiratory distress syndrome (ARDS) | 48
intubation | 48
mechanical ventilation | 48
septic shock | 48
broad-spectrum antimicrobials started | 48
meropenem started | 48
doxycycline started | 48
referred to Intensive Care Unit (ICU) | 48
fever | 48
heart rate 130/min | 48
blood pressure 130/70 mmHg | 48
norepinephrine infusion | 48
sedated with midazolam | 48
sedated with fentanyl | 48
mechanical ventilation | 48
APACHE II 20 | 48
SOFA 12 | 48
improving thrombocytopenia | 48
improving liver function tests | 48
positive dengue IgM | 48
positive scrub typhus serology | 48
elevated procalcitonin | 48
proned | 60
oxygenation status improved | 72
persistent high-grade fever | 72
B. cepacia bacteremia | 0
resistant to amikacin | 0
resistant to aztreonam | 0
resistant to ceftazidime | 0
resistant to cefoperazone–sulbactam | 0
sensitive to levofloxacin | 0
sensitive to meropenem | 0
sensitive to trimethoprim–sulfamethoxazole | 0
methicillin-resistant Staphylococcus aureus | 48
sensitive to linezolid | 48
sensitive to vancomycin | 48
antimicrobials changed | 96
doripenem started | 96
linezolid started | 96
cotrimoxazole started | 96
fever reduced | 120
successful extubation | 144
sterile blood cultures | 168
decreased procalcitonin | 168
cavitatory lesions | 336
bronchiectatic changes | 336
discharged | 504