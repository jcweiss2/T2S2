31 years old | 0
    male | 0
    admitted to the hospital | 0
    presented to the ED | 0
    open sores covering his body | 0
    cigarette burn to left forearm | -336
    sores began at the site of a cigarette burn | -336
    sores spread diffusely over the body | -336
    lesions slightly tender to the touch | 0
    review of systems negative for viral prodrome | 0
    denied fevers | 0
    denied chills | 0
    denied sweats | 0
    denied chest pain | 0
    denied shortness of breath | 0
    denied abdominal pain | 0
    denied nausea | 0
    denied vomiting | 0
    no history of ill contacts | 0
    no animal exposure | 0
    no insect bites | 0
    no recent travel | 0
    denied intravenous drug use | 0
    chronic use of tobacco | 0
    chronic use of alcohol | 0
    chronic use of marijuana | 0
    not taking any medications | 0
    denied known allergies | 0
    denied significant family history | 0
    sought no medical care prior to ED presentation | 0
    arrival to ED via ambulance | 0
    anxious | 0
    avoided unnecessary movement | 0
    temperature 100.1°F | 0
    heart rate 145 bpm | 0
    blood pressure 124/77 mmHg | 0
    respiratory rate 20 breaths per minute | 0
    oxygen saturation 99% on room air | 0
    heart tones regularly tachycardic | 0
    free of murmurs | 0
    free of rubs | 0
    pulmonary exam clear bilaterally | 0
    no crackles | 0
    no wheezes | 0
    no edema of extremities | 0
    no lymphadenopathy | 0
    no hepatosplenomegaly | 0
    skin exam revealed diffuse regions of skin sloughing | 0
    necrosis | 0
    mildly erythematous base along the dermis | 0
    occasional small bullae | 0
    occasional vesicles | 0
    over 50% BSA involved | 0
    back involved | 0
    abdomen involved | 0
    scrotum involved | 0
    perirectal area involved | 0
    forehead spared | 0
    scalp spared | 0
    no purulent discharge | 0
    no pustules | 0
    no purpura | 0
    no ulcerations | 0
    strong foul-smelling odor | 0
    non-affected skin sloughed with lateral traction | 0
    oral mucosa injected | 0
    sloughing apparent | 0
    conjunctivae spared | 0
    temperature increased to 101.7°F | 24
    vancomycin administered | 24
    meropenem administered | 24
    blood cultures sent | 24
    received four liters IV normal saline | 24
    morphine administered | 24
    white blood cell count 12,000/mm | 24
    lactic acid 2.8 mmol/L | 24
    serum bicarbonate 21 mmol/L | 24
    serum glucose 140 mg/dL | 24
    blood urea nitrogen 9 mg/dL | 24
    creatinine 0.9 mg/dL | 24
    anion gap 10 mmol/L | 24
    remained stable | 24
    persistently tachycardic | 24
    admitted to ICU | 24
    developed severe sepsis | 48
    blood cultures positive for oxacillin-sensitive Staphylococcal aureus | 72
    started on steroids | 72
    received IVIG | 72
    cared for in Burn Care Unit | 72
    underwent multiple surgical debridement procedures | 72
    skin biopsy revealed non-specific epidermal necrosis | 72
    discharged home | 168
    over-the-counter NSAID use prior to onset of symptoms | -336
    septicemia | 72
    malodor noted | 0
    biopsy consistent with TEN | 72
    secondary bacterial infection | 72
    TEN diagnosis | 0
    