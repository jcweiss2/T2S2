40 years old | 0
male | 0
HIV-1 infection | -720
high fever | -24
severe malaise | -24
headache | -24
generalized skin rash | -24
sinusitis | -672
symptomatic treatment | -672
fever | 0
shock status | 0
systolic blood pressure 84 mmHg | 0
pulse rate 110 beats/min | 0
mildly altered consciousness | 0
neck stiffness | 0
diminished skin turgor | 0
no focal neurological deficits | 0
no visual disturbances | 0
leukocytosis 11600/µL | 0
elevated C-reactive protein 12.1 mg/L | 0
hyperproteinemia 9.6 g/dL | 0
acute renal dysfunction | 0
creatinine 1.54 mg/dL |
