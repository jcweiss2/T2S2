55 years old | 0
male | 0
admitted to the hospital | 0
ureteral double J stent removal | 0
end-stage renal disease | -8760
compensated chronic renal failure | -8760
ureteroscopic intervention | -720
left ureteric calculus | -720
blood glucose 110 mg/dL | 0
urea 259 mg/dL | 0
creatinin 8.8 mg/dL | 0
uric acid 7.4 mg/dL | 0
sodium 138 mmol/L | 0
potassium 4.93 mmol/L | 0
hemoglobin 7.7 gr/dL | 0
hematocrit 24 (%) | 0
white blood cell count 6000/uL | 0
platelet count 250000/uL | 0
prothrombin time normal | 0
activated partial thromboplastin time normal | 0
bilateral reduced kidney sizes | 0
increased parenchymal echogenicity | 0
creatinin clearance 7.9 mL/min | 0
protein level 2364 mg/day | 0
included in routine hemodialysis program | 0
ureteric catheter removal | 24
abdominal pain | 48
abdominal distension | 48
widespread tenderness | 48
rebound positivity | 48
defense positivity | 48
body temperature 36.5°C | 48
pulse rate 105/min | 48
respiratory rate 20/min | 48
blood pressure 85/50 mm Hg | 48
urea 119 mg/dL | 48
creatinin 4.2 mg/dL | 48
sodium 140 mmol/L | 48
potassium 4.16 mmol/L | 48
hemoglobin 6.7 gr/dL | 48
hematocrit 19.9 (%) | 48
white blood cell count 8000/uL | 48
platelet count 57000/uL | 48
prothrombin time 21.7 s | 48
activated partial thromboplastin time 110 s | 48
INR 1.91 | 48
abdominal tomography | 48
high-density lesion | 48
hematoma | 48
retroperitoneal region | 48
left upper renal pole | 48
subdiaphragmatic area | 48
emergency exploratory operation | 72
free fluid | 72
hemorrhagic character | 72
capsular laceration sites | 72
hematomas | 72
splenectomy | 72
fresh whole blood transfusion | 72
fresh frozen plasma transfusion | 72
thrombocyte suspension transfusion | 72
persistent thrombocytopenia | 96
high INR level | 96
uremic coagulopathy | 96
platelet replacement | 96
fresh frozen plasma replacement | 96
stabilization of blood parameters | 120
pneumococcal vaccine | 120
Haemophilus influenza type B vaccine | 120
meningococcal vaccine | 120
respiratory distress | 240
high fever | 240
pulmonary computed tomography angiography | 240
no thromboembolism | 240
sputum culture positivity | 240
blood culture positivity | 240
Acinetobacter | 240
intravenous colimycin therapy | 240
intensive care unit | 240
progressive deterioration | 240
sepsis | 600
multiorgan failure | 600
death | 600