44 years old | 0
    male | 0
    admitted to Wonkwang University Hospital | 0
    fever | -240
    non-productive cough | -240
    myalgias | -240
    hypertension | -43800
    treated with angiotensin-converting enzyme inhibitor | -43800
    treated with oral quinolone | -216
    resting dyspnea | -48
    productive cough | -48
    fever (before admission) | -48
    admitted to intensive care unit | 96
    mechanically ventilated | 96
    chest CT performed | 120
    fiberoptic bronchoscopy performed | 120
    chest CT scan revealed bilateral peribronchial infiltrates | 120
    bronchoscopy revealed whitish exudative membranes | 120
    endobronchial biopsy specimens revealed Aspergillus species | 120
    bronchial washing fluid revealed Aspergillus species | 120
    high fever persisted | 144
    refractory septic shock | 144
    hypoxemia (persistent) | 144
    IV amphotericin B administered | 144
    supportive care administered | 144
    refractory hypoxemia | 168
    oliguria | 168
    fatal cardiac arrest | 168
    no history of previous respiratory diseases | 0
    no specific family history | 0
    temperature of 38.6℃ | 0
    blood pressure 120/80 mmHg | 0
    heart rate 90 b.p.m | 0
    respiratory rate 30 breaths/min | 0
    bilateral inspiratory coarse crackles | 0
    end-expiratory wheezing | 0
    arterial blood gas: pH 7.343 | 0
    arterial blood gas: PaCO2 41.2 mmHg | 0
    arterial blood gas: PaO2 59.2 mmHg | 0
    arterial blood gas: SaO2 90.7% | 0
    WBC 19,580/mm3 | 0
    neutrophils 82.5% | 0
    ESR 71 mm/h | 0
    C-reactive protein 184.6 mg/L | 0
    hemoglobin A1c 5.8% | 0
    blood urea nitrogen 32.4 mg/dL | 0
    creatinine 1.32 mg/dL | 0
    random glucose 117 mg/dL | 0
    chest X-ray bilateral bronchial wall thickening | 0
    initial sputum stains negative | 0
    sputum cultures negative | 0
    blood cultures negative | 0
    HIV test negative | 0
    empirical therapy with cefoperazone/sulbactam | 0
    empirical therapy with vancomycin | 0
    rapidly deteriorated | 96
    increasing dyspnea | 96
    hypoxemia (initial) | 96
    respiratory failure | 96
    severe CO2 retention | 96
    chest X-ray lesions | 96
    rapidly increasing respiratory acidosis | 120
    hypoxemia (CT time) | 120
    pseudomembranous necrotizing tracheobronchial aspergillosis | 120
    no parenchymal invasion | 120
    no consolidation of the parenchyma | 120
    no post-mortem examination | 168
    refusal of post-mortem examination | 168
    30-pack-a-year ex-smoker | 0
    no invasion of pulmonary parenchyma | 120
    no radiographic abnormalities | 0
    no response to broad-spectrum antibiotics | 96
    no risk factors for immunocompromised state | 0
    no corticosteroid use | 0
    no chronic airway limitation | 0
    no underlying disease | 0
    no T cell dysfunction | 0
    no lymphopenia | 0
    no cutaneous anergy | 0
    no influenza A infection | 0
    no malignancy | 0
    no AIDS | 0
    no bone-marrow transplantation | 0
    no diabetes mellitus | 0
    no chronic liver disease | 0
    no alcoholism | 0
    no diabetic ketoacidosis | 0
    no fungal invasion through bronchial wall | 120
    no pulmonary artery invasion | 120
    no atelectasis | 120
    no parenchymal lung involvement | 120
    no consolidation | 120
    no luminal narrowing | 120
    no patchy atelectasis | 120
    no tracheal narrowing | 120
    no pneumomediastinum | 120
    no parenchymal infiltration on chest X-ray | 0
    no specific radiographic findings | 0
    no response to antibiotics | 96
    no risk factors for immunodeficiency | 0
    no prior respiratory diseases | 0
    no family history of respiratory diseases | 0
    no HIV infection | 0
    no neutropenia | 0
    no exposure to corticosteroids | 0
    no cytotoxic drugs | 0
    no malignancy history | 0
    no bone-marrow transplant history | 0
    no chronic obstructive pulmonary disease | 0
    no asthma | 0
    no fungal invasion into adjacent lung tissue | 120
    no pulmonary parenchyma invasion | 120
    no open-lung biopsy performed | 0
    no microbiological evidence of Aspergillus before bronchoscopy | 0
    no prior antifungal therapy | 0
    no life-saving treatment response | 168
    no alteration of disease course | 168
    no survival | 168