79 years old | 0
woman | 0
surgery on medial collateral ligament of right knee | -175200
TKA for right knee osteoarthritis | -17520
fell from 50 cm height | -72
overstretched right knee at landing | -72
right knee pain | -72
transported to nearby hospital | -72
diagnosed with periprosthetic tibial fracture after TKA | -72
admitted to the hospital | -72
right dorsalis pedis artery not palpable | -72
suspicion of popliteal artery injury | -72
transferred to emergency and critical care center | -72
popliteal artery injury diagnosed by CTA | 0
emergency surgery for revascularization performed | 0
popliteal artery semicircular partial rupture | 0
bifurcation of anterior and posterior tibial arteries injured | 0
anastomosis between popliteal and posterior tibial arteries | 0
popliteal vein damage observed | 0
injured area excised | 0
end-to-end anastomosis performed | 0
external fixation across knee | 0
fracture stabilized | 0
internal fixation on 11th day after injury | 264
Felix classification IIB diagnosis | 264
anatomical locking plates placed | 264
screws inserted forwards and backwards of tibial implant keel | 264
antibiotic treatment started on 5th day after internal fixation | 360
surgical-site sepsis | 360
debridement performed 7 days after internal fixation | 408
exposed plate covered with gastrocnemius muscle flap after 21 days | 504
infection resolved after 50 days | 1200
partial weight-bearing started 3 months after surgery | 2160
bone union confirmed 5 months after surgery | 3600
