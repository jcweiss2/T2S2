48 years old | 0
male | 0
Caucasian | 0
admitted to the hospital | 0
chest pain | -72
dyspnoea | -72
bilateral sensorineural hypacusis | -2880
hearing aids | -2880
cardiac examination | 0
heart rhythm regular | 0
blood pressure similar in both arms | 0
electrocardiogram | 0
short PR interval | 0
narrow QRS complex | 0
inversion of T-waves | 0
non-significant depression of ST segments | 0
elevated high sensitive troponin t | 0
elevated N-terminal proBNP | 0
normal creatinine kinase level | 0
prediabetic metabolic state | 0
slightly elevated ferritin | 0
coronary angiography | 0
excluded coronary artery disease | 0
echocardiography | 0
symmetric non-obstructive HCM | 0
diffuse reduced left ventricular ejection fraction | 0
symmetric increase in myocardial wall thickness | 0
LV wall thickness could not be explained by physical training or valve disease | 0
arterial hypertension excluded | 0
LV intracavitary gradient below 30 mmHg | 0
elevation of LV filling pressure | 0
left ventricular mass index increased | 0
cardiac amyloidosis unlikely | 0
diameter and function of the right ventricle normal | 0
cardiac MRI | 0
mildly reduced LV function | 0
MRI parameters of RV size and function regular | 0
myocardial fibrosis detected by late gadolinium enhancement | 0
endomyocardial biopsy | 0
hypertrophy of cardiomyocytes and diffuse fibrosis | 0
no signs of infiltrative or active inflammatory disease | 0
normal plasma activity of α-D-galactosidase-A | 0
excluded Fabry disease | 0
next-generation sequencing | 0
m.3243A > G mutation | 0
pathogenic variant of mitochondrial DNA | 0
Holter monitoring | 0
no ventricular tachycardia | 0
implantable cardioverter defibrillator therapy not recommended | 0
heart failure medications intended to improve symptoms | 0
follow-up scheduled in 3 months | 0
family history of cardiomyopathy | -10080
mother died of heart failure | -10080
father died of ischemic cardiomyopathy | -10080
half-brother died suddenly | -10080
half-brother diagnosed with HCM | -10080
sister diagnosed with DCM | -10080
m.3243A > G mutation identified in family members | 0
clinical and genetic screening of family members | 0
hearing loss in family members | -10080
diabetes in family members | -10080
kidney disease in family members | -10080
short PQ syndrome in family members | -10080
cardiomyopathy in family members | -10080
MIDD diagnosed in family members | 0
maternally inherited diabetes and deafness | 0
cardiac MRI in 2015 | -1080
cardiac MRI in 2018 | 0
progression of myocardial fibrosis and scarring | 0
LGE in mid-wall pattern | 0
predictor of adverse cardiovascular outcomes | 0
repeated cardiac MRIs recommended | 0
ICD placement not indicated | 0
recommendation for ICD therapy reassessed | 0
intra-familial phenotypic cardiomyopathy variability | 0
heterogeneous spectrum of cardiomyopathies | 0
cardiac hypertrophy more prevalent than dilation | 0
further studies needed | 0