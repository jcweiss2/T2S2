12 years old | 0
female | 0
Thai | 0
admitted to the hospital | 0
behavioural change | -144
fever | -144
headache | -144
bizarre behaviour | -144
conversation with herself | -144
cried or laughed without explaining the reason | -144
alteration of consciousness | -144
abnormal movements of hands | -144
could not write letters | -144
aggressive behaviour | -96
incomprehensive language | -96
intermittent screaming | -96
visual hallucination | -96
received roxithromycin | -144
received fexofenadine | -144
received paracetamol | -144
high-grade fever | -48
intermittent episodes of screaming | -48
aggressive behaviours | -48
computed tomography scan brain | -48
lumbar puncture | -48
received high-dose ceftriaxone | -48
received acyclovir | -48
received azithromycin | -48
received oseltamivir | -48
confusion | 0
disorientation to time | 0
disorientation to place | 0
disorientation to person | 0
low-grade fever | 0
body temperature 38.4°C | 0
pulse rate 110 beats per minute | 0
respiratory rate 24 breaths per minute | 0
Glasgow coma scale E4M5V3 | 0
oromotor dyskinesia | 0
choreoathetosis | 0
reflex 3+ | 0
Babinski's sign equivocal | 0
clonus absent | 0
hemoglobin 123 g/L | 0
white blood cell count 4.83 × 10^9/L | 0
platelet count 310 × 10^9/L | 0
sodium 140 mmol/L | 0
potassium 3.8 mmol/L | 0
chloride 104 mmol/L | 0
bicarbonate 21.4 mmol/L | 0
calcium 2.32 mmol/L | 0
phosphorus 1.12 mmol/L | 0
magnesium 0.97 mmol/L | 0
glucose 5.1 mmol/L | 0
TSH 3.35 µU/mL | 0
FT4 18 ng/L | 0
anti-thyroglobulin < 10 | 0
anti-thyroid peroxidase < 9 IU/mL | 0
C3 1.25 | 0
C4 3.8 g/L | 0
cerebrospinal fluid analysis | 0
colourless fluid | 0
WBC 13 cells/mm^3 | 0
protein 20.1 g/L | 0
glucose 4.2 mmol/L | 0
Gram staining negative | 0
culture from CSF negative | 0
infectious work-ups negative | 0
NMDAR autoantibodies positive | 0
electroencephalogram monitoring | 0
absent sleep-wake pattern | 0
generalized slow waves 1-3 Hertz | 0
delta brush pattern | 0
ictal EEG | 0
generalized rhythmic delta waves | 0
computed tomography scan brain | 0
small hypodense lesions in the left lentiform nucleus | 0
received pulse methylprednisolone | 0
received intravenous immunoglobulin | 0
received plasmapheresis | 0
received phenytoin | 0
received risperidone | 0
developed superrefractory status epilepticus | 336
sent to the paediatric intensive care unit | 336
abdominal bloating | 1008
feeding intolerance | 1008
drooling | 1008
bilious vomiting | 1008
watery diarrhoea | 1008
coffee-ground content | 1008
bilious content | 1008
body temperature 37.8°C | 1008
distended and soft abdomen | 1008
hypoactive bowel sounds | 1008
nasogastric tube inserted | 1008
intravenous fluid infusion | 1008
omeprazole intravenously | 1008
nasogastric fluid content bilious | 1056
drooling | 1056
saliva content | 1056
large volume of stool | 1056
greenish watery stool | 1056
minimally mucous stool | 1056
old blood in stool | 1056
haemoculture from the central line negative | 1056
haemoculture from the arterial line negative | 1056
stool examination | 1056
no white blood cells | 1056
no red blood cells | 1056
no evidence of suspected parasites | 1056
stool culture positive for Pseudomonas aeruginosa | 1056
plain film acute abdomen series | 1056
decreased bowel gas | 1056
CT of the whole abdomen | 1056
circumferential wall thickening | 1056
mucosal hyperenhancement | 1056
drooling inhibited with atropine eye drops | 1056
meropenem | 1056
antidiarrhoeal drugs | 1056
cholestyramine | 1056
octreotide | 1056
lower GI bleeding | 1200
further diagnostic work-up | 1200
serum CMV PCR viral load | 1200
5473 copies/mL | 1200
esophagogastroduodenoscopy | 1200
colonoscopy | 1200
whitish plaque on erythaematous and breaking mucosa | 1200
erythaematous mucosa | 1200
erythaematous friable mucosa | 1200
multiple aphthous ulcers | 1200
multiple small shallow ulcers | 1200
CMV viral load of the colonic tissue | 1200
> 500000 copies/mL | 1200
oesophageal biopsies | 1200
gastric biopsies | 1200
ileal biopsies | 1200
colonic biopsies | 1200
mixed inflammatory cells | 1200
viral-infected cells | 1200
intranuclear and intracytoplasmic inclusions | 1200
immunohistochemistry for CMV positive | 1200
ganciclovir | 1200
pulse methylprednisolone | 1200
unremitting diarrhoea improved | 1344
stool output 1-2 L per day | 1344
no content from the nasogastric tube | 1344
cyclophosphamide | 1344
no serious infection | 1344
no diarrhoea | 1344
neurological status improved | 1344
stable during 10 mo of follow-up | 1344