70 years old | 0
male | 0
admitted to the hospital | 0
consciousness disorder | 0
fever | 0
nausea | 0
vomiting | 0
atopic dermatitis | -8760
colon cancer | -8760
mitral valve stenosis | -8760
ischemic cardiomyopathy | -8760
resection of the sigmoid colon | -2628
adjuvant chemotherapy | -2628
mitral valve replacement | -1752
coronary artery bypass | -1752
local recurrence in the pelvis | -504
totally implantable central venous access device insertion | -504
chemotherapy | -504
impaired consciousness | 0
Glasgow Coma Scale | 0
blood pressure 90/70 mmHg | 0
heart rate 120 beats/min | 0
respiratory rate 24 breaths/min | 0
oxygen saturation 96% | 0
body temperature 38.4℃ | 0
no rash or redness at the site of the totally implantable central venous access device | 0
high inflammation | 0
renal dysfunction | 0
liver dysfunction | 0
disseminated intravascular coagulopathy | 0
high lactate levels | 0
plain computed tomography of the chest and abdominal areas | 0
unremarkable changes | 0
local recurrence at the pelvis showed no change | 0
Gram-positive cluster-forming cocci | 0
antimicrobial therapy with meropenem | 0
antimicrobial therapy with linezolid | 0
intravenous fluids | 0
norepinephrine | 0
mechanical ventilator support | 0
admitted to the intensive-care unit | 0
totally implantable central venous access device removal | 48
no abscess at the surgical site | 48
prosthetic valve endocarditis suspected | 48
transthoracic echocardiograms | 48
MRSA detected in two sets of blood cultures | 72
MRSA detected in urine culture | 72
prolonged state of shock | 72
multiple organ failure | 72
antimicrobial therapy changed to linezolid and clindamycin | 72
intravenous immune globulin | 72
transesophageal echocardiogram | 72
vegetation at the prosthetic mitral valve | 72
diagnosed with PVE caused by MRSA | 72
antimicrobial therapy changed to daptomycin | 96
persistent fever | 144
elevation of CRP | 144
whole-body enhanced CT | 144
multiple cerebral emboli with cerebral abscesses | 144
bilateral renal infarctions with abscesses | 144
spleen infarction | 144
antimicrobial therapy changed to linezolid | 144
recovered from state of persistent shock | 192
weaned off mechanical ventilation | 192
TEE showed enlargement of the vegetation | 264
abscess around the prosthetic valve | 264
surgery for PVE required | 264
mitral valve re-replacement with a bioprosthetic valve | 312
intraoperative valve culture positive for MRSA | 312
antimicrobial therapy with linezolid continued | 312
cerebral infarction | 672
vegetation on the mitral valve | 672
diagnosed with recurrent PVE | 672
antimicrobial therapy changed to vancomycin and rifampicin | 672
all blood cultures obtained after surgery were negative | 672
intravenous antimicrobial therapy continued for four weeks | 672
changed to oral sulfamethoxazole/trimethoprim and rifampicin | 840
became almost permanently bedridden | 840
transferred to a long-term-care sanatorium | 840
antibiotic susceptibility pattern of MRSA | 0
resistance to gentamycin | 0
sensitivity to clindamycin | 0
sensitivity to minocycline | 0
sensitivity to levofloxacin | 0
sensitivity to sulfamethoxazole/trimethoprim | 0
sensitivity to vancomycin | 0
sensitivity to teicoplanin | 0
sensitivity to linezolid | 0
sensitivity to daptomycin | 0
minimum inhibitory concentrations of antimicrobial agents | 0
MLST conducted | 0
ST type obtained | 0
agr typing conducted | 0
Coa typing conducted | 0
SCCmec typing conducted | 0
diagnosis of SCCmecIVl | 0
PCR of various virulence genes | 0
MRSA isolates belonged to ST8 | 0
MRSA isolates belonged to agr l | 0
MRSA isolates belonged to SCCmec type IVl | 0
MRSA isolates belonged to CoaIII | 0
MRSA isolates were negative for PVL | 0
MRSA isolates were negative for ACME-related genes | 0
MRSA isolates were positive for tst-1 | 0
MRSA isolates were positive for sec | 0
MRSA isolates were positive for sel | 0