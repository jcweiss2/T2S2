3 years old | 0 | 0 
female | 0 | 0 
admitted to the hospital | 0 | 0 
fever | -72 | 0 
diarrhea | -72 | 0 
abdominal pain | -72 | 0 
severe dehydration | -72 | 0 
critically ill | 0 | 0 
pediatric intensive care unit admission | 0 | 0 
tachypneic | 0 | 0 
rapid shallow breathing | 0 | 0 
hypotensive | 0 | 0 
evidence of severe dehydration | 0 | 0 
purpuric eruption | 0 | 0 
no organomegaly | 0 | 0 
no lymphadenopathy | 0 | 0 
pancytopenia | 0 | 0 
absolute neutropenia | 0 | 0 
renal impairment | 0 | 0 
electrolyte imbalance | 0 | 0 
hyperuricemia | 0 | 0 
coagulopathy | 0 | 0 
disseminated intravascular coagulation | 0 | 0 
high inflammatory markers | 0 | 0 
gram-negative Bacilli Escherichia coli | 0 | 0 
intravenous fluid therapy | 0 | 168 
blood components transfusion | 0 | 168 
correction of electrolyte disturbance | 0 | 168 
antibiotic therapy | 0 | 168 
provisional diagnosis of acute infectious gastroenteritis | 0 | 0 
sepsis | 0 | 0 
severe dehydration | 0 | 0 
acute renal failure | 0 | 0 
disseminated intravascular coagulation | 0 | 0 
pelvi-abdominal ultrasound | 0 | 0 
bone marrow aspirate | 0 | 0 
hypocellular bone marrow | 0 | 0 
no abnormal cells | 0 | 0 
discharged | 168 | 168 
unexplained irritability | 504 | 504 
abnormal behavior | 504 | 504 
hallucinations | 504 | 504 
failure to recognize parents | 504 | 504 
vital stability | 504 | 504 
well hydrated | 504 | 504 
normal hematological indices | 504 | 504 
normal coagulation parameters | 504 | 504 
normal renal panel | 504 | 504 
normal serum electrolytes | 504 | 504 
brain imaging studies | 504 | 504 
magnetic resonance imaging | 504 | 504 
magnetic resonance arteriography | 504 | 504 
magnetic resonance venography | 504 | 504 
thrombosis in both the left sigmoid and the transverse sinuses | 504 | 504 
workup of thrombophilia | 504 | 504 
no thrombocytosis | 504 | 504 
normal coagulation profile | 504 | 504 
normal protein C and S | 504 | 504 
antithrombin III | 504 | 504 
genetic testing for the thrombophilia mutations panel | 504 | 504 
pediatric cardiologist assessment | 504 | 504 
electrocardiogram | 504 | 504 
echocardiography | 504 | 504 
low molecular weight heparin | 504 | 720 
improved | 504 | 720 
discharged | 720 | 720 
follow-up appointment | 720 | 720 
readmitted | 1008 | 1008 
fever | 1008 | 1008 
pallor | 1008 | 1008 
abdominal enlargement | 1008 | 1008 
leukocytosis | 1008 | 1008 
anemia | 1008 | 1008 
thrombocytopenia | 1008 | 1008 
peripheral smear | 1008 | 1008 
blast cells | 1008 | 1008 
abdominal ultrasonography | 1008 | 1008 
hepatosplenomegaly | 1008 | 1008 
bone marrow examination | 1008 | 1008 
hypercellular bone marrow | 1008 | 1008 
blast cells | 1008 | 1008 
immunophenotyping | 1008 | 1008 
CD10 | 1008 | 1008 
CD20 | 1008 | 1008 
CD79a | 1008 | 1008 
diagnosis of Common ALL | 1008 | 1008 
induction therapy | 1008 | 1008 
consolidation | 1008 | 1008 
thrombophilia mutations panel result | 1056 | 1056 
positive factor XIII V34L | 1056 | 1056 
MTHFR A1298C homozygous mutations | 1056 | 1056 
heterozygous positive factor V Leiden mutation | 1056 | 1056 
follow-up MRV | 1056 | 1056 
complete recanalization of the thrombosed sinuses | 1056 | 1056 
no new thrombi | 1056 | 1056 
complete remission | 1056 | 1056 
regular follow-up | 1056 | 1056 
no other thrombotic events | 1056 | 1056 
no leukemia relapses | 1056 | 1056