18 years old | 0
male | 0
admitted to the hospital | 0
fever | -72
rash | -72
acne | -672
minocycline | -672
increased WBC count | 0
eosinophilia | 0
systemic involvement |?
