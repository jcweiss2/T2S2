83 years old | 0
    female | 0
    chest pain | 0
    abdominal pain | 0
    severe hypotension | 0
    normal ECG | 0
    no change in cardiac enzymes levels | 0
    admitted to intensive care unit | 0
    ileus | 0
    hypovolemic shock | 0
    septic shock | 0
    feculent vomiting | 24
    cardiorespiratory arrest | 24
    resuscitation | 24
    unsuccessful resuscitation | 24
    death | 24
    autopsy | 144
    pallor of entire body skin | 144
    fibrosis of myocardial muscle | 144
    hypertrophy of myocardial muscle | 144
    pulmonary edema | 144
    cerebral edema | 144
    hematoma in left hypochondrium | 144
    liver cyanosis | 144
    fatty changes in liver | 144
    splenic cyanosis | 144
    right kidney cyst | 144
    left kidney surrounded by hematoma | 144
    chronic gastric ulcer | 144
    no acute hemorrhage in gastric ulcer | 144
    severe atherosclerotic changes in arteries | 144
    abdominal aortic rupture | 144
    pulmonary cyanosis | 144
    right lower lobe yellow-brown nodule | 144
    calcified nodule | 144
    mature adipose tissue | 144
    hematopoietic cells | 144
    myeloid cells | 144
    megakaryocytes | 144
    erythroid cells | 144
    mature bony tissue | 144
    no extramedullary hematopoiesis in liver | 144
    no extramedullary hematopoiesis in spleen | 144
    pulmonary myelolipoma | 144
    