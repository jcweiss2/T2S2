61 years old | 0
male | 0
caucasian | 0
admitted to the hospital | 0
shortness of breath | 0
hypoxia | 0
hematemesis | 0
accidental extrication of percutaneous endoscopic gastrostomy (PEG) | -1
type II diabetes mellitus | -672
hypothyroidism | -672
respiratory failure | -672
tracheostomy collar | -672
perforated duodenal ulcer | -4320
septic shock | -4320
ventilator | -4320
tracheostomy | -4320
antibiotics | -4320
PEG placement | -4320
levothyroxine | -4320
insulin | -4320
ipratropium-albuterol nebulizer | -4320
morphine | -4320
intralipid | -4320
clinimix/dextrose amino acid infusion | -4320
scopolamine patch | -4320
pulse oximetry 86% | -1
supplemental oxygen | -1
coffee-ground emesis | -0.5
denies non-steroidal anti-inflammatory drugs use | 0
denies cough | 0
denies fever | 0
denies hemoptysis | 0
denies hematemesis before presentation | 0
supplemental oxygen through trach collar | 0
saturating 96-100% | 0
frail | 0
communicating in complete sentences | 0
blood pressure 113/63 mm Hg | 0
temperature 97.9 F | 0
pulse 110 beats/min | 0
respiratory rate 22 breaths/min | 0
diminished breath sounds | 0
inspiratory wheezing on the right lower base | 0
non-distended | 0
normal bowel sounds | 0
no stigmata of blood or secretions from patent PEG tube insertion site | 0
elevated blood urea nitrogen 54 mg/dl | 0
creatinine 0.9 mg/dl | 0
hemoglobin 10.9 g/dl | 0
leukocytosis 29.4 × 103/mm3 | 0
bandemia (11% of white blood count) | 0
hypoalbuminemia 2.4 g/dl | 0
mildly elevated alanine aspartate (61 u/L) | 0
INR 1.1 | 0
X-ray revealing a possible air-bronchogram on the right lower lobe | 0
pneumonia | 0
intravenous hydration | 1
broad-spectrum intravenous antibiotics | 1
intravenous pantoprazole | 1
esophagogastroduodenoscopy (EGD) | 2
severe esophagitis | 2
diffuse dark mucosal discoloration | 2
erosion | 2
profound ulceration | 2
ischemic necrosis | 2
resolution of gastrointestinal (GI) bleeding | 4
hypoxia | 12
intensive care monitoring | 12
cardiac arrest | 24
death | 24
no obvious signs or symptoms suggesting AEN before experiencing the cardiac arrest | -24