64 years old | 0
female | 0
admitted to intensive care unit | 0
confusion | 0
fever | 0
temperature at 38.8 °C | 0
blood pressure at 105/73 mmHg | 0
heart rate at 129 bpm | 0
agitated behavior | 0
abdominal sensitivity | 0
WBC at 14.000/mm3 | 0
elevated C-reactive protein at 160.6 mg/l | 0
creatinine at 126 μmol/l | 0
all blood cultures were negative | 0
screening for HIV, HCV and HBV was negative | 0
screening for syphilis was negative | 0
MRI of the head showed 4 ring enhancing lesions | 0
cerebral abscesses | 0
cerebellar lesion at 28 mm | 0
frontal right image at 15 mm | 0
parietal lesion at 17 mm | 0
occipital lesion at 15 mm | 0
lumbar puncture found 275/mm3 WBC | 0
4% PNN | 0
89% lymphocytes | 0
no germ was retrieved | 0
total body scan imaging revealed an 11 cm liver abscess | 0
right-sided pleural effusion | 0
negative microbiological cultures from thoracentesis and liver drains | 0
brown purulent liquid recovered | 0
intravenous Ceftriaxone started | 0
oral Metronidazole started | 0
clinical and biological improvement | 120
patient became afebrile | 120
neurological symptoms resolved | 120
transferred to infectious diseases unit | 120
cerebral MRI performed at 3 weeks of treatment | 504
no major difference in the size of the brain abscesses | 504
ultrasound showed stagnation in the size of the liver abscess | 504
craniotomy with drainage of brain abscesses recommended | 504
brain biopsy found a mixed inflammatory reaction | 504
important macrophagic infiltrate and granulomas | 504
no evident pathogenic microorganism | 504
aerobic and anaerobic cultures were negative | 504
PCR product detected with 16S ribosomal DNA from Fusobacterium nucleatum | 504
Ceftriaxone changed to Clindamycine | 504
Metronidazole continued | 504
18F-fludeoxyglucose positron emission tomography (FDG-PET) performed | 504
no other infection site besides the liver, pleura and the brain | 504
MRI of brain performed 12 weeks after the beginning of treatment | 1008
brain abscesses decrease in size | 1008
cerebellar lesion decreased to 8 mm | 1008
frontal right image decreased to 6.5 mm | 1008
parietal and occipital lesions decreased to 6.5 mm | 1008
decrease of ring enhancing intensity and surrounding edema | 1008
treatment with only oral metronidazole continued | 1008
total duration of treatment 20 weeks | 1344
brain, hepatic and pulmonary images performed 6 months after the initial presentation | 2016
stability of brain images | 2016
complete recovery of hepatic abscesses and pleural effusion | 2016
good clinical recovery | 2016
good biological evolution | 2016
CRP at 3.7 mg/l | 2016
no fever | 2016
intra-uterine device removed | -24
culture of device remained negative | -24