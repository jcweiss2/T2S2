65 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
liver cirrhosis | -8760 | 0 | Factual
chronic hepatitis B | -8760 | 0 | Factual
hepatocellular carcinoma | 0 | 0 | Factual
left lobe hepatectomy | 0 | 300 | Factual
intravenous glycopyrrolate | -1 | 0 | Factual
general anesthesia | 0 | 300 | Factual
propofol | 0 | 0 | Factual
rocuronium | 0 | 0 | Factual
remifentanil | 0 | 300 | Factual
sevoflurane | 0 | 300 | Factual
mechanical ventilation | 0 | 300 | Factual
electrocardiography | 0 | 300 | Factual
arterial blood pressure monitoring | 0 | 300 | Factual
central venous pressure monitoring | 0 | 300 | Factual
SpO2 monitoring | 0 | 300 | Factual
stable vital signs | 0 | 60 | Factual
sudden decrease in arterial blood pressure | 60 | 60 | Factual
tachycardia | 60 | 60 | Factual
ST elevation on EKG | 60 | 60 | Factual
resuscitation with colloid and catecholamines | 60 | 120 | Factual
intraoperative ultrasonography | 60 | 120 | Factual
massive air emboli in both heart | 60 | 120 | Factual
diagnosis of VAE and PAE | 60 | 120 | Factual
arterial blood gas analysis | 60 | 60 | Factual
catecholamine administration | 70 | 300 | Factual
systolic blood pressure maintenance | 120 | 300 | Factual
heart rate maintenance | 120 | 300 | Factual
central venous pressure maintenance | 120 | 300 | Factual
end-tidal carbon dioxide restoration | 120 | 300 | Factual
norepinephrine infusion | 120 | 300 | Factual
fluid resuscitation | 120 | 300 | Factual
air emboli disappearance | 130 | 130 | Factual
hepatectomy completion | 130 | 300 | Factual
intensive care unit admission | 300 | 300 | Factual
mechanical ventilation | 300 | 264 | Factual
norepinephrine infusion | 300 | 264 | Factual
abnormal PT/PTT | 300 | 300 | Factual
fibrinogen | 300 | 300 | Factual
d-dimer | 300 | 300 | Factual
antithrombin III | 300 | 300 | Factual
CK-MB | 300 | 300 | Factual
troponin-T | 300 | 300 | Factual
ST elevation on EKG | 300 | 300 | Factual
EKG recovery | 744 | 744 | Factual
trans-thoracic echocardiogram | 744 | 744 | Factual
no patent foramen ovale | 744 | 744 | Factual
vital signs stability | 744 | 744 | Factual
norepinephrine infusion tapering | 744 | 744 | Factual
mental status unchanged | 120 | 264 | Factual
brain CT and MRI | 1200 | 1200 | Factual
multiple acute cerebral infarctions | 1200 | 1200 | Factual
weaning to spontaneous ventilation | 2640 | 2640 | Factual
extubation | 2640 | 2640 | Factual
vital signs instability | 3600 | 3600 | Factual
catecholamine administration | 3600 | 744 | Factual
panperitonitis confirmation | 7440 | 7440 | Factual
cardiac arrest | 7440 | 7440 | Factual
death | 7440 | 7440 | Factual