60 years old | 0
    female | 0
    atrial fibrillation | -8760
    dilated cardiomyopathy | -8760
    implanted biventricular pacing implantable cardioverter defibrillator | -8760
    oral warfarin | -8760
    impaired consciousness | -24
    found lying at home | -24
    transported to hospital by ambulance | -24
    JCS score II-10 | 0
    GCS score 14 (E3V5M6) | 0
    no clear neurological deficits | 0
    non-contrast head CT revealed hemorrhage in third and fourth ventricles | 0
    hemorrhage in bilateral lateral ventricles with left dominance | 0
    hemorrhage confined within ventricles | 0
    brain 3D