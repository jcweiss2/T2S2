54 years old | 0
male | 0
septic shock | 0
malaise | -168
rigors | -168
right upper quadrant pain | -168
flank pain | -168
treated with antibiotics | -168
ceftriaxone | -168
metronidazole | -168
acute cholecystitis | -168
ascending cholangitis | -168
multi-organ failure | 0
oxygen saturations of 80% | 0
haemodynamic compromised | 0
systolic blood pressure of 80 | 0
sinus tachycardia up to 120 beats per minute | 0
bilateral renal angle tenderness | 0
intubated | 0
transferred to the intensive care unit | 0
severe metabolic acidosis | 0
anuric renal failure | 0
thrombocytopenia | 0
dialysis | 0
antibiotics broadened to meropenum | 0
metronidazole | 0
fluconazole | 0
CT scan | 0
bilateral EPN | 0
type two diabetes | 0
referred to the urology service | 0
discussion with the patient's next of kin | 0
decision not to perform bilateral nephrectomies | 0
coagulopathic with an INR of 16 | 24
metabolic acidosis progressed | 24
liver failure | 24
worsening synthetic failure | 24
required maximal inotropic support | 24
case conference | 24
decision to treat medically | 24
supportive care and antibiotics | 24
antibiotics rationalised to ceftriaxone | 72
CT scan on day 3 | 72
no drainable collections | 72
extubated | 144
ongoing dialysis | 144
IV ceftriaxone | 144
transitioned to oral augmentin duo forte | 672
repeat CT after 4 weeks | 672
no significant change in the appearance of the kidneys | 672
afebrile | 672
hemodynamically stable | 672
intermittent hemodialysis | 672
creatinine remained 250 | 672