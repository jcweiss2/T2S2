84 years old | 0
male | 0
admitted to the hospital | 0
febrile | 0
encephalopathic | 0
melanotic stool | 0
stroke with residual left hemiparesis | -8760
gastrointestinal bleed | -8760
heart rate 92 | 0
blood pressure 95/51 | 0
obtunded | 0
dry mucous membranes | 0
non-tender and non-distended abdomen | 0
no evidence of skin changes nor infection | 0
volume resuscitated | 0
initiated on broad spectrum antibiotics | 0
admitted to the intensive care unit (ICU) | 0
presumed diagnoses of gastrointestinal bleed | 0
presumed diagnoses of sepsis of unknown etiology | 0
elevated lactic acid | 0
elevated procalcitonin | 0
hypotension | 0
Gastroenterology consulted | 0
endoscopy deferred | 0
laboratory values normalized | 2
hemodynamics normalized | 2
returned to baseline mental status | 2
no history of weight loss | 0
no history of decreased appetite | 0
no history of recurrent melanotic stool | 0
no history of alterations in bowel habits | 0
right hip erythema | 24
right hip induration | 24
right hip pain | 24
no crepitus | 24
CT of the right hip | 24
concern for necrotizing soft tissue infection | 24
gas involving the right retroperitoneum and upper thigh | 24
no evidence of abscess | 24
General surgery consulted | 24
necrotizing fasciitis | 24
operative intervention declined | 24
clinically improved with non-operative treatment | 56
CT of his abdomen and pelvis | 56
7.1 cm proximal right colon mass | 56
invasion into the retroperitoneum | 56
gas tracking into adjacent soft tissues | 56
concerning for a perforated malignancy | 56
Colorectal surgery consulted | 56
tumor resection with debridement | 56
elected for palliative care | 56
transitioned to hospice care | 56
expired | 240