17 years old | 0
male | 0
admitted to the hospital | 0
past medical history of poorly-controlled persistent asthma | -672
past medical history of obesity | -672
past medical history of hypertension | -672
past medical history of type II diabetes | -672
shortness of breath | 0
febrile | 0
tachycardic | 0
tachypneic | 0
elevated blood pressure | 0
oxygen saturation 98% on room air | 0
weight 122 kg | 0
body mass index (BMI) of 50.1 kg/m2 | 0
skin tenderness and warmth in the gluteal area | -96
2 pack-year history of smoking | -672
non-adherent with metformin | -672
non-adherent with insulin glargine | -672
obese and non-toxic appearing | 0
dry mucous membranes | 0
diminished breath sounds bilaterally without wheezing | 0
soft abdomen without guarding or tenderness | 0
erythematous and indurated left scrotum, left perineum, and bilateral buttocks | 0
sodium of 131 mEq/L | 0
potassium of 3 mEq/L | 0
chloride of 92 mEq/L | 0
phosphate of 2.3 mg/dL | 0
glucose of 320 mg/dL | 0
C-reactive protein (CRP) of 28.6 mg/dL | 0
ultrasound consistent with cellulitis without abscess formation | 0
electrolyte abnormalities | 0
uncontrolled type II diabetes | 0
perineal cellulitis | 0
started on oral clindamycin | 0
started on intravenous (IV) fluids | 0
started on insulin for hyperglycemia | 0
febrile and tachycardic with worsening hypertension | 12
perineal cellulitis progressed to large, fluid-filled blisters | 24
ruptured and drained purulent fluid | 24
broadened antibiotic regimen to cefepime and vancomycin | 24
white blood cell count of 11 K/uL with 35% bands | 24
worsening CRP of 46.4 mg/dL | 24
contrast computed tomography (CT) scan of the pelvis | 24
scrotal wall edema and fluid within the scrotum | 24
extensive fat stranding and air in the subcutaneous tissue | 24
Fournier’s gangrene | 24
general surgery consulted for urgent debridement | 24
IV clindamycin added to vancomycin and cefepime | 24
underwent extensive surgical debridement | 48
intraoperative findings revealed significant necrotic soft tissue | 48
septic shock and diabetic ketoacidosis | 48
transferred to the pediatric intensive care unit | 48
required vasopressors and an insulin infusion | 48
underwent a second debridement | 72
no evidence of ongoing necrotizing infection | 72
vacuum-assisted closure (VAC) performed | 72
wound culture grew Actinomyces species | 72
initial fungal culture and anaerobic cultures had no growth | 72
fungal cultures from a repeat debridement were positive for Candida albicans | 96
blood cultures remained negative | 96
antimicrobial regimen narrowed to piperacillin-tazobactam and fluconazole | 96
underwent a total of 6 surgical debridements | 240
wound VAC changes | 240
diverting colostomy and Foley catheter placement | 240
multiple reconstructive surgeries with split-thickness skin grafts and fasciocutaneous flaps | 240
discharged sixty days after admission | 1440
surgical wounds were healing well at follow-up appointments | 2160
cleared by Plastic Surgery for colostomy takedown | 2160
discharged on a 6-month course of amoxicillin | 2160
no known recurrences | 4320