42 years old | 0
female | 0
anxiety | -8760
obesity | -8760
body mass index 31 kg/m2 | -8760
Roux-en-Y gastric bypass | -8760
dyspepsia | -720
nausea | -720
vomiting | -720
poor oral intake | -720
personality changes | -720
irritability | -720
buspirone | -720
discontinued buspirone | -720
no medications | -2160
confusion | -1440
lethargy | -1440
intermittent confusion and lethargy | -1440
constant confusion and lethargy | -720
sleeping for most of the day | -168
difficulty remembering simple facts | -168
admitted to the emergency department | 0
hyperammonemia | 0
transaminitis | 0
no known liver disease | 0
no alcohol consumption | 0
mild chronic periportal inflammation | -720
moderate macrosteatosis | -720
no cirrhosis | -720
negative acetaminophen level | 0
negative urine drug screen | 0
unremarkable brain computed tomography | 0
fatty liver | 0
no cirrhosis | 0
blood and urine cultures collected | 0
intravenous thiamine | 0
rectal lactulose | 0
admitted to the intensive care unit | 0
excluded Wilson disease | 24
excluded hemochromatosis | 24
excluded viral and autoimmune hepatitis | 24
polymicrobial bacteremia | 24
Escherchia coli | 24
methicillin-sensitive Staphylococcus aureus | 24
Enterococcus faecalis | 24
urine culture grew Enterococcus species | 24
intravenous vancomycin | 72
piperacillin/tazobactam | 72
sodium benzoate/sodium phenylacetate | 72
rifaximin | 72
zinc | 72
arginine | 72
supplemental parenteral lipids | 72
glucose | 72
followed commands | 96
extubated | 120
ammonia and liver enzymes normalized | 168
mentation returned to baseline | 168
discharged home | 240
counseled on a protein-restricted diet | 240
instructed to follow-up with outpatient hepatology | 240
genetic counseling advised | 240