67 years old | 0
male | 0
admitted to the hospital | 0
untreated hypertension | 0
diabetes | 0
acutely increasing chest and back pain | -12
electrocardiogram assessment | 0
ST segment elevation in V1-6 | 0
transthoracic echocardiography | 0
wall motion abnormality in the anterior region | 0
anterior acute STEMI | 0
maximum creatinine kinase level | 0
maximum CK-MB level | 0
coronary angiography | 0
total occlusion at the middle section of the left anterior descending artery | 0
percutaneous coronary intervention | 0
acute strong right subcostal and epigastric pain | 5
abdominal computed tomography | 5
gallstones detected | 5
liver enzyme level did not increase | 5
treated conservatively for biliary colic | 5
symptoms of right heart failure | 5
fatigue | 5
loss of appetite | 5
myocardial enzyme level decreased | 5
no heart murmur | 5
no new ECG abnormalities | 5
daily TTE did not demonstrate new signs of decreased systolic function | 5
myocardial ischemia | 5
mechanical complications | 5
stronger right subcostal and epigastric pain | 120
positive Murphy sign | 120
increase in C-reactive protein | 120
new CT revealed an edematous gallbladder | 120
white blood cell count increased | 120
serum liver and biliary enzymes slightly high | 120
aspartate aminotransferase | 120
alanine aminotransferase | 120
gamma-glutamyl transpeptidase | 120
gallstones vanished | 120
abdominal symptoms suspicious of acute cholecystitis | 120
laparoscopic cholecystectomy | 120
pathological examination revealed chronic cholecystitis | 120
exacerbated pain | 144
admitted to the intensive care unit | 144
restlessness | 144
tachypnea | 144
shock | 144
no new abnormality on TTE and ECG | 144
managed for septic shock | 144
broad-spectrum antibiotics | 144
tracheal intubation | 144
invasive ventilation | 144
continuous renal replacement therapy | 144
norepinephrine administered | 144
dobutamine administered | 144
epinephrine administered | 144
hemodynamic state deteriorated | 144
5th TTE revealed a left-to-right shunt through the ventricular septum | 154
VSR suspected | 154
intra-aortic balloon pumping | 154
venous-artery extracorporeal membrane oxygenation | 154
emergency patch closure of the VSR | 154
perforation at the apical septal region confirmed | 154
intraoperative transesophageal echocardiography | 154
right subcostal pain diminished | 168
hemodynamics improved | 168
left the ICU | 504
transferred | 1776