61 years old | 0
    male | 0
    hypertension | 0
    squamous cell carcinoma of the skin | 0
    cyst removal (unsuccessful) | -1464
    excision of cyst under general anesthesia | -672
    removal of squamous cell skin lesions (left upper arm and central chest) | -672
    TMP-SMX prescribed | -672
    completed TMP-SMX course | -336
    fevers (Tmax 102 F) | -72
    confusion | -72
    admitted to the hospital | 0
    altered mental status | 0
    alert and oriented x1 | 0
    temperature 101.7 F | 0
    BP 120/56 mmHg | 0
    HR 120 beats/min | 0
    RR 22 breaths/min | 0
    O2 saturation 94% on room air | 0
    sinus tachycardia | 0
    mild tenderness in right upper quadrant | 0
    healing excisions (left forearm and central chest) | 0
    sutured wound on upper middle back | 0
    diffuse petechiae | 0
    maculopapular rash (back, chest, abdomen) | 0
    no mucosal/oral involvement | 0
    rash not present on soles/palms | 0
    no bullae or pustules | 0
    WBC 5.1 × 10³/uL | 0
    no eosinophils | 0
    no monocytes | 0
    platelet count 13 × 10³/uL | 0
    sodium 122 mmol/L | 0
    creatinine 2.77 mg/dL | 0
    BUN 50 mg/dL | 0
    AST 238 units/L | 0
    ALT 79 units/L | 0
    PT 12.4 s | 0
    INR 1.1 | 0
    APTT 65 s | 0
    sepsis criteria met | 0
    fluid resuscitation | 0
    blood cultures drawn | 0
    empiric antibiotics (vancomycin, piperacillin/tazobactam) | 0
    platelet transfusion (1 unit) | 0
    transferred to ICU | 0
    consultations (Infectious Disease, Nephrology, Hematology/Oncology) | 0
    peripheral smear (no schistocytes) | 0
    fibrinogen 125 mg/dL | 0
    D-dimer 52,292 ng/mLFEU | 0
    ADAMTS13 activity 34.9% | 0
    G6PD normal | 0
    renal injury (intrinsic) | 0
    hemoglobin 2+ in urine | 0
    trace RBCs in urine | 0
    FeNA 2.79 mEq/L | 0
    diagnosis of delayed hypersensitivity reaction to TMP-SMX | 0
    creatinine worsening | 24
    transaminitis worsening | 24
    hyponatremia worsening | 24
    blood cultures no growth (4 days) | 96
    antibiotics discontinued | 96
    mentation returned to baseline | 72
    maculopapular rash disappeared | 72
    lab values correcting | 96
    transferred out of ICU | 96
    discharged | 120
    advised to avoid TMP-SMX re-challenge | 120
