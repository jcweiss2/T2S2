32 years old | 0
pregnant woman (11 weeks) | 0
previously healthy | 0
hospitalized with hyperemesis | 0
sepsis | 0
disseminated intravascular coagulation | 0
admitted to the intensive care unit | 0
C. albicans cultured from blood | 0
C. albicans cultured from urine | 0
isolate susceptible to all antifungal agents tested | 0
MICs: amphotericin B 0.5 mg/l | 0
MICs: caspofungin 0.125 mg/l | 0
MICs: anidulafungin 0.015 mg/l | 0
MICs: fluconazole ≤0.125 mg/l | 0
MICs: itraconazole ≤0.03 mg/l | 0
MICs: micafungin ≤0.008 | 0
MICs: voriconazole ≤0.03 mg/l | 0
MICs: 5-FC ≤0.125 mg/l | 0
treatment with L-AMB (4 mg/kg) initiated | 0
treatment with caspofungin 70 mg initiated | 0
treatment with broad-spectrum antibiotics initiated | 0
L&AMB dose reduced to 2 mg/kg due to creatinine increase | 0
patient treated with combination for 12 days | 0
L-AMB and antibiotics continued for 9 more days | 0
discharged from intensive care unit | 18
fluctuating C-reactive protein (400–600 mg/l) | 18
slight fever (37.8–38.2 °C) | 18
lost fetus | 18
kidney function never recovered | 18
dependent on hemodialysis | 18
discharged from hospital | 43
no fever | 43
WBC of 7.69×10^9 l−1 | 43
CRP of 188 mg/l | 43
admitted to Department of Infectious Diseases | 77
lumbar back pain | 77
pyrexia | 77
CRP 150 mg/l | 77
bone scintigraphy showed uptake around right hip | 85
bone scintigraphy showed uptake around left sacroiliac joint | 85
bone scintigraphy showed uptake around lower spine | 85
MRI revealed vertebral infection at Th11–12 | 90
MRI revealed vertebral infection at L3–4 | 90
MRI showed no involvement of discs or spinal cavity | 90
fungal etiology suspected | 90
treatment with caspofungin (70 mg loading dose) initiated | 90
treatment with fluconazole (200 mg daily) initiated | 90
biopsy PCR negative | 91
biopsy culture negative | 91
back pain progressed during next 14 days | 90-104
CRP declined from 100 to 60 mg/l | 106
new MRI showed no regression | 106
treatment failure considered | 106
treatment changed to L-AMB 4 mg/kg/day | 106
patient slowly improved during six weeks | 106-148
discharged | 148
asymptomatic | 148
normal CRP (<8 mg/l) | 148
continuous hemodialysis three times a week | 148
fluconazole administered after each HD | 148-228
serum fluconazole concentration 9 mg/L | 228
malaise | 233
vomiting | 233
fluctuating temperature (37–38 °C) | 233
low back pain radiating to right hip | 233
readmitted to hospital | 247
increasing back pain | 247
pyrexia (39.5 °C) | 247
CRP <8 mg/l | 247
CRP increased to 80 mg/l | 248
ESR 50 | 247
L-AMB 4 mg/kg daily initiated | 252
temporal relief of symptoms | 252
pain returned and increased | 280
L-AMB dose increased to 5 mg/kg | 280
MRI showed progression of L3–4 destruction | 293
L-AMB dose increased to 6 mg/kg | 301
combined with 5-FC 3500 mg after each HD | 301
​5-FC treatment discontinued | 378
PET-CT unchanged | 378
MRI showed minimal regression | 378
bone scintigraphy showed regression of Th12-L1 uptake | 378
high dose L-AMB continued for 3 more months | 378-465
leukocyte scintigraphy showed reduced enhancement and edema of L3–4 | 465
MRI showed reduced enhancement and edema of L3–4 | 465
life-long prophylaxis discussed | 465
kidney transplant considered | 465
all anti-fungal treatment discontinued | 465
ESR remained normal | 465-678
bone scintigraphy showed minimal activity | 678
no progression detected on MRI | 678
kidney transplant received | 678
gave birth to healthy child | 678+730
no signs of relapse for 5 years | 678+1825
