hepatitis C-related cirrhosis | -120
recurrent hepatic encephalopathies | -120
chronic portal vein thrombosis | -120
liver transplantation | 0
construction of an end-to-side anastomosis of the donor portal vein to the superior mesenteric vein | 0
end-to-end bile duct anastomosis | 0
massive venous bleeding from local varices | 0
iliac conduit construction | 0
normal liver graft function | 0
stenosis of the bile duct anastomosis | 20
biliary leakage | 20
elevated liver enzymes | 20
pigtail treatment | 20
FCSCEMS insertion | 26
persisting leakage | 26
hepatitis C reinfection | 30
recurrent stenosis of the biliary anastomosis | 30
ERCP | 30
balloon dilatations | 30
placements of pigtails | 30
stent placements | 30
biopsy-proven significant fibrosis | 52
treatment with pegylated interferon and ribavirin | 52
elective ERCP | 104
recovery of 3 plastic double-pigtails | 104
cholangiogram | 104
large portobiliary fistula | 104
hemobilia | 104
FCSEMS placement | 104
prophylactic antibiotic treatment with ciprofloxacin | 104
septic shock | 106
admission to the intensive care unit | 106
hemodynamic support | 106
empiric broad-spectrum antibiotic treatment | 106
computed tomography | 106
angiography | 106
anuric kidney failure | 106
continuous venovenous hemofiltration | 106
intermittent hemodialysis | 110
evaluation for liver re-transplantation | 112
FCSEMS replacement | 136
extraction of the lying FCSEMS | 136
no evidence of persisting leakage | 136
no relevant stenosis | 136
no further endoscopic intervention | 150
no evidence of recurrent stenosis | 150
no evidence of portobiliary fistula | 150