30 years old | 0
female | 0
housewife | 0
ingestion of 15 g of KMnO4 powder | -0.25
ingestion of KMnO4 with a glass of water | -0.25
happily married | 0
no psychiatric illness in the past | 0
reached the hospital within 15 min of ingestion | -0.25
drowsy | 0
hypoxia | 0
stridor | 0
oxygen saturation 85% | 0
arterial blood gas (ABG) revealed pH 7.32/pO252.1/pCO246/HCO322/SpO286.1% | 0
tachycardia | 0
heart rate of 116/min | 0
normal blood pressure (110/70 mmHg) | 0
temperature of 98.2°F | 0
multiple patches of blackish-brown stain on face and hands | 0
oral cavity examination revealed complete brownish black staining | 0
copious secretions | 0
poor differentiation between structures of the oral cavity | 0
vocal cords swollen | 0
almost complete obstruction of airways | 0
percutaneous tracheostomy planned | 0
intubation attempted | 0
difficult intubation | 0
small size (6.5 mm high volume low pressure cuffed) endotracheal tube placed | 0
intermittent positive pressure ventilation initiated | 0
invasive ventilatory support | 0
broad spectrum antibiotics | 0
steroids | 0
proton-pump inhibitor | 0
intravenous fluids started | 0
mechanical ventilation | 0
oxygenation and ABG improved | 12
upper gastrointestinal (GI) endoscopy done on day 1 | 24
diffuse ulceration and necrotic areas in esophagus and fundus of the stomach | 24
bronchoscopy performed | 24
edematous and inflamed mucosa | 24
hemorrhagic patches in entire tracheo-bronchial tree | 24
normal renal and hepatic parameters | 0
normal electrolytes | 0
normal complete hemogram | 0
normal methemoglobin level | 0
liver function test became deranged on 2nd day | 48
rising serum bilirubin | 48
total serum bilirubin increased to 4.5 mg/dl | 48
serum glutamic pyruvic transaminase to 354 IU | 48
coagulation profile deranged | 48
INR of 2.06 | 48
decreased platelet counts (80,000/cumm) | 48
acute hepatic necrosis | 48
coagulation profile started improving on day 4 | 96
serum transaminase levels still elevated | 96
oral cavity examination on day 4 revealed significant reduction in staining of mucosa | 96
edema of upper airway structures reduced | 96
vocal cords swelling reduced | 96
patient extubated | 96
cuff leak check | 96
reintubated | 96
percutaneous tracheostomy done | 96
weaned off the ventilator on day 5 | 120
total parenteral nutrition started | 120
condition gradually improved | 120
started accepting clear liquids orally on day 8 | 192
liver functions and coagulation profile improved slowly | 192
decannulated on day 9 | 216
discharged in good health condition | 216
follow-up after 3 months was normal | 744