63 years old | 0
male | 0
married | 0
smoker | 0
non-drinker | 0
admitted to the hospital | 0
fever | 0
melena | 0
hematemesis | 0
generalized weakness | 0
constant fatigue | 0
shortness of breath | 0
no dysphagia | 0
no dyspepsia | 0
no abdominal pain | 0
no abnormal change of bowel habits | 0
no history of continuous use of NSAIDs | 0
anaemia | -168
juxtarenal abdominal aortic aneurysm | -8760
synthetic grafting aortobifemoral bypass | -8760
hypertension | -8760
type 2 diabetes mellitus | -8760
glaucoma | -8760
lens transplantation | -8760
ischaemic heart disease | -8760
catheterization | -8760
stents | -8760
taking blood pressure medications | -8760
taking diabetes medications | -8760
taking lipid medications | -8760
taking anticoagulant medications | -8760
upper GI endoscopy | 12
CT angiogram | 12
sepsis | 0
transferred to the Surgical ICU | 12
IV antibiotics | 12
referred to the surgical ward | 24
first stage of the operation | 48
exclusion aortic limb graft with endarterectomy | 48
axillofemoral bypass | 48
femoro-femoral bypass | 48
transferred to the ICU | 72
second stage of the operation | 96
intestinal adhesion | 96
aorto-duodenal fistula | 96
aortocecal fistula | 96
infected aortobifemoral graft | 96
infrarenal AAA | 96
infrarenal aortic neck control | 96
removal of old infected aortobifemoral graft | 96
closure of infrarenal abdominal aorta | 96
fistula management | 96
primary repair of the second-third part of the duodenum | 96
right hemicolectomy with primary anastomosis | 96
kept in the SICU post-operation | 120
total parental nutrition | 120
stabilized | 144
transferred to the surgical ward | 168
started on an oral diet | 168
follow-up CT scan | 240
discharged | 288
double secondary aortoenteric fistula | 0
aortoenteric fistula | 0
caecal air bubbles | 12
pus discharge | 12
blood discharge | 12 
GI haemorrhage | 0 
high-grade fever | 0 
aortic graft infection | -168 
aortobifemoral bypass graft infection | -168 
jauxternal AAA reconstruction | -8760 
communication between the aorta and the intestinal wall | 0 
prophylaxis antibiotics | -8760 
recurrence | 0 
continuity of the follow-up | 0 
control and treat any complications | 0 
early stage | 0 
clinicians should suspect AGI and double SAEF | 0 
patients with fever and melena after aneurysm surgery | 0 
intraoperative images | 96 
removal of the jauxternal AAA | 96 
closure of infrarenal abdominal aorta with double layers of protein | 96 
fistula management | 96 
primary repair of the second- third part of the duodenum | 96 
right hemicolectomy with primary anastomosis | 96 
inferior mesenteric vein | 96 
SCARE criteria | 0 
ethical approval | 0 
written informed consent | 0 
source of funding | 0 
author contribution | 0 
conflicts of interest disclosure | 0 
research registration unique identifying number | 0 
data availability statement | 0 
provenance and peer review | 0 
sponsorships or competing interests | 0 
published online | 0