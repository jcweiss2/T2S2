65 years old|0
African American|0
woman|0
BMI 26.5|0
daily smoker|0
peptic ulcer disease|0
omeprazole|0
hysterectomy|0
presented to the Emergency Department|0
worsening left sided abdominal pain|0
nausea|0
emesis|0
hematochezia|-336
denied fevers|0
denied chills|0
anorexia|0
10-pound weight loss|0
afebrile|0
focalized peritoneal signs in the left lower quadrant|0
no generalized peritonitis|0
elevated white blood count (WBC) 15.3|0
potassium 3.0 mmol/L|0
albumin 2.3 g/dL|0
normal CBC|0
normal basic metabolic profile|0
CT abdomen and pelvis showing sigmoid diverticulitis|0
3.8 × 5.5 cm gas containing pericolonic abscess|0
multidisciplinary management initiated|0
treated with intravenous levofloxacin 500 mg|0
metronidazole|0
10 fr drain placed transabdominally|0
20 ccs purulent fluid drained|0
microbial cultures grew streptococcus viridans|0
gram negative rods|0
proteus species|0
continued marked abdominal pain|0
persistent leukocytosis|0
hospital day 3|0
open Hartmann’s operation|0
perforated diverticulitis|0
serositis|0
abscess formation|0
fibrous adhesions|0
fat necrosis|0
granulation tissue|0
negative for malignancy|0
peri-operative antibiotics|0
IV cefepime 2 mg every 12 h|0
IV metronidazole 500 mg every 8 h|0
POD #1|24
mild hypotension|24
tachycardia|24
resolved after epidural infusion temporarily suspended|24
clear liquid diet started|24
minimal intake|24
no evidence of bowel function|24
epidural analgesic catheter removed|96
POD #4|96
Total Parenteral Nutrition started|120
POD #5|120
POD #7|168
continuous hyponatremia|168
hyponatremia ranging 132−134 mmol/L|168
potassium 3.4–3.5 mol/L|168
hypochloremia 95 mmol/L|168
POD #8|192
new onset emesis|192
intermittent periods of hypotension|192
slight sinus tachycardia|192
CT abdomen and pelvis with PO and IV contrast obtained|192
bilateral adrenal enlargement|192
decreased definition consistent with bilateral adrenal gland hemorrhage/infarction|192
random serum cortisol level 2.6 ug/dL|192
no evidence of DVT|192
no evidence of PE|192
serum cardiac troponin level undetectable|192
transthoracic echocardiogram showed EF 60–65%|192
no valvular disease|192
grade 1 diastolic dysfunction|192
endocrinology consulted|192
stress dose hydrocortisone sodium succinate 100 mg started|192
hydrocortisone 100 mg every 8 h|192
clinical status improved within 24 h|216
blood pressure stabilized|216
heart rate stabilized|216
return of bowel function|216
tolerated diet|216
discharged to rehabilitation facility|336
POD#14|336
TPN discontinued|336
antibiotics discontinued|336
steroids tapered down to 5 mg prednisone twice daily|336
5 mg daily thereafter|336
seen in clinic one month after discharge|672
follow up delayed due to transportation issues|672
after four months|2880
continued steroid dependence|2880
no signs of adrenal recovery|2880
continued on hydrocortisone 20 mg in the morning and 10 mg at night|2880
