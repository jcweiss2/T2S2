22 years old | 0
female | 0
admitted to the hospital | 0
upper abdominal pain | 0
LRGB | -2556
lost 50 kg | -2556
gall bladder stones | 0
MRI scan | 0
open cholecystectomy | 24
trans-cystic balloon dilation | 24
cholangiogram | 24
poor drainage | 24
small gallstones | 24
re-operated | 120
cholascos | 120
cystic duct ligation | 120
drainage | 120
endoscopy | 144
hematemesis | 144
blood in the jejunum | 144
severe septicaemia | 216
acute respiratory distress syndrome | 216
transferred to ICU | 216
laparotomy | 312
internal hernia | 312
necrosis of 1 m jejunum | 312
caesarean | 312
premature girl | 312
necrotic intestine removed | 312
second look operation | 336
third look operation | 360
small bowel resections | 360
saliva fistula | 360
jejunostomy | 360
blind closed ileum | 360
infectious complications | 744
pneumothorax | 744
thrombosis of the superior mesenteric vein | 744
thrombosis of the iliac veins | 744
exposed bowel parquet | 744
covered with split skin | 744
transferred to intestinal failure unit | 744
good appetite | 744
no absorption of food | 744
central venous line | 744
Hickmann catheter | 744
received 2200 kcal | 744
SMOF Kabiven | 744
vitamins | 744
trace elements | 744
isotonic saline | 744
fluid balance | 744
complications | 744
Hickmann catheter removed | 744
yeast infection | 744
candida albicans | 744
peripherally inserted central venous catheter | 744
PICCline | 744
discharged | 1200
home parenteral nutrition | 1200
intestinal continuity reconstructed | 1680
defect in the anterior abdominal wall | 1680
closed with bilateral partial component separation | 1680
PICCline occluded | 1848
removed | 1848
trying without parenteral nutrition | 1908
doing well | 1908
weight increased | 1908
bowel movements | 1908
haemoglobin increased | 1908
albumin increased | 1908