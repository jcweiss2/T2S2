32 years old | 0\
    woman | 0\
    presented to the clinic | 0\
    fever of unknown origin | -2160\
    progressively increasing cough | -2160\
    hoarseness of voice | -504\
    odynophagia | -504\
    fever started intermittently | -7200\
    pregnancy | -6480\
    ectopic pregnancy | -6480\
    ruptured ectopic pregnancy | -6480\
    admitted to the hospital | -6480\
    laparoscopic exploration | -6480\
    cultures from fallopian tube positive for Mycobacterium tuberculosis | -6480\
    developed sepsis | -6480\
    adult respiratory distress syndrome | -6480\
    shifted to Intensive Care Unit | -6480\
    central line placed in left subclavian vein | -6480\
    tracheal cultures growth of Pseudomonas aeruginosa | -6480\
    blood cultures presence of Enterobacter cloacae | -6480\
    bronchial lavage confirmed pulmonary tuberculosis | -6480\
    absence of malignancy | -6480\
    antibiotics started | -6480\
    anti-TB medications started | -6480\
    improved | -6480\
    discharged home | -6480\
    mother of two children | 0\
    no comorbidities | 0\
    no family history of TB | 0\
    presented again | -1440\
    vomiting | -1440\
    headache | -1440\
    exertional dyspnea | -1440\
    inability to talk | -1440\
    difficulty opening left eye | -1440\
    significant weight loss | -1440\
    brain MRI revealed disseminated central nervous system TB | -1440\
    anti-TB regimen adjusted | -1440\
    left-sided hemiparesis | -1440\
    gradually recovered | -1440\
    discharged home | -1440\
    presented again | -1440\
    hoarseness of voice | -1440\
    odynophagia | -1440\
    chest radiograph revealed superior mediastinal mass on left | -1440\
    CT scan of chest showed large subclavian artery pseudoaneurysm | -1440\
    CT angiogram confirmed large left subclavian artery pseudoaneurysm | -1440\
    hoarseness attributed to compression effects | -1440\
    odynophagia attributed to compression effects | -1440\
    radial artery blood pressures higher on right than left | -1440\
    preoperative diagnosis of left subclavian artery pseudoaneurysm | -1440\
    repair performed through left posterolateral thoracotomy | -1440\
    fourth intercostal space entered | -1440\
    pleural adhesions excised | -1440\
    large mass visible | -1440\
    distal control achieved | -1440\
    aneurysmal sac opened | -1440\
    pseudoaneurysm confirmed | -1440\
    pericardial patch repair of defect | -1440\
    mediastinal lymph nodes sent for histopathology | -1440\
    excised wall sent for histopathology | -1440\
    lymph nodes showed chronic granulomatous inflammation | -1440\
    no necrosis | -1440\
    negative for fungal hyphae | -1440\
    negative for malignancy | -1440\
    excised wall showed completely necrosed tissue | -1440\
    tolerated procedure well | -1440\
    uneventful recovery | -1440\
    discharged within a week | -1440\
    followed for another 2 months | -1440\
    doing well | -1440\
