42 years old | 0
    woman | 0
    Klatskin tumor | 0
    Bismuth type IV | 0
    acute hepatic failure | -72
    listed for emergency liver transplantation | -72
    elevated liver function profile | 0
    aspartate aminotransferase 170 U/L | 0
    alanine aminotransferase 100 U/L | 0
    hemoglobin decreased from 10.4 g/dl to 4.8 g/dl | 0
    platelet count decreased from 103 × 10³/µl to 60 × 10³/µl | 0
    prothrombin time (INR) 2.03 | 0
    activated partial thrombin time 104.5 seconds | 0
    fibrinogen 97 mg/dl | 0
    fibrin degradation product >5 µg/ml | 0
    D-dimer 3.23 µg/ml | 0
    antithrombin III activity 41% | 0
    plasminogen activity 30% | 0
    protein C activity 43% | 0
    metabolic acidosis pH <7.15 | 0
    base deficit >15 mmol/L | 0
    hypocalcemia <0.8 mmol/L | 0
    hyperglycemia >200 mg/dl | 0
    continuous infusion of calcium gluconate 1 mg/kg/hr | 0
    continuous infusion of 5% albumin | 0
    bicarbonate given intermittently | 0
    insulin given intermittently | 0
    exsanguinating bleeding >1,000 ml/hr | 0
    administration of packed red blood cells 25 units | 0
    administration of fresh frozen plasma 16 units | 0
    administration of cryoprecipitate 16 units | 0
    administration of platelet concentrates 16 units | 0
    continuous infusion of dopamine 10 µg/kg/min | 0
    continuous infusion of norepinephrine 0.35 µg/kg/min | 0
    systolic blood pressure maintained 50-80 mmHg | 0
    diastolic blood pressure maintained 30-65 mmHg | 0
    urine output maintained 20