48 years old | 0
male | 0
high grade urothelial carcinoma | -3360
carcinoma in situ | -3360
radical cystectomy | -3360
orthotopic Studer ileal neobladder | -3360
right laparoscopic nephroureterectomy | -672
upper urinary tract urothelial carcinoma | -672
impaired kidney function | 0
serum creatinine: 3.5 mg/dL | 0
no flank pain | 0
no gross hematuria | 0
no fever | 0
clean intermittent self-catheterization (CIC) | 0
urinary catheter placed | 0
kidney failure | 0
serum creatinine: 4 mg/dL | 0
renal ultrasound | 0
severe hydronephrosis | 0
left solitary kidney | 0
computed tomography (CT) scan | 0
smooth-walled stricture of the distal left ureter | 0
severe dilatation of the urinary tract | 0
empty Studer-type neobladder | 0
benign ureteroileal stricture | 0
percutaneous nephrostomy (PN) tube placed | 0
shaking chills | 1
tachycardia | 1
septic shock | 2
anesthesia consulted | 2
hemodynamic support | 2
discharged from ICU | 48
multifactorial acute kidney failure | 48
elevated serum creatinine: 8 mg/dL | 48
massive hematuria | 168
life-threatening bleeding | 168
bleeding through the PN tube | 168
CT angiography | 168
renal pseudoaneurysm | 168
hyperdense material indicative of blood clots | 168
superselective endovascular embolization | 168
Onyx embolization | 168
exclusion of the pseudoaneurysm | 168
hemoglobin level: 12.8 g/dL | 168
hemoglobin level: 7.2 g/dL | 168
transfusion of 2 red blood cells (RBC) units | 168
hemoglobin level: 9 g/dL | 168
clear urine | 168
renal function improved | 168
creatinine: 3 mg/dL | 168