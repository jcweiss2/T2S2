injuring his leg while working on his farm | -72
trismus | -72
hypertonia | -72
admitted to a local hospital | -72
started treatment with immunoglobulins, tetanus vaccination, and metronidazole | -72
transferred to ICU | -48
tracheostomy | -48
mechanical ventilation | -48
vasoactive support | -48
seizures treated with baclofen, midazolam, and diazepam | -48
electroencephalography revealed severely slow cerebral activity | -48
blood cultures and tracheal secretion samples were sent for laboratory analysis | -24
tracheal secretions tested positive for Klebsiella pneumoniae and methicillin-sensitive Staphylococcus aureus | -24
antibiotic therapy with piperacillin-tazobactam was prescribed | -24
transferred to a geriatric unit in a coma | -24
breathed spontaneously on 4 L/min of supplemental oxygen via a tracheal cannula | -24
antibiotic therapy was switched to linezolid | -18
combined treatment with meropenem | -18
septic shock occurred | -18
patient gradually awoke | -12
feeding tube was removed | -12
developed cholestasis and acute edematous pancreatitis | -12
endoscopic treatment got postponed due to spontaneous recovery | -12
urinary tract infection caused by multidrug-resistant organisms | -12
treated with colistin and amoxicillin-clavulanate | -12
transferred to rehabilitation unit | 0
required tracheal supplemental oxygen | 0
required bladder catheter | 0
developed pressure ulcers | 0
sarcopenic and had low handgrip strength | 0
low appendicular skeletal mass | 0
underwent rehabilitation with good compliance | 1
Clostridioides difficile infection occurred | 1
oral vancomycin was prescribed | 1
presented with AF with a third-degree atrioventricular block | 4
transferred to cardiac ICU | 4
underwent single-chamber pacemaker implantation | 4
presented with hyperkinetic delirium | 6
transferred to hospital | 6
Pseudomonas aeruginosa bloodstream infection | 6
treated with ceftazidime-avibactam and amikacin | 6
tested positive for SARS-CoV-2 | 8
treated with remdesivir | 8
placed on droplet isolation | 8
second recurrence of C. difficile | 10
treated with fidaxomicin | 10
bloodstream infection due to Candida parapsilosis, MSSA, and Candida tropicalis | 14
treated with caspofungin and cefazolin | 14
bloodstream infection caused by P. aeruginosa | 24
antibiotic treatment with piperacillin-tazobactam | 24
antibiotic was shifted to aztreonam and ceftazidime-avibactam | 28
antibiotic was shifted to cefepime | 32
tracheostomy closure was performed | 60
discharged from hospital | 120
able to perform postural transition with assistance | 120
motor and respiratory reconditioning continued | 120 
no shortness of breath | -72
denies chest pain | -72