70 years old | 0
female | 0
admitted to the hospital | 0
pancreatic adenocarcinoma | 0
painless jaundice | 0
jaundice | -4320
weight loss | -4320
poor appetite | -4320
open appendectomy | -4320
appendicitis | -4320
open pancreaticoduodenectomy | 0
nasojejunal feeding tube | 0
enteral nutrition commenced | 6
feed rate increased | 24
transferred to surgical ward | 24
high nasogastric output | 24
osmotic laxative prescribed | 24
nausea | 120
vomiting | 120
increasing central abdominal pain | 120
mild tachycardia | 120
central abdominal tenderness | 120
postoperative anastomotic leak | 120
postoperative collection | 120
small bowel obstruction | 120
internal hernia | 120
computed tomography organized | 120
fluid in distal thoracic esophagus | 120
fluid in stomach | 120
nasojejunal feeding tube tip located appropriately | 120
proximal to mid small bowel obstruction | 120
faecalisation | 120
adhesions postulated | 120
small bowel obstruction caused by enteral nutrition solidification | 120
laparotomy performed | 120
small bowel distension | 120
multiple serosal tears | 120
full thickness enterotomy | 120
faecal contamination | 120
feed contamination | 120
decompression of small bowel | 120
extensive washout | 120
enterotomy repair | 120
nasojejunal feeding tube replaced | 120
standard large bore nasogastric tube | 120
central venous catheter placed | 120
total parenteral nutrition commenced | 120
second admission to ICU | 120
inotropic support | 120
worsening acute kidney injury | 120
antifungal treatment added | 120
wound dehiscence | 144
intra-abdominal collection | 144
percutaneous drains inserted | 144
oral intake resumed | 360
nourishing fluids continued | 360
negative-pressure wound therapy | 360
discharged | 888
wound dehiscence required regular dressing changes | 888
no ongoing issues | 888
full diet resumed | 888
