19 years old | 0
male | 0
admitted to the emergency department | 0
motor vehicle accident | -1
conscious | 0
no abnormal symptoms in airways | 0
normal lung examination | 0
blood pressure 130/85 mmHg | 0
pulse rate 130 beats per minute | 0
no free fluid detected in FAST scan | 0
body mass index (BMI) 36.3 | 0
morbid obesity | 0
no tenderness to palpation on spinal column | 0
no symptoms of laceration in chest and abdomen | 0
no abdominal guarding and tenderness | 0
normal perineal and pelvic examinations | 0
normal distal pulses | 0
deformity in distal third of left forearm | 0
left lower extremity crash injury | 0
left leg nearly amputated below the knee | 0
severe muscle and skin damage | 0
nerves and vessels cut | 0
history of committing suicide | -672
psychological disorders | -672
treated with valproate | -672
nasogastric tube (NGT) inserted | 0
foley catheter inserted | 0
normal chest x-ray | 0
normal pelvic radiograph | 0
normal brain computed tomography (CT) scan | 0
limb amputation planned | 0
below knee amputation performed | 2
aggressive soft-tissue debridement performed | 2
serial examinations and hydration performed | 2
NGT pulled out by patient | 4
tachypnea observed | 4
sinus tachycardia with heart rate 150 beats per minute | 4
complaining of upper abdominal pain | 4
NGT reinsertion | 4
pain alleviation | 4
situation improved | 4
eating despite previous lack of appetite | 4
transferred to operating room | 6
suspicion of gastrointestinal bleeding, ischemia, and necrosis | 6
coffee ground secretions detected | 6
midline laparotomy performed | 6
gastric dilation and discoloration detected | 6
gastric decompression performed | 6
external compression of stomach | 6
discoloration disappeared | 6
suspicious areas necessitated further action | 6
transferred to operating room for second laparotomy | 24
total gastrectomy with Roux-en-Y esophagojejunostomy performed | 24
transferred to intensive care unit (ICU) | 24
condition improved over next three days | 48
infection of amputation stump not controlled | 48
above-knee amputation performed | 72
tachypnea with re-elevated heart rate and anuria | 120
leukocytosis detected | 120
elevated creatinine levels | 120
metabolic acidosis detected | 120
blood culture and urine culture performed | 120
bilateral patchy pulmonary infiltrations detected | 120
infectious disease consultation performed | 120
imipenem, ciprofloxacin, and vancomycin administered | 120
hemodialysis performed | 120
contrast study performed using gastrografin | 144
anastomoses found to be normal with no leakage | 144
patient died due to multi-organ failure | 168