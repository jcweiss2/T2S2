78 years old | 0
male | 0
admitted to Intensive Care Unit | 0
urgent surgical repair | 0
stent-grafting endoleak | 0
aortobronchial fistula | 0
thoracic endovascular repair | -43800
descending thoracic aorta aneurysm | -43800
post-operative course uneventful | 0
acute renal failure | 96
elevated inflammatory markers | 96
bacteremia | 96
refractory shock | 96
broad-spectrum antibiotics | 96
no evidence of bleeding | 96
CT-scan | 96
thickened esophageal wall | 96
small gas bubbles near aortic stent graft | 96
aortoesophageal fistula | 96
upper endoscopy | 96
fistula on posterior surface of esophagus | 96
esophageal stenting | 96
covered self-expanding esophageal stent | 96
Ultraflex Esophageal NG | 96
intravenous proton pump inhibitors | 96
parenteral nutrition | 96
broad-spectrum antibiotics | 96
no signs of hemorrhage | 120
no signs of infection | 120
recovered from shock | 120
suspension of amines | 120
ventilator support | 120
died unexpectedly | 504
rupture of aortic arch | 504