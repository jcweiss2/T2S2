66 years old | 0 | 0 
male | 0 | 0 
diabetes mellitus | 0 | 0 
obesity | 0 | 0 
body mass index 25.3 kg/m2 | 0 | 0 
consumed rice wine | 0 | 0 
colonoscopy | -1 | 0 
positive fecal immunochemical test result | -24 | -24 
glycosylated hemoglobin level 9.1% | -24 | -24 
endoscopic mucosal resection | -1 | 0 
hot snare | -1 | 0 
preventive hemoclips | -1 | 0 
resection of 15 polyps | -1 | 0 
polyps in right colon | -1 | 0 
polyps in left colon and rectum | -1 | 0 
discharged from endoscopy room | 0 | 0 
right abdominal pain | 24 | 24 
tenderness | 24 | 24 
rebound tenderness | 24 | 24 
white blood cell count 21460/mm3 | 24 | 24 
C-reactive protein level 17.8 mg/dL | 24 | 24 
blood urea nitrogen level 28 mg/dL | 24 | 24 
creatinine 2.13 mg/dL | 24 | 24 
lactic acid 2.4 mmol/L | 24 | 24 
total bilirubin 1.7 mg/dL | 24 | 24 
abdominopelvic computed tomography | 24 | 24 
multiple air bubbles in right lateral abdominal muscles | 24 | 24 
broad-spectrum antibiotic therapy | 24 | 48 
piperacillin/tazobactam | 24 | 48 
emergency exploratory laparotomy | 44 | 44 
laparoscopic right hemicolectomy | 44 | 44 
multiple-organ failure | 48 | 48 
metabolic acidosis | 48 | 48 
diagnosis of necrotizing fasciitis | 48 | 48 
surgical debridement and drainage | 72 | 72 
renal replacement therapy | 72 | 72 
intensive care unit | 72 | 72 
imipenem-resistant Acinetobacter baumannii | 96 | 96 
extended spectrum beta-lactamase negative Escherichia coli | 96 | 96 
septic shock | 840 | 840 
multiple-organ failure | 840 | 840 
death | 840 | 840