41 years old | 0
female | 0
severe mitral regurgitation | -52560
mitral valve replacement (MVR) with a high profile bioprosthesis size 31 | -52560
echocardiography showed abnormal position of the bioprosthesis strut | -24
narrowing of the left ventricular outflow tract (LVOT) to 1.7 cm | -24
mean systolic gradient of 35 mmHg | -24
left ventricular (LV) cavity was smallish | -24
intraoperatively noted bioprosthesis strut pressing against the posterior wall of the LVOT | 0
redo MVR with a mechanical valve size 29 Carbomedics | 0
posterior MV leaflet resection due to severe calcification | 0
significant bleeding from chest tubes | 10
hemodynamic instability | 10
surgical re-exploration for bleeding | 10
significant amount of bleeding from the area posterior to the aortic valve annulus | 10
cardiopulmonary bypass instituted | 10
aortic cross clamp | 10
cardioplegia | 10
left atrium opened | 10
no problem with new mechanical mitral valve | 10
no tears identified | 10
tear in posterior wall of LVOT below left coronary cusp | 10
tear opposite to intertrigonal area nearer to left fibrous trigone | 10
tear repaired with multiple pledgeted sutures | 10
patient transferred to intensive care unit | 10
died eight days after | 192
sepsis | 192
disseminated intravascular coagulopathy | 192
