71 years old | 0
male | 0
mild abdominal pain | -72
nausea | -72
profuse diarrhea | -72
pain worsened | -24
diarrhea worsened | -24
became unresponsive | -24
hypotensive | 0
tachycardic | 0
severe pain in lower abdomen | 0
tenderness | 0
no fever | 0
no masses | 0
no lymph nodes | 0
metabolic acidosis | 0
serum lactate level over 6 mmol/L | 0
intravenous fluid reanimation | 0
abdominal CT | 0
whole extent of bowel dilated | 0
no free liquid | 0
no air | 0
abdominal pain worsened | 0
distention worsened | 0
surgical consultation | 0
surgery | 0
intestinal ischemia as differential diagnosis | 0
laparotomy | 0
small bowel purplish color | 0
small bowel edema | 0
no perforation | 0
no necrosis | 0
mesentery engorged | 0
mesentery ecchymosis | 0
bowel visible peristalsis | 0
bowel responded to reanimation maneuvers | 0
second-look laparotomy planned | 0
Bogota bag used | 0
low-molecular-weight heparin initiated | 0
transfer to ICU | 0
angio-3D CT reconstruction | 0
no thrombus | 0
no embolus | 0
celiacomesenteric trunk discovered | 0
superior mesenteric artery and celiac trunk from common trunk | 0
second laparotomy | 24
bowel loops normal color | 24
bowel loops regained mobility | 24
never recovered from acidosis | 24
ventilator-associated pneumonia | 24
sepsis | 24
refractory shock | 24
organ failure | 24
death | 24
