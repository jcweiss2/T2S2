49 years old | 0
female | 0
wheelchair-bound | 0
multiple sclerosis | 0
natalizumab | -120
last dose of natalizumab | -120
encephalopathy | 0
breakthrough seizures | 0
hypothermia | 0
hypotension | 0
tachycardia | 0
tachypnea | 0
hypoxia | 0
mechanical ventilation | 0
elevated white blood cell count | 0
hemoglobin of 10.0 g/dL | 0
platelet count of 511,000/uL | 0
urine toxicology screen | 0
sepsis | 0
pneumonia | 0
cefepime | 0
vancomycin | 0
continuous EEG monitoring | 0
no seizure activity | 0
antiepileptic medication dosing adjusted | 0
mental status unchanged | 0
MRI brain with contrast | 24
lumbar puncture | 24
symmetric marked edema | 24
bilateral basal ganglia | 24
mass effect on lateral ventricles | 24
lymphocytic pleocytosis | 24
low CSF glucose | 24
high protein | 24
viral encephalitis | 24
JC virus testing | 24
negative JC virus testing | 24
herpes encephalitis type 2 | 48
intravenous acyclovir | 48
improvement in mental status | 72
discharged to a rehabilitation center | 168
fever | -24
headache | -24
altered mental status | -24
nausea | -24
vomiting | -24
neurological deficits | -24
receptive aphasia | -24
hemiparesis | -24
seizures | -24
status epilepticus | -24
meningeal signs | -24