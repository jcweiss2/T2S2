45 years old | 0
male | 0
farmer | 0
no significant medical history | 0
presented to the emergency department | 0
chest pain | 0
generalized myalgias | 0
exposed to flood waters | -168
fever | -168
flu-like symptoms | -168
symptoms resolved | -48
nonsmoker | 0
denied alcohol use | 0
denied illicit substance use | 0
blood pressure 86/58 mmHg | 0
heart rate 102 bpm | 0
pulse oximetry 94% | 0
random blood glucose 184 mg/dL | 0
temperature 36.4°C | 0
severely icteric | 0
S3 | 0
no murmurs | 0
decreased air entry | 0
occasional scattered crackles bilaterally | 0
mildly distended abdomen | 0
nontender abdomen | 0
alert and oriented | 0
no neurological deficits | 0
mild pitting edema | 0
chest radiography borderline cardiomegaly | 0
mild interstitial edema | 0
sinus rhythm 94 bpm | 0
no acute dynamic changes | 0
resuscitated with intravenous crystalloid | 0
electrolytes repleted | 0
coronavirus rapid antigen test negative | 0
admitted to medical ICU | 0
intravenous piperacillin-tazobactam | 0
tigecycline | 0
routine management for severe sepsis | 0
respiratory failure | 24
severe hypoxemia | 24
high-flow noninvasive ventilation | 24
moderate global hypokinesis | 24
ejection fraction 30-35% | 24
mild-moderate mitral regurgitation | 24
bilateral air-space disease | 24
serologies positive for leptospirosis | 24
AT | 24
AF | 24
VT | 24
defibrillated | 24
amiodarone infusion 0.5 mg/min | 24
clinically unstable | 24
nonischemic cardiomyopathy | 24
myocarditis | 24
septic shock | 24
cardiogenic shock | 24
inotropic supports | 24
multiorgan failure | 24
succumbed to illness | 24
white cell count 19.6 | 0
hemoglobin 13.4 | 0
platelets 67 | 0
serum sodium 132 | 0
serum potassium 4.4 | 0
serum creatinine 4.3 | 0
blood urea nitrogen 81 | 0
serum calcium 9.2 | 0
serum magnesium 0.9 | 0
fasting blood sugar 84 | 0
ALT 73 | 0
AST 34 | 0
alkaline phosphatase 154 | 0
serum albumin 3.2 | 0
INR 1.2 | 0
PT 14.6 | 0
APTT 34 | 0
total bilirubin 15.5 | 0
conjugated bilirubin 11.1 | 0
troponin I 1.2 | 0
creatine kinase 293 | 0
ESR 55 | 0
CRP 42 | 0
blood cultures negative | 0
urine culture negative | 0
HIV nonreactive | 0
QuantiFERON-TB negative | 0
Biofire respiratory panel negative | 0
COVID-19 test negative | 0
leptospirosis IgM positive | 0
hepatitis B surface antigen negative | 0
hepatitis C IgM negative | 0
hepatitis C IgG negative | 0
dengue IgM negative | 0
dengue IgG negative | 0
malaria negative | 0
urine Legionella antigen negative | 0
jaundice | 0
renal failure | 0
hepatic failure | 0
Weil's syndrome | 0
