18 years old | 0
male | 0
admitted to the hospital | 0
COVID-19 | -720
sore throat | -720
loss of sense of smell | -720
positive COVID-19 PCR | -720
mild COVID-19 illness | -720
full recovery | -720
first dose of inactivated SARS-CoV-2 vaccine | -672
asymptomatic | -672
second dose of inactivated SARS-CoV-2 vaccine | -624
headache | -624
fatigue | -624
fever | -624
sore throat | -624
abdominal pain | -624
high-grade fever | -576
myalgia | -576
nausea | -576
vomiting | -576
diarrhea | -576
faint erythematous non-itchy rash | -576
cough | -576
hypotension | 0
tachycardia | 0
temperature of 39°C | 0
systolic blood pressure of 110 mm Hg | 0
tachycardia, 140 beats per minute | 0
fever persisted | 0
generalised erythematous maculopapular rash | 0
conjunctivitis | 0
proteinuria | 0
WBC (15) | 0
Platelet (122) | 0
Creatinine (115) | 0
AST (53) | 0
ALT (81) | 0
Direct bilirubin (35) | 0
Albumin (16) | 0
C reactive protein (249) | 0
Ferritin (4357) | 0
D-dimer (14) | 0
Procalcitonin (9) | 0
Interleukin-6 (90) | 0
ceftriaxone | 0
levofloxacin | 0
intravenous hydrocortisone | 0
haemodynamic stability | 48
haemodynamic instability | 72
facial puffiness | 72
generalised body oedema | 72
myalgia | 72
anasarca | 72
renal impairment | 72
proteinuria | 72
ECG | 72
sinus tachycardia | 72
non-specific T-wave abnormalities | 72
troponin-I (0.29 ng/mL) | 72
pro-BNP (over 8000 pg/mL) | 72
transthoracic echocardiogram | 72
severe tricuspid regurgitation | 72
pulmonary hypertension | 72
PASP (46 mm Hg) | 72
right atrium and ventricle moderately dilated | 72
pericardial effusion | 72
computed topography scan of the chest | 72
bilateral moderate pleural effusion | 72
basal atelectasis | 72
haemodynamic stability | 120
dexamethasone | 120
normal size of the right atrium and ventricle | 120
trace tricuspid regurgitation | 120
normal pulmonary artery systolic pressure | 120
generalised oedema subsided | 144
skin rash and conjunctivitis resolved | 144
white blood cell count normalised | 144
renal function including albuminuria improved | 144
inflammatory markers came down to normal levels | 144
repeat transthoracic echocardiography | 144
trace tricuspid regurgitation | 144
marked improvement in right ventricular systolic function | 144
normal size of the right atrium and ventricle | 144
normal pulmonary artery systolic pressure | 144
dexamethasone was continued for 8 days | 168
switched to oral prednisolone | 168
discharged home | 168
tapering dose of prednisolone | 168
follow-up | 224
symptoms resolved | 224
general weakness and fatigue | 224
repeat echocardiogram was completely normal | 224