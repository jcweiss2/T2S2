61 years old | 0 | 0 
female | 0 | 0 
non-smoking | 0 | 0 
hypertension | 0 | 0 
chronic cough | -504 | 0 
dyspnea | -504 | 0 
weight loss | -504 | 0 
nausea | -168 | 0 
vomiting | -168 | 0 
cachexia | 0 | 0 
scleral icterus | 0 | 0 
jaundice | 0 | 0 
dry mucous membranes | 0 | 0 
normal bowel sounds | 0 | 0 
decreased breath sounds | 0 | 0 
tachycardia | 0 | 0 
hypotension | 0 | 0 
hyponatremia | 0 | 0 
elevated alkaline phosphatase | 0 | 0 
elevated total bilirubin | 0 | 0 
elevated aspartate aminotransferase | 0 | 0 
elevated alanine aminotransferase | 0 | 0 
pulmonary parenchymal nodules | 0 | 0 
lung mass | 0 | 0 
pleural effusion | 0 | 0 
common bile duct dilation | 0 | 0 
gall bladder distension | 0 | 0 
pancreatic head mass | 0 | 0 
biliary obstruction | 0 | 0 
lung biopsy | 24 | 24 
biliary stenting | 24 | 24 
brain metastases | 48 | 48 
radiation therapy | 48 | 168 
chemotherapy | 48 | 168 
carboplatin treatment | 48 | 168 
pemetrexed treatment | 48 | 168 
pembrolizumab treatment | 48 | 168 
whole brain radiation | 72 | 168 
pneumonia | 120 | 168 
sepsis | 168 | 168 
death | 168 | 168