43 years old | 0
male | 0
admitted to the hospital | 0
left facial swelling | -336
swelling and pain in the left hemifacial area | -336
fever | -240
diabetes mellitus | -6720
uncontrolled diabetes | 0
trismus | 0
thinning of the skin with crepitation | 0
septic shock | 24
tachycardia | 24
hypotension | 24
elevated HbA1C level | 0
high white blood cell count | 0
low hemoglobin level | 0
elevated high-sensitivity C-reactive protein level | 0
high glucose level | 0
low sodium level | 0
cytopenia | 48
seizures | 72
metabolic encephalopathy | 72
renal percutaneous catheter drainage | 168
improvement of clinical symptoms | 168
decrease in abscess size | 600
discharge | 672
no further renal abscesses | 1080
decrease in HbA1C level | 1080
no trismus | 2160
no symptoms suggestive of complications | 2160
lung abscesses | 48
renal abscesses | 48
septic emboli | 48
pneumonia | 48
Klebsiella pneumoniae infection | 0
surgical decompression of CNF | 0
intravenous antibiotics | 0
meropenem | 0
levofloxacin | 0
cefotaxime | 72
metronidazole | 144
ceftriaxone | 168
insulin therapy | 0
blood glucose control | 672
albumin level increase | 168
procalcitonin elevation | 72
LRINEC score | 0
air bubbles in soft tissues | 0
gas-forming air bubbles in the fascia | 0
muscle necrosis invasion | 0
contrast-enhanced CT | 0
facial CT | 0
chest CT | 48
abdominopelvic CT | 72
magnetic resonance imaging | 72
electroencephalography | 72