16 years old | 0
female | 0
weighted 60 kg | 0
lost consciousness | -20
CPR | -20
admitted to the Emergency Department | 0
CPR continuously applied | 0
spontaneous circulation not returned | 0
ECPR performed | 60
ECMO successfully established | 120
heparin administered | 120
spontaneous heart rate returned | 180
transferred to ICU | 240
no history of drug allergy | 0
no history of food allergy | 0
body temperature 35°C (rectal) | 0
heart rate 112 bpm | 0
blood pressure 85/52 mm Hg | 0
deep coma | 0
no pupillary reflex | 0
pupillary size 6 mm | 0
no other abnormalities | 0
balanced salt | 0
lansoprazole | 0
meropenem | 0
vancomycin | 0
no urine output | 0
CRRT used | 0
shivering | 24
left lower extremity edema | 24
ultrasonography indicated arterial blood flow reduction | 24
papaverine administered | 24
thermotherapy applied | 24
pupillary reflex resumed | 24
pupils constricted to 3 mm | 24
sedative stopped | 24
analgesic stopped | 24
painful expression | 24
limb expression | 24
left lower extremity swelling worsened | 48
left lower extremity pale | 48
blood flow completely restricted | 48
echocardiography EF 42% | 48
ECMO stopped | 50
blood flow resumed | 50
no urine output | 50
CRRT performed via right internal jugular vein | 50
enteral nutrition started | 72
anti-infective switched to cefoperazone/sulbactam | 168
spontaneous breathing | 216
shallow coma | 216
diminished coughing | 216
percutaneous dilatation tracheostomy performed | 216
ventilator withdrawn | 240
diarrhea developed | 336
light-yellow stools | 336
high fever (40°C) | 336
shock | 336
sputum culture positive for Acinetobacter baumannii | 336
nasogastric feeding replaced by parenteral nutrition | 336
metronidazole | 336
Smecta | 336
tigecycline | 336
tablets of combined Bifidobacterium, Lactobacillus, Enterococcus, Bacillus cereus | 336
body temperature decreased to 38°C | 336
no significant improvement in diarrhea | 336
vancomycin (0.5g every 6 hours) | 384
metronidazole (0.5g every 6 hours) | 384
diarrhea frequency 20-40 times/day | 384
diarrhea volume 3000#4000 mL | 384
bedside colonoscopy suggested PMC | 432
anti-infectives changed to piperacillin/tazobactam | 432
treatment strategy adjusted | 432
dark red diarrhea | 456
hematochezia | 456
poisoning symptoms | 456
first fecal microbiota transplantation (5 U) | 456
diarrhea volume reduced to 1500#2000 mL | 456
second FMT | 480
third FMT | 528
stool color changed to yellow | 528
nasogastric feeding of lactose-free formula milk | 552
diarrhea reduced to 10 times/day | 552
diarrhea volume 1000 mL | 552
fourth FMT | 624
diarrhea improved to 2-4 times/day | 624
diarrhea volume 300#600 mL | 624
total enteral nutrition started | 648
tracheotomy closed | 672
coronary CTA performed | 864
right coronary artery origin at top of sinus | 864
rehabilitation therapy started | 960
discharged | 1800
grade II brain function | 1800
