22 years old | 0
    gravid | 0
    presented to the Emergency Department | 0
    33 weeks of gestation | 0
    dysuria | -168
    febrile | 0
    body temperature 102.7°F (39.3°C) | 0
    tachycardia | 0
    112 beats per minute | 0
    suprapubic tenderness | 0
    left-sided costovertebral angle tenderness | 0
    blood pressure 105/65 mmHg | 0
    obstetric examination normal | 0
    admitted to the hospital | 0
    sepsis | 0
    acute pyelonephritis | 0
    leukocytosis 15.0×10³/mcl | 0
    urinalysis positive for nitrites | 0
    leucocytes esterase positive | 0
    urine squamous cell 4.8/UL | 0
    urine WBC 566.8/UL | 0
    urine bacteria >10000/UL | 0
    urinary tract infection (UTI) | 0
    urine culture positive for Escherichia coli | 0
    renal ultrasound hyperechoic kidneys | 0
    parenchymal disease renal disease | 0
    intravenous (IV) antibiotics (ceftriaxone 1 g/daily) | 0
    intravenous fluid | 0
    blood culture positive for bacteremia with E. coli | 0
    septic shock | 48
    persistent hypotension | 48
    blood pressures 70/40 mmHg | 48
    unresponsive to 4 liters of crystalloids fluids | 48
    hypoxic | 48
    oxygen saturation 70% on 6 L nasal cannula | 48
    diffused crackles | 48
    extremities warm to touch | 48
    creatinine 1.43 mg/dL | 48
    Hb 10 g/dl | 48
    WBC 20×10³/mcl | 48
    lactic acid 9 mmol/L | 48
    intubated | 48
    acute hypoxic respiratory failure | 48
    norepinephrine infusion started | 48
    norepinephrine titration up to maintain MAP ≥65 | 48
    ABG PH 7.41 | 48
    ABG PCO2 33 mmHg | 48
    ABG PO2 60 mmHg | 48
    pressure-controlled ventilation (PRVC) TV 350 | 48
    RR 18 | 48
    FiO2 100 | 48
    PEEP 10 | 48
    peak pressure 36 cmH₂O | 48
    fetal heart tracings reassuring | 48
    chest x-ray bilateral lung consolidation | 48
    mechanical ventilation with FiO2 100 | 48
    hypoxic | 48
    oxygen saturation 70% | 48
    ABG PO2 50 | 48
    PaO2/FiO2 50 | 48
    severe ARDS | 48
    decision to initiate VV ECMO | 48
    pre8-ECMO vital signs blood pressure 103/72 mmHg | 48
    norepinephrine 6 mcg/min | 48
    oxygen saturation 75% | 48
    RR 18 | 48
    body temp 99.3°F | 48
    pulse rate 102 bpm | 48
    right femoral cannula placed | 48
    right internal jugular vein cannula placed | 48
    23F cannula | 48
    19F cannula | 48
    Amplatz wire used | 48
    ECMO cannulation | 48
    ECMO initiation | 48
    fetal distress | 51
    fetal heart deceleration | 51
    emergency cesarean section | 51
    delivery of viable neonate | 51
    newborn admitted to Neonatal Intensive Care Unit | 51
    5000 Units heparin given | 51
    blood loss 100 ml | 51
    anesthesia with fentanyl | 51
    anesthesia with versed drip | 51
    ECMO circuit Maquet Rotaflow centrifugal pump | 51
    ECMO circuit Maquet oxygenator | 51
    broad-spectrum antibiotics (vancomycin 1250 mg every 12 h) | 51
    broad-spectrum antibiotics (cefepime 1 g every 12 h) | 51
    mechanical ventilation FiO2 0.4 | 51
    ECMO pump speed 1500 RPM | 51
    ECMO pump speed increased to 3000 RPM | 51
    ECMO flow rate 4 LPM | 51
    ECMO sweep 5.5 LPM | 51
    oxygen saturation 96% | 51
    monitored for ECMO chatter | 51
    cannula site examined daily | 51
    anticoagulation with heparin bolus 100 IU/kg | 51
    continuous heparin infusion | 51
    target aPTT 40–60 s | 51
    hemoglobin maintained above 10 g/dl | 51
    received 4 units PRBC | 51
    initial ECHO EF 38% | 51
    mild LV dilatation | 51
    moderate global and diffuse LV hypokinesis | 51
    mild RV dilatation | 51
    mild RV dysfunction | 51
    no pericardial effusion | 51
    daily assessment | 51
    weaning off ECMO support | 51
    safely de-cannulated | 120
    extubated | 168
    chest x-ray marked improvement | 168
    repeat ECHO EF 53% | 168
    no hemodynamically significant valve disease | 168
    no wall motion abnormality | 168
    discharged | 312
    no oxygen requirement | 312
    mother in good health | 312
    child in good health | 312
