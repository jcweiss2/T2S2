20 years old | 0
    male | 0
    presented to accident and emergency department | 0
    headache | -720
    severe | -720
    continuous | -720
    exacerbated with exposure to bright light | -720
    photosensitivity | -720
    nausea | -720
    left eye blurred vision | -720
    generalized body fatigue | -720
    symptoms worsening over a month | -720
    denied history of limb weakness | -720
    denied abnormal movements | -720
    denied seizure | -720
    denied loss of consciousness | -720
    denied sensory manifestations | -720
    managed with analgesia | 0
    MRI brain requested | 0
    MRI showed heterogeneously hyperintense lesion on T2-weighted images | 0
    peripheral hypointensity | 0
    optic chiasm compressed | 0
    optic chiasm displaced superiorly | 0
    cavernous sinuses compressed | 0
    internal carotid artery blood flow spared | 0
    T1 images showed fluid level | 0
    conclusion suggestive of macroadenoma | 0
    mass effect on optic chiasm | 0
    pituitary hormonal assessment done | 0
    history of loss of libido | 0
    failure of erection | 0
    polyuria | 0
    polydipsia | 0
    denied gynaecomastia | 0
    denied change in body part size | 0
    central hypogonadism | 0
    central hypoadrenalism | 0
    normal thyroid function | 0
    mildly elevated prolactin | 0
    commenced on hydrocortisone | 0
    no cranial nerve abnormalities | 0
    no limb abnormalities | 0
    no gait abnormalities | 0
    no thyromegaly | 0
    no signs of acromegaly | 0
    chest X-ray normal | 0
    adrenocorticotropic hormone 4.2 pmol/L | 0
    cortisol 101 nmol/L at zero time | 0
    cortisol 430.53 nmol/L at 30 min | 0
    cortisol 529.60 nmol/L at 60 min | 0
    insulin-like growth factor 1 no reagent available | 0
    thyroxine (T4) free 8.0 pmol/L | 0
    thyroid-stimulating hormone 1.88 mIU/L | 0
    follicle-stimulating hormone 0.1 IU/L | 0
    luteinising hormone 0.6 IU/L | 0
    progesterone 1.32 nmol/L | 0
    prolactin 21.69 ng/mL | 0
    testosterone 0.27 nmol/L | 0
    estradiol 49 pmol/L | 0
    urine osmolality 716 mOsm/kg | 0
    plasma sodium 133 mmol/L | 0
    plasma osmolality 283 mOsm/kg | 0
    differential diagnosis pituitary adenoma | 0
    differential diagnosis pituitary abscess | 0
    differential diagnosis pituitary haemorrhage | 0
    scheduled for trans-sphenoidal removal of pituitary macroadenoma | 0
    trans-sphenoidal surgery | 0
    incision in right nostril | 0
    mucosa separated | 0
    sphenoid sinus mucosa removed | 0
    sellar floor identified | 0
    sellar floor removed | 0
    thick capsule incised | 0
    yellowish pus drained | 0
    cavity cleaned | 0
    cavity irrigated with antibiotics | 0
    cavity irrigated with saline | 0
    pus sent for Gram stain | 0
    pus sent for culture | 0
    pus sent for AFB stain | 0
    pus sent for histopathological evaluation | 0
    pituitary not removed | 0
    histopathology showed inflammatory lesion | 0
    no evidence of pituitary adenoma | 0
    Gram stain showed few WBC | 0
    sterile culture | 0
    AFB stain negative | 0
    shifted to intensive care unit | 24
    overnight observation | 24
    transferred to neurosurgery ward | 24
    commenced on metronidazole | 24
    commenced on ceftriaxone | 24
    commenced on vancomycin | 24
    improvement in symptoms | 24
    normal functional status | 24
    pituitary insufficiency continued | 24
    hydrocortisone continued | 24
    no further headaches | 24
    no other symptoms | 24
    follow-up MRI showed no residual abscess | 24
    complete resolution | 24
    <|eot_id|>
