54 years old | 0
female | 0
soft tissue sarcoma | 0
anaemic | 0
haemoglobin 7.5 mg dL−1 | 0
above-knee amputation | 0
peripheral nerve stimulator-guided psoas compartment block | 0
sciatic nerve block | 0
fentanyl injection 50 μg | 0
lateral decubitus position | 0
insulated 100 mm needle introduction | 0
needle directed towards L4 transverse process | 0
patellar movement seen | 0
current reduced | 0
ropivacaine 25 mL 0.5% injection | 0
negative aspiration for blood and CSF | 0
unresponsive | 2
heart rate decreased to 30 beats min−1 | 2
hypotension 60/40 mm Hg | 2
supine position | 2
ventilation with bag and mask | 2
atropine 0.6 mg administration | 2
mephentermine 6 mg administration | 2
Ringer lactate 1 litre administration | 2
blood pressure improvement | 12
intubation with 7.5 cuffed endotracheal | 12
respiration with 100% oxygen | 12
surgery postponed | 12
shift to ICU | 12
haemodynamically stable | 12
regained consciousness | 14
shallow breathing | 14
fully awake with adequate respiratory effort | 16
extubation | 16
dense bilateral sensory block up to T2 level | 16
sensory block disappearance | 22
full recovery | 22
ICU observation | 24
shift to ward | 48