21 years old | 0
female | 0
Caucasian | 0
admitted to the hospital | 0
severe hypoglycemia | 0
altered mental status | 0
lethargic | 0
plasma glucose 20 mg/dl | 0
dextrose infusion | 0
10% dextrose in water | 0
hypoglycemic | 0
capillary glucose 50-60 mg/dl | 0
transferred to facility | 0
suspected insulinoma | 0
childhood diagnosis of GCK gene mutation | -6336
treated with diazoxide | -6336
treated with octreotide | -6336
repeated episodes of seizures | -4320
syncope | -4320
dizziness | -4320
headaches | -4320
palpitations | -4320
sweating | -4320
seizure-free | -4032
syncopal episode | -4032
extensive inpatient hypoglycemia evaluation | -4032
blood glucose 47 mg/dl | -4032
proinsulin levels 10.4-84.1 pmol/l | -4032
C-peptide level 3.1 ng/ml | -4032
negative insulin antibodies | -4032
negative sulfonylurea screen | -4032
magnetic resonance imaging of abdomen | -4032
no insulinoma | -4032
genetic studies revealed Val452 Leu activating mutation of GCK gene | -4032
treated with diazoxide | -4032
discharged home on oral diazoxide 250 mg daily | -4032
discontinued diazoxide due to side effects | -144
hirsutism | -144
fluid retention | -144
dextrose boluses | 0
continuous infusion of 5% dextrose | 0
low blood glucose level | 0
transferred to intensive care unit | 0
octreotide 200 µg subcutaneously twice daily | 24
diazoxide suspension 100 mg three times a day | 24
neuroglycopenic symptoms improved | 24
hypoglycemia improved | 48
capillary glucose 55-110 mg/dl | 48
discharged | 72