60 years old | 0
male | 0
admitted to the hospital | 0
syncope | 0
received second dose of BNT162b2 COVID-19 vaccine | -48
first dose of BNT162b2 COVID-19 vaccine | -72
fever | -48
malaise | -48
decreased urine output | -24
right leg edema | -24
nausea | -24
dizziness | -24
dyspnea on exertion | -24
lost consciousness | 0
awake and alert | 0
blood pressure 97/50 mmHg | 0
pulse rate 114/min | 0
body temperature 36.0°C | 0
respiratory rate 12 breaths/min | 0
percutaneous oxygen saturation 97% | 0
generalized pitting edema in legs | 0
elevated white blood cell count | 0
hemoglobin 22.2 g/dL | 0
serum creatinine 1.51 mg/dL | 0
urine output increased | 24
blood pressure stabilized | 24
hemoconcentration improved | 24
discharged | 120
first episode of SCLS | -8760
second episode of SCLS | -4380
third episode of SCLS | -2880
fourth episode of SCLS | 0
SCLS diagnosis | 0
IgG-κ-type M-proteinemia | -2880
small JAK2 mutations | -2880
started oral terbutaline and theophylline prophylaxis | 120
no further episodes of SCLS | 8760
received common cold-like symptoms | -8760
nausea and vomiting | -8760
pain and swelling in lower extremities | -8760
oliguria | -8760
hypotension | -8760
hemoconcentration | -8760
sepsis of unknown origin | -8760
fluid and antimicrobial therapy | -8760
discharged after 36 days | -8724
cold-like symptoms | -4380
nausea | -4380
oliguria | -4380
swelling in lower extremities | -4380
acute renal failure of unknown origin | -4380
discharged after 4 days | -4376
left leg swelling | -2880
decrease in urine output | -2880
generalized body edema | -2880
dizziness | -2880
dyspnea on exertion | -2880
hypotension | -2880
strong inflammatory response | -2880
kidney dysfunction | -2880
aggressive fluid therapy | -2880
urine output increased | -2876
blood pressure stabilized | -2876
hemoconcentration improved | -2876
discharged after 9 days | -2871
highly sensitive Troponin I | 0
brain natriuretic peptide | 0
soluble interleukin-2 receptor | 0
C4 and C1 elastase inhibitors | 0
blood culture | 0
anti-streptolysin O antibody | 0
antinuclear antibody | 0
anti-glomerular basement membrane antibody | 0
antineutrophil cytoplasmic antibody | 0
rheumatoid factor | 0
SCLS exacerbation | 0
COVID-19 vaccination | -48
BNT162b2 mRNA COVID-19 vaccine | -48
cytokine storms | -48
IL-2 | -48
IL-11 | -48
tumor necrosis factor | -48
nitric oxide | -48
vasodilation | -48
systemic hypotension | -48
capillary-level water loss | -48
cytotoxic effects on endothelial cells | -48
sepsis-like syndromes | -48
hypovolemic shock | -48
multiple organ failure | -48
death | -48
mortality rate of SCLS | -48
14% | -48
IgG-κ-type monoclonal gammopathy of undetermined significance | -2880
MGUS | -2880
oral terbutaline and theophylline prophylaxis | 120
intravenous immunoglobulin | 0
COVID-19 vaccine administration | -48
SCLS flare-ups | 0
Ad26.COV2-S vaccine | 0
mRNA-1273 vaccine | 0
ChAdOx1 nCoV-19 vaccine | 0
UK Medicines and Healthcare Products Regulatory Agency | 0
MHRA | 0
AstraZeneca vaccine | 0
Moderna vaccine | 0
Pfizer-BioNTech vaccine | -48
Janssen vaccine | 0
Oxford-AstraZeneca vaccine | 0
virus-specific CD4+ and CD8+ T cells | -48
immunomodulatory cytokines | -48
antibodies against SARS-CoV-2 | -48
boosting effect | -48
greater release of cytokines | -48
higher rates of adverse reactions | -48
antibody production | -48
second dose of vaccine | -48
first dose of vaccine | -72
SCLS attack | 0
capillary leakage | 0
hypotension | 0
hemoconcentration | 0
systemic involvement | 0
sepsis | -8760
acute renal failure | -4380
multiple organ failure | -48
death | -48
recovery | 120
discharge | 120
follow-up | 8760
no further episodes | 8760
SCLS exacerbation | 0
COVID-19 vaccination | -48
BNT162b2 mRNA COVID-19 vaccine | -48
SCLS diagnosis | 0
IgG-κ-type M-proteinemia | -2880
small JAK2 mutations | -2880
oral terbutaline and theophylline prophylaxis | 120
intravenous immunoglobulin | 0
COVID-19 vaccine administration | -48
SCLS flare-ups | 0
Ad26.COV2-S vaccine | 0
mRNA-1273 vaccine | 0
ChAdOx1 nCoV-19 vaccine | 0
UK Medicines and Healthcare Products Regulatory Agency | 0
MHRA | 0
AstraZeneca vaccine | 0
Moderna vaccine | 0
Pfizer-BioNTech vaccine | -48
Janssen vaccine | 0
Oxford-AstraZeneca vaccine | 0
virus-specific CD4+ and CD8+ T cells | -48
immunomodulatory cytokines | -48
antibodies against SARS-CoV-2 | -48
boosting effect | -48
greater release of cytokines | -48
higher rates of adverse reactions | -48
antibody production | -48
second dose of vaccine | -48
first dose of vaccine | -72
SCLS attack | 0
capillary leakage | 0
hypotension | 0
hemoconcentration | 0
systemic involvement | 0
sepsis | -8760
acute renal failure | -4380
multiple organ failure | -48
death | -48
recovery | 120
discharge | 120
follow-up | 8760
no further episodes | 8760