37 years old | 0
male | 0
cerebral palsy | 0
multiple enterocutaneous fistulas secondary to a perforated appendix | -175200
perforated appendix | -175200
previous right atrial thrombus | -175200
anticoagulation therapy | -175200
presented to the emergency department | 0
increased enteric drainage from enterocutaneous fistula | -168
occasional rigors | -168
waxing and waning subjective fevers | -168
mechanical fall | -168
long-term indwelling peripherally inserted central catheter (PICC) line | -8760
total parenteral nutrition (TPN) | -8760
enterocutaneous fistula healing well | -168
enterocutaneous fistula opened up after fall | -168
increased output requiring ostomy appliance changes | -168
excellent wound care by caregiver | -168
no signs of infection involving enterocutaneous fistula | -168
afebrile | 0
blood pressure 98/60 mmHg | 0
heart rate within normal limits | 0
respiratory rate within normal limits | 0
serum creatinine 1.88 mg/dL | 0
baseline serum creatinine 0.9 mg/dL | 0
no criteria for systemic inflammatory response syndrome | 0
admitted to general medicine unit | 0
increased enterocutaneous fistula drainage | 0
acute kidney injury | 0
elevated whole blood lactate level 3.4 mmol/L | 24
blood culture samples drawn from PICC line | 24
blood culture samples drawn from peripheral site | 24
broad-spectrum intravenous antibiotics | 24
increasing lactate level | 24
cefepime 2000 mg | 24
metronidazole 500 mg | 24
not hypotensive | 24
lactate level increased to 5.5 mmol/L | 25
hypotensive (blood pressure 91/50 mmHg) | 25
increased temperature 39°C | 25
elevated heart rate 120 beats per min | 25
normal respiratory rate | 25
new diagnosis of severe sepsis | 25
intravenous fluids with normal saline | 25
transferred to medical intensive care unit (MICU) | 25
linezolid 600 mg | 25
vasopressor support with norepinephrine | 25
blood cultures grew lactose fermenting gram-negative rods | 48
linezolid discontinued | 48
PICC line removed | 48
TPN through radiologically inserted jejunostomy tube | 48
continued cefepime and metronidazole | 48
blood culture speciation identified >100 CFU/mL of Rahnella aquatilis | 72
resistance to amoxicillin | 72
resistance to cefazolin | 72
susceptibility to numerous other antibiotics | 72
cefepime and metronidazole de-escalated to ceftriaxone 2000 mg | 72
condition stabilized | 72
transferred back to general medicine unit | 72
PICC line replaced | 72
discharged | 240
outpatient antibiotic therapy with ceftriaxone for 10 days | 240
full recovery from Rahnella aquatilis bacteremia | 240
