67 years old | 0
male | 0
mucosal resection for early gastric cancer | -6720
partial resection for left lung cancer | -6720
collected knee-high wild grass from a riverbed | -240
systemic pain | -168
fatigue | -168
fever | -168
chills | -168
watery diarrhea | -168
loss of appetite | -168
mildly disturbed consciousness | -168
decreased white blood cells (WBC) | -14
decreased platelet counts | -14
elevated hepatic enzyme levels | -14
hospitalized | 0
height of 169.0 cm | 0
body weight of 52.3 kg | 0
Glasgow Coma Scale of 14: E3, V5, M6 | 0
blood pressure of 130/79 mmHg | 0
heart rate (HR) of 96/min | 0
respiratory rate (RR) of 20/min | 0
O2 saturation (SPO2) of 94% | 0
temperature of 38.9°C | 0
crusted skin lesions on the medial surface of the left thigh | 0
freely movable adenopathy of approximately 2 cm in size | 0
aggregated papules in the right inguinal region | 0
no remarkable head-and-neck or chest abnormalities | 0
no remarkable neurological abnormalities | 0
blood count was 1,300 /μL WBC | 0
30,000 /μL platelets | 0
neutrophil count was considerably low at 899 /μL | 0
lymphocyte count was 342 /μL | 0
activated partial thromboplastin time (APTT) of 48.2 seconds | 0
C-reactive protein (CRP) levels at 1.3 mg/dL | 0
elevations in concentrations of aspartate aminotransferase (AST) at 230 U/L | 0
lactate dehydrogenase (LDH) at 760 U/L | 0
creatine kinase (CK) at 746 U/L | 0
sepsis | 24
febrile neutropenia (FN) | 24
hemophagocytosis | 24
administered antibiotics | 24
elevated ferritin levels of 15,165 ng/mL | 48
screened closely for potential antibodies specific for cytomegalovirus and Epstein-Barr virus (EBV) | 48
blood culture was negative | 48
bone marrow biopsy | 48
hemophagocytosis with fewer mature myeloid series cells and more monocytoid and lymphoid cells | 48
immunohistological examination revealed a high number of CD3- and CD4-positive T cells | 48
MUM-1-positive lymphoid cells | 48
CD68, CD163-positive histiomonocytes | 48
no EBV-encoded small RNAs (EBERs)-positive cells | 48
diagnosed with HLH | 48
administered prednisolone (PSL) at 60 mg/day | 48
chest pain | 72
shivering | 72
fever of 39.2°C | 72
blood pressure at 88/52 mmHg | 72
HR at 89/min | 72
RR at 24/min | 72
SPO2 at 94% | 72
elevated CK levels at 953 U/L | 72
elevated LDH at 1,405 U/L | 72
high-sensitivity troponin I (TnI) at 271 pg/mL | 72
severe left ventricular dysfunction [left ventricular ejection fraction (LVEF) of 15%] | 72
electrocardiogram (ECG) showed a slight ST elevation in the V1-2 leads | 72
clinically suspected myocarditis | 72
continued respiratory and circulatory management | 72
infection control in the intensive care unit (ICU) | 72
TnI peaked at 82.6 pg/mL | 96
submitted his serum and urine samples and throat swabs to a responsible public health center | 96
moved him to negative-pressure room | 96
reverse transcription polymerase chain reaction (RT-PCR) analysis of the submitted serum detected 1.77×106 SFTSV RNA copies/mL | 120
submitted pathological sections of his bone marrow to the Division of Virology | 120
infected cells that were stained positively by an anti-SFTSV-nucleoprotein (N) antibody | 120
considered steroid pulse therapy for HLH with SFTS | 120
withdrew from circulatory agonist and ventilator management | 336
ECG showed improvement of ST elevation in the V1-2 leads | 336
re-submitted his serum and confirmed negativity for viremia | 408
released him from quarantine | 408
performed CAG and EMB | 576
no coronary artery stenosis was observed on CAG | 576
pathological evaluation of the EMB specimen revealed that the myocardium was mildly hypertrophic | 576
mild myofibrillar loss and disarrangement | 576
active mononuclear cell infiltration adjacent to the damaged myocardium was not observed | 576
immunohistochemistry revealed increases in the number of CD3-positive T cells | 576
CD68-positive macrophages | 576
tenascin-C expression in the stroma | 576
discharged | 696
follow-up visit 1 month after discharge | 744
transthoracic echocardiography showed a slight improvement with an EF of 52.5% | 744
no heart failure | 744