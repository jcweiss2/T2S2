22 years old | 0
female | 0
type 1 diabetes mellitus | -672
poorly controlled | -672
fever | -120
headache | -120
nausea | -120
vomiting | -120
sumatriptan | -72
Ademalog insulin | -672
insulin glargine | -672
lisinopril | -672
purchased 2 cockatiel birds | -4320
admitted to the hospital | 0
confused | 0
aphasic | 0
nuchal rigidity | 0
right upper-extremity paresis | 0
negative Kernig’s sign | 0
negative Brudzinski’s sign | 0
no papilledema | 0
temperature 39.2°C | 0
pulse 123 beats per minute | 0
respiratory rate 22 per minute | 0
blood pressure 131/75 mmHg | 0
oxygen saturation 100% | 0
WBC count 22 K/µL | 0
hemoglobin 13.8 g/dL | 0
sodium 129 mEq/L | 0
potassium 4 mEq/L | 0
chloride 100 mEq/L | 0
bicarbonate 13 mEq/L | 0
blood urea nitrogen 9 mg/dL | 0
creatinine 0.89 mg/dL | 0
initial creatine phosphokinase 275 U/L | 0
lactic acid 2.5 mmol/L | 0
hemoglobin A1c 13.3% | 0
urine toxicology screen negative | 0
sinus tachycardia | 0
vancomycin | 0
ceftriaxone | 0
acyclovir | 0
isotonic fluids | 0
lumbar puncture | 0
cloudy cerebrospinal fluid | 0
WBC count 2790 cells/µL | 0
total protein 163 mg/dL | 0
glucose 31 mg/dL | 0
Listeria monocytogenes | 7
ampicillin | 7
gentamicin | 7
admitted to MICU | 7
diabetic ketoacidosis | 7
point-of-care ultrasound | 24
hyperdynamic left ventricular function | 24
dilated left ventricle | 48
severely reduced ejection fraction | 48
septic shock | 96
acute respiratory failure | 96
seizure | 96
intubation | 96
invasive mechanical ventilation | 96
vasopressor support | 96
intravenous propofol | 96
levetiracetam | 96
no seizure activity | 96
muscle biopsy deferred | 96
received 49 liters of fluids | 240
vasopressor support with norepinephrine | 264
mental status improved | 336
liberated from mechanical ventilation | 336
transferred to internal medicine ward | 432
tachycardic | 456
short of breath | 456
pulmonary embolism | 456
right atrial thrombus | 456
thrombectomy | 480
heparin infusion | 480
discharged to rehabilitation facility | 552
apixaban | 552
levetiracetam | 552
no residual neurological deficits | 552