68 years old | 0
male | 0
Caucasian | 0
admitted to the Emergency Department | 0
chest pain | -2
vomiting | -2
hypertension | -672
hyperuricemia | -672
Mallory-Weiss syndrome | -672
upper gastrointestinal endoscopy | -672
arterial blood pressure 144/78 mmHg | 0
cardiac frequency 108/min | 0
peripheral oxygen saturation 90% | 0
temperature 37,7 °C | 0
decreased respiratory sounds in both inferior pulmonary areas | 0
pulmonary opacity on the left | 0
mild increase in white blood cell count 10.200/mm3 | 0
electrocardiography normal | 0
high sensitivity troponin I normal | 0
myocardial infarction ruled out | 0
intravenous antibiotic started | 0
oxygen started | 0
deteriorated condition | 48
severe chest pain | 48
respiratory distress | 48
type 1 respiratory failure | 48
increase of white blood cell count | 48
increase of c-reactive protein | 48
increase of d-dimer | 48
chest computed tomographic angiography | 48
pneumomediastinum | 48
hydropneumothorax on the left chest | 48
destruction of the lower esophagus | 48
spontaneous rupture of the esophagus | 48
transhiatal esophagectomy | 72
primary anastomosis | 72
left thoracic drainage | 72
esophageal perforation | 72
pleural effusion | 72
nasojejunal tube | 72
intensive care unit | 80
oral swallow X-ray | 144
clear liquid diet | 144
discharged home | 504
oral contrast esophagogram | 720
no anastomotic leak | 720
no stenosis | 720
asymptomatic | 8760