65 years old | 0
    male | 0
    family history of diabetes mellitus | -672
    prostatic hyperplasia | -672
    umbilical hernia repaired | -672
    admitted to the emergency department | 0
    diffuse abdominal pain | -120
    nausea | -120
    vomiting | -120
    abdominal distension | -120
    inability to pass flatus | -24
    inability to evacuate | -24
    tachycardia | 0
    hypotension | 0
    diffuse abdominal tenderness | 0
    peritoneal irritation | 0
    severe distension | 0
    digital rectal examination | 0
    empty rectum | 0
    leukocytosis | 0
    hemoglobin 18.1 g/dL | 0
    platelet count 207 × 10³ | 0
    acute renal failure | 0
    serum creatinine 3 mg/dL | 0
    blood urea nitrogen 60 mg/dL | 0
    urea 210 mg/dL | 0
    dilated loops | 0
    no signs of gas in the rectum | 0
    bowel obstruction | 0
    no free air | 0
    thick and irregular fibrous capsule | 0
    central low-attenuation necrotic component | 0
    surrounding inflammatory changes | 0
    periappendiceal reactive nodal enlargement | 0
    pneumoperitoneum | 0
    dilated large bowel | 0
    enlarged appendix | 0
    perforation at the tip | 0
    preoperative diagnosis of bowel perforation | 0
    peritonitis | 0
    blood pressure not stabilized | 0
    emergency laparotomy | 0
    massive bowel dilatation | 0
    purulent intraperitoneal fluid | 0
    appendiceal tumor 6 cm × 6 cm | 0
    perforated area 1 cm diameter | 0
    appendectomy | 0
    transfer to surgical intensive care unit | 0
    moderate pain | 24
    oral intake reintroduced | 72
    discharged home | 168
    ambulatory clinic follow-up at 1 month | 720
    ambulatory clinic follow-up at 6 months | 4320
    histological examination | 0
    fibroblastic proliferation | 0
    dense inflammatory infiltrate | 0
    thickened submucosa | 0
    myxoid changes | 0
    spindle cells | 0
    polyclonal plasma cells | 0
    lymphocytes | 0
    perforation lined by fibrinoid exudates | 0
    immunohistochemistry positive for vimentin | 0
    immunohistochemistry positive for smooth muscle actin | 0
    immunohistochemistry negative for ALK | 0
    final diagnosis of inflammatory pseudotumor | 0
    appendiceal perforation | 0
    septic shock | 0
    acute abdomen | 0
    visceral perforation | 0
    tumor-like lesion | 0
    postoperative outcome | 0
    normal renal function | 720
    satisfactory evolution | 4320
<|eot_id|>

