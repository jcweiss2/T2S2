41 years old | 0
    female | 0
    G5P4 | 0
    32 weeks pregnant | 0
    admitted to the hospital | 0
    dry cough | -72
    shortness of breath | -72
    headache | -72
    prenatal care | 0
    no diabetes mellitus | 0
    no hypertension | 0
    no bronchial asthma | 0
    no other comorbidities | 0
    BMI 35.6 | 0
    normal blood pressure | 0
    heart rate 99 bpm | 0
    respiratory rate 24 bpm | 0
    oxygen saturations 93–96% on room air | 0
    chest x-ray diffuse bilateral alveolar infiltrates | 0
    sepsis diagnosis | 0
    community acquired pneumonia | 0
    ceftriaxone | 0
    azithromycin | 0
    COVID-19 PCR positive | 0
    oxygenation worsening | 15
    saturations below 90% | 15
    supplemental oxygen 3 L/min | 15
    desaturations | 24
    high flow nasal cannula (HFNC) 40 L flow with 100% FiO2 | 24
    ABG PaO2 111 mmHg | 24
    moderate ARDS | 24
    transferred to ICU | 24
    repeat ABG PaO2 89 mmHg | 31
    severe ARDS | 31
    furosemide 40 mg | 31
    no effect from furosemide | 31
    intravenous dexamethasone | 31
    intubation decision | 31
    placenta previa | 0
    possible accreta | 0
    high risk for complications | 0
    pregnancy not contributing to condition | 0
    no fetal distress | 0
    no vaginal bleeding | 0
    urgent delivery not indicated | 0
    endotracheal intubation | 35
    emergency cesarean section setup | 35
    sevoflurane | 35
    rocuronium | 35
    succinylcholine | 35
    respiratory instability post-intubation | 35
    PEEP 20 cmH2O | 35
    FiO2 100% | 35
    ABG PaO2 59 mmHg | 35
    fentanyl infusion | 35
    midazolam infusion | 35
    repeat ABG PaO2 150 mmHg | 37
    tidal volume 6 mL/kg | 37
    plateau pressure 39 cmH2O | 37
    PEEP decreased to 15 cmH2O | 37
    vaginal bleeding | 38
    emergency cesarean section | 38
    oxytocin | 38
    phenylephrine | 38
    intravenous bicarbonate | 38
    infant delivered limp | 38
    Apgar score 0 | 38
    Apgar score 5 | 38
    Apgar score 7 | 38
    infant intubated | 38
    infant heart rate drop to 60 | 38
    brief compressions | 38
    no maternal intraoperative respiratory complications | 38
    postoperative ICU transfer | 38
    PEEP 15 cmH2O | 38
    FiO2 100% | 38
    ABG PaO2 438 mmHg | 41
    plateau pressure 25 cmH2O | 41
    convalescent plasma | 41
    oxygenation improvement | 48
    PEEP 10 cmH2O | 48
    FiO2 40% | 48
    ABG PaO2 92 mmHg | 48
    ventilator weaning | 96
    liberated from mechanical ventilation | 168
    transferred out of ICU | 168
    oxygen requirements improvement | 216
    transitioned to room air | 216
    no hypoxemia episodes | 216
    hospital course unremarkable | 264
    discharged | 264
    infant COVID PCR negative at 24 hours | 38
    infant COVID PCR negative at 48 hours | 38
    infant extubated | 86
    infant respiratory stability | 86
    no subsequent COVID PCR tests | 86
    placental tissue no abnormalities | 0
    placental tissue not tested for COVID RNA | 0
    