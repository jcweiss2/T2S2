41 years old | 0
male | 0
admitted to the hospital | 0
found unconscious | 0
signs of multiple trauma | 0
respiratory failure | 0
sepsis | 0
hypotension requiring vasopressors | 0
developed massive hematemesis | -192
drop of hemoglobin from 11.4 to 7.3 g/dL | -192
requiring multiple transfusions | -192
initial upper endoscopy | -168
large cratered 15-mm ulcer | -168
visible bleeding vessel | -168
anterior wall of the duodenal bulb | -168
injection of 12 mL of 1:10,000 epinephrine | -168
blanching of the adjacent mucosa | -168
bipolar cautery applied | -168
oozing pigmented spots | -168
successful hemostasis | -168
vasopressor requirements decreased | -156
hemoglobin 8.5 g/dL | -156
became hypotensive again | -144
hemoglobin dropped to 5.8 g/dL | -144
computed tomography angiogram deferred | -144
transferred to interventional radiology | -144
selective arteriograms showed extravasation | -144
right duodenal branch of the gastroduodenal artery | -144
successful coil embolization | -144
remained in critical condition | -144
active bleeding continued | -144
planned emergent salvage surgery | -144
offered salvage repeat endoscopy | -144
repeat endoscopy | -144
new large >2 cm ulcer | -144
spurting vessel (Forrest type 1a) | -144
posterior-inferior portion of the duodenal bulb | -144
injection of 20 mL of 1:10,000 epinephrine | -144
applications of thermocoagulation | -144
hemostasis grasper | -144
oozing from the ulcer | -144
placement of hemostatic clips not attempted | -144
difficult orientation of the ulcer | -144
risk of perforation | -144
further thermocoagulation risk for perforation | -144
oversew the ulcer with endoscopic sutures | -144
OverStitch endoscopic suture system used | -144
one interrupted suture placed | -144
inferior and superior edges of the ulcer | -144
suture cinched to reduce ulcer size | -144
second running suture placed in parallel | -144
closure of the ulcer bed | -144
hemostasis successful | -144
no further bleeding | -144
hemoglobin 8.1 g/dL at discharge | 0
negative Helicobacter pylori serology | 0
discharged to subacute rehabilitation | 0
no further gastrointestinal bleeding | 0
follow-up telephone call a year after | 8760
developed massive hematemesis | 240
drop of hemoglobin from 11.4 to 7.3 g/dL | 240
requiring multiple transfusions | 240
initial upper endoscopy | 240
large cratered 15-mm ulcer | 240
visible bleeding vessel | 240
anterior wall of the duodenal bulb | 240
injection of 12 mL of 1:10,000 epinephrine | 240
blanching of the adjacent mucosa | 240
bipolar cautery applied | 240
oozing pigmented spots | 240
successful hemostasis | 240
vasopressor requirements decreased | 240
hemoglobin 8.5 g/dL | 240
became hypotensive again | 264
hemoglobin dropped to 5.8 g/dL | 264
computed tomography angiogram deferred | 264
transferred to interventional radiology | 264
selective arteriograms showed extravasation | 264
right duodenal branch of the gastroduodenal artery | 264
successful coil embolization | 264
remained in critical condition | 264
active bleeding continued | 264
planned emergent salvage surgery | 264
offered salvage repeat endoscopy | 264
repeat endoscopy | 264
new large >2 cm ulcer | 264
spurting vessel (Forrest type 1a) | 264
posterior-inferior portion of the duodenal bulb | 264
injection of 20 mL of 1:10,000 epinephrine | 264
applications of thermocoagulation | 264
hemostasis grasper | 264
oozing from the ulcer | 264
placement of hemostatic clips not attempted | 264
difficult orientation of the ulcer | 264
risk of perforation | 264
further thermocoagulation risk for perforation | 264
oversew the ulcer with endoscopic sutures | 264
OverStitch endoscopic suture system used | 264
one interrupted suture placed | 264
inferior and superior edges of the ulcer | 264
suture cinched to reduce ulcer size | 264
second running suture placed in parallel | 264
closure of the ulcer bed | 264
hemostasis successful | 264
no further bleeding | 264
hemoglobin 8.1 g/dL at discharge | 360
negative Helicobacter pylori serology | 360
discharged to subacute rehabilitation | 360
no further gastrointestinal bleeding | 360
