66 years old | 0
male | 0
diabetes mellitus | 0
obesity | 0
colonoscopy | 0
fecal immunochemical test result | 0
no history of trauma | 0
no history of surgery | 0
unknown diabetes mellitus | 0
glycosylated hemoglobin level 9.1% | 0
rice wine consumption | 0
colonoscopic polypectomy | 0
endoscopic mucosal resection | 0
hot snare | 0
preventive hemoclips | 0
right colon polyps | 0
left colon polyps | 0
rectum polyps | 0
cecal intubation | 0
excellent bowel preparation | 0
discharged from endoscopy room | 0
right abdominal pain | 24
tenderness | 24
rebound tenderness | 24
white blood cell count 21460/mm3 | 24
C-reactive protein level 17.8 mg/dL | 24
blood urea nitrogen level 28 mg/dL | 24
creatinine 2.13 mg/dL | 24
lactic acid 2.4 mmol/L | 24
total bilirubin 1.7 mg/dL | 24
abdominopelvic CT | 24
no pneumoperitoneum | 24
no bowel perforation | 24
multiple air bubbles in right lateral abdominal muscles | 24
peritonitis excluded | 24
air bubbles in abdominal muscles | 24
intensive medical treatment | 24
piperacillin/tazobactam | 24
emergency exploratory laparotomy | 44
laparoscopic right hemicolectomy | 44
no perforation found | 44
multiple-organ failure | 44
metabolic acidosis | 44
diagnosis of necrotizing fasciitis | 48
surgical debridement | 48
drainage | 48
extensive broad-spectrum antibiotic therapy | 48
renal replacement therapy | 48
two more surgical debridements | 48
drainages | 48
no bacterial growth in blood cultures | 48
imipenem-resistant Acinetobacter baumannii | 48
extended spectrum beta-lactamase negative Escherichia coli | 48
septic shock | 840
death | 840
