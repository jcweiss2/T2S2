37 years old | 0
female | 0
admitted to the hospital | 0
progressive dyspnea | -72
hypoxia | -72
left lung consolidation | -72
shortness of breath | -72
fever | -72
nonproductive cough | -72
Hepatitis C | -672
intravenous heroin abuse | -672
methadone de-addiction program | -672
smoker | -672
malnourished | 0
dehydrated | 0
multiple skin tattoos | 0
burn marks | 0
temperature 38.2°C | 0
respiratory rate 30/Min | 0
blood pressure 90/50 mmHg | 0
pulse rate 120 beats/min | 0
oxygen saturation 95% | 0
heart sounds dual | 0
no crackles or wheezes | 0
air entry reduced | 0
hemoglobin 99 g/L | 0
white cell count 23.7 × 10^9/L | 0
neutrophil count 22.75 × 10^9/L | 0
lymphocytes 0.79 × 10^9/L | 0
CRP 206 mg/L | 0
ALT 26 U/L | 0
AST 18 U/L | 0
urea 3.5 mmol/L | 0
creatinine 42 μmol/L | 0
CXR showed left-sided consolidation | 0
venous access obtained | 0
resuscitated with normal saline | 0
started on ticaricillin/clavulanate | 0
referred to intensive care unit | 0
hypotensive | 12
noradrenalin infusion initiated | 12
intubated | 12
chest CT performed | 12
consolidation of left lobes | 12
no foreign body described | 12
serology drawn | 12
antibiotic regime augmented | 12
vancomycin added | 12
azythromycin added | 12
transthoracic echocardiogram performed | 12
mild tricuspid regurgitation | 12
no vegetations | 12
normal cardiac function | 12
ventilated on SIMV mode | 12
tidal volume 6 mL/kg | 12
PEEP 10 | 12
FiO2 0.5 | 12
minimal endotracheal aspirate | 24
repeat CXR showed persistence of consolidation | 24
flexible bronchoscopy performed | 48
foreign body revealed | 48
foreign body pulled out | 48
foreign body lodged in ETT | 48
ETT removed | 48
reintubated | 48
foreign body examined | 48
identified as 25G hypodermic needle | 48
CXR showed clearing of consolidation | 96
extubated | 96
transferred to medical ward | 96
sputum culture yielded Pseudomonas aeruginosa | 96
antibiotics de-escalated | 96
discharged | 144
inhaled drugs from same table as drug paraphernalia | -72
inadvertently inhaled hypodermic needle | -72