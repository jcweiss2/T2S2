32 years old | 0
female | 0
admitted to the hospital | 0
fever | 0
rash | 0
diarrhea | 0
cough | -840
cephalosporins cefalexin | -840
itchy rash | -672
fever returned and persisted | -672
diagnosed with erythema multiforme | -672
weight-loss capsule "Likeshou" | -17520
antiallergic treatment prednisone | 0
levofloxacin | 0
cefuroxime | 0
yellowish, watery diarrhea | 0
infectious diarrhea | 0
Bifidobacterium | 0
diarrhea persisted | 0
diarrhea worsened | 0
transferred to ICU | 0
MOF (multiple organ dysfunction syndrome) | 0
fever (38.7°C) | 0
percussion tenderness in left lower quadrant | 0
WBC count 9.94×10^9 cells/L | 0
neutrophil count 8.67×10^9 cells/L | 0
CRP 47 mg/L | 0
ESR 37 mm/h | 0
IL-6 80.93 pg/mL | 0
PCT 1.90 ng/mL | 0
HHV-6 negative | 0
EBV DNA elevated | 0
CMV DNA elevated | 0
abdominal CT thickening small intestine and colon walls | 0
hepatosplenomegaly | 0
normal-sized abdominal lymph nodes | 0
early signs of MOF | 0
diagnosed with DIHS | 0
decreased Bifidobacterium, Lactobacillus, Clostridium | 0
antibiotic treatment stopped | 0
FMT once every week | 0
methylprednisolone pulse therapy | 0
immune globulin pulse therapy | 0
ganciclovir | 0
drop in body temperature (38.9°C to 37.3°C) | 168
recurrent MODS symptoms | 168
sterile blood cultures | 168
stool frequency decline | 216
well-formed stools | 216
normal stool frequency and volume | 264
CRP reduced | 168
PCT reduced | 168
ESR reduced | 168
IL-6 reduced | 168
aspartate aminotransferase normal | 264
alanine aminotransferase normal | 264
improved consciousness | 264
EBV DNA normal | 504
CMV DNA normal | 504
normal stool consistency | 264
normal body temperature | 264
discharged | 1440
