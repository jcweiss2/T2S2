Here is the table of events and timestamps:

7 years old | 0
male | 0
referred to the University Children's Hospital Tuebingen | 0
treatment with a monoclonal bi-specific T-cell engager (blinatumomab) | 0
first relapse of pre-B-ALL | -672
allogeneic HSCT from an unrelated HLA-compatible donor | -672
hemoglobin 8.5 g/dl | 0
thrombocytes 13.000/μl | 0
WBC (white blood cells) 940/μl | 0
50/μl neutrophils | 0
CRP (C-reactive protein) 6.83 mg/dl | 0
ferritin 182 μg/dl | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced general condition | 0
cachexia | 0
chronically reduced