76 years old | 0
    man | 0
    history of poorly controlled diabetes | 0
    HA1c 9.2 | 0
    congestive heart failure | 0
    hypertension | 0
    hyperlipidemia | 0
    sore throat | -18
    negative rapid strep test | -18
    prescription for penicillin | -18
    weakness | -12
    unable to walk | -12
    emergency room presentation | 0
    temperature 102.7°F | 0
    pulse 131 | 0
    respiration 40 | 0
    blood pressure 126/73 | 0
    oxygen saturation 96% | 0
    difficulty swallowing | 0
    hoarseness |!0
    cough | 0
    alert | 0
    no cervical lymphadenopathy | 0
    no tenderness | 0
    pharyngeal erythema | 0
    diminished lung sounds at the bases | 0
    flexible fiber optic laryngoscopy | 0
    mild edema | 0
    erythema of bilateral aryepiglottic folds | 0
    involvement of arytenoids | 0
    involvement of false vocal cords | 0
    mild post-cricoid edema | 0
    bilateral lower extremities edema | 0
    Dexamethasone | 0
    vancomycin hydrochloride 1.5g | 0
    ceftazidime 1g | 0
    Clindamycin 600mg | 0
    rapid strep test negative | 0
    lower respiratory culture beta-hemolytic streptococcus group A | 0
    blood culture beta-hemolytic streptococcus group A | 0
    Centor score 2 | 0
    tonsillar exudates | 0
    temperature > 100.4°F | 0
    net score 1 | 0
    antibiotic regimen narrowed to ceftriaxone | 0
    intravenous ceftriaxone 2g every 24 hours | 0
    responded well to antibiotics | 24
    discharged | 168
    short-term rehabilitation unit | 168
    completed treatment without complications | 168