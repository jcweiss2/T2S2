40 years old | 0
male | 0
admitted to the hospital | 0
polytrauma in a road traffic accident | -48
blunt trauma to the chest | -48
right hemothorax | -48
blunt trauma to the abdomen | -48
right lower lobe liver laceration | -48
fractured right tibia | -48
Injury severity scoring (ISS) of 26 | 0
Sequential Organ Failure Assessment (SOFA) score of 12 | 0
Acute Physiology and Chronic Health Evaluation (APACHE II) score of 18 | 0
required intensive critical care | 0
CECT of the chest and abdomen | 0
deranged renal parameters | 0
coagulopathy | 0
progressively became oliguric | 72
anuric | 72
sepsis | 72
multiorgan failure | 72
respiratory failure | 72
renal failure | 72
metabolic disturbance | 72
required intubation | 144
ventilator support | 144
respiratory distress | 144
heparin-free dialysis | 72
heparin-free dialysis | 96
heparin-free dialysis | 144
no blood products transfused | 0
no active bleeding | 0
GCS decreased from 15 to 6 | 144
noncontrast computed tomography head | 144
massive hemorrhage in parieto-occipital region | 144
intraventricular extension | 144
surgical intervention planned | 144
coagulation profile correction planned | 144
expired | 144
hypovolemia | 0
high lactate | 0
contrast induced nephropathy | 0
inadequate hydration | 0
abdominal compartment syndrome | 0
myoglobinuria | 0
massive intracerebral bleed | 144
no attempt to correct coagulopathy | 0
FFPs recommended for coagulation factor deficiencies | 0
microvascular bleeding | 0
elevated prothrombin time | 0
elevated partial thromboplastin time | 0
platelet transfusions recommended | 0
platelet counts <50000/μL | 0
uremia contributes to platelet dysfunction | 0
uremia contributes to coagulopathy | 0
medications tested for bleeding | 0
conjugated estrogens | 0
desmopressin | 0
cryoprecipitate | 0
thromboelastography (TEG) suggested | 0
