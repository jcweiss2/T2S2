40 years old | 0
male | 0
South Asian | 0
admitted to the hospital | 0
sudden altered consciousness | 0
high fever | 0
progressive shortness of breath | -120
no previous history of any chronic illness | 0
no regular medications | 0
no history of drug allergy | 0
febrile | 0
temperature of 39.6°C | 0
heart rate of 140 beats/minute | 0
oxygen saturation (SpO2) of 72% | 0
thin and cachectic | 0
weighed 62 kg | 0
poor nutritional status | 0
mouth ulcers | 0
scrotal swelling | 0
redness | 0
tenderness | 0
Candida mucositis | 0
emergency admission | 0
test for COVID-19 | 0
real-time polymerase chain reaction (rtPCR) | 0
chest Computed Tomography (CT) | 0
screened for HIV | 0
tested negative for HIV | 0
not tested for T-lymphocyte subsets | 0
high flow nasal cannula (HFNC) therapy | 0
anticoagulation | 0
enoxaparin | 0
remdesivir | 0
broad-spectrum antibiotics | 0
tigecycline | 0
levofloxacin | 0
anidulafungin | 0
insulin sliding scale | 0
insulin glargine | 0
electrolytes replenished | 0
magnesium | 0
potassium | 0
COVID-19 real-time rtPCR test came back as positive | 24
left leg swelling | 24
US Doppler study | 24
iliofemoral deep vein thrombosis (DVT) | 24
enoxaparin increased | 24
regained consciousness | 144
improvement in hemodynamic and ventilatory status | 144
fever gradually subsided | 144
hyperglycemia well-controlled | 144
TLC dropped | 144
oxygenation improved | 144
weaned from HFNC | 144
inflammatory markers improved | 144
anti-cytokine therapy not considered | 144
alternating between supine and self-prone positions | 144
clinical deterioration | 168
GCS dropped | 168
oxygen requirement increased | 168
hypotension | 168
norepinephrine infusion | 168
TLC increased | 168
refractory hypoglycemia | 168
dextrose 50% infusion | 168
remdesivir therapy discontinued | 216
chest X-ray showed worsening bilateral infiltrates | 216
sputum culture | 216
Klebsiella pneumoniae | 216
Candida albicans | 216
hospital-acquired pneumonia (HAP) | 216
invasive mechanical ventilation | 216
antibiotics changed | 216
meropenem | 216
linezolid | 216
anidulafungin therapy continued | 216
gradually improved | 240
fever subsided | 240
TLC counts dropped | 240
euglycemia achieved | 240
vasopressors weaned off | 240
oxygen requirements decreased | 240
extubated | 240
HFNC continued | 240
oxygenation deteriorated | 336
re-intubated | 336
oxygen requirement increased | 336
suspected with pulmonary embolism (PE) | 336
CT angiogram | 336
no evidence of PE | 336
HRCT of chest | 336
large cavitary lesions | 336
pleural effusion | 336
necrotizing pneumonia | 336
lung abscess | 336
right-sided pleural drainage | 336
pleural fluid exudate | 336
no bacterial growth | 336
fiberoptic bronchoscopy | 336
bronchoalveolar lavage (BAL) | 336
Candida albicans | 336
anidulafungin continued | 336
antibiotics continued | 336
clinical signs of gradual improvement | 432
extubated | 456
weaned off HFNC | 504
oxygen support | 576
discharged from the hospital | 1344