48 years old | 0
female | 0
shortness of breath | 0
consciousness disturbance | 0
modified radical mastectomy | -5760
chemotherapy | -5760
radiotherapy | -5760
breast reconstruction | -2880
motorcycle accident | -72
dizziness | -72
cold sweating | -72
right anterior chest pain | -72
disturbed consciousness | 0
blood pressure 74/46 mmHg | 0
heart rate 72/min | 0
respiratory rate 22/min | 0
body temperature 36.7 | 0
white blood cell count 17,100/μL | 0
percentage of neutrophilic segments 92.6% | 0
blood gas pH 7.41 | 0
pCO2 38 mmHg | 0
pO2 62 mmHg | 0
HCO3− 24.1 mmol/L | 0
abdomen- and chest-computed tomography | 0
mass lesion with abscess in the right axillary region | 0
percutaneous abscess drainage | 0
septic shock | 0
resuscitation | 0
fever | 24
bacterial culture | 24
PAD culture | 24
oxacillin-sensitive Staphylococcus aureus | 24
oxacillin | 24
redness and swelling in the upper-outer quadrant of the right breast | 216
fasciectomy and debridement | 216
subcutaneous abscess over the right chest wall | 216
granulation tissue material | 216
foreign body | 216
daily wet dressing | 216
debridement and local flap for the defect reconstruction | 432
postoperative course uneventful | 432
2-month follow-up | 1440
acceptable appearance | 1440
retained surgical sponge | -5760
gossypiboma | -5760
aseptic reaction | -5760
adhesion and encapsulation | -5760
granuloma formation | -5760
right chest contusion | -72
rupture of aseptic encapsulation | -72
inflammation | -72
cytokines release | -72
white blood cells accumulation | -72
pus formation | -72
infectious process | -72
septic shock manifestation | 0
local abscess suspicion | 0
PAD performance | 0
gossypiboma consideration | 24
radiopaque marker | 24
whorl-like pattern | 24
air trapped between surgical sponge fibers | 24