50 years old | 0
male | 0
L5 nerve root radiculopathy | 0
conservative management | - hours not specified, assume -72 
nonsteroidal anti-inflammatory drugs | - hours not specified, assume -72 
physiotherapy | - hours not specified, assume -72 
admission to hospital | 0
planned epidural administration of 80 mg of methylprednisolone | 0
injection of 80 mg of methylprednisolone and 2 ml of 2% lignocaine | 0
dilution with 15% KCl instead of 0.9% NS | 0
severe pain in both lower limbs | 0
pruritus | 0
severe cramps | 0
profuse sweating | 0
progressive weakness of both lower limbs | 5
complete flaccid paraplegia below T11 level | 5
absent reflexes below T11 | 5
high blood pressure | 5
heart rate 124 beats per minute | 5
labetalol administration | 5
refractory hypertension | 5
sweating | 5
agitation | 5
electrocardiography showing hyperkalemia | 5
shift to medicine emergency | 5
review of medication error | 5
shift to Intensive Care Unit | 10
supportive measures | 10
calcium gluconate administration | 10
blood samples showing raised potassium levels | 10
potassium chelating agent administration | 10
return of blood pressure and heart rate to normal | 12
return of sensory modalities | 12
development of spasticity | 12
exaggeration of deep tendon reflexes | 12
extensor plantar reflex | 12
neurological recovery | 14
discharge from Intensive Care Unit | 24