60 years old | 0
male | 0
anxiety disorder | -8760
admitted to hospital | 0
increasing fatigue | -96
weakness | -96
cough | -96
shortness of breath | -96
sharp right-sided pleuritic chest pain | -96
right upper quadrant abdominal pain | -96
denies nausea | -96
denies vomiting | -96
febrile | 0
oral temperature of 39.2°C | 0
hemodynamically stable | 0
edentulous | 0
decreased air entry in the right lower and middle lobes | 0
bronchial breath sounds at the right lung base | 0
crepitations over the rest of the right lung | 0
abdomen tender to palpation in the right upper quadrant | 0
elevated total leukocyte count | 0
neutrophil predominance | 0
blood cultures negative | 0
right-sided pneumothorax | 0
right lower lobe consolidation | 0
pleural fluid | 0
chest tube placed | 0
empirical antimicrobial therapy with levofloxacin and metronidazole | 0
pleural fluid submitted to microbiology laboratory | 0
no polymorphonuclear cells or bacteria on Gram stain | 0
aerobic culture did not demonstrate bacterial growth | 0
anaerobic culture recovered large Gram-positive spore-forming bacillus | 48
organism identified as Clostridium bifermentans | 48
antimicrobial susceptibility testing | 48
isolate susceptible to amoxicillin-clavulanate | 48
isolate susceptible to cefoxitin | 48
isolate susceptible to clindamycin | 48
isolate susceptible to meropenem | 48
isolate susceptible to metronidazole | 48
isolate susceptible to penicillin | 48
continued to complain of significant dyspnea | 72
continued to complain of chest pain | 72
CT scan of chest with contrast | 72
right main pulmonary artery embolus | 72
clinically deteriorated | 72
admitted to intensive care unit | 72
antimicrobial therapy changed to piperacillin-tazobactam and levofloxacin | 72
heparin initiated | 72
thoracotomy and decortication of right lung | 360
empyema fluid submitted to microbiology laboratory | 360
C bifermentans recovered on anaerobic culture | 360
antimicrobial therapy with piperacillin-tazobactam alone | 360
intermittent low-grade fevers | 360
ongoing hypoxia | 360
repeat chest radiography | 360
loculated right-sided pneumothorax | 360
small amount of fluid remaining in empyema cavity | 360
second thoracotomy | 1104
right rib resection | 1104
empyema drainage | 1104
lung tissue obtained for aerobic and anaerobic bacterial culture | 1104
lung tissue found to be sterile | 1104
antimicrobial therapy changed to ceftriaxone and metronidazole | 1104
echocardiogram performed | 1104
no evidence of endocarditis | 1104
no valvular pathology | 1104
gradually improved | 1104
discharged home | 1824
prescription for oral metronidazole | 1824