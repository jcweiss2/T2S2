79 years old | 0
male | 0
admitted to the hospital | 0
fever | -48
unproductive cough | -48
dyspnea on exertion | -48
chronic corticosteroid use | -1344
polymyalgia rheumatica | -1344
gardening | -168
fine crackles of the left lower lobe | 0
anemia | 0
elevated C-reactive protein | 0
elevated creatinine | 0
increased white blood cell count | 0
neutrophilia | 0
lymphopenia | 0
negative pneumococcal urinary antigen test | 0
negative legionella urinary antigen test | 0
initiated antibiotic therapy with ceftriaxone | 0
developed highly productive cough | 24
required cough-assist | 24
rapid progressive respiratory failure | 48
impending hemodynamic instability | 48
intubation | 48
bronchoscopy | 48
minimal left side pleural effusion | 48
changed antibiotic treatment to imipenem-cilastatin and clarithromycin | 48
increased prednisone dosage | 48
transferred to ICU | 72
ventilated on pressure-controlled mode | 72
fraction of inspired oxygen 80% | 72
peak airway pressure <30 cm H2O | 72
positive end-expiratory pressure 8-10 cm H2O | 72
hemodynamic support with norepinephrine | 72
chest computer tomography showed airspace consolidation | 72
bilateral infiltrates | 72
transthoracic echocardiography excluded left ventricular dysfunction | 72
mitral and aortic valves appeared normal | 72
bronchoalveolar lavage sample showed neutrophil predominance | 72
replaced clarithromycin with levofloxacin | 120
Legionella longbeachae grew in bronchial sample culture | 120
definitive diagnosis of L. longbeachae community-acquired pneumonia | 120
acute respiratory distress syndrome | 120
septic shock | 120
progressive improvement | 144
new worsening of respiratory parameters | 216
prone positioning | 216
reduced respiratory support | 240
high fever | 312
worsening respiratory parameters | 312
hemodynamic instability | 312
suspected ventilator-associated pneumonia | 312
withheld further support | 312
died | 312