63 years old | 0
female | 0
diagnosed with papillary thyroid carcinoma | -9
treated by resection and radiotherapy | -9
developed stenosis of the esophagus | -9
repeated aspiration | -9
episodes of respiratory insufficiency due to pneumonia and purulent pleurisy | -9
treated by pleurectomy | -9
developed restrictive ventilation pattern | -9
developed recurrent nerve palsy | -9
treated by percutaneous endoscopic gastrostomy and tracheostoma | -9
put on home ventilation | -9
mobility decreased | -9
secondary depression | -9
nearly stopped talking | -9
mandible nearly fixed | -9
could not open mouth over 20 degrees | -9
left axis vertebralis stented | -6
developed stenosis of the internal axis carotis on both sides | -6
diagnosed with arterial hypertension | -6
diagnosed with secondary lactase deficiency | -6
esophageal stenosis dilated | -6
fistula between the esophagus and tracheal membrane | 0
examined by several chiefs and consultants | 0
deemed too unstable for open surgery | 0
referred to the University of Erlangen | 0
suffering from pneumonia by 4-multiresistente gramnegative Pseudomonas aeruginosa | 0
put on veno-venous extracorporeal membrane oxygenation (vv-ECMO) | 0
ventilated through a tracheostoma with low ventilation forces | 0
thoracic computed tomography confirmed a big fistula of the tracheal membrane | 72
decision to try endobronchial stenting | 72
procedure performed | 96
vv-ECMO began to be partly ineffective | 96
high volume input of physiological saline needed | 96
oral approach would only allow a small flexible bronchoscope | 96
approach for the upper part of the trachea had to be performed through the percutaneous tracheostoma in a retrograde manner | 96
tried different Dumon and one-hybrid self-expanding metalic y-stent | 96
changed to a more floppy Freitag stent (FS) | 96
placed a FS 11 cm in length and an inner diameter of 13 mm | 96
regular tracheal cannula was introduced for ventilation | 96
spontaneous breathing work increased | 120
vv-ECMO support was reduced | 120
lungs became re-aerated again | 120
patient woke up again | 120
could communicate with her family by writing and her eyes | 120
infections continued to be very severe | 120
spontaneous work of breathing never exceeded a tidal ventilation of 170 mL per breath | 120
reduction of intravenous saline injection was limited | 120
patient decided actively to reduce the vv-ECMO support | 120
died on 18 November 2016 due to pulmonary infection | 120