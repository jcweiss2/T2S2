There is no event information in the provided text.