61 years old | 0
male | 0
admitted to the hospital | 0
fever | -192
chills | -192
rigor | -192
hiccup | -192
nausea | -48
breathlessness | -24
administered with arteether | -24
hypertension | -9360
cerebrovascular accident (CVA) | -9360
right-sided hemiparesis | -9360
atenolol | -9360
amlodipine | -9360
amiloride | -9360
aspirin | -9360
confused | 0
temperature 104°F | 0
pulse 110/min | 0
blood pressure 130/80 mmHg | 0
respiration rate 40/min | 0
SPO2 96% | 0
pallor | 0
normal blood sugar | 0
normal ultrasonography (USG) of whole abdomen | 0
increased serum urea | 0
increased serum creatinine | 0
increased serum glutamic oxaloacetic transaminase | 0
increased serum glutamic pyruvic transaminase | 0
increased total leukocytic count | 0
negative Plasmodium vivax | 0
negative Plasmodium falciparum | 0
negative Hepatitis C Virus (HCV) | 0
negative Australian antigen | 0
diagnosed as sepsis with ARF | 0
administered with ceftriaxone | 0
administered with tazobactam | 0
continued arteether | 0
no relief in symptoms | 96
increased serum urea | 96
increased serum creatinine | 96
normal urine output | 96
replaced antibiotics with teicoplanin | 120
replaced antibiotics with meropenem | 120
started hemodialysis | 144
symptoms started abating | 168
increased serum urea | 168
increased serum creatinine | 168
increased total leukocytic count | 168
stopped antibiotics | 240
stopped arteether | 240
administered diuretics | 240
administered cefotaxime | 240
increased total leukocytic count | 288
increased serum urea | 288
increased serum creatinine | 288
added tigecycline | 408
added caspofungin | 576
decreased total leukocytic count | 696
added doripenem | 696
stopped antibiotics | 840
diagnosed as CRF | 840
recommended dialysis | 840
stopped torsemide | 984
stopped metolazone | 984
decreased serum urea | 1008
decreased serum creatinine | 1008
stopped furosemide | 1024
decreased serum urea | 1080
decreased serum creatinine | 1080
normal serum urea | 1440
normal serum creatinine | 1440
normal total leukocytic count | 1440
no dialysis required | 1440