67 years old | 0 | 0 
male | 0 | 0 
admitted to the hospital | 0 | 0 
hypertension | 0 | 0 
degenerative joint disease | 0 | 0 
bilateral knee replacement | -6840 | -6840 
substance abuse | 0 | 0 
trauma to face and chest wall | -24 | -24 
lightheadedness | 0 | 0 
fatigue | 0 | 0 
leukocytosis | 0 | 0 
hemoglobin of 10.2 g | 0 | 0 
venous lactic acid of 2.4 mol/l | 0 | 0 
intramuscular and subpectoral hematoma | 0 | 0 
extrapleural extension into the chest | 0 | 0 
acute right second through fifth anterior rib fractures | 0 | 0 
bilateral lower lobe bronchopneumonia | 0 | 0 
blood cultures obtained | 0 | 0 
empiric antibiotics with intravenous piperacillin–tazobactam | 0 | 48 
afebrile | 0 | 48 
hypotensive | 0 | 48 
vasopressors | 0 | 48 
antibiotics broadened to intravenous vancomycin, cefepime and metronidazole | 48 | 96 
repeat blood, urine and sputum cultures obtained | 48 | 48 
sputum cultures grew methicillin-resistant Staphylococcus aureus | 96 | 96 
antibiotics narrowed to intravenous vancomycin | 96 | 120 
left knee pain | 120 | 120 
swelling on physical exam | 120 | 120 
sterile left knee aspiration | 120 | 120 
synovial fluid cloudy, amber colored | 120 | 120 
white blood cells of 9.28 × 103/mcL | 120 | 120 
calcium pyrophosphate crystals | 120 | 120 
complete washout and debridement of the joint | 144 | 144 
operative note described an infected knee with purulence | 144 | 144 
cultures from the infected area obtained | 144 | 144 
antibiotic regimen transitioned to intravenous cefazolin | 168 | 168 
cultures grew C. bifermentans | 240 | 240 
antibiotic regimen transitioned to intravenous ampicillin–sulbactam | 240 | 336 
contrast computerized tomography scan of the abdomen | 240 | 240 
human immunodeficiency virus screening | 240 | 240 
discharged to a rehabilitation facility | 384 | 384 
follow-up with internal medicine | 744 | 744 
recovered full range of motion of left knee | 744 | 744 
no signs of lingering joint or systemic infection | 744 | 744 
taking Augmentin | 744 | 744 
medication adherence | 744 | 744 
had not yet opted to undergo colonoscopy | 744 | 744