66 years old | 0  
    Japanese woman | 0  
    acute onset of fever | -72  
    systemic fatigue | -72  
    confusion | -72  
    restlessness | -72  
    admitted to the emergency department | 0  
    medical history of depression | 0  
    rectal cancer | 0  
    osteoarthritis of the left knee | 0  
    regular medication with amitriptyline | 0  
    trazodone | 0  
    triazolam | 0  
    flunitrazepam | 0  
    duloxetine | 0  
    aripiprazole | 0  
    no illicit drug use | 0  
    no remarkable family history | 0  
    Glasgow Coma Scale E3V4M5 | 0  
    blood pressure 140/86 mmHg | 0  
    heart rate 130 beats/min | 0  
    body temperature 40.4 °C | 0  
    respiratory rate 26/min | 0  
    SpO2 94% | 0  
    costovertebral angle tenderness | 0  
    neurological examinations unremarkable except for confusion | 0  
    elevated C-reactive protein (16.22 mg/dL) | 0  
    elevated creatine kinase (852 U/L) | 0  
    mild elevation in renal function tests | 0  
    blood urea nitrogen 21 mg/dL | 0  
    serum creatinine 1.37 mg/dL | 0  
    complete blood count within normal range | 0  
    urinary test showing pyuria | 0  
    abdominal CT revealing ureteral stone in the right urinary duct | 0  
    swelling of the right kidney | 0  
    blood pressure gradually decreased | 0  
    continuous intravenous noradrenalin at 0.1 μg/kg/min | 0  
    diagnosed septic shock secondary to obstructive pyelonephritis due to urolithiasis | 0  
    meropenem started | 0  
    intraurethral catheter placed in the right urinary duct | 0  
    haloperidol 5 mg administered via intravenous drip for delirium | 0  
    kept in intensive care unit for general management | 0  
    hemodynamics improved on second day | 48  
    noradrenaline administration ended | 48  
    lucid | 48  
    afebrile | 48  
    consciousness worsened again around noon | 48  
    Glasgow Coma Scale E1VTM2 in the evening | 48  
    hyperthermia (bladder temperature exceeding 40 °C) on third day | 72  
    hyperthermia continued for at least 12 hours | 72  
    head and neck examinations showing roving eye movement | 72  
    no neck stiffness | 72  
    no symptoms of meningeal irritation | 72  
    decreased tonus | 72  
    cogwheel rigidity on fifth day | 120  
    clonic spasms of the face and upper extremities | 120  
    creatine kinase elevated to 9,613 U/L on third day | 72  
    creatine kinase peak of 101,475 U/L on seventh day | 168  
    hepatitis virus antigens negative | 0  
    human immunodeficiency virus antigen negative | 0  
    autoantibodies negative | 0  
    vitamins and trace elements normal | 0  
    contrast-enhanced abdominal CT on third day showed improvement in pyelonephritis | 72  
    brain CT on third day showed no abnormal findings | 72  
    lumbar puncture performed on fourth day | 96  
    cerebrospinal fluid showing albuminocytologic dissociation | 96  
    bacterial culture negative | 96  
    herpes virus PCR negative | 96  
    cytomegalovirus antigen negative | 96  
    lumbar punctures performed at 18th and 26th day | 432, 624  
    albuminocytologic dissociation resolved | 624  
    no evidence of infectious disease | 624  
    electroencephalography showing 5–6 Hz theta rhythm | 0  
    no electrographic seizures | 0  
    diagnosis of NMS | 0  
    dantrolene 160 mg/day administered from fourth day | 96  
    bromocriptine 7.5 mg/day administered from fourth day | 96  
    muscle rigidity eased slowly | 96  
    renal replacement therapy introduced on fourth day | 96  
    anuria | 96  
    renal dysfunction | 96  
    hyperthermia improved after renal replacement therapy | 96  
    elevated creatinine kinase levels improved after renal replacement therapy | 96  
    vital signs recovered gradually | 96  
    laboratory data recovered gradually | 96  
    disturbance of consciousness remained | 96  
    tracheostomy performed | 0  
    brain MRI on 10th day showed diffuse hyperintense signal in cerebellar cortex | 240  
    hyperintense signals in cerebellar dentate nucleus, superior cerebellar peduncle, thalamus | 240  
    brain MRI on 27th day showed hyperintense signals in bilateral substantia nigra and globus pallidus | 648  
    MRI at 3 months showed reduced signal intensities in cerebellum and thalamus | 2160  
    basal ganglia lesions disappeared | 2160  
    transferred to another hospital on 149th day | 3576  
    disturbance of consciousness remained | 3576  
    written consent obtained from patient's daughter | 0  
    NMS diagnosis based on haloperidol exposure | 0  
    hyperthermia | 0  
    rigidity | 0  
    altered mental status | 0  
    creatine kinase elevation | 0  
    unstable hemodynamics | 0  
    negative workup for other disorders | 0  
    cerebellar degeneration | 0  
    multi-organ failure | 0  
    neurogenic degeneration in central nervous system | 0  
    prolonged renal dysfunction | 0  
    severe neurologic sequelae remained | 0  
    brain MRI findings improved | 240  
    neurologic prognosis not reflected by MRI | 240  
    no improvement in disturbance of consciousness | 3576  
    declarations | 0  
    funding statement | 0  
    competing interest statement | 0  
    additional information | 0