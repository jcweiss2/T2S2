70 years old | 0
female | 0
admitted to emergency | 0
acute abdominal pain | 0
type II diabetes | -100000
previous splenectomy | -50400
multiple previous laparotomies | -100000
immunocompromised | 0
CT abdomen | 0
perforated splenic flexure malignancy | 0
laparotomy | 2
grossly dilated large bowel | 2
no obvious perforation | 2
loop colostomy | 2
Intravenous Piperacillin/Tazobactam | 2
vancomycin | 4
fluconazole | 4
admitted to intensive care unit | 4
ongoing shock | 4
high vasopressor | 4
noradrenaline requirement | 4
erythematous patch on left thigh | 14
creatine kinase 19 000 | 14
bedside finger test | 14
dirty dishwater fluid | 14
necrotic fat | 14
lack of bleeding | 14
debridement for suspected NF | 16
Meropenem | 16
Lincomycin | 16
disease progression | 26
gas in muscle compartments | 26
gas throughout the whole left leg | 26
non-contiguous area in right gluteal region | 26
diagnosis of multi-focal non-contiguous necrotising myositis | 26
palliated | 30
swab and tissue microscopy | 30
no pathogen isolated | 30