37 years old | 0
male | 0
cerebral palsy | 0
enterocutaneous fistulas | 0
perforated appendix | -7200
right atrial thrombus | -7200
anticoagulation therapy | -7200
increased enteric drainage | -168
rigors | -168
subjective fevers | -168
mechanical fall | -168
indwelling PICC line | -8760
total parenteral nutrition | -8760
admitted to the hospital | 0
afebrile | 0
blood pressure 98/60 mmHg | 0
heart rate within normal limits | 0
respiratory rate within normal limits | 0
serum creatinine 1.88 mg/dL | 0
elevated whole blood lactate level | 24
blood culture samples drawn | 24
broad-spectrum intravenous antibiotics | 24
cefepime 2000 mg | 24
metronidazole 500 mg | 24
increased lactate level | 25
hypotensive | 25
blood pressure 91/50 mmHg | 25
increased temperature 39°C | 25
elevated heart rate 120 beats per min | 25
normal respiratory rate | 25
severe sepsis | 25
i.v. fluids with normal saline | 25
vasopressor support with norepinephrine | 25
transferred to MICU | 25
linezolid 600 mg | 25
lactose fermenting gram-negative rods | 49
PICC line removed | 49
radiologically inserted jejunostomy tube | 49
TPN through jejunostomy tube | 49
Rahnella aquatilis identified | 60
resistance to amoxicillin | 60
resistance to cefazolin | 60
susceptibility to cefepime | 60
susceptibility to ceftriaxone | 60
de-escalated to ceftriaxone | 60
condition stabilized | 72
transferred back to general medicine unit | 72
PICC line replaced | 72
discharged | 120
outpatient antibiotic therapy with ceftriaxone | 120
full recovery | 240