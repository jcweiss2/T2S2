65 years old | 0
ischemic cardiomyopathy | 0
LVAD implantation | 0
HeartWare HVAD | 0
renal insufficiency | 0
peritoneal dialysis | 0
presented in septic state | -8760
high fever | -8760
elevated inflammatory parameters | -8760
C-reactive protein 16 mg/dL | -8760
leukocytes 17G/L | -8760
Staphylococcus aureus identified in blood cultures | -8760
Staphylococcus aureus identified from peritoneal catheter | -8760
status deteriorated rapidly | -8760
serious right ventricular dysfunction | -8760
requiring inotropic support | -8760
admission to intensive care unit | -8760
driveline infection | -8760
massive swelling of subcutaneous tunnel | -8760
clean entrance site | -8760
driveline tunnel surgically opened | -8760
VAC therapy initiated | -8760
peritoneal catheter explanted | -8760
peritonitis proven laparoscopically | -8760
S. aureus identified at surgical site | -8760
antibiotic treatment with vancomycin | -8760
antibiotic treatment with tigecycline | -8760
antibiotic treatment with meropenem | -8760
VAC dressing changed every third day | -8760
swabs returned sterile | -8760
surgical closure of wound | -528
transfer to normal ward | -432
discharged home | 0
readmitted due to recurrence of driveline infection | 2640
wound reopened | 2640
debrided | 2640
negative pressure therapy initiated again | 2640
evaluation of further surgical options | 2640
does not qualify for heart transplantation | 2640
explantation of assist device not an option | 2640
omentum plasty not an option | 2640
change to VAC Veraflo therapy | 2640
0.04% polyhexanide solution instillation | 2640
vacuum treatment for 3 hours | 2640
changes of dressing | 2640
local debridement | 2640
performed in operation room without general anesthesia | 2640
every 3 days | 2640
surgical closure of wound | 2760
postoperative epicutaneous negative pressure wound therapy | 2760
antibiotic treatment with tazobactam/piperacillin | 2760
antibiotic treatment with rifampicin | 2760
discharged after 31 days hospital stay | 3120
remains free from signs of infection for 12 months | 3120
left ventricular function did not recover | -8760
preceding peritonitis | -8760
lack of space for infection to the pump | -8760
transperitoneal infection | -8760
treatment of recurrent driveline infection | 2640
VAC Veraflo therapy with polyhexanide | 2640
no conflict of interest | 3120
