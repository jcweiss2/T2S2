35 years old | 0
female | 0
mentally disabled | 0
psychiatric history of obsessive behavior in childhood | 0
anxiety disorder | 0
atopic dermatitis | -120
corticoid-based therapy | -120
laterocervical lymphadenopathies | -108
night fever | -108
intense sweating | -108
body computed tomography (CT) | -108
supra- and infra-diaphragmatic lymphadenopathies | -108
abdominal masses | -108
biopsy of a lymphadenopathy | -108
NS classic HL | -108
stage IIIB | -108
International Prognostic Score 2 | -108
ABVD chemotherapy regimen | -96
partial response | -72
early relapse | -24
salvage chemotherapy regimen (ESHAP) | -18
no response | -12
GemOx chemotherapy regimen | -6
neutropenia | -6
thrombocytopenia grade 4 | -6
dose-intensity failures | -6
chemotherapy discontinuation | -6
radiotherapy consolidation | -3
HL progressed | 0
IFE regimen | 3
stable disease | 6
watch-and-wait policy | 24
localized areas of progression | 24
radiotherapy | 24
transient partial responses | 24
new mass appeared in D8–D9 | 48
medullar compression syndrome | 48
biopsy | 48
HL relapse | 48
radiotherapy | 48
GemOx | 48
partial response | 54
new progression | 60
watch-and-wait policy | 60
new clinically symptomatic disease progression | 84
bendamustine | 84
disease stability | 90
HL progressed | 108
significant B symptoms | 108
worsening clinical status | 108
celecoxib | 108
lenalidomide | 108
experimental treatment | 108
compassionate use request | 108
unremarkable toxicity | 120
excellent tolerance | 120
CR | 132
interim CT/PET | 132
final CT/PET | 144
celecoxib maintenance | 144
anemia | 168
gastrointestinal bleeding | 168
celecoxib stopped | 168
new disease relapse | 192
CT/PET | 192
supra- and infra-abdominal adenopathies | 192
hepatic and splenic lesions | 192
biopsies | 192
negative | 192
asymptomatic | 192
celecoxib restarted | 192
disease progressed | 198
ascites | 198
paracentesis | 198
biopsies | 198
negative | 198
final biopsy | 204
HL persistence | 204
brentuximab vedotin | 204
intensive care admission | 210
sepsis | 210
fatal outcome | 210