53 years old | 0
female | 0
presented to the hospital with chest pain | 0
family history noncontributory | 0
social history noncontributory | 0
normal sinus rhythm on EKG | 0
no ischemic changes on EKG | 0
chest pain sudden | previous admission timestamp (assuming previous admission was initial presentation, so timestamp for this event would be before current admission. If current admission is timestamp 0, previous admission events would have negative timestamps. However, the text states "on previous admission", which could be days or weeks before. Assuming previous admission was days prior, let's approximate the time between admissions. The patient had "previous admission" with chest pain, then returned after initial discharge. If she was discharged and returned, the time between could be a few days. Assuming she was discharged after initial admission and returned after a week (168 hours), then the previous admission events would be at -168 hours. However, the case states that blood cultures from the previous admission came back positive during this admission, so the previous admission's events are part of the current admission's history. So the initial chest pain, fever, leukocytosis from previous admission would be at -72 hours (assuming 3 days prior). But the text states "on previous admission, the patient had presented with new-onset chest pain... was discharged on cyclobenzaprine and ibuprofen." Then "the patient’s chest pain did not improve, and she returned after the initial admission to the hospital." So the time between initial admission and return is not specified. Since the exact time isn't given, we need to infer. If the initial admission was a week prior (168 hours), then events from the previous admission would be at -168 hours. However, the current admission's blood cultures from the previous admission came back positive, which took time (e.g., 48 hours after administration of antibiotics). The text says "blood cultures from the previous admission came back positive for Staphylococcus aureus." So the previous admission's blood cultures were taken during that admission, which then came back during the current admission. So the events during the previous admission (chest pain, fever, leukocytosis) would be prior to the current admission. To approximate, let's assign the previous admission's events a timestamp of -72 hours (3 days prior). This is a reasonable approximation.)
chest pain constant | -72
chest pain severe | -72
fever | -72
leukocytosis | -72
viral illness diagnosis | -72
costochondritis diagnosis | -72
discharged on cyclobenzaprine | -72
discharged on ibuprofen | -72
chest pain did not improve | 0
returned to hospital | 0
blood cultures positive for Staphylococcus aureus | 0
leukocytosis 19,000 white blood cells per mL | -72
fever 102°F (39°C) | -72
fever trended down | -72
low-grade fever | 0
no leukocytosis | 0
heart rate above 90 beats per minute | 0
respirations over 20 per minute | 0
septic by criteria | 0
Infectious Disease service contacted | 0
repeat blood cultures recommended | 0
antibiotics administered for 48 hours | 0
switched to IV ceftriaxone 2 g daily | 0
switched from IV vancomycin 1,250 mg twice daily | 0
Staphylococcus sensitive to ceftriaxone | 0
Staphylococcus resistant to penicillins | 0
chest pain | 0
mild murmur | 0
bacteremia | 0
endocarditis suspicion | 0
transthoracic echocardiogram performed | 0
normal ejection fraction | 0
trivial regurgitation of valves | 0
mitral valve mild regurgitation | 0
transesophageal echocardiogram not performed | 0
osteomyelitis treatment | 0
possible endocarditis treatment | 0
no gross abnormalities on echocardiogram | 0
urine cultures no growth | 0
urinalysis no growth | 0
urine collected prior to antibiotics | 0
no sputum production | 0
no cough | 0
good dentition | 0
colonoscopy recommended | 0
no melena | 0
no hematochezia | 0
chest X-ray performed | 0
right pleural effusion | 0
right pleural effusion best visualized on lateral projection | 0
no pleural effusion on first chest X-ray | previous admission timestamp (previous X-ray during previous admission, which we assigned as -72 hours)
CT chest without contrast performed | 0
non-displaced fracture of sternum | 0
osteomyelitis of sternum | 0
MRI chest with and without contrast performed | 0
osteomyelitis involving manubrium and upper sternum body | 0
tender to palpation in manubrium and upper sternum | 0
no overlying erythema | 0
chest pain improved during hospital course | 0
IV antibiotics administered | 0
IV ceftriaxone 2 g once daily for 6 weeks | 0
four complete blood count tests | 0
erythrocyte sedimentation rate tests | 0
C-reactive protein tests | 0
basic metabolic panel tests | 0
ibuprofen provided | 0
oxycodone/acetaminophen provided | 0
erythrocyte sedimentation rate 38 mm/hr | 0
erythrocyte sedimentation rate 18 mm/hr | 0
erythrocyte sedimentation rate 15 mm/hr | 0
erythrocyte sedimentation rate 20 mm/hr | 0
C-reactive protein 9.9 mg/L | 0
C-reactive protein 0.3 mg/L | 0
C-reactive protein 0.1 mg/L | 0
C-reactive protein 2.2 mg/L | 0
no recurrence of infection | 0
chest pain persisted in subsequent months | 0
antinuclear antibody 1:320 centromere pattern | 0
rheumatologic disorder suspicion | 0
HIV test performed | 0
hepatitis panel drawn | 0
hepatitis A negative | 0
hepatitis B core antibody negative | 0
hepatitis B surface antigen negative | 0
hepatitis C antibody negative | 0
urinalysis negative | 0
HIV test negative | 0
elevated liver function tests | 0
aspartate aminotransferase 103 U/L | 0
alanine aminotransferase 180 U/L | 0
alkaline phosphatase 135 U/L | 0
aspartate aminotransferase 76 U/L | 0
alanine aminotransferase 144 U/L | 0
alkaline phosphatase 150 U/L | 0
no abdominal pain | 0
no positive hepatitis panel | 0
no complications from medication | 0
tender to palpation without overlying erythema | 0
no evidence of fracture on MRI | 0
bone marrow edema on T2-weighted images | 0
periosteum enhancement of sternum | 0
increased signal in subcutaneous fat | 0
increased signal in anterior mediastinum fat | 0
no abscess found | 0
infection resolved with IV antibiotics | 0
negative hepatitis panel | 0
negative HIV test | 0
elevated liver function tests trended downward | 0
alkaline phosphatase trended upward | 0
no evidence of endocarditis | 0
no surgical correction needed | 0
no cough or sputum | 0
no abdominal pain or melena | 0
no evidence of fracture | 0
chest pain persisted post-treatment | 0
rheumatologic disorder suspected due to ANA | 0
osteomyelitis diagnosis confirmed | 0
primary osteomyelitis without clear cause | 0
no IV drug abuse | 0
no immunocompromised status | 0
no recent central lines | 0
positive ANA in follow-up | 0
possible rheumatologic disorder | 0
no conflicts of interest reported | 0
chest pain sudden | -72
no leukocytosis |==
- 53 years old | 0
