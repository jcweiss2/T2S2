52 years old | 0
male | 0
admitted to the hospital | 0
swelling in left groin | -120
soreness in left groin | -120
antiviral and antipruritic medications | -120
ineffective treatment | -120
abdominal wall and perineal skin defect | 0
necrosis | 0
suppuration | 0
respiratory rate 20 breaths/min | 0
heart rate 125 beats/min | 0
blood pressure 92/77 mmHg | 0
skin defect in abdomen | 0
exposing rectus abdominus muscle | 0
necrotic tissue | 0
purulent discharge | 0
scrotum and penis with black areas | 0
ulcers | 0
defects | 0
erosion | 0
pus | 0
foul odor | 0
diabetes | -672
no previous record of treatment or complications | -672
normal daily insulin intake | -672
high-sensitivity C-reactive protein 244.34 mg/L | 0
white blood cells 8.79 x 10^9/L | 0
fasting blood glucose 7.64 mmol/L | 0
glycated hemoglobin 6.70% | 0
creatinine 185.0 μmol/L | 0
hemoglobin 118.0 g/L | 0
sodium 130.0 mmol/L | 0
modified LRINEC score 36 | 0
CT scan | 0
contrast-enhanced CT scans | 0
extensive infections in lungs and skin | 0
subcutaneous effusion | 0
gas accumulation | 0
wound debridement | 0
full surgical debridement | 144
general anesthesia | 144
type I respiratory failure | 144
ventilatory support | 144
abdominal tissue pathology | 336
necrosis with infection of adipose tissue | 336
infiltration of numerous neutrophils, lymphocytes, and plasma cells | 336
multinucleated giant cells | 336
acid-fast bacilli | 336
Mycobacterium TB proteins | 336
bronchoscopy | 360
alveolar lavage | 360
NGS testing | 360
pathogenic bacteria | 360
multidrug-resistant Escherichia coli | 360
ornidazole | 0
meropenem | 0
fluid rehydration | 0
daily wound care | 0
daily dressing changes | 0
tigecycline | 360
isoniazid | 360
rifampicin | 360
ethambutol | 360
pyrazinamide | 360
discharged | 408
died | 408