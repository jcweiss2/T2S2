39 years old | 0
    female | 0
    admitted for antibiotic treatment of sepsis | 0
    sepsis of unknown origin | 0
    empirically treated with piperacillin-tazobactam | 0
    diagnosed with renal cell carcinoma | -8760
    clear cell histological features | -8760
    left partial nephrectomy | -8760
    recruited to participate in a clinical trial | -2160
    clinical trial investigating hepatic and pancreatic metastasis | -2160
    received interferon | -2160
    received bevacizumab | -2160
    tomography scan taken | -720
    no indication of pulmonary involvement from cancer | -720
    sudden onset of shortness of breath | 0
    tachypnea | 0
    chest discomfort | 0
    no hemodynamic repercussion | 0
    decreased breath sounds in left hemithorax | 0
    tympanic percussion | 0
    trachea deviation to the right | 0
    bilateral jugular stasis | 0
    saturation 91% | 0
    oxygen given at 10-l/min rate through oxygen mask | 0
    thoracocentesis | 0
    air escape in the second intercostal space | 0
    left-sided hydropneumothorax | 0
    contralateral mediastinal shift | 0
    transferred to ICU | 0
    chest discomfort despite drainage | 0
    chest drain | 0
    odorless, turbid brownish fluid from pleural space | 0
    non-invasive mechanical ventilation | 0
    chest discomfort progressively improved | 0
    both lungs expanded | 0
    discharge from ICU | 0
    liquid resembling nasogastric feed emerged from chest drain | 0
    commencing feeding | 0
    output more than 2300 ml per day | 0
    biochemical analysis of pleural effusion | 0
    neutrophilic exudate | 0
    low pH (6.32) | 0
    low protein (1.5 g/dl) | 0
    normal glucose (103 mg/dl) | 0
    high DHL | 0
    high amylase (873 U/l) | 0
    serum amylase 23 U/l | 0
    cytological exam inconclusive | 0
    suspected esophageal perforation | 0
    methylene blue test performed | 0
    positive result | 0
    leakage in chest drain insertion | 0
    computed tomography with oral contrasted medium | 0
    gastropleural fistula | 0
    originated from greater curvature | 0
    extending to left subphrenic space | 0
    submitted to parenteral nutrition | 0
    sudden bleeding exteriorized by chest tube | 48
    sanguineous pleural effusion | 48
    hypovolemic shock | 48
    transferred to ICU again | 48
    received fluid support | 48
    received blood support | 48
    received vasopressor support | 48
    recovered from shock | 48
    upper gastrointestinal endoscopy | 48
    large blood clot in greater curvature | 48
    large blood clot in fundus | 48
    impeded further exploration | 48
    submitted to embolization of splenic arteries | 48
    successful embolization | 48
    no further bleeding episodes | 48
    transferred to palliative care facility | 48
    died | 360
    death due to shock | 360
    death due to acute respiratory insufficiency | 360