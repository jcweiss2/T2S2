45 years old | 0
female | 0
admitted to the hospital | 0
severe mitral stenosis | 0
left atrial clot | 0
shortness of breath | -168
no cerebral symptoms | -168
conscious | 0
alert | 0
oriented | 0
stable vital signs | 0
blood pressure 110/80 mmHg | 0
diastolic murmur | 0
intact cranial nerves | 0
motor power | 0
sensation | 0
no vasculitis | 0
erythrocyte sedimentation rate (ESR) 4 mm | 0
no leukocytosis | 0
white blood cell (WBC) 10.000 mm3 | 0
electrolytes normal | 0
kidney function normal | 0
liver function normal | 0
chest X-ray showed left cardiac border prominence | 0
electrocardiography no change | 0
two-dimensional echocardiography showed large bulky non-mobile thrombosis | 0
mitral valve area 0.6 cm2 | 0
other cardiac valves normal | 0
negative antinuclear antibodies | 0
negative rheumatoid factor | 0
elevation of C4 & C3 components of complement | 0
negative HBS Antigen | 0
open heart surgery | 0
cardiopulmonary bypass | 0
intraoperative findings | 0
stenotic mitral valve excised | 0
clot excised | 0
left atrial cavity irrigated | 0
valve implanted | 0
left ventricle filled with saline and blood | 0
deaired | 0
weaned off cardiopulmonary bypass | 0
inotropic support commenced | 6
dobutamine | 6
adrenaline | 6
blood pressure dropped | 6
central venous pressure elevated | 6
extremity cool and cyanotic | 6
inotropic drugs tapered | 72
blood pressure stabilized | 72
cyanosis changed to gangrene | 72
acral part of extremity amputated | 288
histopathological examination | 288
non-specific vasculitis with thrombosis | 288
quadriplegic | 24
non-voluntary movements | 24
eyes moved only on vertical plane | 24
pupils small and fixed | 24
responded to questions by blinking or moving eyes vertically | 96
brain MRI showed multiple infarction of brainstem | 96
prolonged ventilatory support | 96
tracheostomy | 96
acute renal failure | 96
anemia | 96
kidneys recovered | 96
locked-in state | 96
no neurological improvement | 672
expired from hepatic failure and generalized sepsis | 672