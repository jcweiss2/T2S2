35 years old | 0
male | 0
school teacher | 0
admitted to the hospital | 0
fever | -360
pain in the right thigh | -360
pain in the right shoulder | -360
pain in the right foot | -336
pain in the left foot | -336
pain in the right index finger | -336
pain in the left ring finger | -336
prescribed oral amoxicillin-clavulanate | -336
prescribed paracetamol | -336
neutrophilic leukocytosis | -168
hyperglycemia | -168
ultrasonography of the right mid arm | -168
ultrasonography of the right forearm | -168
ultrasonography of the right thigh | -168
echogenic intramuscular collections | -168
aspiration of pus | -168
Gram-negative microorganisms | -168
prescribed intravenous antibiotics | -168
prescribed subcutaneous insulin therapy | -168
referred to our hospital | -120
respiratory distress | 0
referred to intensive care unit | 0
encephalopathy | 0
septic shock | 0
impending respiratory failure | 0
diffuse warm and tender swellings | 0
intubated | 0
ventilated | 0
vasopressor support | 0
norepinephrine | 0
repeat ultrasound | 0
inflamed muscle membranes | 0
fibrillary pattern of muscle lost | 0
Doppler screen of limbs | 0
no venous thrombosis | 0
two-dimensional-echocardiogram | 0
no infective endocarditis | 0
empirical antimicrobials | 0
meropenem | 0
vancomycin | 0
admission blood cultures | 0
B. cepacia | 0
pancytopenia | 0
hyperferritinemia | 0
hypertriglyceridemia | 0
hepatosplenomegaly | 0
secondary hemophagocytic lymphohistiocytosis | 0
bone marrow examination | 0
hemophagocytosis | 0
growth of B. cepacia | 0
resistant to amikacin | 0
resistant to gentamicin | 0
resistant to piperacillin tazobactam | 0
sensitive to meropenem | 0
sensitive to cotrimoxazole | 0
sensitive to levofloxacin | 0
no granuloma | 0
no necrosis | 0
no fungal elements | 0
cotrimoxazole added to therapy | 0
shock improved | 120
hypoxemia improved | 120
febrile | 0
afebrile | 240
meropenem stopped | 168
vancomycin stopped | 168
cotrimoxazole continued | 168
transferred to ward | 360
discharged home | 360