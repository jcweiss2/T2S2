84 years old | 0
male | 0
admitted to the hospital | 0
edema on both legs | -720
diabetes mellitus | -13140
hypertension | -8760
idiopathic Parkinsons disease | -50400
abdominal ultrasound examination | 0
alcoholic liver cirrhosis | 0
small ascites around the liver | 0
serum albumin concentration 2.5 g/dL | 0
serum bilirubin concentration 2.4 mg/dL | 0
prothrombin time 88% | 0
thrombocytopenia | 0
diabetic chronic renal failure | 0
mild cardiomegaly | 0
brain natriuretic peptide 193 pg/mL | 0
left ventricle ejection fraction 55% | 0
leg edema improved | 48
diuretics administration | 48
albumin administration | 48
dyspnea | 192
tachycardia | 192
tachypnea | 192
hypoxemia | 192
oxygen supplementation | 192
septic shock | 192
endotracheal intubation | 192
hypotension | 216
exacerbated tachycardia | 216
hypothermia | 216
WBC 700/mm3 | 216
Hb 9.7 g/dL | 216
platelet count 59,000/mm3 | 216
BUN/Cr 57/2.2 mg/dL | 216
C-reactive protein 8.3 mg/dL | 216
lactic acid concentration 4.4 mmol/L | 216
urinalysis | 216
urine culture | 216
chest radiograph | 216
piperacillin/tazobactam administration | 216
ciprofloxacin administration | 216
intravenous fluid administration | 216
central venous pressure 12 mmHg | 216
dobutamine administration | 216
dopamine administration | 216
norepinephrine administration | 216
continuous veno-venous hemodialysis | 216
anuria | 216
azotemia | 216
vasopressin administration | 242
skin necrosis | 246
purpura on both wrists and both lower legs | 246
necrotic skin lesions expanded | 250
discontinued vasopressin infusion | 268
Escherichia Coli growth | 268
hemodynamic instability | 268
death | 268