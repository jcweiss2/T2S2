syncope | -12
leg ecchymosis | -12
sepsis due to acute prostatitis | -12
anuria | 0
rhabdomyolysis-induced AKI | 0
increased urea | 0
increased creatinine | 0
increased myoglobin | 0
increased CPK | 0
increased LDH | 0
increased CRP | 0
increased PCT | 0
increased total bilirubin | 0
increased direct bilirubin | 0
increased AST | 0
increased ALT | 0
increased PSA | 0
increased white blood cell count | 0
no hydronephrosis | 0
empty bladder | 0
traces of blood in bladder catheter | 0
no indications to urologic surgery | 0
volume expansion started | 0
diuretic treatment started | 0
antibiotic treatment started | 0
femoral central venous catheter placed | 0
HFR-Supra treatment started | 0
furosemide administered | 0
low molecular weight heparin administered | 0
urea decreased | 96
creatinine decreased | 96
myoglobin decreased | 96
CPK decreased | 96
LDH decreased | 96
CRP decreased | 96
PCT decreased | 96
urine output increased | 96
furosemide tapered | 192
antibiotic therapy switched | 192
HFR-Supra sessions continued | 120
significant reduction in myoglobin | 120
significant reduction in CPK | 120
significant reduction in LDH | 120
significant reduction in CRP | 120
significant reduction in PCT | 120
femoral hemodialysis catheter removed | 168
right jugular central venous catheter placed | 168
on-line hemodiafiltration started | 168
high-flux hemodialysis started | 168
dialysis therapy prolonged | 168
urea decreased | 504
creatinine decreased | 504
CRP decreased | 504
total bilirubin decreased | 504
ASL decreased | 504
ALT decreased | 504
PSA decreased | 504
white blood cells count decreased | 504
urine output increased | 504
dialysis no longer required | 504
urea decreased | 1008
creatinine decreased | 1008
GFR increased | 1008