35 years old | 0
male | 0
admitted to the hospital | 0
coughing | -168
respiratory distress | -24
no fever | -168
no nasal discharge | -168
no chest pain | -168
no hemoptysis | -168
no hematuria | -168
no passage of worms in stool | -168
no atopy | -168
no recent travel | -168
no exposure to pets | -168
no exposure to birds | -168
no exposure to cotton | -168
no exposure to dust | -168
no exposure to metal fumes | -168
pallor | 0
use of accessory muscles of respiration | 0
no lymphadenopathy | 0
no cyanosis | 0
no clubbing | 0
no pedal edema | 0
no palpable purpura | 0
no elevated jugular venous pressure | 0
bilateral rhonchi | 0
bilateral crackles | 0
liver palpable | 0
spleen palpable | 0
normal cardiovascular examination | 0
normal neurological examination | 0
hemoglobin level of 8.3 g/dL | 0
white cell count of 27.6×10^9/L | 0
differential count of 39% polymorphs | 0
differential count of 11% lymphocytes | 0
differential count of 2% monocytes | 0
differential count of 48% eosinophils | 0
absolute eosinophil count of 13.2×10^9/L | 0
platelet count of 420×10^9/L | 0
erythrocyte sedimentation rate of 24 mm/hour | 0
lactate dehydrogenase level of 1,000 U/L | 0
uric acid level of 565 µmol/L | 0
normal renal function | 0
normal liver function | 0
type-1 respiratory failure | 0
pH of 7.38 | 0
partial pressure of oxygen of 67 mmHg | 0
partial pressure of carbon dioxide of 35.5 mmHg | 0
oxygen saturation of 85% | 0
bilateral fluffy alveolar opacities on chest X-ray | 0
normal cardiac size and contour on chest X-ray | 0
confluent symmetrical central airspace opacities on computed tomography | 0
negative troponin I expression | 0
pulmonary capillary wedge pressure of 5 mmHg | 0
normal serum procalcitonin level | 0
sterile blood cultures | 0
negative leptospira serology | 0
negative mycoplasma serology | 0
negative legionella serology | 0
negative filariasis serology | 0
negative strongyloides stercoralis serology | 0
negative legionella urine antigen | 0
negative anti-nuclear antibody | 0
negative anti-neutrophil cytoplasmic antibody | 0
no cysts/ova on stool examination | 0
serum immunoglobulin E level of 708 IU/mL | 0
normal nerve conduction | 0
diethylcarbamazine administration | 0
glucocorticoid administration | 0
no improvement in symptoms | 24
worsening type-1 respiratory failure | 24
bronchoscopy | 24
eosinophil-rich infiltrate on bronchoalveolar lavage | 24
fibroblastic proliferation with formation of Masson bodies on histopathological examination | 24
granulocytic hyperplasia on bone marrow examination | 24
marked increase in eosinophils on bone marrow examination | 24
FIP1L1-PDGFRA mRNA detected | 24
no BCR-ABL1 mRNA detected | 24
myeloid neoplasm associated with eosinophilia and PDGFRA gene rearrangement diagnosis | 24
imatinib administration | 24
marked clinical improvement | 168
marked radiological improvement | 168
marked hematological improvement | 168
complete hematological remission | 336
discharged in stable condition | 336