56 years old| 0
male | 0
admitted to the hospital | 0
external hemorrhoids | -175200
thrombosed external protruding hemorrhoid | 0
severe anal pain | -24
bleeding | -24
hemorrhoidectomy | 0
post-operation day 1 | 24
temperature 36.4 oC | 24
blood pressure 85/50 mmHg | 24
pulse 83 beats per minute | 24
moderate wound pain | 24
mild swelling | 24
no pus or bloody discharge | 24
mefenamic acid 250mg QID PO | 24
pethidine 50mg PRN | 24
post-operation day 2 | 48
pulse 108 beats per minute | 48
blood pressure 76/54 mmHg | 48
no dizziness | 48
no chills | 48
no weakness | 48
no poor appetite | 48
no low urine output | 48
no tarry stool | 48
no epigastric discomfort | 48
post-operation day 3 | 72
fever 38.6 oC | 72
chills | 72
blood pressure 70/42 mmHg | 72
pulse 124 beats per minute | 72
oxygen saturation 97% | 72
leukocytosis 13100/µL | 72
elevated C-reactive protein 33.12 mg/dL | 72
blood urea nitrogen 40.6 mg/dL | 72
creatinine 2.6 mg/dL | 72
decreased platelets 81000/µL | 72
intravenous fluid | 72
cefmetazole 1g Q8H | 72
blood pressure 155/110 mmHg | 74
pulse 88 beats per minute | 74
oxygen saturation 95% | 74
general soreness | 74
discomfort | 74
consciousness change | 78
temperature 36.1 oC | 78
blood pressure 68/51 mmHg | 78
pulse 144 beats per minute | 78
respiratory rate 27 per minute | 78
oxygen saturation 95% | 78
artery blood gas analysis pH 7.32 | 78
pCO2 16.9 mmHg | 78
pO2 118.9 mmHg | 78
HCO3 8.5 mmol/L | 78
intensive care unit admission | 78
endotracheal tube placement | 78
sodium bicarbonate | 78
continuous venous-venous hemofiltration | 78
cardiac arrest | 78
cardiopulmonary resuscitation | 78
extracorporeal membrane oxygenation (ECMO) | 78
no significant swelling | 78
no pus discharge | 78
swab culture from deep wound | 78
second cardiac arrest | 80
expired | 80
Streptococcus pyogenes culture | 80
Streptococcal toxic shock syndrome (STSS) | 80
metabolic acidosis | 78
acute respiratory distress syndrome | 78
renal impairment | 72
coagulopathy | 72
abnormal liver function | 72
septic shock | 72
multiorgan failure | 78
persistent hypotension | 48
leukocytosis | 72
elevated C-reactive protein | 72
blood urea nitrogen elevation | 72
creatinine elevation | 72
decreased platelets | 72
tachypnea | 78
low oxygen saturation | 78
generalized edema | 78
pleural effusion | 78
peritoneal effusion | 78
hypoalbuminemia | 78
soft tissue necrosis | 78
gangrene | 78
skin rash | 78
severe sepsis | 72
stress ulcer induced gastrointestinal bleeding | 48
dehydration | 48
Streptococcus pyogenes induced necrotizing fasciitis | 80
invasive GAS disease | 78
persistent metabolic acidosis | 78
tissue perfusion | 78
life threatening sepsis | 78
fecal impaction | 0
infection | 0
urinary retention | 0
bleeding | 0
anus stenosis | 0
septic complication | 0
Escherichia coli | 0
Bacteroides | 0
necrotizing soft tissue infection | 80
postpartum endometritis | 0
puerperal sepsis | 0
tonsillitis | 0
skin infections | 0
soft tissue infections | 0
toxic shock syndrome (TSS) | 80
invasive group A streptococcal disease | 78
streptococcal TSS | 80
necrotizing fasciitis | 80
myositis | 80
high mortality | 80
morbidity | 80
septic complications | 0
portal of entry for GAS | 0
local sepsis | 78
distant sepsis | 78
predominant organisms Escherichia coli | 0
Bacteroides fragilis | 0
Staphylococcus aureus | 0
Streptococcus pyogenes induced STSS | 80
aggressive intervention | 78
high mortality rate | 80
morbidity rate | 80
catastrophic complications | 0
GAS infection following hemorrhoidectomy | 78
presenting features of STSS | 0
early diagnosis | 78
effective therapeutic drugs | 78
informed consent | 0
conflict of interest | 0
CARE Checklist | 0
peer review | 0
provenance | 0
grade B review | 0
