64 years old | 0
male | 0
Caribbean | 0
admitted to the hospital | 0
diabetes | -672
skin lesions | -168
sepsis | -168
tachycardia | 0
pustules | 0
crusted papules | 0
atrophic cribriform plaques | 0
slit-like ulcerations | 0
axillary lymphadenopathy | 0
jagged red to purplish ulcerations | 0
vancomycin | 0
piperacillin-tazobactam | 0
intravenous fluids | 0
leukocytosis | 0
neutrophilic predominance | 0
elevated inflammatory markers | 0
high sensitivity C-reactive protein | 0
lactate dehydrogenase | 0
mild transaminitis | 0
blood cultures | 0
punch biopsy | 0
bacterial cultures | 0
fungal cultures | 0
viral cultures | 0
ulcerative dermatitis | 0
sub-adjacent neutrophilic infiltrate | 0
pyoderma gangrenosum | 0
prednisone | 24
clobetasol | 24
doxycycline | 24
discharged | 24
biopsy results | 48
intraepidermal vesicular dermatitis | 48
atypical lymphoid infiltrate | 48
CD25 positivity | 48
CD2 positivity | 48
CD3 positivity | 48
CD5 positivity | 48
ALK1 negativity | 48
CD8 negativity | 48
CD20 negativity | 48
CD34 negativity | 48
flow-cytometry | 72
HTLV1/2 levels | 72
autoimmune panel | 72
human immunodeficiency virus | 72
rapid plasma reagin | 72
hepatitis serologies | 72
Quantiferon assay | 72
urine and protein electrophoresis | 72
polyclonal gammopathy | 72
HTLV1/2 serology | 72
elevated interleukin-2 receptor levels | 72
ATLL | 72
altered mental status | 120
severe hypercalcemia | 120
corrected calcium | 120
aggressive hydration | 120
calcitonin | 120
zoledronic acid | 144
hypoxic respiratory failure | 168
disseminated intravascular coagulopathy | 168
emergent intubation | 168
PET/CT scan | 168
organ-system lymphomatous involvement | 168
lungs | 168
spleen | 168
kidneys | 168
diaphragm | 168
scalp | 168
multi-level lymphadenopathy | 168
axillary/chest wall | 168
retroperitoneal | 168
pelvic | 168
cervical chains | 168
goals of care discussion | 192
full comfort care | 192
passed away | 216