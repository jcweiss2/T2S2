68 years old | 0
    female | 0
    hypothyroidism | 0
    bipolar disorder | 0
    sodium valproate | -17520
    clozapine | -17520
    risperidone | -17520
    trihexyphenidyl | -17520
    drowsy | -24
    no limb weakness | -24
    hypothermic | 0
    pulse 50/min | 0
    blood pressure 90/60 mmHg | 0
    respiratory rate 24/min | 0
    bilateral mute plantars | 0
    crepitations over right lower lung fields | 0
    pancytopenia | 0
    normal renal function | 0
    normal liver function | 0
    right lower lobe consolidation | 0
    right middle lobe consolidation | 0
    crystalloids | 0
    antibiotics | 0
    hydrocortisone | 0
    sepsis | 0
    right lower zone pneumonia | 0
    withheld sodium valproate | 0
    withheld clozapine | 0
    withheld risperidone | 0
    withheld trihexyphenidyl | 0
    TSH 22.86 mIU/L | 0
    normal FT4 | 0
    normal FT3 | 0
    anti-thyroid peroxidase antibodies negative | 0
    thyroxine dose escalated to 100 mcg/day | 0
    respiratory distress worsened | 72
    more drowsy | 72
    intubated | 72
    mechanical ventilation | 72
    vasopressors | 72
    sedatives tapered | 168
    infection controlled | 168
    vasopressors stopped | 168
    lethargic | 168
    poor respiratory efforts | 168
    percutaneous tracheostomy | 240
    MRI brain normal | 240
    CSF examination normal | 240
    total creatine kinase levels normal | 240
    electroencephalography normal | 240
    lethargic | 240
    fixed gaze | 240
    limited blinking | 240
    fixed flexor posturing | 240
    increased muscle tone in all limbs | 240
    psychiatry consultation | 240
    provisional diagnosis of catatonia | 240
    lorazepam test performed | 240
    limb rigidity improved | 240
    IV lorazepam 2 mg q8h | 240
    fully conscious | 288
    weaned off ventilator | 576
    neuromuscular power improved | 576
    tracheostomy tube removed | 576
    stoma strapped | 576
    discharged | 840
    