50 years old | 0
male | 0
admitted to the hospital | 0
fever | -120
acute respiratory failure | -120
shortness of breath | -24
dry cough | -24
unremarkable medical history | 0
bilateral multifocal involvement of the lungs | 0
diffuse interstitial pattern | 0
mildly elevated white blood cells | 0
increased C-reactive protein | 0
low procalcitonin | 0
tachypnea | 0
hypotension | 0
tachycardia | 0
diminished vesicular breath sounds | 0
cigarette smoke | -120
unprotected heterosexual intercourse | -120
denies recent travel history | 0
denies close contacts with animals | 0
denies contacts with sick people | 0
denies intravenous drugs use | 0
Pneumocystis jirovecii pneumonia | 0
positive HIV-1 antibody-antigen test | 0
positive pneumococcal urinary antigen | 0
arterial blood gas analysis | 0
severe hypoxemia | 0
empirical therapy with piperacillin-tazobactam | 0
empirical therapy with levofloxacin | 0
empirical therapy with cotrimoxazole | 0
mechanical ventilation | 0
bronchoscopy | 96
Gram stain of bronchoalveolar lavage negative | 96
no bacterial or fungal growth on BAL cultures | 96
no P jirovecii on BAL | 96
cotrimoxazole ceased | 96
no acid-fast bacteria on Ziehl-Neelsen staining | 96
negative Mycobacterium tuberculosis-complex PCR | 96
negative cytomegalovirus | 96
negative Epstein-Barr virus | 96
negative herpes simplex virus 1/2 | 96
negative adenovirus | 96
negative influenza A/B | 96
negative Aspergillus galactomannan antigen | 96
BAL cytology showed macrophages | 96
BAL cytology showed neutrophils | 96
BAL cytology showed lymphocytes | 96
no neoplastic cells on BAL cytology | 96
negative pneumococcal urinary antigen | 96
negative blood cultures | 0
negative Legionella urinary antigen | 0
negative serology for intracellular bacteria | 0
repeated bronchoscopy | 144
repeated Gram stain negative | 144
repeated Ziehl-Neelsen stain negative | 144
no bacterial or fungal growth on repeated BAL cultures | 144
negative Pneumocystis jirovecii IFA | 144
negative PCR-mediated tests for viruses | 144
repeated procalcitonin | 144
no substantial clinical or radiological improvement | 144
persistently febrile | 144
severe respiratory distress | 144
control chest x-rays showed marked interstitial bilateral pattern | 144
control chest x-rays showed acute respiratory distress syndrome radiological signs | 144
confirmatory HIV Western blot | 120
positive HIV Western blot | 120
plasma HIV-ribonucleic acid above 10000000 copies | 120
CD4+ T-cell count 571 cells/mm3 | 120
CD8+ T-cell count 234 cells/mm3 | 120
CD4+/CD8+ ratio 2.44 | 120
previous negative HIV test | -432
HIV-RNA on BAL 206647 cps/mL | 120
antiretroviral treatment introduced | 192
tenofovir disoproxil fumarate/emtricitabine | 192
darunavir/ritonavir | 192
raltegravir | 192
worsening respiratory failure | 192
onset of septic shock | 192
noradrenaline | 192
neutrophilia | 192
increased CRP | 192
positive Klebsiella pneumoniae carbapenemase-producing K. pneumoniae | 192
high-dose meropenem | 216
gentamicin | 216
tygeclicine | 216
negative blood cultures | 192
negative blood cultures | 216
hemodynamically stable | 216
progressive improvement of respiratory distress | 216
radiological improvement on control chest x-rays | 336
extubated | 336
transferred to pneumology ward | 432
transferred to infectious diseases unit | 432
oxygen supply de-escalated | 432
remarkable clinical improvement | 432
follow-up bronchoscopy | 648
BAL cultures still positive for KPC-Kp | 648
HIV-RNA on BAL diminished | 648
antiretroviral treatment well tolerated | 648
complete clinical recovery | 816
discharged | 816
plasma HIV-RNA after 8 weeks of ART decreased | 1344
plasma HIV-RNA after 12 weeks of ART decreased | 2016