67 years old | 0
female | 0
admitted to the hospital | 0
right-sided headaches | -336
visual disturbance | -336
acute confusion | -168
fever | -168
vomiting | -168
photophobia | -168
right-sided radicular leg pain | -168
extreme lethargy | -168
thirst | -168
weight loss | -168
loss of appetite | -168
new onset nocturia | -168
hyponatraemia | -168
primary breast carcinoma | -8760
wide local excision | -8760
post-operative radiotherapy | -8760
adjuvant pharmacological treatment with letrozole | -8760
brain MRI | -336
partly solid, partly cystic suprasellar tumour | -336
compression of the optic apparatus | -336
repeat MRI | -168
progression of the tumour | -168
widespread metastatic lesions in the ventricular system | -168
MRI spine | -168
intradural extramedullary lesion at the level of L1 | -168
equivocal pial nodules of enhancement | -168
lumbar puncture | 672
squamous cells compatible with papillary craniopharyngioma | 672
BRAF V600K mutation | 672
atypical papillary craniopharyngioma | 0
stealth-guided endoscopic resection | 0
CSF cytology | 0
BRAF inhibitors | 672
discharged | not mentioned