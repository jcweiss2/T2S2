87 years old | 0
female | 0
Caucasian | 0
admitted to the hospital | 0
left knee septic arthritis | -96
bilateral conjunctivitis | -96
swelling in hand joint | -96
swelling in first metatarsophalangeal joint of left foot | -96
fevers | -96
episodic altered mental status | -96
denied sore throat | 0
denied dysphagia | 0
denied odynophagia | 0
denied hoarseness | 0
denied other esophageal symptoms | 0
hypertension | 0
paroxysmal atrial fibrillation | 0
diabetes mellitus type I | 0
hypothyroidism | 0
sick sinus syndrome | 0
status post pacemaker placement | 0
total abdominal hysterectomy | 0
multiple caesarean deliveries | 0
cholecystectomy | 0
hernia repair | 0
bilateral conjunctival erythema | 0
mild mucopurulent discharge | 0
irregular heart rhythm | 0
left knee swollen | 0
left knee erythematous | 0
left knee tender | 0
elevated white blood cell count | 0
elevated erythrocyte sedimentation rate | 0
elevated C-reactive protein | 0
transthoracic echocardiography | 0
TEE performed | 0
intravenous sedation with midazolam | 0
pharyngeal local anesthesia with benzocaine | 0
nausea | 1
vomiting | 1
severe chest pain | 1
severe back pain | 1
urgent chest radiography | 1
Gastrografin study | 1
esophageal perforation | 1
contrast seen above gastroesophageal junction | 1
esophagogastroduodenoscopy | 2
mucosal tear | 2
moderate to severe inflammation throughout esophagus | 2
no obvious bleeding | 2
WallFlex stent placement | 2
transferred to intensive care unit | 2
Diflucan started | 2
broad-spectrum antibiotics started | 2
repeat Gastrografin esophagram | 48
no leakage | 48
liquid diet started | 48
respiratory failure | 72
multiorgan failure | 72
palliative care | 120
expired | 168