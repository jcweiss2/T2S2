61 years old | 0
    female | 0
    peripheral arterial disease | 0
    hyperlipidemia | 0
    previous tobacco use | 0
    presented to the emergency department | 0
    midsternal chest pain | -48
    acute occlusion of the right anterior artery | -34560
    right common iliac artery stenting | -34560
    stenting in the right tibial artery | -34560
    stent occluded in the right tibial artery | 0
    unvaccinated for COVID-19 | 0
    no respiratory symptoms | 0
    no nausea | 0
    no vomiting | 0
    admitted to the hospital | 0
    ruled out acute coronary syndrome | 0
    seen by cardiology service | 0
    initial laboratory tests | 0
    troponins | 0
    D-dimer | 0
    results not significant | 0
    normal vitals | 0
    heart rate in the 60s | 0
    COVID-19 antigen test | 0
    COVID-19 PCR test | 0
    both COVID-19 tests positive | 0
    evaluated by infectious disease service | 0
    started on dexamethasone 6 mg IV daily | 0
    started on NMV/r | 0
    risk factors for severe COVID&minus;19 | 0
    medication list reviewed | 0
    apixaban 5 mg oral daily | 0
    atorvastatin 40 mg oral at bedtime | 0
    clopidogrel 75 mg oral daily | 0
    atorvastatin held | 0
    apixaban dose adjusted to 2.5 mg twice daily | 0
    nirmatrelvir 300 mg | 0
    ritonavir 100 mg twice daily | 0
    planned duration of 5 days | 0
    heart rate progressively declined | 0
    sinus bradycardia on telemetry | 0
    heart rate in mid 30s | 0
    NMV/r discontinued | 0
    ECG showing sinus bradycardia | 0
    no contributing medications | 0
    denied chest pain | 0
    denied headache | 0
    denied dizziness | 0
    denied blurry vision | 0
    electrolytes within normal limits | 0
    administered atropine 0.5 mg IV twice | 0
    placed on transcutaneous pacer | 0
    transferred to ICU | 0
    blood pressure 90/45 mmHg | 0
    heart rate 33 bpm | 0
    MAP 60 | 0
    dobutamine drip started | 0
    dobutamine titrated up to 5 µg/kg/min | 0
    palpitations | 0
    drip titrated back down | 0
    dobutamine discontinued after 10 hours | 0
    terbutaline tablet 5 mg ordered | 0
    terbutaline discontinued | 0
    no hypoxemia | 0
    no elevated inflammatory markers | 0
    low cortisol levels | 0
    appropriate cosyntropin stimulation tests | 0
    MRI of the brain | 0
    MRI negative | 0
    remained asymptomatic from COVID-19 | 0
    medication-induced bradycardia | 0
    discharged | 0
    