17 years old | 0
girl | 0
admitted to the hospital | 0
headache | -720
occupying lesion located in bilateral and third ventricles | 0
neuronavigation-assisted IVT tumor excision | 0
external ventricular drainage | 0
perioperative i.v. antibiotic prophylaxis with cefazolin | 0
vancomycin | -24
ceftriaxone | -144
marked leucocytosis | -24
abnormal laboratory examination of CSF | -24
fever | -48
body temperature 38.4°C | -48
nausea | -48
emesis | -48
apathy | -48
CSF cultures showed carbapenem-resistant Enterobacter cloacae infection | -12
blood culture positive | -12
removed drainage tube of external ventricular | -12
catheter cultured | -12
tigecycline i.v. | -12
amikacin i.v. | -12
cardiac arrest | -12
respiratory arrest | -12
herniation of the brain | -12
placed another EVD | -12
adjusted antibiotics | 0
meropenem i.v. | 0
cotrimoxazole | 0
allergic to cotrimoxazole | 0
fever persisted | 0
highest temperature 38.8°C | 0
state of consciousness deteriorated into lethargy | 0
CSF cultures still showed carbapenem-resistant Enterobacter cloacae infection | 0
IVT amikacin | 24
elevated WBC count in CSF | 72
CSF culture persistently positive | 72
EVD on left side | 192
EVD on right side | 264
CSF culture negative | 408
IVT amikacin discontinued | 432
ventricular drainages removed | 480
CSF culture continuously negative | 624
stopped meropenem | 624
stopped amikacin | 624
mental status improved | 624
fever subsided | 624
meningitis effectively treated | 624
no nephrotoxicity | 624
no seizures | 624
no focal deficits | 624
central neurocytoma confirmed | 624
transferred to receive radiotherapy | 624
third ventriculostomy | 624
septostomy of the septum pellucidum | 624
obstructive hydrocephalus | 624
full recovery | 624
normal life | 624
