70 years old | 0
male | 0
laboratory-confirmed diagnosis of COVID-19 | -72
respiratory symptoms (dyspnea, tachypnea) | 0
dyspnea | 0
tachypnea | 0
PaO2 68.2 mmHg | 0
FiO2 0.4 | 0
transferred to ICU | 0
dyspnea worsened | 0
PaO2 60.5 mmHg | 0
FiO2 0.9 | 0
intubation | 480
ventilator for 8 days | 480
extubation | 672
unable to breathe properly | 720
re-intubation | 720
planned tracheostomy | 768
preoperative chest X-ray | 768
reposition ET tube balloon below second tracheal ring | 768
confirm balloon position with X-ray | 768
thrombocytopenia | 0
septic shock | 0
platelet transfusion | 768
surgical tracheostomy | 768
FiO2 lowered to=0.4 | 768
balloon overinflated | 768
ET tube withdrawal | 768
transparent film dressing applied | 768
tracheostomy tube insertion | 768
check tracheostomy tube patency | 768
ventilator connected | 768
ET tube removed | 768
oxygen saturation maintained above 98% | 768
medical staff asymptomatic after 14 days | 768 + (14 × 24) = 768 + 336 = 1104
discharged | 2520
