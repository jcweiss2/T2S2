59 years old | 0
female | 0
blood type O | 0
Rh positive | 0
admitted to the hospital | 0
segment-V space-occupying lesion | -365
liver cancer | -365
transarterial embolization | -365
sorafenib | -304
dizziness | -91
skin ulcers | -91
computed tomography scan | -30
radiation therapy | -14
Piggyback LT | 0
hepatitis B | 0
entecavir | 0
HBV serology test | 0
hepatitis B virus | 0
human immunodeficiency virus | 0
hepatitis A | 0
hepatitis C | 0
donor | 0
brain death | 0
car accident | 0
HLA class-I | 0
HLA class-II | 0
blood products | 0
irradiated | 0
filtered | 0
transplantation process | 0
acute renal failure | 0
hematoma | 0
hepatitis B immunoglobulin | 24
immunosuppressive drugs | 24
steroids | 24
tacrolimus | 24
hemodialysis | 24
fresh frozen plasma | 24
leukocyte-depleted red blood cells | 24
pathological analyses | 240
HCC | 240
massive tumor necrosis | 240
liver function | 240
improvement | 240
aspartate aminotransferase | 240
alanine aminotransferase | 240
gamma-glutamyl transpeptidase | 240
alkaline phosphatase | 240
fever | 240
procalcitonin | 240
PCT levels | 240
blood cultures | 312
cytomegalovirus | 312
Epstein-Barr virus | 312
rash | 312
obscure red spots | 312
chest | 312
tacrolimus administration | 408
sirolimus | 408
mycophenolate mofetil | 408
immune suppression | 408
sputum culture | 432
Acinetobacter baumannii | 432
methicillin-resistant Staphylococcus aureus | 432
infections | 432
rash advanced | 456
erythematous macules | 456
papules | 456
limbs | 456
palms | 456
neck | 456
face | 456
oral examination | 456
white ulcers | 456
buccal mucosa | 456
lips | 456
bone marrow suppression | 456
white blood cell count | 456
platelet count | 456
hemoglobin level | 456
intensive care unit | 456
dermatologist | 456
gamma globulin administration | 456
skin biopsy | 456
fluorescence in situ hybridization | 456
peripheral blood | 456
abdominal incision | 696
sutured | 696
bone marrow aspiration | 768
bone marrow pathology | 768
granulocytes | 768
red blood cells | 768
megakaryocytes | 768
macrophages | 768
neutrophils | 768
platelets | 768
bone marrow cell morphology | 768
megakaryocyte production | 768
platelet levels | 768
FISH analysis | 792
donor lymphocytes | 792
skin biopsy specimens | 792
epidermal dyskeratosis | 792
basic vacuolization | 792
lymphocytic infiltrates | 792
grade-1 acute lt-GVHD | 792
multidisciplinary team | 816
steroids | 816
tacrolimus | 816
granulocyte colony-stimulating factor | 816
meropenem | 816
voriconazole | 816
anti-infective therapy | 816
rash reduced | 816
general condition | 816
deteriorate | 816
serum ferritin levels | 816
esophageal ulcers | 816
oral ulcers | 816
eating | 816
temperature | 1128
hallucinations | 1128
septic shock | 1320
multiple organ dysfunction syndrome | 1320
death | 1320