65 years old | 0
male | 0
diabetic | 0
transhiatal oesophagectomy | -264
gastric resection | -264
adenocarcinoma of the gastro-oesophageal junction | -264
progressive breathlessness | 240
severe breathlessness | 264
reduced air entry on left hemithorax | 264
chest X-ray revealing large bowel loops in left hemithorax | 264
diaphragmatic hernia | 264
emergency thoracolaparotomy | 264
severe respiratory distress | 264
inability to lie down | 264
nasal flaring | 264
active accessory muscles | 264
sweating | 264
dilated neck veins | 264
respiratory rate 40/min | 264
thready pulse | 264
pulse rate 180/min | 264
blood pressure 90/60 mmHg | 264
oxygen saturation 85-90% | 264
supplemental oxygen 6 l/min | 264
preoxygenation | 264
induction in sitting position | 264
fluid resuscitation | 264
rapid sequence induction technique | 264
haemodynamic instability | 264
noradrenaline infusion initiated | 264
airway pressures up to 42 cm H2O | 264
improvement in haemodynamic parameters | 264
resolution of high airway pressures | 264
noradrenaline infusion weaned off | 264
transfer to intensive care unit | 288
ventilatory support | 288
severe mixed acidosis | 288
weaned off ventilator | 312
extubation | 312
succumbed to septic shock | 384
anastomotic leak | 384
