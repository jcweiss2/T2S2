53 years old | 0
female | 0
liposculpture surgery | 0
wide liposuction of the dorsal region | 0
wide liposuction of the flanks | 0
wide liposuction of the thighs | 0
fat graft insertion into the gluteal area | 0
fever | -168
disabling pain at the surgical site | -168
extensive bullae formation | -168
signs of septic shock | -72
vasopressor support | -72
mechanical ventilation | -72
acute renal failure | -72
admitted to the intensive care unit | -72
air transportation | 0
septic shock | 0
multiple and extensive lesions | 0
subcutaneous emphysema | 0
leakage of purulent material | 0
erythema | 0
necrosis at the wound edges | 0
CT scan of the abdomen | 0
cutaneous dehiscence towards the left flank | 0
cutaneous dehiscence towards the right flank | 0
extension to the iliac crests | 0
extension to the left gluteal region | 0
extension to the perineal region | 0
extensive generalized soft tissue emphysema | 0
air dissected some of the muscular planes | 0
striation of subcutaneous fatty tissue | 0
diagnosis of necrotizing soft tissue infection | 0
surgical wound cleansing | 0
mechanical scrubbing | 0
debridement | 0
use of prophylactic antibiotics | 0
correct identification of the pathogen involved | 0
surgical intervention for drainage | 0
placement of a negative pressure therapy system | 0
metabolic acidosis | 0
hyperlactatemia | 0
leukocytosis with a left shift | 0
thrombocytopenia | 0
elevated CRP | 0
elevated ESR | 0
hyperglycemia | 0
remained in the intensive care unit for 7 days | 168
source of infection controlled | 168
hemodynamic stabilization achieved | 168
hospitalized for 42 days | 1008
15 surgical interventions performed | 0
multiple wound cleansing | 0
advancement of flaps | 0
lesions reconstruction | 0
procurement and placement of grafts | 0
secretion cultures | 0
E. Coli found | 0
Finegoldia magna found | 0
Streptococcus mitis found | 0
antibiotic management with Vancomycin | 0
antibiotic management with Meropenem | 0
antibiotic management with Clindamycin | 0
discharged | 1008
intensive rehabilitation program | 1008
no further complications | 1008
