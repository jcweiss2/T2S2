68 years old | 0
female | 0
admitted to the hospital | 0
jaundice | -72
general weakness | -72
fatigue | -72
decreased appetite | -72
icteric sclera | 0
acute bronchitis | 0
tranexamic acid | -168
N-acetylcysteine | -168
dihydrocodeine | -168
azithromycin | -168
normal vital signs | 0
CT scan | 0
bronchoscopy | 0
no history of allergic diseases | 0
denies alcohol consumption | 0
denies smoking | 0
white blood cell count | 0
hemoglobin level | 0
platelet count | 0
aspartate aminotransferase level | 0
alanine aminotransferase level | 0
total bilirubin level | 0
direct bilirubin level | 0
alkaline phosphatase level | 0
gamma-glutamyl transferase level | 0
total protein concentration | 0
albumin level | 0
blood urea nitrogen level | 0
creatinine level | 0
sodium concentration | 0
potassium concentration | 0
amylase level | 0
lipase level | 0
ammonia concentration | 0
prothrombin time | 0
partial thromboplastin time | 0
high sensitivity C-reactive protein level | 0
hepatitis A virus immunoglobulin M antibody | 0
hepatitis B surface antigen | 0
anti-HCV | 0
Epstein-Barr virus viral capsid antigen-IgM | 0
Epstein-Barr virus early antigen-diffuse restrict IgM | 0
cytomegalovirus IgM | 0
cytomegalovirus real-time polymerase chain reaction | 0
herpes simplex virus-IgM | 0
herpes simplex virus-immunoglobulin G | 0
toxoplasma IgM | 0
human immunodeficiency virus serum | 0
antinuclear antibody | 0
anti-mitochondrial antibody | 0
anti-smooth muscle antibody | 0
liver kidney microsomal antibody | 0
IgG serum level | 0
CT image | -168
periportal edema | 0
gallbladder wall edema | 0
ascites | 0
azithromycin-induced liver injury | 0
discontinuation of medications | 0
Roussel Uclaf Causality Assessment Method | 0
RUCAM score for azithromycin | 0
RUCAM score for tranexamic acid | 0
RUCAM score for N-acetylcysteine | 0
RUCAM score for dihydrocodeine | 0
hepatocellular type | 0
diagnosis of azithromycin-induced liver injury | 0
diagnosis of acute liver failure | 0
medical treatment | 0
worsening laboratory test values | 24
flapping tremor | 72
decreased level of consciousness | 72
hepatic encephalopathy | 72
semi-coma | 72
living donor liver transplantation | 192
recovery of consciousness | 192
recovery of liver function | 192
discharge from hospital | 240
histological examination of explanted liver | 240
fulminant hepatitis | 240
zone 3 necrosis | 240
extensive hepatocyte death | 240