9 years old | 0
male | 0
admitted to the hospital | 0
painful skin eruption | -720
fever | -720
generalized malaise | -720
erythematous macules | 0
papules | 0
necrotic plaques | 0
hemorrhagic crusts | 0
mucous membrane involvement | 0
oral mucosa involvement | 0
small painful ulcers on the tongue | 0
small painful ulcers on the inner lip | 0
mild leukocytosis | 0
elevated erythrocyte sedimentation rate | 0
elevated C-reactive protein | 0
anemia | 0
skin biopsy | 0
focal full-thickness epidermal necrosis | 0
exocytosis | 0
vacuolar interface dermatitis | 0
prominent superficial and deep perivascular lymphocytic infiltrate | 0
focal hemorrhage | 0
diagnosis of FUMHD | 0
systemic antibiotics | 0
azithromycin | 0
systemic steroids | 0
left the hospital | 240
treated at another hospital | 240
intravenous immunoglobulins | 240
cyclosporine | 240
returned to the hospital | 504
ulceronecrotic papules increased in number and size | 504
ulceronecrotic plaques became confluent | 504
Pseudomonas aeruginosa infection | 504
gangrenous ulcers | 504
central black eschars | 504
erythematous borders | 504
ecthyma gangrenosum | 504
systemic vancomycin | 504
gentamycin | 504
systemic inflammatory response syndrome | 504
tachypnea | 504
tachycardia | 504
hypothermia | 504
supportive measures | 504
intravenous fluids | 504
refractory hypotension | 504
myocardial dysfunction | 504
generalized edema | 504
fulminant sepsis | 504
multiple organ failure | 504
death | 528