72 years old | 0
female | 0
admitted to the hospital | 0
fever | -24
pain in bilateral big toes | -24
no history of trauma | 0
no insect bites recently | 0
episodes of fever and pain happen twice a year | 0
resolves spontaneously | 0
used to take Traditional Chinese Medicine | 0
drug toxicology screen was negative | 0
no diagnosis of joint problem | 0
no autoimmune problem | 0
vasculitis screen was negative | 0
borderline positive anti-nuclear antibody | 0
no risk factors for peripheral vascular disease | 0
pain on bilateral big toes | 0
bilateral podagra | 0
minimal swelling | 0
full range of motion | 0
pulses were well felt | 0
diagnosis of streptococcal septicaemia | 0
growth of Streptococcus pneumoniae in blood culture | 0
broad spectrum antibiotics started | 0
hypotension | 0
urine output of <20 ml/h | 0
dopamine used | 0
noradrenaline used | 48
vital signs normalized | 48
extremities were noted to be dusky | 48
livedo reticularis | 48
patches of ecchymosis | 72
mottled skin | 72
necrotic terminal digits | 120
necrotic tip of nose | 120
signs of dry gangrene | 120
ecchymotic bullae | 168
plantar gangrene | 168
dorsalis pedis and posterior tibial pulses were not palpable | 168
radial pulses were not palpable | 168
dry gangrene involved all digits | 168
referral to vascular surgeon | 168
diagnosis of microvascular spasm | 168
inotropes resulting in peripheral gangrene | 168
arterial occlusion test | 168
moderate calcification of bilateral lower limb arteries | 168
referral to plastic surgery | 168
plan to await dry gangrene to demarcate | 168
dry gangrene progressed to bilateral ankles and wrists | 720
dry gangrene demarcated | 720
elective 4 limb amputations | 1440
bilateral below knee amputations | 1440
bilateral above elbow amputations | 1440
recovery was smooth post-operatively | 1440
rehabilitation started | 1440
ambulatory with bilateral lower limb prosthesis | 2160
utilizes bilateral upper limb prosthesis | 2160