71 years old | 0
female | 0
mRCC | -672
mixed papillary and clear cell type | -672
retroperitoneal lymph node metastases | -672
right ovarian metastases | -672
liver metastases | -672
ipilimumab | -672
nivolumab | -672
maintenance single-agent nivolumab | -336
immune-related primary hypoadrenalism | -336
hypopituitarism | -336
secondary hypoadrenalism | -336
secondary hypothyroidism | -336
exogenous hydrocortisone | -336
fludrocortisone | -336
thyroxine replacement | -336
short synacthen test | -336
MRI pituitary | -336
disease progression | 0
sunitinib | 0
admitted to the hospital | 14
presumed sepsis | 14
fever | 14
hypotension | 14
tachycardia | 14
broad-spectrum antibiotics | 14
intravenous stress dose steroids | 14
inotropes | 14
septic screen | 14
discharged from the hospital | 21
steroid replacement adjusted | 21
sunitinib restarted | 21
re-presented with the same symptoms | 26
broad-spectrum antibiotics | 26
intravenous stress dose steroids | 26
inotropes | 26
septic screen | 26
baseline steroid dose reviewed | 26
reduced dose of sunitinib | 26
re-presented with the same symptoms | 27
ICU admission | 27
stress dose steroids | 27
inotropes | 27
broad-spectrum antibiotics | 27
septic screen | 27
tunnelled venous access catheter removed | 27
baseline steroid dose revised | 27
elective admission for a trial of sunitinib | 28
sunitinib administration | 28
profoundly hypotensive | 29
tachycardic | 29
aggressive intravenous fluid replacement | 29
intravenous steroids | 29
inotropes | 29
haemodynamic parameters normalized | 30
transitioned back to oral steroids | 30
sunitinib therapy permanently discontinued | 30