64 years old | 0
male | 0
hypertension | -672
tobacco consumption | -672
moderate obesity | -672
alcohol consumption | -672
hepatocellular carcinoma | -672
abdominal pain | -672
appendicular syndrome | -672
liver steatosis | -672
liver fibrosis | -672
liver cirrhosis | 0
portal hypertension | 0
normal liver function | 0
prothrombin time | 0
bilirubinemia | 0
albuminemia | 0
creatininemia | 0
platelet count | 0
tumor in right liver | -672
extended right hepatectomy | 0
perioperative Doppler ultrasound | 0
vascular patency | 0
intermittent portal clamping | 0
caval clamping | 0
hemodynamic insufficiency | 0
crystalloids administration | 0
red blood cells transfusions | 0
R0 resection | 0
hepatocellular carcinoma resection | 0
non-severe pulmonary embolism | 48
post-operative day 2 | 48
remnant liver volume measurement | 48
PHLF | 120
hyperbilirubinemia | 120
ascites | 120
sepsis | 120
antibiotic treatment | 120
intensive care | 120
remnant liver volume measurement | 216
left hepatic vein stenosis | 432
DUS | 432
cavography | 432
pressure gradient measurement | 432
percutaneous transluminal angioplasty | 432
metallic stent placement | 432
LHV-IVC gradient measurement | 432
post-intervention recovery | 432
bilirubinemia reduction | 432
discharge | 720
bilirubin level measurement | 1440
PT measurement | 1440
liver function tests | 2880
morphological imaging | 2880
liver regeneration | 2880
metallic stent permeability | 2880