12 years old | 0
male | 0
stung by numerous (around 500 stings) African bee | -1
stung on the face | -1
stung on the upper limbs | -1
stung on the trunk | -1
admitted to a local hospital | 0
IV fluids | 0
hydrocortisone | 0
diclofenac IM for pain | 0
facial edema progressive | 28
decrease in urine output | 28
furosemide (2 mg/kg) | 28
BP 100/70 mmHg | 28
HR 68 beat/min | 28
RR 35 breath/min | 28
referred to tertiary hospital | 28
conscious | 28
could not see well | 28
facial swelling | 28
peri-orbital edema | 28
erythema stings marks on face | 28
erythema stings marks on trunk | 28
erythema stings marks on upper limbs | 28
saturating in room air at 97% | 28
RR 28 breath/min | 28
HR 94 beat/min | 28
BP 118/70 mmHg (90th percentile) | 28
broad spectrum antibiotic (ceftriaxone) | 28
fluid restriction | 28
creatinine 116 mmol/l | 28
urea 15.4 mmol/l | 28
hyperkalemia 6.9 mmol/l | 28
D10% plus Insulin | 28
calcium gluconate | 28
hyponatremia 128mmol/l | 28
catheter inserted | 28
urine dipstick RBC+++ | 28
muddy brown cast | 28
leucocytosis 25 | 28
neutrophils 89.7% | 28
hemoglobin 13.8 g/dl | 28
normocytic normochromic | 28
platelet count 269 | 28
K 5.15 mmol/l | 28
Na 128 mmol/l | 28
urine output 200 ml | 28
amber colored urine | 28
creatinine 248 mmol/l | 28
urea 22.52 mmol/l | 28
fluid input 700 ml | 28
urine output 100 ml | 28
creatinine 402 mmol/l | 28
urea 29.83 mmol/l | 28
potassium 5.4 mmol/l | 28
sodium 127 mmol/l | 28
transferred to PICU | 28
hemodialysis considered inevitable | 28
potassium 5.99 mmol/l | 28
creatinine 462 mmol/l | 28
urea 34.65 mmol/l | 28
five dialysis sessions | 28
high grade fever 38.6°C | 28
blood cultures collected | 28
vancomycin every third day for 1 month | 28
cultures negative on Day 7 | 28
urine output raised to 1.8 ml/kg/h | 28
creatinine 172 mmol/l | 28
urea 11 mmol/l | 28
K+ 4.6 mmol/l | 28
Na+ 138mmol/l | 28
hospital stay 2 weeks | 336
creatinine 52 mmol/l | 504
urea 2.96 mmol/l | 504
electrolytes normal | 504
facial swelling disappeared | 28
creatinine recovered to normal | 28
urine output recovered to normal | 28
blood in urine | 28
acute kidney injury | 28
acute tubular necrosis | 28
acute tubular interstitial nephritis | 28
rhabdomyolysis | 28
pigment tubulopathy | 28
erythema on skin | 28
skin healed leaving black spots | 28
anaphylaxis | 28
hypotension | 28
hemodialysis | 28
fluid retention | 28
metabolic worsening | 28
hematocrit 43.7% | 28
MCV 85.8 fl | 28
MCH 27.1 pg | 28
MCHC 31.6 g/dl | 28
leukocyte 25 × 10^9 cells/ml | 28
lymphocytes 5.3% | 28
monocytes 2.7% | 28
eosinophils 2.1% | 28
basophils 0.2% | 28
platelet 550 × 10^9/ml | 28
Hepatitis B surface antigen Negative | 28
Hepatitis C antigen Negative | 28
blood cultures no bacterial growth | 28
