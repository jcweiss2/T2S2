27 years old| 0
male| 0
admitted to the hospital (psychiatric department)| 0
acute psychiatric syndrome| 0
personality change| 0
behavioral change| 0
friendly behavior| 0
focused attention| 0
clear consciousness| 0
slow response to questions| 0
emotional instability| 0
interruption of thinking| 0
thinking burst| 0
absence of hallucination| 0
absence of delusion| 0
absence of impulsive aggression| 0
psychotropic drugs use| 0
no response to psychotropic drugs| 0
rigidity emerged| 168
transferred to neurology department| 288
suspected viral encephalitis| 288
neurological impairment| 288
abnormal movements| 288
tachycardia| 288
progressed to status epilepticus| 288
insomnia| 288
confusion of consciousness| 288
memory deficits| 288
absence of fever| 288
EEG showed diffuse slowing| 288
EEG showed general slowing| 288
MRI brain normal| 288
CSF protein elevation (90 mg/dL)| 288
CSF karyocyte count elevation (50 × 106/L)| 288
CSF glucose normal| 288
NMDAR antibodies detected in CSF (1/100)| 288
NMDAR antibodies detected in serum (1/10)| 288
tumor screening negative| 288
ANMDARE diagnosis| 288
anti-epileptic drugs| 288
corticosteroids (methylprednisolone 1 g/d for 5 days)| 288
tapered oral prednisolone| 288
IVIG (400 mg/kg daily for 5 days)| 288
discharge from hospital| 288
clear mind at discharge| 288
normal behaviors at discharge| 288
readmission to EICU| 720
hyperpyrexia (39.0°C)| 720
dyspnea| 720
severe status epilepticus| 720
decreased level of consciousness| 720
limb convulsions| 720
supplemental oxygen therapy| 720
perspiration| 720
cutaneous pallor| 720
tachypnea (35 bpm)| 720
hypoxemia (SaO2 86%)| 720
scattered crackles| 720
diffuse crackles| 720
rhonchi| 720
CRP elevation (75 mg/L)| 720
PCT elevation (22 ng/mL)| 720
chest CT showing acute lung inflammation| 720
CSF NMDAR antibodies positive (1/80)| 720
HSV DNA PCR negative| 720
Acinetobacter baumannii in sputum culture| 720
ANMDARE relapse diagnosis| 720
acinetobacter baumannii pneumonia diagnosis| 720
steroid pulse therapy| 720
IVIG pulse therapy| 720
antibacterial agents| 720
supportive therapies| 720
no tumor detection| 720
gradual recovery| 720
mild psychiatric sequelae| 720
