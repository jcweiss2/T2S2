72 years old | 0
    man | 0
    referred to emergency department | 0
    fever | -168
    non-productive cough | -168
    shortness of breath | -168
    gradual onset | -168
    increasing severity | -168
    history of malignancy | 0
    no malignancy | 0
    history of diabetes | 0
    no diabetes | 0
    history of cardiovascular disease | 0
    no cardiovascular disease | 0
    PCR-based test for SARS-CoV-2 | -168
    positive SARS-CoV-2 | -168
    respiratory rate 55 breaths per minute | 0
    peripheral oxygen saturation 74% | 0
    15 L/min oxygen | 0
    non-rebreather mask | 0
    blood pressure 144/91 mmHg | 0
    heart rate 145 beats per minute | 0
    body temperature 36.8°C | 0
    increased white cell count 15,840 cells/μL | 0
    8% lymphocytes | 0
    normal platelet count 192,000 platelets/μL | 0
    blood gas analysis pH 7.42 | 0
    pCO2 23 mmHg | 0
    pO2 43 mmHg | 0
    HCO3 15 mmol/L | 0
    base deficit -9 mmol/L | 0
    lactic acid 7.46 mmol/L | 0
    BUN 36 mg/dL | 0
    creatinine 1.4 mg/dL | 0
    ALT 169 U/L | 0
    AST 238 U/L | 0
    increased procalcitonin 51.36 ng/mL | 0
    hs-CRP 391 mg/L | 0
    elevated D-dimer >50,000 ng/mL FEU | 0
    increased fibrinogen 439 mg/dL | 0
    CKMB 31.8 ng/mL | 0
    troponin I 0.61 ng/mL | 0
    sinus tachycardia | 0
    chest X-ray heterogenous consolidation | 0
    blood culture negative | 0
    initiated HFNO therapy | 0
    oxygen flow 40 liters/minute | 0
    100% FiO2 | 0
    oxygen saturation improved to 92% | 0
    respiratory rate improved to 26 breaths per minute | 0
    blood pressure improved to 130/80 mmHg | 0
    heart rate improved to 120 beats per minute | 0
    informed consent | 0
    central venous catheter placement | 0
    arterial catheter placement | 0
    treated with aspirin | 0
    treated with clopidogrel | 0
    infusion with UFH | 0
    aPTT checked every 6 hours | 0
    target aPTT 2 to 2.5 times control value | 0
    transferred to ICU | 0
    management in ICU | 0
    meropenem 1 gram every 8 hours | 0
    levofloxacin 750 mg/day | 0
    dexamethasone 5 mg every 12 hours | 0
    famotidine 20 mg/day | 0
    vitamin D 400 IU/day | 0
    ascorbic acid 500 mg every 8 hours | 0
    zinc 100 mg/day | 0
    atorvastatin 40 mg/day | 0
    NAC 200 mg every 8 hours | 0
    nebulized lidocaine | 0
    average UFH dose 25,191 units/day | 0
    mean aPTT 64.35 seconds | 0
    condition improved | 0
    oxygen down-titrated to simple face mask | 264
    blood gas analysis pH 7.41 | 264
    pCO2 37 mmHg | 264
    pO2 74 mmHg | 264
    HCO3 24 mmol/L | 264
    base deficit -1 mmol/L | 264
    lactic acid 1.36 mmol/L | 264
    procalcitonin decreased to 7.4 ng/mL | 264
    hs-CRP decreased to 0.13 mg/dL | 264
    D-dimer decreased to 5,308 ng/mL FEU | 264
    increased fibrinogen 523 mg/dL | 264
    ALT decreased to 153 U/L | 264
    AST decreased to 62 U/L | 264
    sudden clinical deterioration | 264
    labored breathing | 264
    desaturation | 264
    hypotension | 264
    altered mental status | 264
    endotracheal intubation | 264
    inotropic agents | 264
    vasopressor agents | 264
    CTPA revealed bilateral pulmonary artery thrombosis | 288
    multiple pulmonary vein thrombosis | 288
    brain CT scan infarct left parietal lobe | 288
    infarct pons | 288
    infarct left cerebellum | 288
    rescue thrombolytic therapy | 288
    streptokinase loading dose 250,000 IU | 288
    streptokinase 100,000 IU/hour over 12 hours | 288
    critical condition | 336
    no improvement after thrombolytic therapy | 336
    hs-CRP 221.1 mg/dL | 336
    ferritin >15,000 μg/L | 336
    D-dimer 2,597 ng/mL FEU | 336
    fibrinogen 634 mg/dL | 336
    tocilizumab 600 mg infusion | 336
    died due to multiple end-organ failure | 432
    