18 years old| 0
male | 0
admitted to the hospital | 0
fever | -72
rash | -72
acne |  -672
minocycline |  -672
increased WBC count | 0
eosinophilia| 0
systemic involvement| 0
diffuse erythematous or maculopapular eruption| 0
pruritis | 0
DRESS syndrome | 0
fever persisted | 0
rash persisted | 0
discharged | 24
Separate conjunctive phrases into its component events and assign them the same timestamp (for example, the separation of 'fever and rash' into 2 events: 'fever' and 'rash')  If the event has duration, assign the event time as the start of the time interval. Attempt to use the text span without modifications except 'history of' where applicable. Include all patient events, even if they appear in the discussion; do not omit any events; include termination/discontinuation events; include the pertinent negative findings, like 'no shortness of breath' and 'denies chest pain'.  Show the events and timestamps in rows, each row has two columns: one column for the event, the other column for the timestamp.  The time is a numeric value in hour unit. The two columns are separated by a pipe '|' as a bar-separated file. Skip the title of the table. Reply with the table only. Create a table from the following case:
17 years old| 0
female | 0
admitted with fever | -504
productive cough | -504
right pleuritic chest pain | -504
crepitations bilaterally | 0
reduced breath sounds at right lower hemithorax | 0
stony dullness on percussion | 0
hemoglobin 9.0 g/dL | 0
platelet count 386,000/μL | 0
white blood cell count 12,140/μL | 0
coagulation profile normal | 0
chest radiograph showing large right loculated pleural effusion | 0
28-French chest tube inserted | 0
drained 1.2 L of pus | 0
diagnosed with right loculated empyema thoracis | 0
started on intravenous co-amoxiclav | 0
vital signs returned to normal | 48
chest tube replaced due to blockage | 72
chest tube drainage remained poor | 72
persistent pleural effusion | 72
flushing with normal saline | 72
started on intrapleural streptokinase | 72
complained of palpitations | 108
sweating | 108
giddiness | 108
respiratory rate 25 breaths/minute | 108
blood pressure 70/50 mm Hg | 108
pulse rate 140 beats/minute | 108
temperature 38.3°C | 108
hemoglobin dropped to 6.5 g/dL | 108
platelet count 209,000/μL | 108
white cell count 18,600/μL | 108
International Normalized Ratio 1.5 | 108
activated partial thromboplastin time normal | 108
chest radiograph showing right massive hemothorax | 108
diagnosed with right massive hemothorax | 108
thoracic surgical consult sought | 108
chest tube replaced again | 108
drained 1.1 L of altered blood | 144
transfused 7 units of packed red blood cells | 144
hemoglobin level 9.6 g/dL post-transfusion | 144
coagulation profile normalized | 144
transferred to cardiothoracic center | 336
underwent right lung decortications | 336
recovered uneventfully | 336
