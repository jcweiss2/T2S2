19 years old | 0
male | 0
presented with a two-day history of fever | -48
presented with a two-day history of malaise | -48
presented with a two-day history of headache | -48
presented with a two-day history of vomiting | -48
presented with a two-day history of an episode of near-syncope | -48
no relevant medical history | 0
confused | 0
fever of 39.3 °C | 0
blood pressure of 124/66 mmHg | 0
pulse rate of 126 bpm | 0
oxygen saturation of 100% on ambient air | 0
maculopapular rash spread in the legs and thigh | 0
tender, solid, non-fluctuant, mobile nodule in the left armpit | 0
developed a few days back | -72
normal breath sounds bilaterally | 0
no lymphadenopathy | 0
white count of 26.9 k/mm³ | 0
neutrophils of 91% with bands | 0
procalcitonin of 0.42 ng/mL | 0
lactic acid of 3.1 mmol/L | 0
chest radiography showed no acute pulmonary disease | 0
negative urine analysis | 0
negative SARS-CoV-2 RT-PCR | 0
negative Legionella urinary antigen | 0
negative pneumococcus urinary antigen | 0
started on ceftriaxone | 0
started on doxycycline | 0
admitted to the general medical ward | 0
lumbar puncture performed | 0
cerebrospinal fluid analysis showed no evidence of infection | 0
transthoracic echocardiogram done | 0
no evidence of vegetations | 0
day 2 admission developed persistent hypotension | 48
day 2 admission developed tachycardia | 48
day 2 admission developed fever to 40 °C | 48
day 2 admission developed profound upper and lower extremities weakness | 48
transferred to the ICU | 48
white count increased to 41.7 k/mm³ | 48
AST 113 IU/L | 48
ALT 151 IU/L | 48
CK 319 IU/L | 48
high sensitivity troponin 27 pg/mL | 48
D-dimer 1067 ng/mL FEU | 48
C-reactive protein 18 mg/dL | 48
erythrocyte sedimentation rate 42 mm/h | 48
interleukin-6 1620 pg/mL | 48
fibrinogen 625 mg/dL | 48
repeat SARS-CoV-2 RT-PCR negative | 48
IgG antibodies negative | 48
respiratory viral panel negative | 48
MRSA PCR screen positive | 48
negative gonococcus DNA probe | 48
negative Chlamydia DNA probe | 48
negative HSV1 and 2 antigen/antibodies | 48
negative hepatitis panel | 48
negative Rickettsia antibody agglutination | 48
negative Brucella antibody agglutination | 48
negative EBV IgM and IgG VCA antibodies | 48
negative EBV PCR | 48
negative CMV antibodies | 48
negative West Nile Virus antibody panel | 48
negative Lyme IgM and IgG antibodies Western Blot | 48
negative Syphilis screen | 48
negative interferon release assay for tuberculosis | 48
negative malarial smear | 48
negative Histoplasma galactomannan urine antigen | 48
normal C3 complement levels | 48
normal C4 complement levels | 48
negative ANA | 48
negative P2-ANCA | 48
negative C-ANCA | 48
negative rheumatoid factor | 48
MRI spine ruled out spinal abscess | 48
MRI spine ruled out paravertebral abscess | 48
CT head ruled out intracranial infections | 48
CT chest ruled out new lung involvement | 48
CT abdomen ruled out intraabdominal infection | 48
started on IV vancomycin | 48
day 4 white count trending down | 96
day 4 lactic acid trending down | 96
day 4 fever decreased | 96
day 4 vitals became stable | 96
discharged from the ICU | 96
left armpit pain | 96
nodule evolved into an abscess with fluctuance | 96
flushed | 96
nonspecific erythrasma on the lower limbs | 96
deep palmar erythema | 96
suspicion for staphylococcal TSS | 96
incision and drainage of the abscess performed | 96
culture sent | 96
gradually improved | 96
rashes started to have central clearance | 96
flaky skin in the palms | 96
monitored for possible generalized desquamation | 96
discharged in stable condition | 96
oral amoxicillin-clavulanate for 14 days | 96
diffuse erythroderma nearly resolved except palms and soles | 96
flakiness with pinkish coloration in the palms | 96
rash started to improve on vancomycin | 96
vancomycin-induced rash deemed unlikely | 96
wound cultures showed methicillin-susceptible Staphylococcus aureus | 96
definitive diagnosis of staphylococcal TSS secondary to abscess | 96
