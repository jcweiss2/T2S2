78 years old | 0
male | 0
leg edema | -24
ruptured abdominal aortic aneurysm | -8760
aorto-bi-iliac graft | -8760
smoking history | -87600
widowed | 0
retired public school employee | 0
new onset atrial fibrillation | 0
warfarin | 0
digoxin | 0
diuretic therapy | 0
shortness of breath | -48
leg edema (persisted) | -72
nonproductive cough | -168
malaise | -504
fatigue | -504
weakness | -504
denied fever | 0
denied chills | 0
denied sweats | 0
temperature 36.8oC | 0
pulse 132/minute | 0
blood pressure 105/56 mmHg | 0
respirations 28/minute | 0
jugular venous distension | 0
irregularly irregular pulse | 0
left-sided rhonchi | 0
bibasilar pulmonary crackles | 0
left lower pulmonary infiltrate | 0
left pleural effusion | 0
cardiomegaly | 0
atrial fibrillation | 0
no ischemic changes | 0
creatine phosphokinase 2205 U/L | 0
AST 128 U/L |
