77 years old | 0
female | 0
uncontrolled diabetes | 0
hypertension | 0
chronic obstructive airway disease | 0
admitted to ICU | 0
bilateral pneumonia | 0
acute kidney injury | 0
intubated | 0
subclavian central line inserted | 0
vasopressors started | 0
injection piperacillin and tazobactum combination started | 0
injection clindamycin started | 0
injection meropenem started | 0
injection teicoplanin started | 0
injection colistin started | 0
injection Fluconazole started | 120
watery diarrhea | 168
injection racecadotril started | 168
injection metronidazole started | 168
Saccharomyces containing sachet started | 168
stool routine/microscopy done | 168
stool culture done | 168
stool toxin for C. difficile done | 168
diarrhea settled | 168
hypotension | 216
diarrhea again | 216
injection fluconazole changed to injection caspofungin | 216
blood culture done | 216
blood culture report sterile | 264
blood culture report showed growth of yeast | 336
yeast reported as Saccharomyces cerevisiae | 336
injection caspofungin stopped | 336
injection amphotericin B started | 336
Saccharomyces containing probiotic stopped | 336
central line removed | 336
repeat blood cultures done | 360
repeat blood cultures showed no fungal growth | 432
patient died | 576