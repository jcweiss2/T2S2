19 years old | 0
male | 0
Han nationality | 0
student | 0
unmarried | 0
admitted to the hospital | 0
chest pain | -240
oliguria | -240
phlegm | -168
Nuss surgery 4 years ago | -34560
pectus excavatum | -34560
metal bar removed | -1440
no special medical history | 0
no family history | 0
nausea after drinking milk | -240
violent vomiting | -240
sent to local hospital | -240
emergent electrocardiogram | -240
ST-segment elevation | -240
coronary angiogram | -240
midsection anterior descending branch | -240
acute myocardial infarction suspected | -240
myocarditis suspected | -240
admitted to cardiology department | -240
chest pain improved | -216
nausea persisted | -216
vomiting persisted | -216
anuria | -216
acute liver failure considered | -216
acute renal failure considered | -216
transferred to ICU | -216
emergency blood tests | -216
WBC 18.3×109/L | -216
neutrophiles granulocyte 87.5% | -216
glutamic-pyruvic transaminase 3469 U | -216
glutamic oxalacetic transaminase 3815 U/L | -216
total bilirubin 54.2 μmol/L | -216
creatinine 217 mmol/L | -216
urea nitrogen 10.8 mmol/L | -216
serum potassium 7.47 mmol/L | -216
creatine kinase 541 U/L | -216
creatine kinase 50.4 U/L | -216
lactate dehydrogenase 4138 U/L | -216
procalcitonin 0.13 ng/mL | -216
C-reactive protein 22.8 mg/L | -216
complement and protein 148 | -216
anti-infection | -216
continuous renal replacement treatment | -216
symptomatic treatments | -216
specimens collected | -216
etiological examination | -216
toxicological examination | -216
vital signs stabilized | -216
sudden shock | -168
decreasing heart rate | -168
emergency endotracheal intubation | -168
mechanical ventilation | -168
cardiopulmonary resuscitation | -168
fluid resuscitation | -168
low blood pressure | -168
vasopressors | -168
Dopamine 10 μg/kg/min | -168
Norepinephrine 0.1 μg/kg/min | -168
vital signs stabilized again | -168
vasopressors stopped | -72
endotracheal intubation removed | -48
transferred to our hospital | 0
admitted to ICU | 0
temperature 36°C | 0
respiration rate 24 breaths/min | 0
pulse rate 102 beats/min | 0
blood pressure 154/98 mmHg | 0
clear consciousness | 0
poor spirits | 0
skin and mucosa slightly yellow | 0
scattered bleeding points | 0
subcutaneous ecchymosis | 0
soft neck | 0
no resistance | 0
thoracic deformity funnelform | 0
old surgical scar | 0
increased respiratory mobility | 0
increased respiratory frequency | 0
coarse breath sounds | 0
moist rales | 0
sputum sounds | 0
neat heart rhythm | 0
low-pitched heart sounds | 0
weakened muscle strength | 0
weakened muscle tension | 0
edema in lower extremities | 0
no other abnormalities | 0
WBC 8.36×109/L | 0
Grn% 95.4% | 0
platelet 65 g/L | 0
Troponin T 0.182 ng/mL | 0
creatine kinase 7.590 ng/mL | 0
myoglobin 835.3 ng/mL | 0
brain natriuretic peptide 6265 pg/mL | 0
chest radiograph lung infection | 0
left pleural effusion | 0
pericardial effusion | 0
pulmonary infection diagnosis | 0
renal failure diagnosis | 0
liver failure diagnosis | 0
acute cardiac insufficiency diagnosis | 0
acute myocardial infarction diagnosis | 0
myocarditis diagnosis | 0
poisoning suspected | 0
vital signs stable | 0
abundant sputum | 0
difficulty in sputum expectoration | 0
CT scan | 0
echocardiography | 0
palpitation | 24
dyspnea | 24
defecating 400 mL yellow mucous stools | 24
sweating | 24
cyanosis | 24
heart rate 130–140 bpm | 24
blood pressure 120–130/70-80 mmHg | 24
oxygen saturation 85%–90% | 24
heart rate continued to rise | 24
intubation | 24
mechanical ventilation | 24
oxygen saturation 92%–94% | 24
arterial blood gas oxygenation index 86.6 mmHg | 24
lactic acid 4.3 mmol/L | 24
emergency echocardiography | 24
restricted ventricular diastole | 24
stroke volume 17 mL | 24
diastolic pericardial fluid sonolucent area | 24
anechoic area post pericardium 1.8 cm | 24
anechoic area left ventricular lateral 1.0 cm | 24
anechoic area subcostal four chamber 1.4 cm | 24
apical pericardium 2.8 cm | 24
right ventricular lateral pericardium 4.1 cm | 24
flocculent echo | 24
no abnormal blood flow | 24
thorax puncture and drainage | 24
tawny turbid effusion | 24
pericardiocentesis | 24
drainage tube indwelled | 24
ultrasonography confirmed drainage tube | 24
200 mL dark red fluid drained | 24
symptoms slightly relieved | 24
vital signs more stable | 24
pericardiocentesis guided by ultrasonography | 48
bloody fluid extracted | 48
coagulation function disorder | 48
low prothrombin complex | 48
low fibrinogen | 48
coagulation factors added | 48
coagulation corrected | 48
stable for one day | 48
fraction of inspired oxygen decreased | 48
toxicology tests negative | 48
etiology tests negative | 48
oxygen saturation declined | 72
echocardiography reexamination | 72
effusion in right ventricle inferior wall | 72
active bleeding suspected | 72
no improvement after adjusting tube | 72
consultation with cardiologist | 72
consultation with thoracic surgeon | 72
consultation with radiologist | 72
chest CT showed sharp osteophyte | 72
osteophyte caused by Nuss surgery | 72
osteophyte damaged pericardium | 72
pericardial effusion | 72
acute cardiac tamponage | 72
repeated shock symptoms | 72
multiple organ dysfunction | 72
coagulation dysfunction | 72
surgical risk high | 72
communication with family | 72
thoracotomy under general anesthesia | 168
atelectasis lower left lobe | 168
partial consolidation | 168
thoracic hydrothorax 500 mL | 168
pericardium adhered to chest wall | 168
300 mL blood fluid extracted | 168
damage to left ventricle anterior wall | 168
fibrinoid material | 168
local blood exudation | 168
scar formation 3 cm | 168
horizontal mattress suture | 168
osteophytes trimmed | 168
bone wax applied | 168
returned to ward | 168
drainage tube bloody fluid | 168
fluid resuscitation | 168
vasopressor needed | 168
active bleeding | 168
hemoglobin 51 g/L | 168
emergency surgical exploration | 168
diffuse extravasation | 168
extensive hemostasis | 168
coagulation factors supplied | 168
second operation | 168
mechanical ventilation | 168
anti-infection | 168
CRRT | 168
tracheotomy | 312
intermittent blood supplementing | 312
ventilator parameters turned down | 312
antibiotics stopped | 408
renal function recovered | 600
CRRT stopped | 600
rehabilitation exercise | 600
ventilator removed | 1272
tracheal tube removed | 1272
discharged | 2592
