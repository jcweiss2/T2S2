37 years old | 0
male | 0
admitted to the hospital | 0
pain in left hemithorax | -168
pain in left upper abdomen | -168
fever | -168
body temperature of 39.1°C | -168
severe cough | -168
purulent greenish sputum | -168
alcohol abuser | -13140
tobacco smoker | -13140
periodic upper abdominal pain | -8760
shortness of breath | -168
dyspnea | -168
cough with increased sputum volume | -168
inability to remain in a prone position | -168
blood pressure of 140/90 mmHg | 0
heart rate of 98 beats per minute | 0
temperature of 38.2°C | 0
respiratory rate of 23 breaths per minute | 0
absent breath sound in the lower half of the left hemithorax | 0
reduced breath sounds with wheezing under the upper half of the left hemithorax | 0
hemoglobin of 12.5 g/dL | 0
white blood cells of 16 800/mm3 | 0
platelets of 590 000/mm3 | 0
elevated serum amylase | 0
elevated lipase | 0
elevated C-reactive protein | 0
positive for hepatitis C | 0
negative for human immunodeficiency virus (HIV) | 0
left pleural effusion | 0
structural changes of the pancreas | 0
chronic gastric and duodenal inflammation | 0
diagnosed with left-sided pneumonia | 0
diagnosed with pleural effusion | 0
diagnosed with acute onset of chronic alcoholic pancreatitis | 0
thoracentesis | 0
antibiotic treatment | 0
analgesics | 0
intravenous hydration | 0
pleural fluid and sputum cultures showed no bacterial growth | 24
sputum analysis for mycobacterium tuberculosis was negative | 24
repeated chest radiographs showed infiltration in the left lower lobe | 48
persisting pleural effusion | 48
abdominal computed tomography (CT) scans showed cystic changes of the pancreatic head and body | 48
fluid in the subhepatic space | 48
antibiotic treatment scheme was changed | 72
repeated x-rays showed 2 left lung abscesses | 96
left pleural cavity was drained | 96
measurement of the pleural fluid enzymes was undertaken | 96
high concentrations of amylase and lipase in pleural fluid | 96
suspected PPF | 96
abdominal magnetic resonance imaging (MRI) revealed a slightly dilated pancreatic duct | 96
cystic transformation of the pancreatic head | 96
pseudocyst in the body of the gland | 96
transferred to Mariinsky Hospital | 168
dyspnea | 168
cough with purulent sputum | 168
fever | 168
unable to sleep in a supine position | 168
chest CT showed multiple left lung abscesses | 168
lung abscesses were drained under radiologic guidance | 216
additional abscess cavity was drained | 216
pancreatic body pseudocyst was externally drained | 216
amylase level in pseudocyst fluid was 13 200 IU/L | 216
condition slowly improved | 240
fluid outflow from pseudocyst drain remained stable | 240
fluid outflow from pleural drains remained stable | 240
stenting of the pancreatic duct | 360
transcutaneous external-internal stenting with 14 Fr pancreatic stent | 360
puncture of slightly dilated duct was done | 360
fistula track from the pancreatic body pseudocyst was found | 360
ductal stricture was found in the head of the gland | 360
guide-wire and stent were pushed through it into the duodenum | 360
postoperative period was uneventful | 360
octreotide injections | 360
serum amylase level dropped to 150 IU/L | 384
pseudocyst drain outflow was stopped | 384
pseudocyst drain was removed | 384
pleural drains were removed | 504
symptoms quickly improved | 504
normalization of body temperature | 504
decrease of dyspnea | 504
disappearance of cough and sputum | 504
follow-up CT scan revealed small localized hydropneumothorax | 504
abdominal MRI showed diffuse parenchymal changes | 504
ductal hypertension | 504
PPF track was still visible | 504
discharged | 720
readmitted | 840
pancreatic surgery | 840
Bern modification of duodenum-preserving pancreatic head resection | 840
pancreatowirsungojejunal anastomosis with Roux-en-Y retrocolic jejunal loop | 840
postoperative period was uncomplicated | 840
discharged | 1008
outpatient ultrasound examination | 2160
signs of CP | 2160
no pseudocysts and ductal dilatation | 2160
telephone survey | 8760
no complaints | 8760
works as a builder | 8760
smokes 5 to 8 cigarettes per day | 8760
consumes strong alcoholic beverages in small doses | 8760
no clinical signs of exocrine and endocrine pancreatic insufficiency | 8760
does not use pancreatic enzyme supplementation | 8760