25 years old | 0
African American | 0
female | 0
admitted to the hospital | 0
found on the floor at home | -96
verbally incomprehensible | -96
complete bilateral vision loss | -96
altered mental status | -96
not eating well | -96
not taking medications | -96
systemic hypertension | -672
stage 4 chronic kidney disease | -672
idiopathic intracranial hypertension | -672
ventriculoperitoneal shunt | -672
hypertensive retinopathy | -672
optic neuropathy | -672
loss of peripheral vision in right eye | -672
loss of central vision in left eye | -672
medication non-compliance | -672
carvedilol | -672
nifedipine | -672
blood pressure 168/98 mmHg | 0
pulse 100 beats per minute | 0
incomprehensible | 0
minimally verbal | 0
obtunded | 0
total bilateral vision loss | 0
altered mental status | 0
left sided rib pain | 0
coughing | 0
head CT | 0
hypodensities in the cerebellum | 0
hyperdensities in the posterior occipital lobe | 0
brain MRI | 2
T2/FLAIR hyperintensity | 2
T1 hypointensity | 2
no restricted diffusion | 2
vasogenic edema | 2
cerebellum involvement | 2
posterior parietal and occipital lobes involvement | 2
blood urea nitrogen 92.0 mg/dL | 2
creatinine 17.56 mg/dL | 2
echocardiogram | 2
right-sided atrial septum vegetation | 2
culture-negative endocarditis | 2
blood cultures negative | 2
PRES diagnosis | 4
labetalol | 4
hydralazine | 4
clevidipine | 10
blood pressure control | 10
neurological examination checks | 10
VP shunt interrogation | 10
tunneled catheter | 12
dialysis treatment | 12
sevelamer carbonate | 12
vancomycin | 12
ceftazidime | 12
empiric antibiotic regimen | 12
regained baseline cognition | 24
regained vision | 24
cerebral metamorphopsia | 24
visual distortion | 24
cartoon-like vision | 24
no hallucinations | 24
resolved metamorphopsia | 168
follow-up MRI | 168
resolution of vasogenic edema | 168
discharged | 168