43 years old | 0
female | 0
admitted to the hospital | 0
behavioral abnormalities | -32400
depressed mood | -32400
dysphoria | -32400
easy irritability | -32400
difficulty to gain weight | -32400
sleep disorders | -32400
insomnia | -32400
increased prolactin levels | -32400
bradycardia | -32400
hypotension | -32400
hypoglycemia | -32400
sudden death of sister | -129600
behavioral problems in children | -129600
carbolithium treatment | -720
abnormal thinking | -720
personality changes | -720
poor concentration | -720
confusion | -720
memory impairment | -720
anxiety | -720
poor judgment | -720
on carbolithium treatment | -720
acute onset of permanent dystonic posture | -216
numbness | -216
tingling | -216
diplopia | -216
low potassium levels | -216
admitted to neurology unit | -216
treated with muscle relaxants | -216
treated with potassium | -216
neurological bladder | -192
catheterized | -192
discharged | -192
olanzapine treatment | -168
psychosis worsening | -168
difficulty in walking | -168
confined to bed | -168
sacral decubitus | -168
fever | -168
increased difficulty in movements | -168
low potassium levels | -168
admitted to neurology unit | -168
marked bradycardia | -168
atrial fibrillation | -168
ventricular fibrillation | -168
lost consciousness | -168
orotracheal intubation | -168
transferred to intensive care unit | -168
involuntary parossistic eye movements | 0
involuntary parossistic head movements | 0
bilateral ptosis | 0
oculogyric crises | 0
dystonia of the head | 0
generalized muscle hypotrophy | 0
absent deep tendon reflexes | 0
no pathological reflexes | 0
hemocromocytometric test | 0
biochemical parameters | 0
urine analysis | 0
electroencephalography | 0
diffuse theta mixed to paroxysmal activities | 0
brain MRI | 0
symmetric hyperintense lesions | 0
restricted diffusion | 0
globus pallidus | 0
untreatable bradycardia | 24
fever | 24
blood tests | 24
white blood count | 24
pancytopenia | 48
procalcitonin increase | 48
hemocultures | 48
Enterococcus faecalis | 48
Acinetobacter baumanii | 48
tigecycline | 48
colistin | 48
sedation | 72
whole exome sequencing | 72
p.Ser250Phe mutation | 72
DDC gene | 72
heterozygous state | 72
pyridoxine treatment | 96
pramipexole treatment | 96
death | 120
autopsy | 120
sepsis | 120
no macro- and microscopic brain abnormalities | 120