7 years old | 0
male | 0
admitted to the hospital | 0
non-productive cough | -720
asthma | -720
albuterol inhaler use | -720
non-bloody emesis | -672
non-bilious emesis | -672
temperature of 104 | -672
decreased appetite | 0
4 pound weight loss | 0
denial of pets | 0
denial of recent travel | 0
denial of sick contacts | 0
denial of foreign or new foods |#0
denial of animal or insect bites | 0
denial of fevers | 0
denial of diarrhea | 0
denial of constipation | 0
denial of chills | 0
well-controlled asthma | -2160
albuterol as needed | -2160
last albuterol use over three months ago | -2160
fully immunized | 0
no allergies to medications | 0
unremarkable family history | 0
previous normal growth and development | 0
no surgical history | 0
non-tender lymphadenopathy | 0
palpable lymphadenopathy | 0
mobile lymphadenopathy | 0
right submental lymph node (1 cm) | 0
anterior cervical lymph node (0.7 cm) | 0
bilateral supraclavicular lymph nodes (0.5 cm) | 0
clear lung auscultation | 0
para-tracheal mass on chest radiograph | 0
transfer to higher level of care | 0
CT scan showing paratracheal mass | 0
supraclavicular lymph nodes | 0
differential diagnosis: teratoma | 0
differential diagnosis: thymoma | 0
differential diagnosis: lymphoma | 0
differential diagnosis: thyroid related tumor | 0
differential diagnosis: granulomatous process | 0
transfer to hematology/oncology service | 0
extensive laboratory evaluation | 0
ceftriaxone started | 0
pediatric surgery consultation | 0
infectious disease consultation | 0
white blood cell count 6.8 ×10³/mL | 0
hemoglobin 11.5 g/dL | 0
platelets 307 ×10³/mL | 0
neutrophil 23% | 0
lymphocytes 46% | 0
monocytes 12% | 0
eosinophils 18% | 0
ESR 30 mm/hr | 0
CRP <0.012 mg/dL | 0
LDH 197 U/L | 0
uric acid 2.7 mg/dL | 0
unremarkable comprehensive metabolic panel | 0
unremarkable glucose | 0
unremarkable bilirubin | 0
unremarkable urinalysis | 0
unremarkable TSH/T4 | 0
unremarkable HIV | 0
unremarkable PPD | 0
unremarkable homovanillic acid | 0
unremarkable vanillylmandelic acid | 0
unremarkable angiotensin converting enzyme | 0
unremarkable ANCA | 0
MRI of the brain normal | 0
blood cultures negative | 0
stool cultures negative | 0
serum cryptococcal antigen positive (1:20) | 0
repeat cryptococcal antigen undetectable | 72
histoplasmosis H band negative | 0
histoplasmosis M band antibody present | 0
chronic infection with histoplasmosis (last 6 months to 3 years) | 0
thoracotomy performed | 0
purulent fluid obtained | 0
cultures sent | 0
mediastinal lymph node biopsies | 0
right upper lung lobe biopsy | 0
mediastinal nodule biopsy | 0
mediastinal mass biopsy | 0
post-op pneumothorax | 0
right-sided chest tube | 0
transfer to pediatric intensive care unit | 0
return to OR for spinal tap | 0
cerebral spinal fluid analysis: colorless clear fluid | 0
cerebral spinal fluid: one red blood cell | 0
cerebral spinal fluid: one white blood cell | 0
cerebral spinal fluid: 85 lymphocytes | 0
cerebral spinal fluid: 15 monocytes | 0
cerebral spinal fluid: negative Indian ink stain | 0
cerebral spinal fluid: negative bacterial culture | 0
cerebral spinal fluid: negative fungal culture | 0
biopsy results unclear | 0
confirmation of histoplasmosis | 0
necrotizing granulomatous inflammation | 0
calcification | 0
histoplasmosis mediastinal granuloma diagnosis | 0
start of itraconazole course | 0
pain control with Hydrocodone/Acetaminophen | 0
pain control with Ketorolac | 0
incentive spirometry | 0
serial chest x-rays showing improvement | 0
chest tube set to water seal | 0
chest tube removal | 288
intermittent fevers | 0
cultures negative at discharge | 0
afebrile >24 hours prior to discharge | 0
exposure to dirt | 0
possible histoplasma inoculation | 0
denial of living near demolition or construction sites | 0
lack of H bands | 0
calcifications on biopsy | 0
mass size 3.1×2.7×3.7 cm | 0
discharge after 12 days | 288
repeat serum cryptococcal antigen test at one week post discharge | 360
compliant to itraconazole course | 288
itraconazole level monitoring | 336
itraconazole dose adjustment | 336
