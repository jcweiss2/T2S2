81 years old | 0
male | 0
admitted to the hospital | 0
inginoscrotal hernia | -672
auricular fibrillation | -672
chronic heart failure | -672
chronic renal dysfunction | -672
upper abdominal pain | 0
temperature 36.1 °C | 0
abdominal distention | 0
tenderness of the epigastric area | 0
bilateral giant inguinoscrotal hernia | 0
white blood cell count 4900/mm2 | 0
C-reactive protein 1.2 mg/dl | 0
creatinin 1.71 mg/dl | 0
prothrombin 18.7 s | 0
PT-INR 1.61 | 0
computed tomography scan | 0
slightly dilated stomach | 0
dilated jejunum | 0
large bilateral inguinoscrotal hernia | 0
small bowel in hernia sac | 0
cecum in hernia sac | 0
ascending colon in hernia sac | 0
sigmoid colon in hernia sac | 0
acute entire abdominal pain | 48
decreased blood pressure | 48
free air in the right inguinal hernia sac | 48
much ascites | 48
emergency operation | 48
diagnosis of acute generalized peritonitis | 48
small bowel perforation in the inguinal hernia sac | 48
general anesthesia | 48
mid-lower median abdominal incision | 48
transverse incision at the right inguinal area | 48
dirty ascites in the inguinal sac | 48
perforated cecum | 48
necrotic terminal ileum | 48
rupture of the inferior duodenum angle | 48
right hemicolectomy | 48
side-to-side anastomosis of duodenum and jejunum | 48
primary closure of the peritoneum at the hernia gate | 48
transferred to intensive care unit | 48
septic shock | 72
leakage of the duodenum–jejunum anastomosis | 72
antibiotic agents | 72
vasopressure agent | 72
continuous hemodiafiltration | 72
death | 432