39 years old | 0
female | 0
ingested caffeine tablets | -1
generalized tonic–clonic seizure | -1
broad complex tachycardia | -1
cardiopulmonary resuscitation | -1
defibrillations | -1
epinephrine | -1
amiodarone | -1
intubated | 0
sinus rhythm | 0
blood pressure 62/33 mmHg | 0
heart rate 140/min | 0
activated charcoal | 0
multiple ventricular extrasystoles | 0
intravenous magnesium | 0
intravenous calcium | 0
hypotension | 0
crystalloids | 0
epinephrine boluses | 0
continuous infusion | 0
lactic acidosis | 0
intravenous sodium bicarbonate | 0
haemodialysis | 5
blood samples drawn | 5
serum caffeine concentrations measured | 5
recurrent cardiovascular instability | 5
concomitant lactic acidosis | 5
dobutamine | 5
hypotension | 5
rhabdomyolysis | 5
acute renal failure | 48
creatinine kinase max 69 885 U/L | 48
aspartate transaminase max 1908 U/L | 48
volume overload | 48
persistent haemodynamic instability | 48
chronic veno-venous haemodiafiltration (CVVHDF) | 48
pending serum caffeine concentration measurements reported | 72
daily haemodialysis therapy recommenced | 72
pulmonary failure | 120
tricuspid endocarditis | 120
line sepsis | 120
renal function improved | 336
haemodialysis therapy stopped | 336
total of 14 haemodialysis sessions | 336