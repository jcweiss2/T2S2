33 years old | 0
female | 0
admitted at 19 wk gestation | 0
fever | -504
chills | -504
hospitalized at 14 wk gestation | -1176
dry cough | -1176
empirical antibiotic treatment (ceftriaxone, azithromycin) | -1176
intermittent mild fever (37.5C-38.0C) | -672
contact dermatitis of both hands | -?
steroid ointment application | -?
blister on contact dermatitis | -1176
antibiotic ointment application | -1176
healed blisters | -1176
anesthesiology resident | -?
worked in intensive care units | -?
rounding patients | -?
endotracheal intubation | -?
central venous catheterization | -?
physical examination unremarkable | 0
no abdominal pain | 0
no urinary symptoms | 0
vaginal examination showed no leaking amniotic fluid | 0
increased white blood cell count | 0
high CRP (15.8 mg/dL) | 0
elevated procalcitonin (0.503 ng/mL) | 0
normal thyroid function | 0
normal liver function | 0
normal renal function | 0
normal coagulation profile | 0
normal electrolytes | 0
normal lactate levels | 0
normal vaginal PCR for STDs | 0
normal rheumatological studies | 0
blood cultures grew S. marcescens | 48
abdominal ultrasonography nonspecific | 0
gallbladder polyp | 0
normal fetus | 0
normal placenta | 0
normal obstetric ultrasonography | 0
normal abdominal MRI | 0
normal pelvic MRI | 0
S. marcescens bacteremia diagnosis | 48
chorioamnionitis diagnosis | 336
empirical cefepime IV | 0
ceftriaxone IV | 48
fever recurrence | 96
cefepime resumed | 96
watery discharge | 552
PPROM diagnosis | 552
cefepime IV | 552
clarithromycin PO | 552
induced labor | 552
delivered dead fetus | 552
afebrile | 768
normalized leukocytosis | 768
normalized CRP | 768
discharged | 768
placenta culture grew S. marcescens | 768
chorioamnionitis with focal infarct | 768
miscarriage | 552
