61 years old | 0
male | 0
admitted to the hospital | 0
persistent productive cough | -360
chills | -360
fever | -360
aminophylline | -360
deflazacort | -360
formoterol + budesonide fumarate | -360
amoxicillin + clavulanate potassium | -240
clarithromycin | -196
blood tests | 0
computed tomography scan of the chest | 0
elevation of C-reactive protein | 0
leukocytosis | 0
lymphopenia | 0
BSR elevation | 0
centrilobular nodular opacities | 0
bronchi with thickened walls | 0
facial glass nodular opacities | 0
non-calcified nodular opacities | 0
opacity in a fibroatelectasic range | 0
absence of lymphadenomegaly | 0
absence of pleural effusion | 0
sputum examination | 0
Stenotrophomonas maltophilia identified | 0
sensitivity to levofloxacin | 0
sensitivity to sulfamethoxazole/trimethoprim | 0
treatment with levofloxacin | 0
resolution of cough | 360 
no shortness of breath | 0
no comorbidities | 0 
no malignancy | 0
no organ transplantation | 0
no HIV infection | 0
no chronic obstructive pulmonary disease | 0
no cystic fibrosis | 0
no prolonged hospital stay | 0
no intensive care unit admission | 0
no mechanical ventilation | 0
no permanent catheter therapy | 0
no corticosteroid or immunosuppressive therapy | 0 
no recent antibiotic treatment | 0