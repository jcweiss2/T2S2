20 years old | 0
male | 0
arrived at the emergency department | 0
fever | -336
productive cough | -336
night sweats | -336
malaise | -336
myalgia | -336
non-smoker | 0
occupational smoke exposure | 0
policeman in region with domestic waste burning | 0
treated with roxithromycin | -168
temperature 38.4°C | 0
blood pressure 130/70 mmHg | 0
pulse 88 bpm | 0
oxygen saturation 97% | 0
dyspnoea | 0
tachypnoea |0
bronchial breathing sounds |0
crackles over right lung |0
white blood cells 11.54×10³/μl |0
total eosinophils 92×10⁴/μl |0
haemoglobin 13.7 g/dl |0
creatinine 1.1 mg/dl |0
C-reactive protein 11 mg/dl |0
elevated liver enzymes |0
ALP 524 |0
GGT 320 |0
ALT 406 |0
AST 137 |0
normal abdominal ultrasound |0
chest radiograph infiltrates right lung |0
IV cefuroxime initiated |0
negative blood cultures |48
negative sputum cultures |48
negative urine Legionella antigen test |48
persistent high-grade fever |48
antibiotic treatment changed to moxifloxacin |48
sterile blood cultures |48
respiratory distress |96
persistent fever |96
oxygen saturation 88% |96
PaO2 67 mmHg |96
CRP 14 mg/dl |96
elevated liver enzymes |96
leucocytosis 12.8×10³/μl |96
eosinophil count 1.33×10³/μl |96
chest radiogram bilateral infiltrates |96
respiratory distress worsened |120
intubated |120
mechanically ventilated |120
transferred to intensive care unit |120
broncho-alveolar lavage 30% eosinophils |144
diagnosis of AEP |144
IV glucocorticoids administered |144
prompt improvement |144
resolution of fever |144
successful extubation |168
chest radiogram regression infiltrates |168
eosinophil count 260/μl |168
discharged |192
oral prednisone 60 mg/day |192
tapering over 3 months |192
elevated eosinophil count during deterioration |96
rapid decrease eosinophil count after glucocorticoids |144
no long-term pulmonary complications |192
