48 years old | 0
male | 0
seizure disorder | -8760
antiepileptics | -8760
valproic acid | -8760
carbamazepine | -8760
clobazam | -8760
type-2 diabetes mellitus | -8760
hypertension | -4380
impaired level of consciousness | -24
admitted to critical care unit | 0
blood pressure 160/100 mmHg | 0
heart rate 96/min | 0
respiratory rate 22/min | 0
Glasgow coma score 11 | 0
poor coughing | 0
coarse crepts on right base | 0
intubated | 0
mechanical ventilation | 0
antiepileptics stopped | 0
intravenous infusion of propofol | 0
elevated creatinine | 0
BUN 40 mg/dl | 0
blood sugar 176 mg/dl | 0
total leukocyte count 11,400 | 0
liver function test | 0
ultrasound abdomen | 0
medical renal disease | 0
serum creatinine 2.1 mg/dl | -2160
MRI head | 0
cerebrospinal fluid analysis | 0
electroencephalogram | 0
continuous generalized slowing | 0
uremic encephalopathy | 0
hemodialysis | 0
BUN level 68 mg/dl | 0
BUN level 21 mg/dl | 24
ammonia level 274 μmol/L | 24
valproate-induced hyperammonemic encephalopathy | 24
L-carnitine | 24
refractory septic shock | 168
ICU-acquired multidrug resistant infection | 168
death | 168