43 years old | 0
female | 0
weight gain | -720
leg edema | -720
nephrotic syndrome | -720
admitted to hospital | 0
minimal change nephrotic syndrome | 0
steroid therapy | 0
steroid pulse | 0
prednisolone | 0
fever | 168
acute kidney injury | 168
drowsy | 168
blood pressure 121/93 mmHg | 168
pulse rate 80/min | 168
body temperature 36.8°C | 168
bilateral lower extremity edema | 168
no chest pain | 168
no abdominal tenderness | 168
high inflammation | 168
abnormal cardiac biomarkers | 168
renal dysfunction | 168
CRP 48.93 mg/dL | 168
Alb 1.4 g/dL | 168
CK 2529 mg/dL | 168
CK-MB 196 mg/dL | 168
Cr 3.75 mg/dL | 168
troponin-T 14.19 ng/mL | 168
PCT 100 ng/mL | 168
marked proteinuria | 168
ST-elevation | 168
pleural effusion | 168
reduced wall motion of the left ventricle | 168
ejection fraction 30% | 168
hypokynesis | 168
severe respiratory distress | 192
pulmonary congestion | 192
anuria | 192
non-invasive positive pressure ventilation | 192
continuous hemodiafiltration | 192
Meropenem | 192
Levofloxacin | 192
Escherichia coli | 192
sepsis | 192
calcification | 216
Warfarin | 336
remission of MCNS | 720
reduction in prednisolone | 720
discharged | 912
follow-up with CT | 912
calcification | 912
impaired cardiac function | 912
EF 46% | 912
MRI | 912
wall motion impaired | 912
Late Gadolinium Enhancement | 912
myofiber fibrosis | 912
follow-up with CT | 8760
calcification | 8760
improved cardiac function | 8760
EF 60.6% | 8760
wall motion not fully recovered | 8760