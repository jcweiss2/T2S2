39 years old | 0
male | 0
ulcerative colitis | -87600
sclerosing cholangitis | -87600
admitted to the hospital | 0
elective liver transplantation |DISCUSSION
azathioprine | -87600
ursacol | -87600
prednisone | -87600
simvastatin | -87600
spironolactone | -87600
folic acid | -87600
calcium carbonate | -87600
general condition good | 0
healthy skin tone | 0
well hydrated | 0
feverless | 0
jaundiced +++/IV | 0
stable vital signs | 0
target painless hepatomegaly | 0
spider veins | 0
lower limb edema | 0
high fever | 12
tachycardia | 12
myalgia in the calves | 12
anuria | 12
ceftriaxone | 12
lesions resembling purplish erythematous plaques | 12
rapid growth | 12
proximal progression | 12
recent trip to the coastal area of Paraná | -24
samples for leptospirosis | 12
samples for dengue | 12
samples for yellow fever | 12
samples for spotted fever | 12
samples for meningococcemia | 12
negative test results | 12
unresponsive to volume | 24
dyspnea | 24
respiratory distress | 24
transferred to the ICU | 24
vasoactive drugs | 24
mechanical ventilation | 24
clinical condition progressively worsened | 24
increased need for vasoactive drugs | 24
skin lesions became confluent | 24
blisters | 24
sero-sanguineous fluids discharge | 24
ceftriaxone changed to meropenem | 24
ceftriaxone changed to oxacillin | 24
blood cultures growth of gram-negative bacillus | 24
Vibrio vulnificus identified | 24
died | 30
gram-negative bacilli in subepidermal space | 12
gram-negative bacilli in splenic small vessels | 12
Vibrio vulnificus infection | 12
sepsis | 12
disseminated intravascular coagulation | 24
septic shock | 24
bullous cellulitis | 12
pain and swelling in affected limb | 12
rash | 12
bullous lesions with seroDISCUSSIONhemorrhagic fluids | 24
necrotizing fasciitis | 24
leukocytosis | 24
major shift to the left |
