12 years old | 0
male | 0
Tanzanian | 0
admitted to the hospital | 0
stung by numerous African bees | -1
stung on the face, upper limbs and trunk | -1
given IV fluids | 0
given hydrocortisone | 0
given diclofenac IM for pain | 0
facial edema | 0
decrease in urine output | 28
given furosemide | 28
referred to tertiary hospital | 28
conscious | 28
could not see well | 28
facial swelling | 28
peri-orbital edema | 28
erythema stings marks on face, trunk and upper limbs | 28
treated with broad spectrum antibiotic | 28
fluid restriction | 28
initial laboratory investigations | 28
creatinine 116 mmol/l | 28
urea 15.4 mmol/l | 28
hyperkalemia 6.9 mmol/l | 28
hyponatremia 128 mmol/l | 28
catheter inserted | 28
urine for dipstick showed RBC+++ | 28
microscopy examination revealed muddy brown cast | 28
leucocytosis 25 | 28
neutrophils 89.7% | 28
hemoglobin 13.8 g/dl | 28
platelet count 269 | 28
correction control electrolytes | 28
potassium 5.15 mmol/l | 28
sodium 128 mmol/l | 28
urine output 200 ml | 48
amber colored urine | 48
creatinine 248 mmol/l | 48
urea 22.52 mmol/l | 48
fluid input restricted to 700 ml | 48
close monitoring of input and output | 48
produced only 100 ml of urine | 60
creatinine 402 mmol/l | 60
urea 29.83 mmol/l | 60
potassium 5.4 mmol/l | 60
sodium 127 mmol/l | 60
transferred to pediatric intensive care unit | 60
hemodialysis considered | 60
initiation of hemodialysis | 72
potassium 5.99 mmol/l | 72
creatinine 462 mmol/l | 72
urea 34.65 mmol/l | 72
five sessions of hemodialysis | 72
high grade fever 38.6°C | 96
blood cultures collected | 96
vancomycin administered | 96
cultures were all negative | 168
urine output raised to 1.8 ml/kg/h | 168
creatinine 172 mmol/l | 168
urea 11 mmol/l | 168
electrolytes normal | 168
discharged | 336
follow-up after discharge | 504
biochemistry back to normal | 504
creatinine 52 mmol/l | 504
urea 2.96 mmol/l | 504
electrolytes normal | 504