65 years old | 0
male | 0
hypertension | 0
depression | 0
fever | -168
malaise | -168
chest x-ray | -168
COVID swab | -168
dental work | -192
presented to ambulatory respiratory care unit | 0
referred to emergency department | 0
temperature 97.7 Fahrenheit | 0
heart rate 63 beats per minute | 0
blood pressure 74/44 mmHg | 0
respiratory rate 20 breaths per minute | 0
oxygen saturation 99% | 0
crackles at the right lung base | 0
holosystolic murmur | 0
AST 89 IU/L | 0
ALT 103 IU/L | 0
proBNP 16093 pg/mL | 0
Troponin-T 0.79 ng/mL | 0
CRP > 300 mg/L | 0
creatinine 2.6 mg/dL | 0
lactate 3.4 mmol/L | 0
atrial fibrillation | 0
intraventricular conduction delay | 0
ST elevation | 0
preserved LVEF | 0
tricuspid regurgitation | 0
no pericardial effusion | 0
gram-positive cocci | 0
coagulase-negative staphylococcus | 0
CT angiogram negative for pulmonary embolism | 0
negative urine antigens | 0
LVEF 54% | 24
dilated right ventricle | 24
RV systolic dysfunction | 24
TAPSE 1.3 cm | 24
leftward interventricular septal shift | 24
tricuspid regurgitation | 24
no significant left-sided valvular disease | 24
no pericardial effusion | 24
admitted to medical ICU | 24
administered IV fluids | 24
vasopressors | 24
empiric antibiotics | 24
vancomycin | 24
ceftriaxone | 24
doxycycline | 24
unfractionated heparin | 24
fever abated | 32
blood pressure stabilized | 32
vasopressors weaned | 32
renal function improved | 32
peak troponin-T 1.24 | 36
peak CK-MB 57 | 36
coronary angiography | 96
no obstructive coronary artery disease | 96
CMR imaging myopericarditis | 120
pericardial effusion | 120
sub-epicardial late gadolinium enhancement | 120
anaplasma serology positive | 144
anaplasma PCR positive | 144
discharged | 144
doxycycline | 144
followed up with infectious disease | 336
stopped antibiotics | 336
repeat CMR | 336
followed up with heart failure | 672
sinus rhythm | 672
no atrial fibrillation | 672
no high-grade heart block | 672
LVEF 59% | 672
normal RV size | 672
resolution of pericardial effusion | 672
normal T2 signal | 672
no dyspnoea | 672
no chest pain | 672
