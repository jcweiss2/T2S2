57 years old | 0 | 0 
Hispanic | 0 | 0 
male | 0 | 0 
admitted to the hospital | 0 | 0 
history of coronary artery disease | -6336 | 0 
history of myocardial infarction | -6336 | 0 
history of ischemic dilated cardiomyopathy | -6336 | 0 
pocket infection of his cardiac resynchronization therapy defibrillator | -48 | 0 
erythema around his left upper chest implant site | -144 | -48 
discomfort around his left upper chest implant site | -144 | -48 
edema around his left upper chest implant site | -48 | -48 
serosanguinous drainage around his left upper chest implant site | -48 | -48 
oral amoxicillin treatment | -48 | 0 
nonbacteremic | 0 | 0 
afebrile | 0 | 0 
laboratory investigations within normal limits | 0 | 0 
severely reduced left ventricular systolic function | 0 | 0 
ejection fraction of 20%–25% | 0 | 0 
global hypokinesis of the left ventricle | 0 | 0 
no evidence of vegetations | 0 | 0 
leads scarred to the lateral wall of the superior vena cava | 0 | 0 
transvenous lead extraction | 0 | 24 
cardiac resynchronization therapy defibrillator pocket capsule dissected out | 0 | 1 
device removed | 0 | 1 
coronary sinus and right atrial leads extracted | 0 | 2 
right ventricular lead extracted | 0 | 2 
hypotensive | 2 | 2 
transesophageal echocardiography revealed a large pericardial effusion | 2 | 2 
emergency midsternotomy | 2 | 3 
pericardium opened | 2 | 3 
significant amount of blood seen | 2 | 3 
bleeding manually controlled with pressure | 2 | 4 
cardiopulmonary bypass instituted | 4 | 24 
5-mm tear in the superior cavoatrial junction | 4 | 4 
perforation in the right atrium | 4 | 4 
oozing hematoma at the level of the innominate vein | 4 | 4 
lesions repaired with multiple 4-0 polypropylene sutures | 4 | 6 
right ventricular lead capped and abandoned | 6 | 6 
intra-aortic balloon pump placed | 6 | 168 
coagulopathy | 6 | 24 
transfusions of cryoprecipitate, platelets, fresh frozen plasma, and factor VII | 6 | 24 
chest closed | 24 | 24 
transferred to the intensive care unit | 24 | 24 
severe cardiogenic shock | 24 | 168 
multiorgan failure | 24 | 168 
hypotensive | 24 | 168 
required large doses of vasopressin, epinephrine, and norepinephrine | 24 | 168 
hypoxic respiratory failure | 24 | 168 
mechanical ventilation | 24 | 168 
liver failure | 24 | 168 
albumin | 24 | 168 
blood products given | 24 | 168 
broad-spectrum antibiotics | 24 | 168 
oliguric | 24 | 168 
continuous venovenous hemodialysis | 24 | 408 
bilateral, symmetrical cyanotic changes to all 5 digits of his upper and lower extremities | 48 | 216 
vasopressor administration stopped | 48 | 48 
upper- and lower-digit ischemia progressed to dry gangrene | 216 | 216 
dull pain | 216 | 216 
no ability to move his fingers and toes | 216 | 216 
bilateral stiffness | 216 | 216 
2+ pitting edema | 216 | 216 
nonexistent capillary refill time | 216 | 216 
palpable 2+ peripheral pulses | 216 | 216 
Doppler study showed flat waveforms on all digits and toes bilaterally | 216 | 216 
no proximal occlusion or stenosis | 216 | 216 
intra-aortic balloon pump removed | 168 | 168 
endotracheal tube removed | 168 | 168 
albumin discontinued | 240 | 240 
liver enzymes returned to normal limits | 240 | 240 
kidney function gradually improved | 240 | 408 
hemodialysis stopped | 408 | 408 
mental status improved | 240 | 408 
necrotic lesions treated conservatively with povidone-iodine dressings | 240 | 408 
debridement | 312 | 312 
negative-pressure wound therapy | 312 | 408 
purulent, foul-smelling material from his left infraclavicular operative site | 408 | 408 
transferred to our facility | 408 | 408 
preoperative transesophageal echocardiography | 408 | 408 
diminished ejection fraction of 10%–15% | 408 | 408 
laser extraction of his retained lead | 432 | 432 
pus drained from the subfascial area | 432 | 432 
antibiotic regimen | 432 | 432 
microbial cultures grew Enterobacter cloacae and Staphylococcus epidermidis | 432 | 432 
transvenous implantable cardioverter-defibrillator system implanted | 448 | 448 
evaluation of his hands and feet | 448 | 448 
no signs of local infection or wet gangrene | 448 | 448 
black skin changes and demarcation lines | 448 | 448 
frank mummification of his digits and toes | 448 | 448 
discharged to home health services | 552 | 552 
amputation and debridement of his necrotic feet | 760 | 760 
amputation of his fingers scheduled | 760 | 760