63 years old | 0
man | 0
history of smoking | 0
hypertension | 0
vascular disease | 0
diagnosis of clinically T3 | -2160
diagnosis of N3 | -2160
diagnosis of M0 | -2160
diagnosis of poorly differentiated adenocarcinoma | -2160
right upper lobe | -2160
stage IIIB | -2160
concurrent chemoradiation | -2160
3 courses carboplatin/etoposide chemotherapy | -2160
60 Gy radiation therapy | -2160
dysphagia grade 3 | -1680
weight loss | -1680
gastroscopy | -1680
radiation esophagitis | -1680
stenosis | -1680
nasogastric tube placement | -1680
tube feeding | -1680
presented at emergency room | -1680
sepsis | -1680
acute dyspnea | -1680
right sided thoracic pain | -1680
reduced right sided airflow | -1680
tachycardia | -1680
hypotension | -1680
saturation of 85% | -1680
C-reactive protein of 348 mg/L | -1680
leukocytosis of 24.8 × 10^9/L | -1680
chest x-ray showing atelectasis | -1680
right sided pleural effusion | -1680
CT scan showing mediastinal air configuration | -1680
admitted to intensive care unit | -1680
acute respiratory failure | -1680
sepsis due to pneumonia | -1680
empyema | -1680
noninvasive ventilation | -1680
intravenous broad-spectrum antibiotics | -1680
fluid resuscitation | -1680
bronchoscopy revealing bronchopleural fistula | -1680
20 French chest tube placement | -1680
repeated CT scan after 10 days | -1680
decrease of empyema | -1680
consolidations | -1680
mediastinal air configuration unchanged | -1680
no signs of cancer recurrence | -1680
multidisciplinary consultation | -1680
enteral feeding | -1680
antibiotics for intrapulmonary consolidations | -1680
surgical coverage with latissimus dorsi flap | -1680
no respiratory support required | -1680
no fever | -1680
low infection parameters | -1680
improved nutritional status | -1680
operation performed | 0
latissimus dorsi muscle flap harvested | 0
thoracotomy in fifth intercostal space | 0
lung adhesive to thoracic wall | 0
inflammation | 0
fibrosis of mediastinum | 0
salvage pneumonectomy considered | 0
latissimus dorsi flap fixated dorsally to bronchus | 0
insignificant air leak | 0
full coverage of defect | 0
28 French intrathoracic chest tube placement | 0
lung reinsufflated | 0
no air leakage | 0
wound closure | 0
recovery after 6 days | 168
transferred to surgical ward | 168
limited air leakage for 8 days | 192
drain removed | 240
dismissed to rehabilitation center | 360
readmitted after 10 weeks | 1680
hemoptysis | 1680
pneumonia | 1680
anemia | 1680
bronchoscopy showing large defect | 1680
palliative care started | 1680
died | 2400
