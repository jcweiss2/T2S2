21 years old | 0
female | 0
admitted to the hospital | 0
dyspnea | -48
fever | -48
malaise | -48
lymphadenopathy | -48
axillary lymphadenopathy | 0
cervical lymphadenopathy | 0
inguinal lymphadenopathy | 0
multifocal pneumonia | 0
treatment for community-acquired pneumonia | 0
ceftriaxone | 0
azithromycin | 0
oxygen therapy | 0
mechanical ventilation | 24
computerized tomography chest | 24
bilateral lung consolidation | 24
pericardial effusion | 24
HIV test | 24
streptococcus pneumonia test | 24
legionella test | 24
histoplasma test | 24
brucella test | 24
aspergillus test | 24
tuberculosis test | 24
influenza test | 24
respiratory syncytial virus test | 24
mycoplasma IgM test | 24
chlamydia antibody titer test | 24
bronchoscopy | 48
bronchoalveolar lavage | 48
transthoracic echocardiogram | 48
cervical lymph node biopsy | 72
histopathology | 72
septic work up | 72
blood cultures | 72
sputum cultures | 72
urine cultures | 72
high dose steroids | 96
intravenous immune globulin | 96
hemolytic work up | 120
haptogobin test | 120
schistocytes test | 120
thrombocytopenia | 120
partial thromboplastin time test | 120
prothrombin time test | 120
D-dimer test | 120
fresh frozen plasma | 144
disseminated intravascular coagulopathy | 168
death | 168
Kikuchi-Fujimoto disease | 0 
lymphoma | 0 
tumor necrosis factor-alpha | 0 
interleukin-1 | 0 
interleukin-6 | 0 
cytokine release | 0 
hydroxychloroquine | 0 
relapse | 0 
sepsis | 0 
acute myeloid leukemia | 0 
verbal consent | -24 
informed consent | -24 
conflict-of-interest statement | -24 
institutional review board statement | -24 
peer-review report classification | -24 
peer-review started | -744 
first decision | -624 
article in press | -408 
P- Reviewer | -24 
S- Editor | -24 
L- Editor | -24 
E- Editor | -24