22 years old | 0
male | 0
Hispanic | 0
admitted to the hospital | 0
intermittent fevers | -336
headache | -336
fatigue | -336
malaise | -336
nausea | -336
vomiting | -336
diarrhea | -336
nosebleeds | -336
non-productive cough | -336
sore throat | -336
light sensitivity | -336
rash | -72
petechial rash | 0
no shortness of breath | 0
no chest pain | 0
no bloody stools | 0
no neck stiffness | 0
worked as a taxidermist | -72
had a cat | -672
had two dogs | -672
fleas in home | -672
seen rats in home | -672
afebrile | 0
blood pressure 97/47 | 0
pulse rate 136 | 0
respiratory rate 22 | 0
hyponatremic | 0
elevated BUN | 0
elevated creatinine | 0
elevated AST | 0
elevated ALT | 0
elevated ALP | 0
elevated D-dimer | 0
low fibrinogen | 0
elevated lactic acid | 0
thrombocytopenia | 0
elevated WBC | 0
diagnosed with severe sepsis | 0
diagnosed with DIC | 0
treated with vancomycin | 0
treated with ceftriaxone | 0
lumbar puncture not performed | 0
seen by infectious diseases specialist | 24
diagnosed with murine typhus | 24
treated with doxycycline | 24
Rickettsia typhi titers positive | 24
cryoprecipitate administered | 24
fever resolved | 48
transferred out of MICU | 72
repeat infection work-up | 120
Rickettsia typhi serum antibody titers high | 120
discharged | 120
improvement in symptoms | 120