65 years old | 0
female | 0
admitted to the hospital | 0
fever | -744
nausea | -168
vomiting | -168
neutrophil count 6.96×10^9/L ↑ | 0
monocyte count 0.86×10^9/L ↑ | 0
lymphocyte percentage 14.9% ↓ | 0
red blood cell count 3.17×10^12/L ↓ | 0
hemoglobin content 87 g/L ↓ | 0
hematocrit 0.28 L/L ↓ | 0
average red blood cell hemoglobin concentration 312 g/L ↓ | 0
platelet count 363×10^9/L ↑ | 0
platelet distribution width 8.3 fl ↓ | 0
C-reactive protein (CRP) 52.01 mg/L ↑ | 0
secondary infectious thrombocytopenia | 0
gram-negative bacilli septicemia (Klebsiella pneumoniae) | 0
liver abscess | 0
bilateral lung inflammation | 0
type 2 diabetes | 0
hypertension grade 3 (extremely high risk) | 0
vancomycin | 0
caspofungin | 0
dexamethasone | 0
posaconazole oral suspension | 0
liver abscess puncture and drainage treatment | 0
light perception disappeared in the left eye | 72
eyelid redness and pain | 72
purulent secretion | 72
repeated fever | 72
left-sided headache | 72
endogenous endophthalmitis (left) | 72
orbital cellulitis (left) | 72
rubeosis iridis (left) | 72
exudative retinal detachment (left) | 72
diabetic retinopathy (right) | 72
intravitreal injection with vancomycin and ceftazidime | 72
left eyeball enucleation | 336
fever | 336
moxifloxacin | 336
sulperazon | 336
inflammation of both lungs | 432
pericardial effusion | 432
bilateral pleural thickening and effusion | 432
atelectasis in right inferior lobe | 432
liver cyst | 432
liver abscess | 432
right renal cyst | 432
myoma of the uterus | 432
convulsion with unconsciousness | 480
lacunar infarction | 480
encephalomalacia | 480
bilateral pleural effusion | 480
intracranial infection | 480
lumbar puncture | 480
cerebrospinal fluid (CSF) biochemistry analysis | 480
microbial metagenomic next-generation sequencing (mNGS) | 480
glucose <1.1 mmol/L ↓ | 480
chlorine 108 mmol/L ↓ | 480
CSF protein >3,000 mg/L ↑ | 480
Klebsiella pneumoniae with drug-resistant gene blaSHV | 480
meropenem | 480
pulmonary edema | 744
pleural effusion | 744
discharged from the hospital | 744