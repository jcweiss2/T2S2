55 years old | 0
man | 0
resection of a right adrenal tumor | -87600
right adrenal tumor | -87600
excessive secretion of aldosterone | 0
excessive secretion of cortisol |D0
excessive secretion of catecholamines |D0
excessive secretion of sexual hormones |D0
monoclonal gammapathy |D0
mass (diameter 10.6 cm) |D-87600
post-traumatic hematuria |D-87600
normal blood pressure |D-87600
stage II tumor (> 5 cm) |D-87600
anesthetic procedure |D-87600
surgical procedure |D-87600
annual follow-up (computed tomography and PET) |D-87600
asymptomatic until January 2019 |0
liver enzymes disturbances |0
large intrahepatic mass (14.4 × 12.6 cm) |0
FDG-18 PET-scan |0
liver biopsy |0
molecular research assay |0
surgical resection of intrahepatic tumor |0
pre-anesthetic visit |0
normal arterial blood pressure (133/73 mmHg) |0
normal heart rate (58/min) |0
laboratory investigations for abnormal endocrine hormonal secretion |0
biomarkers of liver cancer |0
induction of anesthesia |0
maintenance with sevoflurane |0
mobilization of the right liver |0
severe adhesions between liver and vena cava |0
bleeding at hepatico-caval small vessels |0
hypotension |0
blood transfusions (1347 mL) |0
norepinephrine infusion (up to 0.65 μg/kg/min) |0
parenchymal transection |0
portal vein not opened |0
hepatic vein not opened |0
residual bleeding not present |0
cristalloids (6000 mL) |0
colloids (2000 mL) |0
oxygen saturation no changes |0
end-tidal carbon dioxide no changes |0
arrival in ICU |0
norepinephrine infusion rate (2 μg/kg/min) |0
arterial blood pressure dependent on fluid replacement |0
cristalloids (16000 mL over 8 hours) |0
hemoglobin concentration (8.4 g/dL to 11.5 g/dL) |0
total plasma protein concentration (14 g/L) |0
refractory vasoplegic shock |0
transthoracic echocardiography |0
well preserved left ventricular function |0
low filling pressures |0
fluids received (47000 mL over first postoperative day) |0
vasopressors (norepinephrine up to 5 μg/kg/min) |0
methylprednisolone |0
ventilation with 1.0 FiO2 |0
generalized edema |0
anuric renal failure |0
lactic acidosis |0
four-limb ischemia |0
rhabdomyolysis |0
abdominal compartment syndrome (ACS) |0
bladder pressure >20 mm Hg |0
multiple organ dysfunction |0
second laparotomy for ACS decompression |0
no acute liver failure |0
no intestinal ischemia |0
postoperative day 7 |168
hemodynamic improvement |168
decrease of vasopressors |168
decrease of lactic acidosis |168
blood cultures positive for Escherichia coli |168
no evidence of intestinal ischemia |168
no evidence of perforation |168
refractory septic shock |168
acute respiratory distress syndrome |168
died on postoperative day 9 |216
determination of catecholamines impossible |0
determination of cortisol concentration impossible |0
immunohistochemical features of intrahepatic tumor similar to primary adrenal tumor |0
Ki67 index >30% |0
metastatic adrenocortical carcinoma |0
postmortem examination findings |216
acute tubular necrosis |216
centrilobular liver necrosis |216
hemorrhagic necrosis of the spleen |216
lung congestion |216
diffuse intra-alveolar hemorrhage |216
inflammatory cell infiltration |216
normal coronary arteries |216
no inflammatory or ischemic injury in myocardium |216
