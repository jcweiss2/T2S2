56 years old | 0
male | 0
Chinese | 0
admitted to the hospital | 0
diarrhea | -480
yellow loose stools | -480
diarrhea 6-8 times a day | -480
aggravated diarrhea | -240
dark green watery stool | -240
diarrhea up to 10 times a day | -240
palpitations | -240
shortness of breath | -240
dizziness | -240
dry mouth | -240
dry skin | -240
sunken eye socket symptoms | -240
no history of fevering | -168
no abdominal pain | -168
no travelling | -168
liver cancer | -720
hepatitis B cirrhosis | -720
allograft | -720
immunosuppressive therapy | -720
tacrolimus | -720
mycophenolic acid | -720
sirolimus | -720
septic shock | 0
metabolic acidosis | 0
intubated | 0
transferred to the intensive care unit | 0
oliguria | 0
serum creatinine 170 μmol/L | 0
continuous renal replacement treatment | 0
white blood cell count 13.46×10^9/L | 0
neutrophil ratio 87.9% | 0
procalcitonin 3.32 ng/mL | 0
C-reactive protein 190 mg/L | 0
Troponin-T 191.2 ng/L | 0
possible abdominal or lung infection | 0
myocardial injury | 0
no significant changes in liver function test | 0
no significant changes in blood coagulation test | 0
no significant changes in platelet count | 0
tacrolimus concentration within the target treatment range | 0
temperature continued to rise to 38.5°C | 24
empirical treatment with piperacillin/tazobactam | 24
no significant improvement | 48
bronchoalveolar lavage solution for culture | 48
Aspergillus fumigatus | 48
carbapenem-resistant Klebsiella pneumoniae | 48
antibacterial agents replaced by meropenem and voriconazole | 48
tacrolimus and sirolimus discontinued | 48
stool for detection | 48
intestinal bacterial culture negative | 48
microscopic examination of parasite negative | 48
clostridium difficile antigen negative | 48
compound berberine | 48
electrolyte balance and acid-base balance corrected | 48
diarrhea significantly mitigated | 72
enteral nutrition solution | 72
probiotics | 72
high frequency diarrhea | 96
fever | 96
temperature fluctuating around 39 °C | 96
parasitic examination of stool negative | 96
fecal bacterial cultures negative | 96
blood sample for PACEseq mNGS analysis | 96
Klebsiella pneumoniae | 120
Cryptosporidium parvum | 120
oval bodies in stool samples | 120
Cryptosporidium oocysts | 120
azithromycin | 120
cyclosporine | 120
trough concentration of cyclosporine 194.00 μg/L | 144
cyclosporine dose adjusted | 144
diarrhea did not improve | 168
azithromycin stopped | 168
nitazoxanide | 168
diarrhea frequency reduced | 192
diarrhea subsided | 336
fecal samples collected again | 336
no Cryptosporidium oocysts | 336
nitazoxanide stopped | 336
systemic infection controlled | 960
disconnected from the ventilator intermittently | 960
creatinine decreased to normal baseline level | 960
liver function gradually recovered | 960
transferred to the general ward | 1128
rehabilitation treatment | 1128