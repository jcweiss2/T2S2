34 years old | 0
woman | 0
gravida 4 | 0
para 3 | 0
presented to the Obstetric Department for labor induction | 0
suspected macrosomic fetus | 0
39th gestational week | 0
periodic depression | 0
whiplash | 0
overweight (BMI 34) | 0
active phase of labor | 6
amniotomy | 6
clear amnion fluid | 6
oxytocin use | 6
spontaneous birth | 10
male infant | 10
4230 g | 10
Apgar score 7 | 10
Apgar score 10 | 10
discharge | 14
readmission | 24
pain | 24
chills | 24
hypotension (96/72 mmHg) | 24
tachycardia (112) | 24
fever | 24
oliguria | 24
generalized abdominal tenderness | 24
guarding | 24
peritoneal signs | 24
enlarged uterus | 24
abdominal ultrasound examination | 24
transvaginal ultrasound examination | 24
empty uterus | 24
no intraabdominal fluid | 24
culture samples collected | 24
intravenous antibiotic therapy with metronidazole | 24
intravenous antibiotic therapy with cefuroxime | 24
elevated CRP | 24
elevated creatinine | 24
normal white blood cell counts | 24
normal hemoglobin | 24
normal platelets | 24
abdominal CT-scan with intravenous contrast | 36
enlarged uterus | 36
ascites | 36
circulatory instability | 36
transfer to ICU | 36
tentative diagnosis of severe puerperal endometritis | 36
circulatory stabilization | 38
operation theater | 38
manual exploration of the uterus | 38
progressive elevation of CRP | 38
leucocytosis | 38
no retained placental tissue | 38
no uncontrolled hemorrhage | 38
antibiotic therapy changed to meropenem | 38
antibiotic therapy changed to metronidazole | 38
fulminate circulatory shock | 38
fluid resuscitation | 38
heavy vasopressor therapy | 38
cardiac arrest | 38
cardiopulmonary resuscitation | 38
intravenous adrenaline | 38
sinus rhythm | 38
transthoracic echocardiography | 38
right ventricular heart failure | 38
left ventricular heart failure | 38
lowered ejection fraction | 38
transfer to TICU | 38
invasive cardiopulmonary support | 38
cardiac failure reversed | 38
kidney function improved | 38
Group A streptococcus in urine sample | 38
Group A streptococcus in vaginal culture | 38
negative blood cultures | 38
allergy to penicillin | 38
meropenem continued | 38
metronidazole continued | 38
return to regional ICU | 168
stable condition | 168
intubated | 168
sedated | 168
circulatory instability | 168
temperature increased above 42°C | 168
active cooling | 168
CVVHDF | 168
new CT scan | 168
necrosis in uterus suspicion | 168
thrombosis in right uterine artery suspicion | 168
explorative laparotomy | 168
total abdominal hysterectomy | 168
necrotic uterus | 168
enlarged uterus | 168
thromboembolus in right uterine artery | 168
microscopic examination of acute necrotizing inflammation | 168
microscopic examination of reactive endometrial changes | 168
septic thromboemboli in uterine artery | 168
intensive care management | 168
resuscitative efforts | 168
respiratory assistance | 168
dialysis | 168
altered consciousness | 168
paralysis of all four extremities | 168
absent tendon reflexes | 168
preserved eye movements | 168
preserved oculus reflex | 168
MRI-scan | 168
EEG | 168
lumbar puncture | 168
no obvious explanation found | 168
severe Critical Illness Polyneuropathy (CIP) | 168
transfer to neurorehabilitation department | 2880
still patient at the center (4 months postpartum) | 2880
condition improving | 2880
