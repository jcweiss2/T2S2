665 g | 0
male | 0
emergency cesarean section | 0
severe preeclampsia | 0
intubated | 0
transferred to neonatal intensive care unit | 0
mechanical ventilation | 0
total parenteral nutrition | 0
minimal enteral nutrition with breast milk | 0
delayed meconium passage | 0
abdominal distension | 0
increased gastric residuals | 0
NEC | 0
minimal enteral feeding discontinued | 0
gastric free drainage | 0
broad-spectrum antibiotic therapy | 0
operated | 6
perforated NEC | 6
multiple areas of perforation | 6
circulatory disturbances in the intestinal wall | 6
long segment including jejunum and ileum resected | 6
stoma formed | 6
distal end left closed | 6
TPN until postoperative seventh day | 7
minimal enteral feeding started | 7
enteral nutrition alone insufficient | 7
short bowel syndrome | 7
thyroid screening tests | 14
fT4: 0.87 ng/dL | 14
TSH: 0.061 mIU/L | 14
cortisol: 5.75 µg/dL | 14
serum total bilirubin: 12.12 mg/dL | 14
direct reacting bilirubin: 11.48 mg/dL | 14
fT4 level decreasing | 21
close to lower limit of normal | 21
enteral levothyroxine 5 µg/kg/day | 21
no response to treatment | 21
enteral dose increased to 10 µg/kg/day | 21
no increase in fT4 levels | 21
poor absorption | 21
main site of oral thyroxine absorption incomplete | 21
rectal levothyroxine tablet | 21
ground and diluted with saline | 21
administered rectally | 21
dose 10 µg/kg/day | 21
fT4 levels increased | 30
bilirubin levels decreased | 30
died | 77
severe bronchopulmonary dysplasia | 77
surgical NEC | 77
short bowel syndrome | 77
sepsis | 77
