59 years old | 0
    man | 0
    admitted to the hospital | 0
    ascending aortic aneurysm | 0
    atrial fibrillation | 0
    congestive heart failure | 0
    reduced ejection fraction | 0
    bilateral lower extremity venous stasis ulcers | 0
    stage 3 chronic kidney disease | 0
    multinodular goiter | 0
    ground-level fall | 0
    ambulating | 0
    heart racing | 0
    denied dyspnea | 0
    denied chest pain | 0
    denied loss of consciousness | 0
    deterioration of health | -720
    unable to properly care for bilateral lower extremity wounds | -720
    clean wounds with water and washcloth daily | -720
    septic shock | 0
    blood pressure 84/53 mm Hg | 0
    heart rate 124 beats per minute | 0
    lactate 3 mg/dL | 0
    lower extremity ulcers below the knee | 0
    right extremity medial ulcers 8 × 5 cm (depth to muscle tissue) | 0
    right extremity medial ulcers 6 × 3 cm | 0
    left extremity medial ulcer 8 × 5 cm (depth to muscle tissue) | 0
    necrotic skin | 0
    subcutaneous tissue | 0
    maggots | 0
    C-reactive protein 6.97 mg/L | 0
    creatinine 3.54 mg/dL |6 0
    elevated troponin 0.06 ng/mL | 0
    elevated white blood cell count 14.8 × 10³ cells per mL | 0
    83.6% neutrophils | 0
    atrial fibrillation with rapid ventricular rate | 0
    enlarged heart | 0
    tortuous aorta | 0
    negative osteomyelitis | 0
    bilateral subcutaneous gas formation | 0
    admitted to ICU | 0
    treatment of septic shock | 0
    non-ST elevation myocardial infarction | 0
    sepsis bundle initiated | 0
    fluid resuscitation | 0
    vasopressor support with norepinephrine | 0
    blood cultures obtained | 0
    urine culture obtained | 0
    initiated on vancomycin | 0
    initiated on piperacillin/tazobactam | 0
    acute coronary syndrome protocol initiated | 0
    elevated troponins | 0
    amiodarone initiated | 0
    digoxin refractory | 0
    debridement of bilateral lower extremity necrotic skin and soft tissue | 0
    muscle tissue not involved | 0
    blood cultures grew S. fonticola | 0
    blood cultures grew MSSA | 0
    S. fonticola resistant to amoxicillin/clavulanate | 0
    vancomycin discontinued | 96
    piperacillin/tazobactam de-escalated to ceftriaxone | 96
    dilation of all cardiac chambers | 0
    mild concentric left ventricular hypertrophy | 0
    left ventricular systolic function severely depressed | 0
    ejection fraction 15% to 20% | 0
    diastolic function unable to be assessed | 0
    abnormal septal motion | 0
    bundle branch block | 0
    abnormal regional wall motion | 0
    underlying coronary acute disease | 0
    myocardial infarction | 0
    right ventricle moderately dilated | 0
    mild to moderate reduced right ventricular systolic function | 0
    systolic pressure 45 mm Hg | 0
    moderate tricuspid regurgitation | 0
    TEE performed | 0
    severe left ventricular systolic dysfunction | 0
    severe low-flow low-gradient aortic valve stenosis | 0
    mitral valve vegetation less than 1 cm | 0
    mobile echo density 0.8 × 1.6 cm | 0
    left atrium thrombus | 0
    source of infection determined | 0
    chronic bilateral lower extremity skin infection | 0
    severe 2 vessel coronary artery disease | 0
    ceftriaxone changed to cefepime | 96
    infective endocarditis | 0
    Amp-C beta-lactamase production concern | 0
    duration of cefepime treatment 6 weeks | 0
    discharged to skilled nursing facility | 0
    uneventful recovery | 0
    completed 6 weeks antibiotic therapy | 1008
    outpatient management | 1008
    multidisciplinary approach | 1008
    cardiology follow-up | 1008
    nephrology follow-up | 1008
    infectious disease follow-up | 1008
    primary care follow-up | 1008
    S. fonticola bacteremia | 0
    endocarditis | 0
    colonization | 0
    local infection | 0
    hematogenous spread | 0
    β-Lactamase producing S. fonticola | 0
    susceptible organism | 0
    coinfection with MSSA | 0
    mitral valve endocarditis | 0
    