66 years old | 0
female | 0
admitted to the emergency department | 0
general weakness | -168
poor oral intake | -168
diabetes | -8760
hypertension | -8760
metformin | -8760
glimepiride | -8760
hydrochlorothiazide | -8760
losartan | -8760
atorvastatin | -8760
severe osteoarthritis | -8760
steroid injections | -336
urinary tract infection | -336
blood culture | -336
urine culture | -336
Escherichia coli | -336
ceftriaxone | -336
tazobactam | -336
no antihypertensive medication | -336
height 152 cm | 0
body weight 57 kg | 0
blood pressure 70/50 mmHg | 0
heart rate 70 beats per minute | 0
respiratory rate 20 per minute | 0
body temperature 36.5°C | 0
decreased skin turgor | 0
decreased tongue turgor | 0
pulmonary examination unremarkable | 0
cardiac examination unremarkable | 0
abdominal examination unremarkable | 0
neurologic examination unremarkable | 0
pyuria | 0
hypotension | 0
UTI sepsis | 0
antibiotics | 0
massive hydration | 0
stabilization of vital signs | 24
normalization of inflammatory signs | 48
normalization of blood pressure | 48
elevated serum calcium | 0
elevated serum creatinine | 0
poor oral intake | 0
general weakness | 0
administration of saline | 72
administration of calcitonin | 72
decrease in serum calcium | 96
increase in serum calcium | 120
contrast-enhanced computed tomography | 120
whole body bone scintigraphy | 120
no evidence of malignancy | 120
serum protein electrophoresis | 120
urine protein electrophoresis | 120
anti-neutrophil cytoplasmic antibody titers | 120
tumor marker studies | 120
thyroid function profile | 120
normal thyroid stimulating hormone | 120
normal free thyroxine | 120
bone mineral density T-score | 120
osteopenia | 120
suppressed PTH-vitamin D axis | 120
intact parathyroid hormone | 120
PTH-related peptide | 120
serum 25-hydroxy vitamin D | 120
adrenocortical function assessment | 120
low serum cortisol | 120
elevated adrenocorticotropic hormone | 120
ACTH stimulation test | 120
inadequate cortisol response | 120
diagnosis of secondary adrenal insufficiency | 120
hydrocortisone administration | 240
normalization of serum calcium | 264
improvement of general weakness | 264
improvement of anorexia | 264
normalization of magnesium level | 264
follow-up | 336
loss to follow-up | 672