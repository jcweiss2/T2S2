75 years old | 0
female | 0
admitted to the hospital | 0
mildly itching skin rash | -48
fever | -48
shivering | -48
weakness | -48
self-medication with cetirizine | -48
no improvement | -48
no signs of respiratory disorders | -48
no signs of gastrointestinal disorders | -48
SARS-CoV-2 polymerase chain reaction test negative | -48
chest X-ray did not show pulmonary infiltrates | -48
prescribed allopurinol for hyperuricemia | -504
antihypertensive drugs (amlodipine, valsartan) | -504
maculopapulous exanthema | 0
oral lesions not apparent | 0
skin lesions caused by viral infection | 0
adverse drug reaction induced by allopurinol | 0
allopurinol discontinued | 0
oral prednisolone prescribed | 0
cetirizine prescribed | 0
treatment on an outpatient basis | 0
worsening exanthema | 48
hospital admission | 48
highly painful widespread blistering and skin peeling | 48
oral involvement | 48
mucosal ulceration and erythema of the conjunctiva | 48
diagnosis of TEN | 48
prednisolone intravenously | 48
cyclosporine | 48
skin biopsy for histopathological examination | 48
typical signs of TEN | 48
transferred to Intensive Care Unit (ICU) | 48
multidisciplinary supportive team | 48
SCORTEN predicted hospital mortality of 90% | 48
fluid replacement | 48
conservative approach for skin management | 48
large blisters decompressed | 48
warm sterile lotions of polyhexanide and octenidine | 48
nonadhesive gauze, antiseptic gel, and sterile compresses | 48
metalline foil to prevent shearing forces | 48
oral lesions rinsed with saline and antiseptic lotions | 48
intensive analgesia including opiates | 48
patient-controlled analgesia | 48
nasogastric feeding | 48
prophylactic anticoagulation | 48
bacteriuria treated with antibiotics | 48
ophthalmologic consultations | 48
gynecological consultations | 48
signs of involvement with superficial necrolysis at the labia minora and introitus | 48
no evidence of superinfection | 48
skin lesions and general condition improved | 168
laboratory findings showed regression of renal failure and inflammatory markers | 168
transferred to the Dermatology Department | 168
recovered completely | 1008
discharged | 1008