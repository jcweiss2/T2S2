55 years old | 0 | 0 
male | 0 | 0 
nonalcoholic steatohepatitis | -672 | 0 
alpha 1 antitrypsin deficiency | -672 | 0 
orthotopic liver transplant | 0 | 0 
incarcerated inguinal hernia | 0 | 24 
hernia repair | 0 | 24 
cytomegalovirus viremia | 0 | 168 
valganciclovir | 0 | 168 
mycophenolate mofetil | 168 | 720 
tacrolimus | 168 | 720 
prednisone | 168 | 720 
encephalopathy | 720 | 744 
increasing home oxygen requirements | 720 | 744 
oxygen saturation <92% | 720 | 744 
sparse speech | 744 | 744 
disorientation | 744 | 744 
nonfocal neurologic examination | 744 | 744 
white blood cell count 9.3 × 10^9/L | 744 | 744 
creatinine 2.12 mg/dL | 744 | 744 
blood urea nitrogen 53 mg/dL | 744 | 744 
arterial ammonia 204 µmol/L | 744 | 744 
intravenous ganciclovir | 744 | 768 
vancomycin | 744 | 768 
meropenem | 744 | 768 
micafungin | 744 | 768 
intravenous micronutrient supplementation | 744 | 768 
lumbar puncture | 744 | 744 
encapsulated yeast suspicious for Cryptococcus | 744 | 744 
liposomal amphotericin B | 744 | 768 
flucytosine | 744 | 768 
continuous renal replacement therapy | 744 | 768 
rifaximin | 744 | 768 
zinc | 744 | 768 
lactulose | 744 | 768 
ammonia 692 µmol/L | 768 | 768 
mechanical ventilation | 768 | 840 
empiric intravenous doxycycline | 768 | 840 
urine and bronchial aspirate for Mycoplasma and Ureaplasma PCR | 768 | 768 
ammonia <100 µmol/L | 840 | 840 
Cryptococcal serum and cerebrospinal fluid antigen titers >1:2560 | 840 | 840 
cultures from bronchoalveolar lavage, CSF, and blood revealed cryptococcal growth | 840 | 840 
repeat lumbar punctures | 840 | 1008 
thrombocytopenia | 840 | 1008 
tracheostomy | 1008 | 1008 
splenectomy | 1008 | 1008 
sepsis | 1008 | 1008 
duodenal leak | 1008 | 1008 
renal failure | 1008 | 1008 
failure to thrive | 1008 | 1008 
comfort care in hospice | 1008 | 1008 
urea cycle disorder screening studies | 1008 | 1008 
low urine orotic level | 1008 | 1008 
normal serum citrulline and arginine level | 1008 | 1008 
weight loss 15 lb | -720 | 0 
hyperammonemia | 744 | 840 
cerebral edema | 840 | 840 
brain herniation | 840 | 840 
urease production | 840 | 840 
acetohydroxamic acid | 1008 | 1008 
inborn error of metabolism | 1008 | 1008 
ornithine transcarbamylase deficiency | 1008 | 1008 
ureaplasma | 1008 | 1008 
valproic acid overdose | 1008 | 1008 
ackee fruit | 1008 | 1008 
magnetic resonance imaging of the brain | 840 | 840 
cytotoxic edema | 840 | 840 
hydrocephalus | 1008 | 1008 
splenic infarcts | 1008 | 1008 
necrosis | 1008 | 1008 
oliguric renal failure | 1008 | 1008 
persistent thrombocytopenia | 840 | 1008 
large volume drainage | 840 | 1008 
permanent CSF diversion | 840 | 840 
altered mental status | 720 | 840 
central nervous system cryptococcosis | 840 | 840 
disseminated cryptococcal infection | 840 | 840 
urease-producing organisms | 840 | 840 
cryptococcal infection | 840 | 840 
hyperammonemia caused by urease-producing organisms | 840 | 840 
adjunctive treatment | 1008 | 1008 
control of plasma ammonia levels | 840 | 1008 
combination antifungal therapy | 840 | 1008 
early consultation with nephrology | 840 | 840 
initiation of CRRT | 840 | 840 
critical intervention | 840 | 840 
neurological outcome | 1008 | 1008 
transient improvement | 840 | 840 
normal brain MRI | 840 | 840 
slow neurological improvement | 1008 | 1008 
complete recovery | 1008 | 1008 
genetic analysis | 1008 | 1008 
informed consent | 0 | 0 
ethics approval | 0 | 0 
funding | 0 | 0 
conflicts of interest | 0 | 0 
ORCID iD | 0 | 0 
anonymized patient information | 0 | 0 
publication | 0 | 0 
research | 0 | 0 
authorship | 0 | 0 
article | 0 | 0 
institution | 0 | 0 
representative | 0 | 0 
case reports | 1008 | 1008 
cryptococcal infection | 840 | 1008 
hyperammonemia | 744 | 1008 
liver transplant | 0 | 1008 
urease production | 840 | 1008 
cryptococcal infections | 840 | 1008 
therapeutic target | 1008 | 1008 
acetohydroxamic acid | 1008 | 1008 
FDA-approved | 1008 | 1008 
irreversible enzyme inhibitor | 1008 | 1008 
struvite stones | 1008 | 1008 
in vitro | 1008 | 1008 
adjunctive treatment | 1008 | 1008 
control of plasma ammonia levels | 840 | 1008 
CRRT | 840 | 1008 
nephrology | 840 | 840 
initiation of CRRT | 840 | 840 
critical intervention | 840 | 840 
neurological outcome | 1008 | 1008 
transient improvement | 840 | 840 
normal brain MRI | 840 | 840 
slow neurological improvement | 1008 | 1008 
complete recovery | 1008 | 1008 
genetic analysis | 1008 | 1008 
informed consent | 0 | 0 
ethics approval | 0 | 0 
funding | 0 | 0 
conflicts of interest | 0 | 0 
ORCID iD | 0 | 0 
anonymized patient information | 0 | 0 
publication | 0 | 0 
research | 0 | 0 
authorship | 0 | 0 
article | 0 | 0 
institution | 0 | 0 
representative | 0 | 0 
case reports | 1008 | 1008 
cryptococcal infection | 840 | 1008 
hyperammonemia | 744 | 1008 
liver transplant | 0 | 1008 
urease production | 840 | 1008 
cryptococcal infections | 840 | 1008 
therapeutic target | 1008 | 1008 
acetohydroxamic acid | 1008 | 1008 
FDA-approved | 1008 | 1008 
irreversible enzyme inhibitor | 1008 | 1008 
struvite stones | 1008 | 1008 
in vitro | 1008 | 1008 
adjunctive treatment | 1008 | 1008 
control of plasma ammonia levels | 840 | 1008 
CRRT | 840 | 1008 
nephrology | 840 | 840 
initiation of CRRT | 840 | 840 
critical intervention | 840 | 840 
neurological outcome | 1008 | 1008 
transient improvement | 840 | 840 
normal brain MRI | 840 | 840 
slow neurological improvement | 1008 | 1008 
complete recovery | 1008 | 1008 
genetic analysis | 1008 | 1008 
informed consent | 0 | 0 
ethics approval | 0 | 0 
funding | 0 | 0 
conflicts of interest | 0 | 0 
ORCID iD | 0 | 0 
anonymized patient information | 0 | 0 
publication | 0 | 0 
research | 0 | 0 
authorship | 0 | 0 
article | 0 | 0 
institution | 0 | 0 
representative | 0 | 0 
case reports | 1008 | 1008 
cryptococcal infection | 840 | 1008 
hyperammonemia | 744 | 1008 
liver transplant | 0 | 1008 
urease production | 840 | 1008 
cryptococcal infections | 840 | 1008 
therapeutic target | 1008 | 1008 
acetohydroxamic acid | 1008 | 1008 
FDA-approved | 1008 | 1008 
irreversible enzyme inhibitor | 1008 | 1008 
struvite stones | 1008 | 1008 
in vitro | 1008 | 1008 
adjunctive treatment | 1008 | 1008 
control of plasma ammonia levels | 840 | 1008 
CRRT | 840 | 1008 
nephrology | 840 | 840 
initiation of CRRT | 840 | 840 
critical intervention | 840 | 840 
neurological outcome | 1008 | 1008 
transient improvement | 840 | 840 
normal brain MRI | 840 | 840 
slow neurological improvement | 1008 | 1008 
complete recovery | 1008 | 1008 
genetic analysis | 1008 | 1008 
informed consent | 0 | 0 
ethics approval | 0 | 0 
funding | 0 | 0 
conflicts of interest | 0 | 0 
ORCID iD | 0 | 0 
anonymized patient information | 0 | 0 
publication | 0 | 0 
research | 0 | 0 
authorship | 0 | 0 
article | 0 | 0 
institution | 0 | 0 
representative | 0 | 0 
case reports | 1008 | 1008 
cryptococcal infection | 840 | 1008 
hyperammonemia | 744 | 1008 
liver transplant | 0 | 1008 
urease production | 840 | 1008 
cryptococcal infections | 840 | 1008 
therapeutic target | 1008 | 1008 
acetohydroxamic acid | 1008 | 1008 
FDA-approved | 1008 | 1008 
irreversible enzyme inhibitor | 1008 | 1008 
struvite stones | 1008 | 1008 
in vitro | 1008 | 1008 
adjunctive treatment | 1008 | 1008 
control of plasma ammonia levels | 840 | 1008 
CRRT | 840 | 1008 
nephrology | 840 | 840 
initiation of CRRT | 840 | 840 
critical intervention | 840 | 840 
neurological outcome | 1008 | 1008 
transient improvement | 840 | 840 
normal brain MRI | 840 | 840 
slow neurological improvement | 1008 | 1008 
complete recovery | 1008 | 1008 
genetic analysis | 1008 | 1008 
informed consent | 0 | 0 
ethics approval | 0 | 0 
funding | 0 | 0 
conflicts of interest | 0 | 0 
ORCID iD | 0 | 0 
anonymized patient information | 0 | 0 
publication | 0 | 0 
research | 0 | 0 
authorship | 0 | 0 
article | 0 | 0 
institution | 0 | 0 
representative | 0 | 0 
case reports | 1008 | 1008 
cryptococcal infection | 840 | 1008 
hyperammonemia | 744 | 1008 
liver transplant | 0 | 1008 
urease production | 840 | 1008 
cryptococcal infections | 840 | 1008 
therapeutic target | 1008 | 1008 
acetohydroxamic acid | 1008 | 1008 
FDA-approved | 1008 | 1008 
irreversible enzyme inhibitor | 1008 | 1008 
struvite stones | 1008 | 1008 
in vitro | 1008 | 1008 
adjunctive treatment | 1008 | 1008 
control of plasma ammonia levels | 840 | 1008 
CRRT | 840 | 1008 
nephrology | 840 | 840 
initiation of CRRT | 840 | 840 
critical intervention | 840 | 840 
neurological outcome | 1008 | 1008 
transient improvement | 840 | 840 
normal brain MRI | 840 | 840 
slow neurological improvement | 1008 | 1008 
complete recovery | 1008 | 1008 
genetic analysis | 1008 | 1008 
informed consent | 0 | 0 
ethics approval | 0 | 0 
funding | 0 | 0 
conflicts of interest | 0 | 0 
ORCID iD | 0 | 0 
anonymized patient information | 0 | 0 
publication | 0 | 0 
research | 0 | 0 
authorship | 0 | 0 
article | 0 | 0 
institution | 0 | 0 
representative | 0 | 0 
case reports | 1008 | 1008 
cryptococcal infection | 840 | 1008 
hyperammonemia | 744 | 1008 
liver transplant | 0 | 1008 
urease production | 840 | 1008 
cryptococcal infections | 840 | 1008 
therapeutic target | 1008 | 1008 
acetohydroxamic acid | 1008 | 1008 
FDA-approved | 1008 | 1008 
irreversible enzyme inhibitor | 1008 | 1008 
struvite stones | 1008 | 1008 
in vitro | 1008 | 1008 
adjunctive treatment | 1008 | 1008 
control of plasma ammonia levels | 840 | 1008 
CRRT | 840 | 1008 
nephrology | 840 | 840 
initiation of CRRT | 840 | 840 
critical intervention | 840 | 840 
neurological outcome | 1008 | 1008 
transient improvement | 840 | 840 
normal brain MRI | 840 | 840 
slow neurological improvement | 1008 | 1008 
complete recovery | 1008 | 1008 
genetic analysis | 1008 | 1008 
informed consent | 0 | 0 
ethics approval | 0 | 0 
funding | 0 | 0 
conflicts of interest | 0 | 0 
ORCID iD | 0 | 0 
anonymized patient information | 0 | 0 
publication | 0 | 0 
research | 0 | 0 
authorship | 0 | 0 
article | 0 | 0 
institution | 0 | 0 
representative | 0 | 0 
case reports | 1008 | 1008 
cryptococcal infection | 840 | 1008 
hyperammonemia | 744 | 1008 
liver transplant | 0 | 1008 
urease production | 840 | 1008 
cryptococcal infections | 840 | 1008 
therapeutic target | 1008 | 1008 
acetohydroxamic acid | 1008 | 1008 
FDA-approved | 1008 | 1008 
irreversible enzyme inhibitor | 1008 | 1008 
struvite stones | 1008 | 1008 
in vitro | 1008 | 1008 
adjunctive treatment | 1008 | 1008 
control of plasma ammonia levels | 840 | 1008 
CRRT | 840 | 1008 
nephrology | 840 | 840 
initiation of CRRT | 840 | 840 
critical intervention | 840 | 840 
neurological outcome | 1008 | 1008 
transient improvement | 840 | 840 
normal brain MRI | 840 | 840 
slow neurological improvement | 1008 | 1008 
complete recovery | 1008 | 1008 
genetic analysis | 1008 | 1008 
informed consent | 0 | 0 
ethics approval | 0 | 0 
funding | 0 | 0 
conflicts of interest | 0 | 0 
ORCID iD | 0 | 0 
anonymized patient information | 0 | 0 
publication | 0 | 0 
research | 0 | 0 
authorship | 0 | 0 
article | 0 | 0 
institution | 0 | 0 
representative | 0 | 0 
case reports | 1008 | 1008 
cryptococcal infection | 840 | 1008 
hyperammonemia | 744 | 1008 
liver transplant | 0 | 1008 
urease production | 840 | 1008 
cryptococcal infections | 840 | 1008 
therapeutic target | 1008 | 1008 
acetohydroxamic acid | 1008 | 1008 
FDA-approved | 1008 | 1008 
irreversible enzyme inhibitor | 1008 | 1008 
struvite stones | 1008 | 1008 
in vitro | 1008 | 1008 
adjunctive treatment | 1008 | 1008 
control of plasma ammonia levels | 840 | 1008 
CRRT | 840 | 1008 
nephrology | 840 | 840 
initiation of CRRT | 840 | 840 
critical intervention | 840 | 840 
neurological outcome | 1008 | 1008 
transient improvement | 840 | 840 
normal brain MRI | 840 | 840 
slow neurological improvement | 1008 | 1008 
complete recovery | 1008 | 1008 
genetic analysis | 1008 | 1008 
informed consent | 0 | 0 
ethics approval | 0 | 0 
funding | 0 | 0 
conflicts of interest | 0 | 0 
ORCID iD | 0 | 0 
anonymized patient information | 0 | 0 
publication | 0 | 0 
research | 0 | 0 
authorship | 0 | 0 
article | 0 | 0 
institution | 0 | 0 
representative | 0 | 0 
case reports | 1008 | 1008 
cryptococcal infection | 840 | 1008 
hyperammonemia | 744 | 1008 
liver transplant | 0 | 1008 
urease production | 840 | 1008 
cryptococcal infections | 840 | 1008 
therapeutic target | 1008 | 1008 
acetohydroxamic acid | 1008 | 1008 
FDA-approved | 1008 | 1008 
irreversible enzyme inhibitor | 1008 | 1008 
struvite stones | 1008 | 1008 
in vitro | 1008 | 1008 
adjunctive treatment | 1008 | 1008 
control of plasma ammonia levels | 840 | 1008 
CRRT | 840 | 1008 
nephrology | 840 | 840 
initiation of CRRT | 840 | 840 
critical intervention | 840 | 840 
neurological outcome | 1008 | 1008 
transient improvement | 840 | 840 
normal brain MRI | 840 | 840 
slow neurological improvement | 1008 | 1008 
complete recovery | 1008 | 1008 
genetic analysis | 1008 | 1008 
informed consent | 0 | 0 
ethics approval | 0 | 0 
funding | 0 | 0 
conflicts of interest | 0 | 0 
ORCID iD | 0 | 0 
anonymized patient information | 0 | 0 
publication | 0 | 0 
research | 0 | 0 
authorship | 0 | 0 
article | 0 | 0 
institution | 0 | 0 
representative | 0 | 0 
case reports | 1008 | 1008 
cryptococcal infection | 840 | 1008 
hyperammonemia | 744 | 1008 
liver transplant | 0 | 1008 
urease production | 840 | 1008 
cryptococcal infections | 840 | 1008 
therapeutic target | 1008 | 1008 
acetohydroxamic acid | 1008 | 1008 
FDA-approved | 1008 | 1008 
irreversible enzyme inhibitor | 1008 | 1008 
struvite stones | 1008 | 1008 
in vitro | 1008 | 1008 
adjunctive treatment | 1008 | 1008 
control of plasma ammonia levels | 840 | 1008 
CRRT | 840 | 1008 
nephrology | 840 | 840 
initiation of CRRT | 840 | 840 
critical intervention | 840 | 840 
neurological outcome | 1008 | 1008 
transient improvement | 840 | 840 
normal brain MRI | 840 | 840 
slow neurological improvement | 1008 | 1008 
complete recovery | 1008 | 1008 
genetic analysis | 1008 | 1008 
informed consent | 0 | 0 
ethics approval | 0 | 0 
funding | 0 | 0 
conflicts of interest | 0 | 0 
ORCID iD | 0 | 0 
anonymized patient information | 0 | 0 
publication | 0 | 0 
research | 0 | 0 
authorship | 0 | 0 
article | 0 | 0 
institution | 0 | 0 
representative | 0 | 0 
case reports | 1008 | 1008 
cryptococcal infection | 840 | 1008 
hyperammonemia | 744 | 1008 
liver transplant | 0 | 1008 
urease production | 840 | 1008 
cryptococcal infections | 840 | 1008 
therapeutic target | 1008 | 1008 
acetohydroxamic acid | 1008 | 1008 
FDA-approved | 1008 | 1008 
irreversible enzyme inhibitor | 1008 | 1008 
struvite stones | 1008 | 1008 
in vitro | 1008 | 1008 
adjunctive treatment | 1008 | 1008 
control of plasma ammonia levels | 840 | 1008 
CRRT | 840 | 1008 
nephrology | 840 | 840 
initiation of CRRT | 840 | 840 
critical intervention | 840 | 840 
neurological outcome | 1008 | 1008 
transient improvement | 840 | 840 
normal brain MRI | 840 | 840 
slow neurological improvement | 1008 | 1008 
complete recovery | 1008 | 1008 
genetic analysis | 1008 | 1008 
informed consent | 0 | 0 
ethics approval | 0 | 0 
funding | 0 | 0 
conflicts of interest | 0 | 0 
ORCID iD | 0 | 0 
anonymized patient information | 0 | 0 
publication | 0 | 0 
research | 0 | 0 
authorship | 0 | 0 
article | 0 | 0 
institution | 0 | 0 
representative | 0 | 0 
case reports | 1008 | 1008 
cryptococcal infection | 840 | 1008 
hyperammonemia | 744 | 1008 
liver transplant | 0 | 1008 
urease production | 840 | 1008 
cryptococcal infections | 840 | 1008 
therapeutic target | 1008 | 1008 
acetohydroxamic acid | 1008 | 1008 
FDA-approved | 1008 | 1008 
irreversible enzyme inhibitor | 1008 | 1008 
struvite stones | 1008 | 1008 
in vitro | 1008 | 1008 
adjunctive treatment | 1008 | 1008 
control of plasma ammonia levels | 840 | 1008 
CRRT | 840 | 1008 
nephrology | 840 | 840 
initiation of CRRT | 840 | 840 
critical intervention | 840 | 840 
neurological outcome | 1008 | 1008 
transient improvement | 840 | 840 
normal brain MRI | 840 | 840 
slow neurological improvement | 1008 | 1008 
complete recovery | 1008 | 1008 
genetic analysis | 1008 | 1008 
informed consent | 0 | 0 
ethics approval | 0 | 0 
funding | 0 | 0 
conflicts of interest | 0 | 0 
ORCID iD | 0 | 0 
anonymized patient information | 0 | 0 
publication | 0 | 0 
research | 0 | 0 
authorship | 0 | 0 
article | 0 | 0 
institution | 0 | 0 
representative | 0 | 0 
case reports | 1008 | 1008 
cryptococcal infection | 840 | 1008 
hyperammonemia | 744 | 1008 
liver transplant | 0 | 1008 
urease production | 840 | 1008 
cryptococcal infections | 840 | 1008 
therapeutic target | 1008 | 1008 
acetohydroxamic acid | 1008 | 1008 
FDA-approved | 1008 | 1008 
irreversible enzyme inhibitor | 1008 | 1008 
struvite stones | 1008 | 1008 
in vitro | 1008 | 1008 
adjunctive treatment | 1008 | 1008 
control of plasma ammonia levels | 840 | 1008 
CRRT | 840 | 1008 
nephrology | 840 | 840 
initiation of CRRT | 840 | 840 
critical intervention | 840 | 840 
neurological outcome | 1008 | 1008 
transient improvement | 840 | 840 
normal brain MRI | 840 | 840 
slow neurological improvement | 1008 | 1008 
complete recovery | 1008 | 1008 
genetic analysis | 1008 | 1008 
informed consent | 0 | 0 
ethics approval | 0 | 0 
funding | 0 | 0 
conflicts of interest | 0 | 0 
ORCID iD | 0 | 0 
anonymized patient information | 0 | 0 
publication | 0 | 0 
research | 0 | 0 
authorship | 0 | 0 
article | 0 | 0 
institution | 0 | 0 
representative | 0 | 0 
case reports | 1008 | 1008 
cryptococcal infection | 840 | 1008 
hyperammonemia | 744 | 1008 
liver transplant | 0 | 1008 
urease production | 840 | 1008 
cryptococcal infections | 840 | 1008 
therapeutic target | 1008 | 1008 
acetohydroxamic acid | 1008 | 1008 
FDA-approved | 1008 | 1008 
irreversible enzyme inhibitor | 1008 | 1008 
struvite stones | 1008 | 1008 
in vitro | 1008 | 1008 
adjunctive treatment | 1008 | 1008 
control of plasma ammonia levels | 840 | 1008 
CRRT | 840 | 1008 
nephrology | 840 | 840 
initiation of CRRT | 840 | 840 
critical intervention | 840 | 840 
neurological outcome | 1008 | 1008 
transient improvement | 840 | 840 
normal brain MRI | 840 | 840 
slow neurological improvement | 1008 | 1008 
complete recovery | 1008 | 1008 
genetic analysis | 1008 | 1008 
informed consent | 0 | 0 
ethics approval | 0 | 0 
funding | 0 | 0 
conflicts of interest | 0 | 0 
ORCID iD | 0 | 0 
anonymized patient information | 0 | 0 
publication | 0 | 0 
research | 0 | 0 
authorship | 0 | 0 
article | 0 | 0 
institution | 0 | 0 
representative | 0 | 0 
case reports | 1008 | 1008 
cryptococcal infection | 840 | 1008 
hyperammonemia | 744 | 1008 
liver transplant | 0 | 1008 
urease production | 840 | 1008 
cryptococcal infections | 840 | 1008 
therapeutic target | 1008 | 1008 
acetohydroxamic acid | 1008 | 1008 
FDA-approved | 1008 | 1008 
irreversible enzyme inhibitor | 1008 | 1008 
struvite stones | 1008 | 1008 
in vitro | 1008 | 1008 
adjunctive treatment | 1008 | 1008 
control of plasma ammonia levels | 840 | 1008 
CRRT | 840 | 1008 
nephrology | 840 | 840 
initiation of CRRT | 840 | 840 
critical intervention | 840 | 840 
neurological outcome | 1008 | 1008 
transient improvement | 840 | 840 
normal brain MRI | 840 | 840 
slow neurological improvement | 1008 | 1008 
complete recovery | 1008 | 1008 
genetic analysis | 1008 | 1008 
informed consent | 0 | 0 
ethics approval | 0 | 0 
funding | 0 | 0 
conflicts of interest | 0 | 0 
ORCID iD | 0 | 0 
anonymized patient information | 0 | 0 
publication | 0 | 0 
research | 0 | 0 
authorship | 0 | 0 
article | 0 | 0 
institution | 0 | 0 
representative | 0 | 0 
case reports | 1008 | 1008 
cryptococcal infection | 840 | 1008 
hyperammonemia | 744 | 1008 
liver transplant | 0 | 1008 
urease production | 840 | 1008 
cryptococcal infections | 840 | 1008 
therapeutic target | 1008 | 1008 
acetohydroxamic acid | 1008 | 1008 
FDA-approved | 1008 | 1008 
irreversible enzyme inhibitor | 1008 | 1008 
struvite stones | 1008 | 1008 
in vitro | 1008 | 1008 
adjunctive treatment | 1008 | 1008 
control of plasma ammonia levels | 840 | 1008 
CRRT | 840 | 1008 
nephrology | 840 | 840 
initiation of CRRT | 840 | 840 
critical intervention | 840 | 840 
neurological outcome | 1008 | 1008 
transient improvement | 840 | 840 
normal brain MRI | 840 | 840 
slow neurological improvement | 1008 | 1008 
complete recovery | 1008 | 1008 
genetic analysis | 1008 | 1008 
informed consent | 0 | 0 
ethics approval | 0 | 0 
funding | 0 | 0 
conflicts of interest | 0 | 0 
ORCID iD | 0 | 0 
anonymized patient information | 0 | 0 
publication | 0 | 0 
research | 0 | 0 
authorship | 0 | 0 
article | 0 | 0 
institution | 0 | 0 
representative | 0 | 0 
case reports | 1008 | 1008 
cryptococcal infection | 840 | 1008 
hyperammonemia | 744 | 1008 
liver transplant | 0 | 1008 
urease production | 840 | 1008 
cryptococcal infections | 840 | 1008 
therapeutic target | 1008 | 1008 
acetohydroxamic acid | 1008 | 1008 
FDA-approved | 1008 | 1008 
irreversible enzyme inhibitor | 1008 | 1008 
struvite stones | 1008 | 1008 
in vitro | 1008 | 1008 
adjunctive treatment | 1008 | 1008 
control of plasma ammonia levels | 840 | 1008 
CRRT | 840 | 1008 
nephrology | 840 | 840 
initiation of CRRT | 840 | 840 
critical intervention | 840 | 840 
neurological outcome | 1008 | 1008 
transient improvement | 840 | 840 
normal brain MRI | 840 | 840 
slow neurological improvement | 1008 | 1008 
complete recovery | 1008 | 1008 
genetic analysis | 1008 | 1008 
informed consent | 0 | 0 
ethics approval | 0 | 0 
funding | 0 | 0 
conflicts of interest | 0 | 0 
ORCID iD | 0 | 0 
anonymized patient information | 0 | 0 
publication | 0 | 0 
research | 0 | 0 
authorship | 0 | 0 
article | 0 | 0 
institution | 0 | 0 
representative | 0 | 0 
case reports | 1008 | 1008 
cryptococcal infection | 840 | 1008 
hyperam