48 years old|0
male|0
born with spina bifida|0
paraplegia waist downward|0
long-term indurethral catheter|0
temperature of 39°C|0
urine microbiology revealed Pseudomonas aeruginosa|0
prescribed ciprofloxacin 500 mg twice a day|0
ultrasound examination of urinary tract|0
bilateral renal calculi|0
largest calculus in the right kidney measuring 1 cm|0
large staghorn calculus in the left kidney|0
no hydronephrosis|0
isotope renogram|0
divided renal function of 70% for the right kidney|0
divided renal function of 30% for the left kidney|0
persistent obstructive pattern in the left kidney|0
slightly reduced tracer uptake in the left upper moiety|0
left upper moiety accounted for 11% of function|0
left lower moiety accounted for 18% of function|0
left upper moiety appeared obstructed for 30 minutes|0
persistent retention of tracer|0
CT revealed large staghorn calculus in the left kidney|0
moderately severe left hydronephrosis|0
pronounced in the upper pole|0
left staghorn calculus measured ~4 cm at its maximum diameter|0
13 mm calculus in the left upper ureter|0
left kidney measured 9.5 cm|0
diffuse mid> and upper-pole cortical thinning|0
multiple calculi in the mid and lower poles of the right kidney|0
no bladder calculi|0
flexible uretero-renoscopy was performed|0
preoperative discussion|0
left ureteroscopy with laser lithotripsy| -624
insertion of left ureteric stent| -624
very tight stricture at the left ureteropelvic junction| -624
stricture was dilated sequentially| -624
access sheath of size 12/14 French was used| -624
laser lithotripsy| -624
40%–50% of stones were fragmented| -624
large amounts of stones left behind| -624
ureter was clear| -624
stented with 8-French stent| -624
repeat left ureterorenoscopy and laser lithotripsy| -504
flexible ureteroscope| -504
time taken was 3 hours| -504
majority of stone fragments were retrieved| -504
some fragments were left to pass| -504
fragments were left in lower pole| -504
ureter was clear| -504
4.8-French stent inserted in the left ureter| -504
no intraoperative complications| -504
no postoperative complications| -504
CT of kidney, ureters, bladder performed 3 weeks after the second ureteroscopy| -504
generalized shrinkage of left kidney| -504
multifocal scarring| -504
irregularity of its outline| -504
ureteric stent in situ| -504
three lower pole stones in individual calyces| -504
two of them quite large| -504
largest measuring about 19 mm in diameter| -504
some dilatation of the upper pole pelvicalyceal system| -504
presence of the ureteric stent| -504
no stones in the left ureter| -504
calcification in the prostate| -504
small stone fragments in the base of the bladder| -504
right kidney of normal size| -504
small area of upper pole cortical scarring| -504
cortical thickness otherwise reasonably maintained| -504
multiple upper and lower pole calyceal stones| -504
largest at the lower pole measuring about 14 mm| -504
1 cm stone in the renal pelvis| -504
left JJ stent removed| -504
stone analysis revealed struvite| -504
blood pressure recorded as 143/97 mmHg|0
recording of 24-hour blood pressure not done|0
no treatment instituted|0
urine sample sent for microbiology|0
report was “mixed growth”|0
antibiotic sensitivity not reported|0
left rigid ureterorenoscopy performed|0
patient received gentamicin 240 mg intravenously|0
ureter was normal|0
size 13/15, 46 cm access sheath used|0
flexible ureteroscopy|0
laser lithotripsy|0
fragments removed with a basket|0
difficult to negotiate the scope into calyceal diverticulum|0
vision was poor because of bleeding|0
some fragments remained|0
right rigid ureteroscopy performed|0
possible intrarenal mucosal perforation|0
4.8-Fr, 26 cm, JJ stent inserted in both ureters|0
surgery lasted for 2 hours and 40 minutes|0
blood pressure during surgery: 80/40 mmHg|0
blood pressure remained stable at 90/50 mmHg|0
frank hematuria|0
sinus tachycardia|0
admitted to the critical care unit|0
hemodynamically stable|0
hemoglobin: 116 g/L|0
white blood cell count: 24.5×109/L|0
neutrophils: 22.6×109/L|0
INR: 1.2|0
APTT: 32 seconds|0
APTT ratio: 1.3|0
C-reactive protein: 137 mg/L|0
creatinine: 64 μmol/L|0
prescribed cefuroxime intravenously|0
transferred to the spinal unit the following day|24
temperature of 38°C|24
urine was dark red|24
blood tests: INR: 1.1|24
hemoglobin: 120 g/L|24
white blood cell count: 20×109|24
neutrophils: 17.9×109|24
C-reactive protein: 168.1 mg/L|24
prescribed gentamicin for 5 days|24
hematuria subsided|24
discharged home|24
both ureteric stents removed|168
gentamicin 160 mg administered|168
three days later developed temperature|168
CT of kidneys requested|168
hemoglobin: 128 g/L|168
white blood cell count: 9.6×109|168
C-reactive protein: 133.4 mg/L|168
urine culture: P. aeruginosa|168
prescribed ciprofloxacin 500 mg twice a day|168
CT of urinary tract performed 4 weeks after ureteroscopy|672
9×7 cm subcapsular collection on the left kidney|672
minor perinephric fat stranding|672
few residual stones/fragments in the lower pole calyces|672
largest measuring 19 mm|672
multiple residual stones in the mid and lower pole calyces of the right kidney|672
largest about 9 mm|672
no ureteric or bladder stones|672
chest X-ray revealed elevated left hemidiaphragm|672
minimal atelectasis in the left lower zone|672
percutaneous drainage not carried out|672
managed conservatively|672
monitoring body temperature|672
monitoring C-reactive protein|672
monitoring white blood cell count|672
prescribed ciprofloxacin 500 mg twice a day for 5 days|672
urine sample showed growth of Pseudomonas aeruginosa resistant to gentamicin and ciprofloxacin|672
ciprofloxacin discontinued|672
remained well in himself|672
prescribed ferrous sulfate 200 mg daily|672
isotope renogram performed 8 weeks after ureterorenoscopy|1344
deterioration in the left renal function|1344
left kidney contributed only 17%|1344
right kidney contributed 83%|1344
renographic analysis showed both kidneys draining spontaneously without obstruction|1344
renographic drainage curve normal on the right|1344
good drainage on the left|1344
ultrasound scan of left kidney performed 9 weeks after ureterorenoscopy|1512
residual hematoma 3.3 cm in depth|1512
CT of kidney, ureters, bladder performed 14 weeks after ureterorenoscopy|2352
left renal subcapsular collection reduced to 3×2 cm|2352
some inflammatory stranding in the left perinephric fat|2352
no hydronephrosis|2352
several residual calculi in both kidneys|2352
blood pressure was 146/93 mmHg|2352
24-hour mean blood pressure: 130/91 mmHg|2352
prescribed ramipril 1.25 mg daily|2352
four months after the third ureteroscopy|2688
hemoglobin increased to 157 g/L|2688
ethical approval not necessary|0
