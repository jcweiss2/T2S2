47 years old | 0
male | 0
admitted to hospital | 0
COVID-19 infection | -48
fever | -48
sweats | -48
cough | -48
shortness of breath | -48
nasopharyngeal swab | 0
diagnosis of COVID-19 | 0
CXR | 0
right basal atelectasis | 0
inpatient duration | 0
ventilatory support | 0
dexamethasone | 0
discharged | 504
represented with chest pain | 336
shortness of breath | 336
COVID-19 tests negative | 336
CTPA | 336
large left hydropneumothorax | 336
air fluid levels | 336
empirical antimicrobial therapy | 336
clarithromycin | 336
piperacillin/tazobactam | 336
antibiotics escalated to meropenem | 336
intercostal drain inserted | 336
pleural fluid sampling | 336
pH of 7.1 | 336
microbiology cultures reported negative | 336
broad spectrum antibiotics | 336
failed to drain pleural cavity | 336
left uniportal video-assisted thoracoscopy | 1008
left pleural washout and decortication | 1008
necrotic lung | 1008
left lower lobectomy | 1008
antibiotics continued | 1008
fall in white cell count | 1008
C reactive protein | 1008
sinus tachycardia | 1008
resolved by the time of discharge | 1056
antibiotics discontinued | 1056
mobile and independent | 1056
no subsequent readmission | 1056
CXR at discharge | 1056
clear pleural spaces | 1056
loss of volume in left hemithorax | 1056
macroscopic inspection of lung | 1008
microscopic evaluation | 1008
bronchial oedema | 1008
organising pneumonia | 1008
airway oedema | 1008
pulmonary haemorrhage | 1008
acute fibrinous pneumonia | 1008