39 years old | 0
female | 0
height 155 cm | 0
weight 44.5 kg | 0
mild dyspnea | 0
adenoid cystic carcinoma in the carina | 0
carinal resection and reconstruction | 0
chest computed tomography | -24
bronchoscopy | -24
mass almost totally obstructed the left mainstem bronchus | -24
mass extended to the carina and right mainstem bronchus | -24
internal diameter of the RMB 11 mm | -24
length of the RMB 12 mm | -24
length of the distal LMB not involved by the mass 20 mm | -24
preoperative examinations were normal findings | -24
moderate obstructive pattern of the pulmonary function test | -24
forced expiratory volume in one second of 1.88 liter | -24
forced vital capacity of 2.81 liter | -24
ratio of 67% | -24
general anesthesia induced | 0
target-controlled infusion of propofol | 0
remifentanil | 0
rocuronium | 0
tracheal intubation | 0
right-sided double-lumen tube | 0
patient moved to the right lateral position | 0
left bronchi and vasculature dissected | 0
thoracoscopic surgery under right OLV | 0
arterial oxygen tension 462 mmHg | 20
inspired oxygen fraction 1.0 | 20
right-sided double-lumen tube replaced | 20
single-lumen endotracheal tube | 20
bronchial blocker | 20
left lateral position | 20
right thoracotomy | 20
peak airway pressure 28 cmH2O | 40
tidal volume 300 ml | 40
PaO2 110 mmHg | 40
FIO2 1.0 | 40
carinal resection | 40
LMB resected | 40
sterile reinforced endotracheal tube | 40
left OLV | 40
airway pressure increased to 35 cmH2O | 40
oxygen saturation by pulse oximetry decreased to 70% | 40
RMB resected | 40
additional sterile endotracheal tube | 40
differential bilateral lung ventilation | 40
SpO2 restored to 100% | 42
carina removed | 42
lower trachea resected | 42
separated RMB anastomosed with the resected trachea | 42
no air leak in the anastomotic site | 42
left lung removed | 42
left endobronchial tube removed | 42
non-dependent right lung ventilated | 42
low tidal volume of 200-250 ml | 42
airway pressure lower than 20 cmH2O | 42
SpO2 decreased below 80% | 42
tube reinserted into the LMB | 42
both lungs ventilated | 42
sufficient two-lung ventilation | 47
FIO2 1.0 | 47
right OLV reattempted | 47
SpO2 decreased below 90% | 50
left pulmonary artery clamped | 50
right OLV attempted | 50
SpO2 maintained 100% | 55
left main pulmonary artery ligated | 55
silicone vascular loop | 55
ligating clip | 55
left endobronchial tube removed | 55
right thoracotomy closed | 55
PaO2 360 mmHg | 115
FIO2 1.0 | 115
patient moved to the right lateral position | 115
left thoracotomy | 115
left pulmonary artery and veins resected | 115
left pneumonectomy completed | 115
patient shifted to the supine position | 115
chin tightly sutured to the chest | 115
tracheal extubation | 115
patient transferred to the intensive care unit | 115
discharged on the 13th postoperative day | 318
no complications | 318