85 years old | 0
male | 0
admitted to the hospital | 0
dog bite | -360
fever | -48
aggressive behavior | -120
mental confusion | -120
psychomotor agitation | -120
impaired consciousness | -120
healing wound | 0
nuchal rigidity | 0
Brudzinski’s sign | 0
leukocytosis | 0
low platelet cell count | 0
elevated C-reactive protein | 0
normal liver function tests | 0
normal renal function tests | 0
normal glycosylated hemoglobin level | 0
negative Anti-HIV 1/2 Western blot | 0
negative blood cultures | 0
positive RT-PCR for SARS-CoV-2 | 0
normal cranial computed tomography | 0
cerebrospinal fluid analysis | 0
glucose levels of 9 mg/dL | 0
protein concentration of 171.3 mg/dL | 0
white blood cell count of 727 cells/mm3 | 0
CSF Gram stain with gram-negative bacilli | 0
CSF culture | 48
translucent, spotty and flat colonies | 48
identification of C. canimorsus | 48
treatment with ceftriaxone | 0
no clinical improvement | 120
treatment with meropenem | 120
clinical response | 120
admitted to ICU | 0
discharged from ICU | 120
discharged from hospital | 336
full clinical resolution of symptoms | 336
no sequelae at six-month follow-up | 4320