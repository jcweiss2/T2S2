57 years old | 0
female | 0
diabetes | 0
hypertension | 0
transferred to our facility | 0
high-grade fever | -72
fall | -336
initial treatment at a primary health center | -336
ambulating well at home | -336
conscious | 0
oriented | 0
febrile | 0
hypotensive | 0
minimal respiratory distress | 0
sepsis due to unknown source | 0
managed with fluid resuscitation | 0
cultures | 0
imaging to identify potential source | 0
broad-spectrum antibiotics | 0
leukocytosis | 0
toxic neutrophil granulation | 0
normal renal panel | 0
normal liver panel | 0
normal coagulation panel | 0
electrocardiogram: right axis deviation | 0
electrocardiogram: S1Q3T3 pattern | 0
echocardiography: no right heart strain | 0
lower limb venous Doppler: no DVT | 0
compression ultrasound: no DVT | 0
CT pulmonary angiogram ruled out PE | 0
initiated on unfractionated heparin | 0
blood cultures grew MSSA | 0
antibiotic de-escalated | 0
patient gradually improving | 0
rest of cultures negative | 0
tropical infections screening negative | 0
CT abdomen revealed D8 vertebral fracture | 0
transesophageal echocardiography: no infective endocarditis | 0
acute left lower limb swelling | 24
left lower limb pain | 24
left lower limb redness | 24
repeat venous Doppler: acute DVT | 24
DVT extending from left internal iliac to popliteal vein | 24
normal coagulation profile | 24
normal platelet count | 24
peripheral smear normal | 24
connective tissue workup negative | 24
vasculitis workup negative | 24
therapeutic anticoagulation with heparin | 24
MRI spine: T8 and T11 wedging | 24
MRI spine: no cord edema | 24
MRI spine: no cord mass | 24
compression of left common iliac vein by right common iliac artery | 24
acute thrombus in left common iliac vein | 24
May-Thurner syndrome diagnosis | 24
catheter-based thrombolysis suggested | 24
venous stenting suggested | 24
IVC filter placement | 24
long-term anticoagulation with rivaroxaban | 24
afebrile at discharge | 168
stable at discharge | 168
asymptomatic during follow-up | 672
