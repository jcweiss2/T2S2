male | 0
born | 0
uncomplicated pregnancy | 0
cesarean section | 0
gestational weeks | 0
birth weight | 0
height | 0
head circumference | 0
no history of consanguinity | 0
no known genetic disorders | 0
admitted to pediatric intensive care unit | -84
RSV infection | -84
failure to thrive | -84
bulging of the anterior fontanel | -84
lumbar puncture | -84
severe intracranial hypertension | -84
CSF analysis | -84
negative for central nervous system infection | -84
extensive external hydrocephalus | -84
need for ventriculoperitoneal shunt placement | -84
rapid improvement of the clinical condition | -84
deflection of the growth curve | -84
radiographs of the entire skeleton | -84
generalized sclerosis of the bone | -84
diagnosis of infantile osteopetrosis | -84
bone marrow biopsy | -84
osteoclast-poor osteopetrosis | -84
genetic testing | -84
homozygous TCIRG1 mutation | -84
allogeneic HSCT | -35
conditioning with busulphan | -35
conditioning with fludarabin | -35
conditioning with melphalan | -35
conditioning with anti-thymocyte globulin | -35
referred to the department of Otorhinolaryngology | -35
clinical and audiological evaluation | -35
newborn hearing screening | -168
brainstem audiometric testing | -35
normal hearing | -35
neurologic and ophthalmologic evaluation | -35
normal cranial nerve functions | -35
impaired vision of the right eye | -35
recurrent episodes of acute otitis media | 108
recurrent episodes of otitis media with effusion | 108
bilateral tympanostomy tubes | 108
persistent OME | 108
impact on hearing acuity | 108
free-field audiometry preoperative | 108
bluish mass behind the right tympanic membrane | 108
dehiscent jugular bulb | 108
middle ear effusion | 108
placement of tympanostomy tubes | 108
hearing test postoperatively | 108
low frequency | 108
severe conductive hearing loss | 108
cone beam CT scan | 108
small tympanic cavity | 108
thickened superstructures | 108
thickened footplates | 108
upward and medial angulation of the petrous bone apex | 108
rehabilitation with a conventional or bone-anchored hearing aid | 108
no recurrence of otitis media | 240
no need for replacing tympanostomy tubes | 240
audiometric thresholds remain stable | 240
good functional results | 240
monocular blindness | 240
good general health | 240
favorable development | 240
stable blood values | 240
since allogeneic HSCT | 240