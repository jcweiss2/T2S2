84 years old|0
    hip joint endoprosthesis|0
    increased bleeding during operation|0
    postoperative anemia|0
    hemodynamic instability|0
    received 3 units of packed red blood cells|0
    fever|312
    antibiosis with piperacillin-tazobactam|312
    diarrhea|312
    deterioration|312
    intensive care unit admission|384
    severe septic shock|384
    circulatory failure|384
    lactic acidosis|384
    blood smear ordered|384
    high concentration of plasmodia detected|384
    rapid test positive for Plasmodium falciparum|384
    artesunate administration|384
    ventilation|408
    hemodynamic support|408
    death|432
    no travel history|0
    Plasmodium falciparum transmission via packed red blood cells|0
    look back process initiated|0
    donor with multiple donations|0
    recent travel to malaria endemic country|0
    malaria contracted without symptoms|0
    blood donation 2 weeks after return from endemic area|0
    donor did not mention recent return from endemic area|0
    donor did not report intake of malaria prophylaxis drugs|0
    donor released to donate whole blood|0
    donor had general symptoms of illness|408
    donor had fever|408
    donor did not report symptoms|408
    donor diagnosed with malaria|408
    no information passed to blood transfusion service|408
    donor took malaria prophylaxis|408
    negligent manslaughter|432
    donor confronted with legal consequences|432
    indictment by public prosecutor|432
    sentenced to criminal fine|432
    heirs sued for damages|432
    donor convicted under civil law|432
    bereavement compensation|432
    funeral expenses|432
    judgment not legally binding|432
    
    <|eot_id|>
    84 years old|0
    hip joint endoprosthesis|0
    increased bleeding during operation|0
    postoperative anemia|0
    hemodynamic instability|0
    received 3 units of packed red blood cells|0
    fever|312
    antibiosis with piperacillin-tazobactam|312
    diarrhea|312
    deterioration|312
    intensive care unit admission|384
    severe septic shock|384
    circulatory failure|384
    lactic acidosis|384
    blood smear ordered|384
    high concentration of plasmodia detected|384
    rapid test positive for Plasmodium falciparum|384
    artesunate administration|384
    ventilation|408
    hemodynamic support|408
    death|432
    no travel history|0
    Plasmodium falciparum transmission via packed red blood cells|0
    look back process initiated|0
    donor with multiple donations|0
    recent travel to malaria endemic country|0
    malaria contracted without symptoms|0
    blood donation 2 weeks after return from endemic area|0
    donor did not mention recent return from endemic area|0
    donor did not report intake of malaria prophylaxis drugs|0
    donor released to donate whole blood|0
    donor had general symptoms of illness|408
    donor had fever|408
    donor did not report symptoms|408
    donor diagnosed with malaria|408
    no information passed to blood transfusion service|408
    donor took malaria prophylaxis|408
    negligent manslaughter|432
    donor confronted with legal consequences|432
    indictment by public prosecutor|432
    sentenced to criminal fine|432
    heirs sued for damages|432
    donor convicted under civil law|432
    bereavement compensation|432
    funeral expenses|432
    judgment not legally binding|432