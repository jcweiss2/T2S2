65 years old | 0
male | 0
no history of smoking | 0
no underlying pulmonary diseases | 0
admitted to the hospital | 0
4-day history of shortness of breath | -96
fever | -96
dry cough | -96
fatigue | -96
breath sounds were reduced | 0
oxygen saturation (SpO2) was 93% | 0
bilateral peripheral ground-glass attenuation | 0
patchy consolidation | 0
lung involvement was 60%-70% | 0
nasopharyngeal SARS-CoV-2 RT-PCR test was positive | 0
symptoms gradually worsened | 0
increased temperature | 0
saturation with free breathing decreased to 90% | 0
white cell count: 7.93 х 109/ L | 0
hemoglobin 159 g/l | 0
platelet count: 468 х 109/l | 0
Westergren ESR 41 mm/h | 0
interleukine 6 102 pg/ml | 0
С-reactive protein 142 mg/l | 0
ferritin 939.92 μg/ml | 0
D-dimer 609 ng/ml | 0
procalcitonin 0,11 ng/ml | 0
treatment of SARS-CoV-2 infection included dexamethason | 0
heparin | 0
tocilizumab | 0
acetylcysteine | 0
pantoprazole | 0
nadroparin calcium | 0
oxygen supplementation | 0
air and pleural effusion in the right pleural cavity | 360
collapse of the right lung | 360
thoracentesis | 360
thoracostomy | 360
1400 ml of a yellowish opaque liquid was evacuated | 360
linezolid and imipenem/cilastatin therapy | 360
daily drainage volume was from 300 to 1000 ml of fluid | 384
pleural effusion with gas bubbles | 432
focal area of subpleural infiltration | 432
central cavity of destruction | 432
air layer up to 47 mm of anteroposterior thickness | 432
radiological sings of the left side hydropneumothorax | 432
pleural fluid analysis confirmed an exudative lymphocytic-rich effusion | 432
Acinetobacter baumannii and Pseudomonas aeruginosa were cultured | 432
urine culture was positive for Klebsiella pneumonia | 432
needle thoracocentesis and new pleural drainage | 504
air and creamy purulent mass have been aspirated | 504
200 to 800 ml of serofibrinous hemorrhagic fluid was drawn daily | 504
diagnosis of pleural empyema | 540
transferred to the Surgical Department | 540
right pleural space was daily irrigated with antiseptic solutions | 540
lung expansion was achieved by continuous vacuum aspiration technique | 540
encapsulated pleural effusion located in the upper anterior area of the right hemithorax | 624
ultrasound-guided puncture of this effusion was performed | 624
new drainage of the pleural cavity was installed | 624
4-week antibiotic therapy | 672
discharged from the hospital | 744
oxygen saturation (SpO2) was 97% on room air | 744
chest CT after chest tube removing showed the presence of a small amount of fluid | 744
lab test scores came back to normal range | 744
level of С-reactive protein was 11.7 mg/l | 744
procalcitonin < 0,1 ng/ml | 744