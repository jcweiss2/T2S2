40 years old | 0
female | 0
vomiting | -24
diarrhea | -24
loss of consciousness | -24
common cold treatment | -24
garenoxacin | -24
hypothyroidism | -6720
admitted to the hospital | 0
fever | -24
shock | 0
dopamine | 0
noradrenaline | 0
antibiotics | 0
referred to the Critical Care Center | 24
body temperature 38.6°C | 24
blood pressure 62/46 mmHg | 24
heart rate 100-110 beats/min | 24
respiratory rate 20 breaths/min | 24
oxygen saturation 100% | 24
Glasgow Coma Scale 15/15 | 24
elevated white blood cell count | 24
elevated C-reactive protein | 24
elevated procalcitonin | 24
sepsis-induced disseminated intravascular coagulation | 24
elevated creatinine kinase | 24
elevated creatinine kinase MB | 24
elevated troponin T | 24
sequential organ failure assessment score 8 | 24
septic shock with unknown focus | 24
antibiotics (meropenem, vancomycin, clindamycin) | 24
intravenous immunoglobulin | 24
vasoactive agents (noradrenaline and arginine vasopressin) | 24
hydrocortisone | 24
dobutamine | 24
pulse-induced contour cardiac output monitoring | 24
low cardiac output | 24
intubated | 24
mechanical ventilation | 24
circulatory status not improved | 120
electrocardiography revealed widespread ST elevation | 120
echocardiography revealed reduced left ventricular ejection fraction | 120
cardiogenic shock with concomitant septic shock | 120
coronary angiography | 120
Swan-Ganz catheter measurements | 120
intra-aortic balloon pumping (IABP) | 216
circulatory status stable | 216
improved left ventricle motion | 270
initiated CRRT | 270
reduced doses of noradrenaline and dobutamine | 600
discontinued dobutamine | 864
reduced IABP assist ratio | 960
discontinued IABP | 1728
discontinued vasoactive agents | 1728
fever resolved | 144
discontinued CRRT | 168
discontinued mechanical ventilation | 264
echocardiography showed improved LVEF | 168
inflammatory markers improved | 168
discontinued antibiotics | 336
posttreatment investigation for pathogens | 408
returned to the previous hospital for rehabilitation | 528
thyroid function normal | 1368