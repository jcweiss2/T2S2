39 years old | 0
male | 0
admitted to the hospital | 0
intermittent fever | -720
moderate exertion dyspnoea | -168
orthopnoea | -24
systolic murmurs in aortic and pulmonary areas | 0
elevated C-reactive protein | 0
leucocytosis | 0
neutrophilia | 0
anaemia | 0
empiric antibiotic therapy started | 0
piperacillin–tazobactam | 0
transoesophageal echocardiography | 24
vegetation attached to the non-coronary cusp of the aortic valve | 24
severe aortic regurgitation | 24
aortic root abscess | 24
left ventricle-to-right atrium fistula | 24
blood cultures | 24
Capnocytophaga canimorsus | 24
ceftriaxone | 48
surgery | 72
aortic valve replacement | 72
closure of the fistula | 72
worsening of patient’s general condition | 360
acute mediastinitis | 360
pericardial abscess | 360
cardiac tamponade | 360
emergency surgery | 360
pericardial abscess culture | 480
Enterococcus faecalis | 480
ampicillin | 480
patient exits intensive care unit | 480
discharged | 912
antibiotic therapy | 912
metronidazole | 912
linezolid | 912
dog bite | -1440
owned a pet dog | -1440