2 years old | 0
male | 0
admitted to pediatric polyclinic | 0
fever | 0
fever one week before | -168
treated for upper respiratory tract infection | -168
developed fever again | -7
cesarean section | -730
birth weight 3450 g | -730
length 50 cm | -730
head circumference 35 cm | -730
hospitalized at the newborn intensive care unit | -730
hyperbilirubinemia | -730
neonatal sepsis | -730
no reproduction in the blood and urinary cultures | -730
physical examination normal | 0
body temperature 37.2 oC | 0
body weight 12.5 kg | 0
height 87 cm | 0
WBC 19.2x103/µL | 0
neutrophil 52.6% | 0
lymphocyte 37% | 0
Hb 10.7 g/dL | 0
HTC 31.9% | 0
MCV 74 fL | 0
RDW 16.8 | 0
Plt 332000x103/µL | 0
C-reactive protein 3.04 mg/dL | 0
biochemical parameters normal | 0
urine dipstick positive for leukocytes | 0
urine dipstick negative for blood/hemoglobin | 0
urine dipstick negative for nitrite | 0
leukocytes in urinary sediment | 0
amorphous crystals in urinary sediment | 0
urinary system ultrasound | 0
7.5-mm stone in the left ureter | 0
grade 2 hydronephrosis | 0
R. ornithinolytica in urinary culture | 0
antibiotic sensitivity report | 0
sensitive to trimethoprim/sulfamethoxazole | 0
sensitive to amoxicillin/clavulanic acid | 0
sensitive to gentamicin | 0
sensitive to cefuroxime axetil | 0
resistant to ampicillin | 0
urine sample and culture obtained with a catheter | 24
oral cefuroxime axetil started | 24
urinary culture taken with the catheter | 48
105 CFU/mL R. ornithinolytica reproduced | 48
antibiotic sensitivity report same as former one | 48
immunoglobulins normal | 48
tests for stone etiology ordered | 48
calcium/creatinine normal | 48
oxalate normal | 48
citrate normal | 48
magnesium normal | 48
uric acid normal | 48
endoscopic stone removal | 72
double J catheter introduced | 72
follow-up of the patient | 120
remission of hydronephrosis | 120
cefuroxime therapy for 10 days | 120
follow-up urine culture negative | 240