32 years old | 0  
    male | 0  
    admitted to the hospital | 0  
    fever | -48  
    cough | -48  
    shortness of breath | -48  
    diarrhea | -96  
    denied diarrhea on admission | 0  
    denied chest pain | 0  
    denied abdominal pain | 0  
    denied nausea | 0  
    denied vomiting | 0  
    exposure to father with similar symptoms | -48  
    father admitted to hospital to rule out SARS-CoV-2 | -48  
    no known sick contacts | 0  
    admitted to rule out community acquired pneumonia | 0  
    admitted to rule out viral syndrome secondary to SARS-CoV-2 | 0  
    admitted to rule out viral syndrome secondary to influenza | 0  
    regular heart rate | 0  
    regular heart rhythm | 0  
    no murmurs | 0  
    no rubs | 0  
    no gallops | 0  
    no jugular venous distension | 0  
    lungs clear to auscultation bilaterally | 0  
    ecchymosis from cupping marks on back | 0  
    normotensive | 0  
    no tachycardia | 0  
    respiratory rate 18 breaths per min | 0  
    oxygen saturation 95% on room air | 0  
    unremarkable complete blood count | 0  
    hyperglycemia 282 mg/dL | 0  
    hemoglobin A1c 14% | 0  
    elevated lactate dehydrogenase 792 U/L | 0  
    elevated C-reactive protein 126.61 mg/L | 0  
    mild acidemia | 0  
    normal sinus rhythm on electrocardiogram | 0  
    no QTc prolongation | 0  
    chest X-ray showing peripheral patchy opacities | 0  
    started on IV ceftriaxone | 0  
    started on IV azithromycin | 0  
    started on IV hydroxychloroquine | 0  
    started on oral zinc supplementation | 0  
    SARS-CoV-2 RNA nasal swab sent for RT-PCR | 0  
    influenza A and B antigen nasal swab sent for RT-PCR | 0  
    desaturated to 79% SpO2 | 0  
    required 6 L/min supplemental oxygen | 0  
    switched to high-flow nasal cannula | 0  
    IV linezolid added | 0  
    insulin regimen started | 0  
    SARS-CoV-2 RNA positive | 24  
    influenza A positive | 24  
    oseltamivir added | 24  
    chest CT showing bilateral ground-glass opacities | 24  
    continuous fever spikes | 0  
    stable until hospital day 5 | 120  
    worsening tachypnea | 120  
    increased FiO2 requirement | 120  
    worsening PaO2/FiO2 ratio | 120  
    SpO2 87% on HFNC | 120  
    respiratory rate 28-32 breaths per min | 120  
    repeat chest X-ray showing worsening opacities | 120  
    elevated ferritin 884 ng/mL | 120  
    persistently elevated LDH 870 U/L | 120  
    arterial blood gas showing hypoxia | 120  
    elevated bicarbonate level | 120  
    ARDS secondary to sepsis | 120  
    sepsis secondary to coinfection with SARS-CoV-2 | 120  
    sepsis secondary to coinfection with influenza A | 120  
    intubated | 120  
    mechanical ventilation | 120  
    upgraded to ICU | 120  
    IV tocilizumab | 120  
    acute kidney injury | 120  
    anuric | 120  
    hemodialysis started | 120  
    linezolid discontinued | 120  
    IV meropenem started | 120  
    IV lopinavir and ritonavir started | 120  
    self-extubated | 120  
    transitioned to BIPAP | 120  
    transitioned to HFNC | 120  
    downgraded to medical floor | 120  
    found hypoxic | 120  
    repeat chest X-ray showing worsening opacities | 120  
    BIPAP placed again | 120  
    respiratory distress | 120  
    re-intubated | 120  
    placed back in ICU | 120  
    died | 120  
    
    