79 years old | 0
female | 0
on a ventilator | 0
biliary sepsis | -168
treated with antibiotics | -168
treated with supportive treatment | -168
jaundiced | 0
heart problems | 0
hypothyroidism | 0
diabetes mellitus | 0
high total bilirubin | 0
high direct bilirubin | 0
high CRP | 0
abdominal ultrasound | -168
MRI evaluation | -168
large cyst | -168
gastric compression | -168
bile duct obstruction | -168
large stone | -168
piperacillin-tazobactam | 0
amikacin | 0
levothyroxine | 0
insulin therapy | 0
supportive treatments | 0
abdominal MRI review | 0
pancreatic pseudocyst | 0
biliary drainage | 0
bedside biliary drainage procedure | 24
transabdominal US guidance | 24
dilated bile duct | 24
bile fluid aspiration | 24
guide wire insertion | 24
PTBD pigtail catheter insertion | 24
cyst evaluation | 48
infected cyst | 48
cyst fluid analysis | 48
amylase | 48
lipase | 48
CEA | 48
decreased bilirubin | 72
decreased CRP | 72
breathing improvement | 72
ventilator mode change | 72
pigtail catheter dislodged | 144
ERCP procedure | 144
cholangiogram | 144
large stone | 144
7-Fr double-pigtail stent | 144
EUS procedure | 144
cyst evaluation | 144
cyst puncture | 144
guide wire insertion | 144
cystotome | 144
7-Fr double-pigtail stent insertion | 144
improved condition | 168
spontaneous breathing | 168
discharged from ICU | 168
discharged from hospital | 240
repeat ERCP procedure | 2160
CBD stone crushing | 2160
pancreatic cyst reduction | 2160
pancreatic cyst stent maintenance | 2160