57 years old | 0
female | 0
right lateral ankle pain | -12
ankle injury | -12
swelling on lateral aspect | -12
physical exam: swelling | 0
2 cm round ecchymotic lesion | 0
limited range of motion | 0
intact pulses | 0
no other skin findings | 0
right leg x-ray | 0
lateral malleolar edema | 0
no acute osseous findings | 0
discharged | 0
worsening swelling | 6
ecchymotic lesion expansion | 6
increased pain | 6
shortness of breath | 6
cardiac arrest | 6
hypoxic respiratory failure | 6
intubated | 6
hypotension | 6
sinus tachycardia | 6
mechanically ventilated | 6
extensive hemorrhagic lesion | 6
bullous formation | 6
white blood cell count 3.3 K/mm3 | 6
hemoglobin 8.9 g/dL | 6
mean corpuscular volume 112.8 fL | 6
platelet count 36 K/mm3 | 6
potassium 5.1 mmol/L | 6
carbon dioxide 11 mmol/L | 6
anion gap 33 mEq/L | 6
creatinine 2.9 mg/dL | 6
lactic acid 21.4 mmol/L | 6
total bilirubin 1.7 mg/dL | 6
aspartate transaminase 327 U/L | 6
alanine transaminase 164 U/L | 6
troponin 0.110 ng/mL | 6
prothrombin time 25.9 seconds | 6
INR 2.25 | 6
fibrinogen 318 mg/dL | 6
d-dimer 5200 ng/mL | 6
creatinine kinase 3197 U/L | 6
arterial blood gas: pH 6.69 | 6
pCO2 69.1 mmHg | 6
HCO3 8.3 mmol/L | 6
chest x-ray clear | 6
endotracheal tube | 6
head CT: subarachnoid hemorrhage | 6
chest CT angiography: no pulmonary embolism | 6
admitted to ICU | 6
intravenous fluids | 6
blood cultures obtained | 6
general surgery consulted | 6
intravenous vancomycin | 6
intravenous meropenem | 6
intravenous clindamycin | 6
bedside fasciotomy | 6
bedside below knee guillotine amputation | 6
tissue cultures obtained | 6
second blood cultures | 6
progression of acidosis | 6
nephrology consulted | 6
continuous renal replacement therapy | 6
worsening acidosis | 24
multiple pressors | 24
clinical deterioration | 24
expired | 24
blood cultures: P. fluorescens | 24
tissue cultures: P. putida | 24
