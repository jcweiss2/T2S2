55 years old | 0
male | 0
admitted to the intensive care unit | 0
ingestion of sodium chlorite | -24
ingestion of whiskey | -24
ingestion of ibuprofen | -24
attempted hanging | -24
found lying on the floor | -24
cyanotic | -24
lowered consciousness | -24
inadequate response to verbal stimulus | -24
vomiting | -24
transported to the emergency department | -24
Glasgow Coma Scale score 13 | 0
body temperature 33.6°C | 0
heart rate 110/min | 0
blood pressure 150/80 mmHg | 0
respiratory rate 28/min | 0
pulse oximetry 65% | 0
generalized skin cyanosis | 0
neck markings after strangulation | 0
silent abdomen | 0
incontinence for urine and feces | 0
chocolate brown serum | 0
no abnormalities on further physical examination | 0
depression | 0
previous suicide attempt | 0
alcohol abuse | 0
no regular medication | 0
sedated | 0
intubated | 0
mechanically ventilated | 0
hemoglobin 179 g/L | 0
erythrocytes 5.45 × 10^12/L | 0
hematocrit 0.54 | 0
leukocytes 28.5 × 10^9/L | 0
platelet count 279 × 10^9/L | 0
BUN 5.5 mg/dL | 0
creatinine 142 μmol/L | 0
potassium 7.5 mM | 0
osmolality 351 mosm/L | 0
arterial lactate 6.5 mM | 0
myoglobin 433 ng/mL | 0
bilirubin 28 mM | 0
normal liver enzymes | 0
normal coagulation factors | 0
arterial blood gas pH 7.25 | 0
PaCO2 4.45 kPa | 0
PaO2 52.45 kPa | 0
BE −12.2 mmol/L | 0
HCO3 14.1 mmol/L | 0
SaO2 99% | 0
lactate 6.48 mmol/L | 0
MetHb 40.1% | 0
alcohol in blood 2 mg/g | 0
ibuprofen in gastric content | 0
ibuprofen in urine | 0
gastric fibroscopy | 0
superficial necrotic spots in antrum, stomach body, duodenum | 0
edema of pylorus | 0
ulcérations in upper esophagus, stomach, duodenum after 3 days | 72
electrocardiogram showed peaked T waves | 0
normal chest x ray | 0
normal CT scan of brain | 0
methylene blue therapy | 2
continuous venovenous hemodiafiltration initiated | 4.5
hyperkalemia | 4.5
metabolic acidosis | 4.5
hemodialysis for hyperkalemia | 4.5
lactate dropped to 2.55 mmol/L | 14
MetHb decreased to 15.2% | 14
MetHb decreased to 10.2% | 29
hemolytic anemia | 24
disseminated intravascular coagulation | 24
hemoglobin dropped from 179 to 116 g/L | 24
thrombocytes dropped from 279 to 164 × 10^9/L | 24
D dimer 29.1 mg/mL | 24
INR 1.8 | 24
APTT ratio 1.4 | 24
hemoglobin dropped to 59 g/L | 120
platelet count dropped to 77 × 10^9/L | 120
packed red blood cells transfused | 120
norepinephrine drip instituted | 20
hypotension 80/60 mmHg | 20
bronchopneumonia | 192
sepsis | 192
body temperature 39°C | 192
antibiotics initiated | 192
gastric ulceration improved | 240
esophageal ulceration improved | 240
weaned from mechanical ventilation | 312
intermittent hemodialysis every second day | 408
started urinating 2500 mL/24h | 408
blood urea 12 mg/dL | 408
creatinine 428 μmol/L | 408
estimated GFR 15.6 mL/min | 408
transferred to medium care facility | 528
no further need of hemodialysis | 528
discharged from hospital | 1536
written informed consent | 1536
