32 years old | 0
    woman | 0
    history of intravenous drug use | 0
    attention deficit/hyperactivity disorder | 0
    presented for evaluation of fevers | -24
    presented for evaluation of chills | -24
    presented for evaluation of shortness of breath | -24
    fever | -168
    chills | -168
    generalized weakness | -168
    shortness of breath | -72
    non-smoker | 0
    did not consume alcohol | 0
    abusing fentanyl intravenously | -168
    on dextroamphetamine/amphetamine | 0
    denied exposure to other medications | 0
    denied exposure to chemicals | 0
    temperature 102.7 °Fahrenheit | 0
    blood pressure 102/56 mmHg | 0
    pulse 136 beats per minute | 0
    respiratory rate 38 breaths per minute | 0
    oxygen saturation 94% on room air | 0
    well-developed female | 0
    moderate respiratory distress | 0
    bilateral rhonchi | 0
    regular heart rhythm | 0
    tachycardia | 0
    no murmur | 0
    no rub | 0
    no gallop | 0
    WBC 12,200/mm³ | 0
    hemoglobin 10.9 g/dL | 0
    platelet count 85,000/mm³ | 0
    ESR 60 mm/hr | 0
    hyponatremia (sodium 124 mmol/L) | 0
    creatinine 2.8 mg/dL | 0
    BUN 98 mg/dL | 0
    NT-proBNP 1028 pg/mL | 0
    ECG sinus tachycardia | 0
    chest radiograph bilateral lower lobe infiltrates | 0
    chest radiograph small pleural effusions | 0
    IV fluids | 0
    levofloxacin | 0
    clinical deterioration | 24
    transferred to ICU | 24
    septic shock | 24
    acute respiratory failure | 24
    pressor support | 24
    mechanical ventilation | 24
    blood cultures gram-positive cocci | 24
    vancomycin therapy | 24
    transthoracic echocardiogram vegetation at tricuspid valve | 24
    moderate-to-severe tricuspid regurgitation | 24
    cardiothoracic surgery consulted | 24
    transesophageal echocardiogram patent foramen ovale | 24
    CT chest multiple cavitary peripheral lung nodules | 24
    septic emboli | 24
    non-oliguric AKI | 24
    renal replacement therapy | 24
    acute tubular necrosis | 24
    perfusion-related kidney injury | 24
    MSSA | 72
    oxacillin initiated | 72
    pressors weaned off | 336
    extubated | 336
    renal function recovery | 336
    bilateral nontender purpuric papules | 408
    bullous lesions | 432
    anterior knee lesions | 432
    lateral thigh lesions | 432
    no mucosal involvement | 408
    no palmar involvement | 408
    no abdominal pain | 408
    no arthralgias | 408
    no paresthesia | 408
    no fever | 408
    no chills | 408
    HIV negative | 408
    hepatitis B negative | 408
    p2-ANCA negative | 408
    c2-ANCA negative | 408
    cryoglobulin negative | 408
    rheumatoid factor negative | 408
    ANA weakly positive (1:40) | 408
    anti-ds DNA negative | 408
    complement C3 low (14 mg/dL) | 408
    complement C4 normal (28 mg/dL) | 408
    anti-HCV positive | 408
    HCV viral load 4.16 × 10⁵ IU/mL | 408
    no significant RBC changes | 408
    no significant leukocyte count changes | 408
    no significant kidney function changes | 408
    eosinophil count normal | 408
    bullous fluid no bacteria | 408
    gram staining negative | 408
    punch biopsies leukocytoclastic vasculitis | 408
    perivascular neutrophil infiltration | 408
    fibrinoid necrosis of small vessels | 408
    no bacteria | 408
    no fungi | 408
    no viral inclusions | 408
    oxacillin-associated LCV diagnosis | 408
    vancomycin started | 408
    oxacillin discontinued | 408
    skin lesion resolution | 408
    no scar formation | 408
    tricuspid valve replacement surgery | 720
    no perioperative complications | 720
    no recurrence of skin lesions | 720
    isolated cutaneous LCV | 0
    oxacillin-induced cutaneous LCV | 0
    