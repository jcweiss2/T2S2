23 years old | 0
female | 0
admitted to the regional hospital | 0
hypogastric pain | -168
vomiting | -168
expressive aphasia | 0
vertigo | 0
unsteady gait | 0
severe metabolic acidosis | 0
hyperlactataemia | 0
brain computed tomography | 0
lumbar puncture | 0
treated with i.v. bicarbonate | 0
treated with infusions | 0
treated with antipyretics | 0
pyrexia | 0
toxicology screening | 0
ethylene glycol in urine | 0
glycolic acid in urine | 0
treated with i.v. ethanol | 0
lost consciousness | 16
developed convulsions | 16
intubated | 16
admitted to the intensive care unit | 16
aspiration pneumonia | 16
sepsis | 16
renal failure | 16
treated with antibiotics | 16
treated with continuous haemodiafiltration | 16
CRRT used bicarbonate-buffered solutions | 16
citrate-calcium module | 16
estimated citrate level | 16
improvement of consciousness | 120
extubation attempt | 168
failed extubation | 192
reintubation | 192
dilatation tracheostomy | 288
bleeding from tracheostomy | 288
referred to the tertiary hospital | 384
intractable metabolic alkalosis | 384
two organ failures | 384
initial bronchoscopy | 384
atelectasis eliminated | 384
open bronchial tree | 384
microbiology specimens | 384
ceased antibiotics | 432
echocardiography | 384
mildly globally reduced ejection fraction | 384
thrombus in the right internal jugular vein | 384
chest X-ray | 384
infiltration of the right lower lobe | 384
metabolic alkalosis | 384
hypernatraemia | 384
elevation of the renal parameters | 384
urea | 384
serum creatinine | 384
total to ionised calcium ratio | 384
citrate accumulation | 384
high total plasma protein | 384
electrophoresis | 384
immunoassay on the free light chains | 504
free kappa | 504
free lambda | 504
kappa/lambda ratio | 504
treated with CRRT | 384
treated with RCA | 384
trisodium citrate | 384
calcium chloride replacement | 384
calcium-free lactate-buffered solution | 384
plasmatic natrium lowered | 408
normal acid-base parameters | 480
restored consciousness | 480
weaning of the respiratory support | 528
decannulated | 528
CRRT ceased | 552
restoration of diuresis | 552
transferred back to the regional hospital | 552
discharged home | 1152
good performance status | 1152
healed tracheostomy | 1152
normal renal functions | 1152