50 years old | 0
    male | 0
    fever | -336
    loss of appetite | -336
    watery diarrhea (more than 10 times per day) | -336
    heavy drinker for about 10 years | 0
    consumed approximately 250 g of alcohol per day in the previous 6 mo | -4320
    admission | 0
    increased WBC count (17280/μL) | 0
    increased neutrophils (82.4%) | 0
    increased C-reactive protein level (3.97 mg/dL) | 0
    increased total bilirubin level (8.0 mg/dL) | 0
    increased prothrombin time (55%) | 0
    hepatomegaly with severe steatosis | 0
    splenomegaly | 0
    diffuse, edematous colon | 0
    diagnosed with acute alcoholic hepatitis | 0
    diagnosed with infectious enteritis | 0
    alcohol abstinence | 0
    prescribed antibiotics | 0
    WBC count increased to 43650/μL | 0
    neutrophils increased to 85.7% | 0
    total bilirubin increased to 20.8 mg/dL | 0
    prothrombin time decreased to 34% | 0
    renal failure progressed | 0
    hyporesis | 0
    creatinine increased to 3.26 mg/dL | 0
    transferred to our hospital | 0
    fever | 0
    jaundice | 0
    anuria | 0
    ascites | 0
    pretibial edema | 0
    hepatomegaly | 0
    hepatic encephalopathy | 0
    flapping tremor | 0
    WBC count increased to 54000/μL | 0
    neutrophils increased to 85.7% | 0
    total bilirubin increased to 26.8 mg/dL | 0
    aspartate aminotransferase increased to 99 IU/L | 0
    alanine aminotransferase increased to 48 IU/L | 0
    NH3 increased to 92 μg/dL | 0
    albumin decreased to 4 g/dL | 0
    blood urea nitrogen increased to 71 mg/dL | 0
    creatinine increased to 3.26 mg/dL | 0
    CRP increased to 6.73 mg/dL | 0
    procalcitonin increased to 8.53 ng/mL | 0
    prothrombin time decreased to 32% | 0
    interleukin-6 increased to 116.09 pg/mL | 0
    tumor necrosis factor-α increased to 5.4 pg/mL | 0
    diagnosis of severe alcoholic hepatitis with multiple organ failure | 0
    diagnosis of severe infectious enteritis | 0
    Maddrey discriminant function score 66 | 0
    Glasgow alcoholic hepatitis score 11 | 0
    infection with multidrug resistance Pseudomonas aeruginosa | 0
    intensive care | 0
    plasma exchange | 0
    hemodialysis | 0
    antibiotics administration | 0
    no improvement of liver failure | 0
    granulocytapheresis (GCAP) performed | 336
    WBC count decreased to 46450/μL | 336
    total bilirubin improved to 15.8 mg/dL | 336
    GCAP performed three times within 1 week | 336
    WBC count improved to 35000/μL | 336
    interleukin-6 improved | 336
    tumor necrosis factor1-α improved | 336
    meropenem administered | 336
    levofloxacin administered | 336
    diarrhea improved | 336
    fever improved | 336
    laboratory parameters improved | 336
    disappearance of Pseudomonas aeruginosa | 336
    renal failure improved | 336
    transferred to previous hospital | 1680
    no steroids administered | 0
    