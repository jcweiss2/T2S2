40 years old | 0
female | 0
admitted to the hospital | 0
lower abdominal pain | -168
nonbilious vomiting | -168
loose stools | -168
breathlessness | -168
decreased urine output | -168
fever | -72
history of fever | -72
afebrile | 0
thin patient | 0
dry tongue | 0
no pedal edema | 0
no generalized lymphadenopathy | 0
pulse rate of 130/min | 0
blood pressure 96/80 mmHg | 0
oxygen saturation 90% | 0
respiratory rate 34/min | 0
body temperature 98.4°F | 0
tenderness in the right iliac fossa | 0
no palpable mass | 0
audible bowel sounds | 0
hemoglobin 98 g/L | 0
high total leukocyte count | 0
platelet count 263.4 × 10^9/L | 0
deranged renal function | 0
urea 42.83 mmol/L | 0
creatinine 159.12 mmol/L | 0
electrolyte tests within normal limits | 0
liver function profile abnormal | 0
total bilirubin 12.65 mmol/L | 0
direct bilirubin 6.15 mmol/L | 0
alanine aminotransferase 8.2 mkat/L | 0
aspartate aminotransferase 50.9 mkat/L | 0
alkaline phosphatase 247.6 U/L | 0
gamma-glutamyl transferase 25.2 U/L | 0
total protein 57 g/L | 0
albumin 30.8 g/L | 0
hepatitis C virus positive | 0
bilateral moderate pleural effusion | 0
plain chest X-ray | 0
screening two-dimensional echocardiography | 0
no abnormality on echocardiography | 0
intravenous normal saline | 0
pain management | 0
supplemental oxygen | 0
empirical intravenous antibiotic therapy | 0
ceftriaxone 1 g every 12 h | 0
metronidazole 500 mg every 8 h | 0
ultrasound-guided thoracic paracentesis | 2
purulent aspirate | 2
pleural fluid sent for analysis | 2
lactate dehydrogenase level raised | 2
serum procalcitonin elevated | 2
abdominal ultrasound scan | 2
intrabdominal collection | 2
contrast-enhanced computed tomography scan | 4
bilateral pleural effusion | 4
multiple subcentimetric ground-glass centrilobular nodules | 4
acute appendicitis with rupture | 4
adjacent collection extending in the right posterior pararenal and perihepatic spaces | 4
suspicious communication between the peritoneal and pleural cavities | 4
COVID-19 pneumonia in differential diagnosis | 0
hollow viscus perforation with acute respiratory distress syndrome in differential diagnosis | 0
disseminated tuberculosis in differential diagnosis | 0
non-Hodgkin lymphoma with chylothorax in differential diagnosis | 0
RT-PCR test negative for COVID-19 | 4
erect chest X-ray | 4
no free air under the right dome of the diaphragm | 4
pleural fluid analysis favoring infective nature | 4
adenosine deaminase level high | 4
triglyceride levels in pleural fluid within normal limits | 4
bilateral intercostal tube drainage | 6
ultrasound guidance | 6
local anesthesia | 6
evacuation of purulent content | 6
urgent exploratory laparotomy | 12
appendectomy | 12
retroperitoneal collection | 12
gangrenous appendix | 12
injection noradrenaline 8 mg at 2 ml/h | 12
inotrope | 12
hypotension | 12
patient not extubated | 12
ionotropic support | 12
ventilatory support | 12
ICU admission | 12
mean arterial pressure | 12
noradrenaline support increased | 72
injection vasopressin at 2 units/h | 72
postoperative evolution satisfactory | 72
average urine output maintained | 72
kidney function tests within normal limits | 72
urea 6.7 mmol/L | 72
creatinine 97 mmol/L | 72
tracheostomy | 168
total parenteral nutrition | 168
ionotropic support tapered | 240
cessation of ionotropic support | 240
bilateral ICD outputs monitored | 240
bilateral ICD removed | 264
Klebsiella pneumoniae on culture medium | 240
pleural fluid culture revealed K. pneumoniae | 240
antibiotics adjusted | 240
blood culture negative | 240
pus evacuated from pleural cavity | 240
no AFB on Ziehl-Neelsen staining | 240
cartridge-based nucleic acid amplification test negative for tuberculosis | 240
histopathological examination of the appendix | 240
transmural necrosis of the appendicular wall | 240
dense acute inflammatory infiltrates | 240
bacterial colonies | 240
right-sided ICD removal | 216
left-sided ICD removal | 264
Ryle’s tube feeding | 264
oral feeds | 408
decannulation | 408
weaned off ventilator | 432
shifted out of ICU | 432
healing laparotomy wound | 432
suture removal | 504
monitored in high-dependency unit | 504
discharged | 504
follow-up visit | 720
no fresh complaints | 720
able to carry out daily activities | 720