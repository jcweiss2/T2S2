31 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
SLE | -8760 | 0 | Factual
lupus nephritis | -8760 | 0 | Factual
prior stroke | -8760 | 0 | Factual
intravenous drug use | -8760 | 0 | Factual
cardiogenic shock | 0 | 0 | Factual
mental status changes | 0 | 0 | Factual
elevated jugular venous pressure | 0 | 0 | Factual
prominent v wave | 0 | 0 | Factual
body temperature 36.3°C | 0 | 0 | Factual
blood pressure 95/66 mm Hg | 0 | 0 | Factual
heart rate 94 beats/min | 0 | 0 | Factual
hemoglobin 10.3 g/dL | 0 | 0 | Factual
white blood cell count 18.9 × 10^9/L | 0 | 0 | Factual
platelet count 64 × 10^9/L | 0 | 0 | Factual
international normalized ratio 3.6 | 0 | 0 | Factual
creatinine level 1.7 mg/dL | 0 | 0 | Factual
drug studies positive for narcotics | 0 | 0 | Factual
drug studies positive for cannabis | 0 | 0 | Factual
antiphospholipid serology normal | 0 | 0 | Factual
blood cultures negative | 0 | 0 | Factual
infectious endocarditis considered | 0 | 0 | Possible
broad-spectrum intravenous antibiotics | 0 | 24 | Factual
mitral valve replacements | -720 | -168 | Factual
NBTE | -720 | 0 | Factual
mitral valve prosthesis dehiscence | 0 | 0 | Factual
severe perivalvular regurgitation | 0 | 0 | Factual
annular pseudoaneurysm | 0 | 0 | Factual
fourth sternotomy | 24 | 24 | Factual
mitral valve annulus reconstruction | 24 | 24 | Factual
bioprosthesis integration | 24 | 24 | Factual
left atrial dome reconstruction | 24 | 24 | Factual
interatrial septal incision reconstruction | 24 | 24 | Factual
postoperative TEE | 24 | 24 | Factual
well-seated mitral valve bioprosthesis | 24 | 24 | Factual
mean gradient 3 mm Hg | 24 | 24 | Factual
no regurgitation | 24 | 24 | Factual
extracorporeal membrane oxygenation | 24 | 120 | Factual
multiple blood product transfusions | 24 | 120 | Factual
layered thrombus in left atrium | 120 | 120 | Factual
surgical clot removal | 120 | 120 | Factual
thrombus reaccumulation | 120 | 120 | Factual
extracorporeal membrane oxygenation withdrawn | 120 | 120 | Factual
patient died | 120 | 120 | Factual
autopsy declined | 120 | 120 | Factual