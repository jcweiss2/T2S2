66 years old|0
male|0
intense abdominal pain|0
acute renal failure|0
urea 178 mg/dL|0
serum creatinin 7.92 mg/dL|0
erroneous receipt of high dose amphotericin B deoxycholate|0
nasal leishmaniasis|0
HIV infection|-120
non-adherent to treatment|-120
gastroesophageal reflux disease|-120
former smoker|-120
HIV viral load 92,494 copies/ml|-120
CD4 count 5 cells/mm3|-120
CD4/CD8 ratio 0.08|-120
pancytopaenic|0
haemoglobin 6.0 g/dL|0
leucocytes 1,620 cells/μL|0
lymphocytes 142 cells/μL|0
platelets 64,000 cells/μL|0
afebrile|0
emaciated|0
severe nasal lesion|0
ulcer in the hard palate|0
extensive necrotic lesion involving left nasal ala and septum|0
dysphonic|0
chest computed tomography scan revealed consolidative lesions in both lungs|0
small bilateral pleural effusions|0
no treatment started for the lungs lesions|0
haemodialysis required during hospitalization|0
worsening renal failure after receiving treatment for nasal leishmaniasis|0
received 16 days of amphotericin B treatment|0
first 3 days received 5 mg/kg/day d-AmB|0
switched to L-AmB 4 mg/kg/day|3
remained stable until episode of acute respiratory distress|16
pulmonary sepsis by P. aeruginosa|16
admission to the intensive care unit (ICU)|16
melena|16
severe blood dyscrasia|16
partial response to nasal lesion following treatment|16
testicular mass discovered|16
local swelling|16
hyperemia|16
ultrasound diagnosed multiseptate fluid collection on right scrotal testicle|16
thick walls measuring 3.2 × 2.5 cm|16
contact with the epididymis on the same side|16
diagnostic orchiectomy required|16
swollen testicle|16
areas of necrosis|16
fluid accumulation|16
unfavourable clinical outcome|16
died|25
genitourinary histoplasmosis diagnosed post-mortem|27
disseminated histoplasmosis|0
lack of awareness of this condition|0
testicular histoplasmosis|0
granulomatous inflammation|0
histopathology|0
culture of testicular sample analysis|27
misdiagnosis of nasal lesion as leishmaniasis|0
confusion between amastigotes and yeast structures|0
drug toxicity leading to paused antifungal therapy|0
testicular tuberculosis (TB)|0
granulomatous diseases|0
bilateral disease|0
unilateral disease|0
lack of common clinical presentation|0
diagnosis confirmed post-mortem|27
