61 years old | 0
    male | 0
    presented to the emergency department | 0
    diarrhea | -24
    hematochezia | -24
    melena | -24
    nausea | 0
    foul-smelling belching | 0
    vomiting | 0
    hematemesis | 0
    stabbing epigastric pain | 0
    radiation | 0
    intermittent chills | 0
    dizziness | 0
    fever | 0
    headache | 0
    recent travel | 0
    sick contacts | 0
    unusual food intake | 0
    ulcerative colitis | -168
    total proctocolectomy with ileal-anal anastomosis | -168
    remission of ulcerative colitis | 0
    bowel movements | 0
    diabetes mellitus | 0
    hypercholesterolemia | 0
    hypertension | 0
    sitagliptin-metformin | 0
    atorvastatin | 0
    enalapril | 0
    metoprolol tartrate | 0
    excessive NSAID consumption | 0
    smoking | 0
    alcohol abuse | 0
    hypotension | 0
    blood pressure 80/56 mmHg | 0
    pulse 60 | 0
    respiratory rate 16 | 0
    temperature 36°C | 0
    soft abdomen | 0
    non-distended abdomen | 0
    mild epigastric tenderness | 0
    rebound tenderness | 0
    guarding | 0
    leukocytosis | 0
    white blood cell count 20.9×10^9/L | 0
    elevated lactate | 0
    anion gap metabolic acidosis | 0
    bicarbonate 14.6 mEq/L | 0
    gap 14 mEq/L | 0
    sodium 135 mEq/L | 0
    potassium 3.9 mEq/L | 0
    acute kidney injury | 0
    creatinine 299 µmol/L | 0
    non-contrast CT findings of gastric emphysema | 0
    portal venous gas in liver | 0
    left adrenal nodule | 0
    intravenous fluids | 0
    piperacillin/tazobactam | 0
    intravenous pantoprazole | 0
    admission to intensive care unit | 0
    rapid resolution of symptoms | 0
    negative stool studies for Clostridium difficile | 0
    negative stool studies for Salmonella spp. | 0
    negative stool studies for Shigella spp. | 0
    negative stool studies for Campylobacter spp. | 0
    negative stool studies for Escherichia coli | 0
    diet advancement | 72
    improved renal function | 72
    follow-up CT abdomen with contrast | 72
    resolution of emphysematous gastritis | 72
    discharge home | 72
    oral pantoprazole | 72
    ciprofloxacin | 72
    metronidazole | 72
    follow-up with gastroenterology | 72
    upper endoscopy | 72
    follow-up CT abdomen in 6 months | 72
    stability of adrenal nodule | 72<|eot_id|>
    