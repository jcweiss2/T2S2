42 years old | 0
female | 0
granular dystrophy | 0
DALK | 0
big bubble technique | 0
8 mm recipient stromal flap partially dissected | 0
air injected into the substance of the remaining stroma | 0
donor button cut 8.25 mm | 0
DM peeled off | 0
donor button placed over the recipient DM | 0
sutured with recipient rim | 0
age of donor cornea 36 years | 0
in situ cornea excision | 0
surgery gone quite well | 0
whitish infiltrates along the graft-host junction | 24
severe anterior chamber reaction | 24
postoperative keratitis | 24
graft removed | 24
another stromal graft placed | 24
corneal scrapings sent for microbiology | 24
host DM clear and intact | 24
topical vancomycin started | 27
topical ceftazidime started | 27
Gram-stain showed Gram-negative Bacilli | 48
infiltrates along the entire graft host junction | 48
hypopyon | 48
topical antibiotics increased | 48
corneal scrapings revealed Klebsiella pneumoniae | 72
Klebsiella pneumoniae resistant to multiple antibiotics | 72
sensitive to imipenem, tigecycline, and partially sensitive to gatifloxacin | 72
imipenem drops started | 72
infiltration extended toward center of graft | 96
hypopyon persisted | 96
therapeutic penetrating keratoplasty | 120
infiltrates observed in host DM | 120
graft clear without infiltrates or hypopyon | 144
imipenem continued | 144
gatifloxacin drops added | 144
prednisolone drops added | 192
unaided vision 6/60 | 1008
vision improved to 6/18 with pin hole | 1008
graft clear | 1008
anterior segment quiet | 1008
intraocular pressure normal | 1008
pathogen eradicated | 1008