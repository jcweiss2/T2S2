26 years old | 0
male | 0
admitted to the acute surgical unit | 0
folliculitis | 0
multiple carbuncles |! 0
ulcerative colitis | -672
