47 years old | 0
male | 0
motor vehicle collision | -168
subarachnoid hemorrhage | -168
bilateral lung contusions | -168
rib fractures | -168
blunt abdominal injury | -168
lumbar fractures | -168
open-book pelvic fracture | -168
abdominal CT scan | -168
no ascites | -168
no free gas | -168
injury severity score 48 | -168
FAST | -96
presence of ascites | -96
diagnostic paracentesis | -96
dark green ascites | -96
emergency exploratory laparotomy | -96
mass intestinal fluid | -96
severe edema of the intestinal wall | -96
complete rupture of the jejunum | -96
primary anastomosis | -96
debridement of the injured area | -96
removal of the ruptured jejunum | -96
postoperative Gram-negative sepsis | -96
hypotension | -96
multiple vasopressors | -96
MODS | -96
AKI | -96
acute gastrointestinal injury | -96
hyperbilirubinemia | -96
hepatic dysfunction | -96
transfer to trauma referral center | 0
coma | 0
Glasgow coma scale score 2T1 | 0
shock | 0
heart rate 125 beats/min | 0
mean arterial pressure < 70 mmHg | 0
norepinephrine 1.2 mg·kg−1·min−1 | 0
acidosis | 0
pH 7.25 | 0
base excess −6.55 mEq/L | 0
lactic acid 3.92 mmol/L | 0
peritonitic | 0
jaundice | 0
admitted to TICU | 0
salvage resuscitation | 0
hemodynamic monitoring | 0
abdominal examinations | 0
serial laboratories | 0
imaging | 0
organ support | 0
digestive juice-like fluid drainage | 0
hemoglobin 78 g/L | 0
red-cell count 2.7 × 1012/L | 0
white-cell count 17.3 × 109/L | 0
platelet count 190 × 109/L | 0
prothrombin time 20 s | 0
activated partial thromboplastin time 50 s | 0
international normalized ratio 3.12 | 0
C-reaction protein 289.3 mg/L | 0
procalcitonin 10.7 ng/mL | 0
interleukin-6 826 ng/L | 0
albumin 26 g/L | 0
total bilirubin 391.5 μmol/L | 0
direct bilirubin 284.1 μmol/L | 0
indirect bilirubin 58.7 μmol/L | 0
alanine aminotransferase 35 U/L | 0
aspartate aminotransferase 58 U/L | 0
FAST ascites | 0
CT exudation | 0
dilated proximal jejunum | 0
DCS initiation | 24
hemodynamic instability | 24
MODS | 24
continuous renal replacement therapy | 24
bilirubin adsorption | 24
AKI | 24
hyperbilirubinemia | 24
hyperkalemia | 24
negative pressure irrigation tubes | 24
passive drainage to gravity | 24
broad-spectrum antibiotic therapy | 24
transfer to operating room | 48
intestinal fluid in abdominal cavity | 48
small intestinal edema | 48
complete rupture of primary anastomosis | 48
DCL | 48
temporary abdominal closure | 48
TDE creation | 48
postoperative transfer to TICU | 48
hemodynamic stability | 96
bioelectrical impedance analysis-directed fluid restriction | 96
ultrafiltration rate | 96
net negative fluid balance | 96
bedside dressing change | 96
split-thickness skin grafting | 1752
high risk of malnutrition | 0
Nutrition Risk Screening 2002 score 6 | 0
EN initiation | 96
glucose sodium chloride EN | 96
nasogastric tube | 96
proximal portion EN | 96
short peptide formula EN | 120
cholestatic cholecystitis | 96
percutaneous gallbladder puncture and drainage | 96
tracheostomy tube | 96
oral diet | 96
jejunal feeding tube insertion | 168
chyme reinfusion | 168
separation of intestinal adhesions | 168
clear abdominal drainage | 168
methylene blue injection | 168
chyme drainage | 168
chyme filtration | 168
chyme injection to distal TDE | 168
hermetic device | 168
trained nursing staff | 168
bilirubin adsorption | 168
bilirubin level decrease | 168
jaundice relief | 168
distal portion EN initiation | 192
short peptide formula | 192
supplemental enteral glutamine | 192
EN dosage increase | 192
protein increase | 192
standard EN formula | 432
weight gain | 432
laboratory normalization | 432
discharge to orthopedic department | 2280
home EN | 2280
home CR | 2280
staged reconstruction | 2280
jejunal feeding tube removal | 2280
anastomosis of TDE | 2280
abdominal wall reconstruction | 2280
regular diet | 2280
discharge | 2280
