51 years old | 0
man | 0
abdominal pain | 0
vomiting | 0
admitted | 0
suspected diagnosis of intestinal obstruction | 0
eaten uncertain quantities of persimmon | -several days
previous abdominal operation to repair small bowel perforation | -20 years
leukocytosis (19,240/µL) | 0
hemoglobin concentration of 18.3 g/dL | 0
normal C-reactive protein (0.07 mg/dL) | 0
body temperature 36.5℃ | 0
abdominal distension | 0
mild tenderness over epigastric area | 0
HIV antibody negative | 0
abdominal CT scan revealed mechanical obstruction in ileum | 0
ovoid bezoar 5.5 × 2.5 cm | 0
mild splenomegaly | 0
decrease of leukocytosis (7,690/µL) | 96
increase of C-reactive protein (4.02 mg/dL) | 96
symptoms not resolved by day 5 of hospitalization | 120
bezoar removal operation | 120
small bowel dilatation | 120
no signs of small bowel ischemia | 120
bezoar extracted through enterotomy | 120
decompression of dilated bowel | 120
postoperative recurrent fever >38℃ | 48
postoperative atelectasis | 48
passing flatus | 120
progressive diet started | 120
dyspnea | 168
chest radiography showed diffuse ground glass opacity | 168
ARDS diagnosed | 168
mechanical ventilation | 168
blood cultures collected postoperative day 4 | 96
started empiric fluconazole | 96
C. famata in blood cultures | 96
C. parapsilosis in blood cultures | 144
fluconazole treatment for 4 days | 96
fever persisted | 96
leukocytosis persisted | 96
history of antifungal treatment for tinea pedis 3 years ago | -three years
changed to amphotericin B | 96
methylprednisolone administered | 96
stool culture grew C. glabrata | 288
amphotericin-associated nephrotoxicity | 432
changed to caspofugin | 432
afebrile | 168
clinical improvement | 168
sterile blood cultures days 7, 10, 14 after antifungal therapy | 168
30-day antifungal therapy | 888
discharged | 888
ARDS caused by C. parapsilosis and C. famata | 168
no urinary or central venous catheters used | 0
Candida species other than C. albicans increased | 0
mucosal breakdown | 0
no immunocompromised state | 0
no self-administering illicit IV drugs | 0
reduced susceptibility to echinocandins and azoles | 0
initiation of liposomal amphotericin B | 96
small bowel bezoar as cause of candidemia | 0
