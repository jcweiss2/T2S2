49 years old | 0
male | 0
previously fit and well | 0
admitted to the emergency department | 0
swollen and painful scrotum and penis | -168
infective episode of balanitis | -672
Ciprofloxacin | -672
pyrexial | 0
temperature of 39°C | 0
swollen tender scrotum and penis | 0
scrotal oedema | 0
no gangrenous patches | 0
no skin breaks | 0
raised white cell count | 0
C-reactive protein of 269mg/L | 0
unremarkable urine dipstick | 0
blood cultures taken | 0
empirical antibiotics commenced | 0
intravenous Gentamicin | 0
Co-amoxiclav | 0
scrotal ultrasound scan | 0
scrotal cellulitis | 0
oedema | 0
lymphadenopathy | 0
CT thorax, abdomen and pelvis | 0
no intra-abdominal pathology | 0
echocardiogram | 0
bilateral lower limb doppler study | 0
no infective endocarditis | 0
no deep vein thrombosis | 0
Streptococcus Anginosus | 24
antibiotics rationalised | 24
Benzylpenicillin | 24
Clindamycin | 24
repeat ultrasound scan | 72
skin cellulitis | 72
abscess in the root of the penis | 72
reactive hydroceles | 72
MRI | 72
10×6cm abscess | 72
abscess abutting the ventral aspect of the root of the penis | 72
abscess extending to perineum and base of scrotum | 72
displacing but not invading the urethra | 72
incision and drainage of the abscess | 96
wound exploration and washout | 120
necrotic corpus cavernosum | 144
possible ischiorectal involvement | 144
flexible sigmoidoscopy | 144
normal recto-sigmoid colon | 144
suprapubic catheter | 144
comprehensive debridement | 144
further operative attempts at debridement | 192
wound washouts | 192
antibiotic therapy continued | 0
discharged | 1008
declined to attend follow up | 1008