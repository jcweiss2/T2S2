male | 0
40 + 2 weeks’ gestation | 0
primigravida mother | 0
25 years old | 0
uncomplicated pregnancy | -672
spontaneous onset of labor | -1
fetal distress | -1
ventouse-assisted delivery | 0
birth weight 3940 grams | 0
resuscitation with mask ventilation | 0
intubated | 0.13
transferred to NICU | 0.13
synchronized intermittent positive pressure ventilation | 0.13
gentamicin | 0.13
benzyl penicillin | 0.13
neutropenia | 18
left shift | 18
elevated C-reactive protein | 18
elevated procalcitonin | 18
lumbar puncture | 23
normal cell count | 23
negative for pathogens | 23
placental surface eSwab | 23
Gram-negative diplococci | 23
Neisseria meningitidis | 23
molecular testing | 23
blood cultures negative | 0.48
heel-prick blood | 5.5
N. meningitidis genogroup W DNA | 5.5
benzylpenicillin dosage decreased | 13.5
cefotaxime | 13.5
maternal bloods | -2.5
elevated leucocyte count | -2.5
neutrophil count | -2.5
mother remained well | 0
baby improved | 13.5
discharged home | 192
contact tracing | 192
chemoprophylaxis | 192
vaccination | 192
quadrivalent conjugate meningococcal vaccine | 192
counseling | 192 
funisitis | -1
chorioamnionitis | -1 
maternal and fetal inflammatory response | -1 
extubated | 13.5