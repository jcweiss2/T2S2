4 years old | 0
female | 0
admitted to the hospital | 0
fever | -96
generalized edema | -48
oliguria | -48
erythematous rash | -24
vomiting | -24
tachycardia | 0
hypotension | 0
poor peripheral perfusion | 0
macular erythematous rash | 0
cervical lymphadenopathy | 0
oral cheilosis | 0
tender hepatomegaly | 0
splenomegaly | 0
dengue considered | 0
leptospirosis considered | 0
sepsis considered | 0
Kawasaki's disease considered | 0
hemoglobin 8.7 gm% | 0
white cell count 10,000/cu.mm | 0
platelets 430,000 cells/cu.mm | 0
ESR 4 mm | 0
blood culture negative | 0
peripheral smear no malarial parasites | 0
liver function tests deranged | 0
SGPT 155 IU/L | 0
total proteins 4.8 g/dL | 0
albumin 2 g/dL | 0
dengue IgM negative | 0
leptospira IgM negative | 0
Cardioscope monitoring no arrhythmia | 0
serum creatinine normal | 0
CPK normal | 0
IV Ceftriaxone started | 0
normal saline bolus started | 0
Dopamine started | 0
fever persisted | 24
red lips developed | 24
strawberry tongue developed | 24
rash disappeared | 48
Dopamine stopped | 96
platelet count 477,000/cu.mm | 120
ESR 135 mm | 120
mild pericardial effusion | 120
dilated coronary arteries | 120
IVIG started | 120
edema subsided | 216
inotropic support omitted | 216
ESR decreased to 40 mm | 216
ESR decreased to 20 mm | 360
desquamation of the soles and palms | 504
Aspirin started | 504