49 years old| 0
male | 0
bronchiectasis | 0
fibrosis of the middle lobe | 0
dyspnea | 0
recurrent hemoptysis | 0
nonproductive cough |8
conservative management | 0
progressive decrease in physical endurance | 0
deterioration of the quality of life | 0
computerized tomography (CT) scan of the chest | 0
fibroatelectasis of the right middle lobe (RML) | 0
echocardiography | 0
large atrial septal defect (ASD) | 0
biventricular enlargement | 0
severe mitral regurgitation | 0
severe tricuspid regurgitation | 0
mitral prolapse | 0
moderate pulmonary artery hypertension | 0
multidisciplinary evaluation | 0
simultaneous procedure | 0
thoracoscopic uniportal cardiac intervention | 0
lobectomy | 0
femoral artery cannulation | 0
femoral vein cannulation | 0
cardiopulmonary bypass (CPB) | 0
transesophageal echocardiography | 0
cross-clamping of the aorta | 0
Chitwood clamp | 0
antegrade cardioplegia | 0
right atriotomy | 0
mitral valve ring annuloplasty | 0
De Vega annuloplasty of the tricuspid valve | 0
closure of the interatrial septal defect | 0
bovine pericardial patch | 0
heparin reversal | 0
isolation of the middle lobe vein | 0
transection of the middle lobe vein | 0
division of the middle lobe bronchus | 0
division of the middle lobe artery | 0
division of the parenchymal bridge | 0
endoscopic gastrointestinal anastomosis (endo GIA) stapler | 0
extubated | 72
transfer from the intensive care unit | 24
chest tube removal | 96
discharged | 192
improved exercise tolerance | 7392
resolution of hemoptysis | 7392
normalization of the cardiac chamber dimensions | 7392
absence of regurgitation | 7392
