75 years old | 0
male | 0
admitted to the hospital | 0
fever | -96
myalgia | -96
dyspnoea | -96
quit smoking | -131040
hypertension | 0
valsartan | 0
amlodipine | 0
travelled recently | -168
stayed in a motel | -168
temperature 38.7°C | 0
blood pressure 132/67 mmHg | 0
heart rate 102 beats per min | 0
respiratory rate 24 breaths per min | 0
severe hypoxaemia | 0
arterial oxygen tension 47.1 mmHg | 0
arterial carbon dioxide tension 40.9 mmHg | 0
pH 7.464 | 0
HCO3− 28.4 mmol·L−1 | 0
arterial oxygen saturation 84.2% | 0
anaemia | 0
haemoglobin 10.7 g·dL−1 | 0
elevated white blood cells | 0
elevated C-reactive protein | 0
hyponatraemia | 0
serum Na+ 127 mmol·L−1 | 0
infiltrates in both lungs | 0
antibiotic therapy with ampicillin/sulbactam | 0
antiviral therapy with oseltamivir | 0
Legionella urinary antigen test positive | 12
antibiotic therapy changed to moxifloxacin | 12
haemoptysis | 24
haemodynamic instability | 24
type I respiratory failure | 24
intubated | 24
transferred to the respiratory failure unit | 24
chest computed tomography | 24
extensive bilateral infiltrates | 24
blood in the bronchial secretions | 24
high oxygenation index | 24
increased need for haemodynamic support | 24
renal function deteriorated | 24
creatinine 4.75 mg·dL−1 | 24
haemoglobin 6.7 g·dL−1 | 24
many red blood cells in urine | 24
severe morphological deterioration | 24
bronchoscopy | 24
bloody secretions | 24
iron-laden macrophages | 24
microbiology results negative | 24
transfused with fresh frozen plasma and red blood cells | 24
samples for ANCA and anti-GBM antibodies | 24
positive C-ANCA | 24
negative anti-GBM | 24
methylprednisolone 1 g per 24 h i.v. | 24
cyclophosphamide 15 mg·kg−1 | 24
severe diffuse alveolar haemorrhage | 48
respiratory and haemodynamic instability | 48
unresponsive to mechanical ventilation | 48
plasma and blood transfusion | 48
vasopressor therapy | 48