55 years old | 0
male | 0
non-insulin dependent diabetes mellitus | 0
ingestion of methidathion | 0
semi-comatose | 0
myoclonus-like movements | 0
intubated | 0
mechanical ventilation | 0
intravenous infusion of atropine | 0
intravenous infusion of norepinephrine | 0
intravenous infusion of vasopressin | 0
intravenous infusion of dobutamine | 0
intravenous infusion of epinephrine | 0
intravenous infusion of PAM-A | 0
intravascular volume expansion | 0
gastric lavage | 0
midazolam | 0
remifentanyl | 0
vecuronium | 0
arterial blood gas analysis | 0
ethanol level in blood | 0
albumin | 0
glucose | 0
Hemoglobin A1c | 0
total CO2 content | 0
leukocyte count | 0
hemoglobin | 0
hematocrit | 0
platelets | 0
transferred to intensive care unit | 24
tests for hepatitis A, B, and C | 24
human immunodeficiency virus test | 24
free T4 level | 24
arterial blood gases | 24
blood cultures | 24
intravenous infusion of vecuronium discontinued | 48
intravenous infusion of epinephrine tapered off | 48
norepinephrine reduced | 48
vasopressin reduced | 48
dobutamine reduced | 48
metabolic acidosis resolved | 48
urine output decreased | 48
intravenous infusion of atropine discontinued | 96
glycopyrrolate given | 96
urine output decreased | 96
sputum culture | 96
piperacillin/tazobactam started | 96
doses of vasopressors and inotropic not reduced | 120
interleukin-6 | 120
procalcitonin | 120
intravenous infusion of remifentanil and midazolam maintained | 120
lactate level | 144
fibrinogen | 144
d-dimer | 144
ultrasonography | 144
transthoracic echocardiography | 144
total parenteral nutrition started | 144
enteral feeding not considered | 144
intravenous midazolam infusion discontinued | 216
vasopressors and inotropic reduced | 216
ulnar nerve stimulation test | 288
sputum culture | 288
vancomycin started | 288
arterial blood gas analysis | 408
leukocyte count | 408
platelet count | 408
ultrasonography of abdomen | 408
CT scan of abdomen | 408
exploratory laparotomy | 408
pulmonary artery catheter inserted | 408
laparotomy | 408
bowel resected | 408
peritoneum closed | 408
vasopressors and inotropic required | 408
urine output | 408
arterial blood gases | 408
lactate | 408
creatinine | 408
leukocyte count | 408
platelet count | 408
fibrinogen level | 408
glycopyrrolate given for the last time | 480
cultures from peritoneal drain and blood | 480
procalcitonin | 480
interleukin-6 | 480
C-reactive protein | 480
fibrinogen | 480
platelet count | 480
ulnar nerve stimulation test | 480
pathologic report | 480
voriconazole started | 480
culture of peritoneal drain fluid | 648
blood culture | 648
second laparotomy | 744
total colectomy | 744
septic shock | 744
vasopressors and inotropic required | 744
intravascular volume expansion | 744
thermodilution cardiac output | 744
metabolic acidosis | 744
lactate level | 744
galactomannan test | 744
cardiac arrest | 912
cardiopulmonary resuscitation | 912