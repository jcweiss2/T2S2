70 years old | 0
female | 0
admitted to intensive care unit | 0
altered sensorium | 0
hypotension | 0
fever | -48
diabetes mellitus type 2 | -672
essential hypertension | -672
chronic kidney disease | -672
hemodialysis | -672
hospitalized 1 month ago | -672
volume overload | -672
worsening renal parameters | -672
tender swellings over inner thighs | -672
tender swellings over buttocks | -672
punch biopsies advised | -672
punch biopsies declined | -672
awake | 0
confused | 0
disoriented to time | 0
disoriented to place | 0
disoriented to person | 0
no focal neurological deficit | 0
pulse rate 110/min | 0
blood pressure 70/50 mm Hg | 0
SPO2 98% | 0
afebrile | 0
bilateral basal crepitations | 0
violaceous nodules | 0
indurations | 0
extremely tender to palpation | 0
retiform purpura | 0
hemoglobin 6.6 g/dl | 0
total leucocyte count 25.0 thou/cumm | 0
neutrophilic leukocytosis | 0
erythrocyte sedimentation rate 119 mm/1st hour | 0
c-reactive protein 247 mg/L | 0
serum albumin 1.01 g/dl | 0
corrected serum calcium 11.08 mg/dl | 0
serum phosphate 4.95 mg/dl | 0
calcium phosphate product 54.8 | 0
creatine phosphokinase 57 U/L | 0
subcutaneous edema | 0
no deep vein thrombosis | 0
subcutaneous fat reticulation | 0
edema | 0
soft tissue changes related to lipodermatosclerosis | 0
metabolically inactive subcutaneous fat stranding | 0
panniculitis | 0
no evidence of metabolically active disease | 0
ANA profile negative | 0
p ANCA negative | 0
c ANCA negative | 0
APLA IgM negative | 0
IgG kappa monoclonal band | 0
plasma cell <10% | 0
monoclonal gammopathy of uncertain significance | 0
calciphylaxis | 0
empirical IV antibiotics (meropenem) | 0
empirical IV antibiotics (vancomycin) | 0
antifungal agent micafungin | 0
worsening sepsis | 0
persistent hypotension | 0
intravenous colistin | 0
blood cultures sterile | 0
urine cultures sterile | 0
calcitonin | 0
zoledronic acid | 0
alternate-day hemodialysis | 0
low calcium dialysate | 0
intravenous vitamin K | 0
no improvement in symptoms | 0
punch biopsies | 0
vasculopathic lymphoid infiltrate | 0
focal panniculitis | 0
no specific deposits on diffuse immunofluorescence | 0
intravascular lymphoma | 0
refractory septic shock | 0
intravenous hydrocortisone 50 mg 6-hourly | 0
no escalation of therapy | 0
deterioration of sensorium | 24
expired | 48
