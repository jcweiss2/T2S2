28 years old | 0
male | 0
admitted to the hospital | 0
abdominal pain | 0
persistent diarrhea | -48
dissection of the basilar artery | -216
dissection of the right common iliac artery | -240
retroperitoneal hematoma | -240
dissection and embolism of the renal artery | -144
definitively diagnosed as having vEDS | -216
genetic testing | -216
missense variants in COL3A1 | -216
panperitonitis | 0
rebound tenderness | 0
muscular defensiveness | 0
blood pressure 152/92 mmHg | 0
pulse rate 110 bpm | 0
peripheral arterial oxygen saturation 92% | 0
body temperature 37.8°C | 0
WBC 3100/μL | 0
TP 6.1 g/dL | 0
CK 903 U/L | 0
RBC 448×10^4/μL | 0
Alb 4.0 g/dL | 0
CRP 0.44 mg/dL | 0
Hb 13.3 g/dL | 0
BUN 11.2 mg/dL | 0
Glucose 111 mg/dL | 0
Ht 38.3% | 0
Cre 0.62 mg/dL | 0
HbA1c 6.4% | 0
Plt 19.1×10^4/μL | 0
Na 139 mmol/L | 0
K 4.2 mmol/L | 0
PT-INR 1.01 | 0
APTT 30.9 sec | 0
T-Bil 0.89 mg/dL | 0
D-dimer 1.2 ug/mL | 0
AST 39 U/L | 0
ALT 56 U/L | 0
LDH 224 U/L | 0
non-localized intraabdominal free air | 0
enlargement of a right common iliac arterial aneurysm | 0
intestinal perforation | 0
laparotomy | 0
perforation of the sigmoid colon | 0
intestinal tract wall fragile | 0
mesentery fragile | 0
mesenteric vessels fragile | 0
resection of the sigmoid colon | 0
end-colostomy | 0
pathological findings | 0
thinning of muscular layer | 0
tear of the muscular layer | 0
infiltration of inflammatory cells | 0
septic shock | 0
ventilator management | 0
analgesic agents | 0
fentanyl | 0
acetaminophen | 0
discharged | 696
follow-up with CT imaging | 696
no events after 18 months | 1092