50 years old | 0
    female | 0
    severe lower abdominal pain | -120
    lower abdominal pain irradiating to the lumbar region | -120
    nausea | -120
    vomiting | -120
    fever | -120
    constipation | -120
    generalized abdominal pain | -1344
    diarrhea | -1344
    hypertension | -1344
    dyslipidemia | -1344
    heart failure | -1344
    rheumatologic disease | -1344
    furosemide | -1344
    captopril | -1344
    spironolactone | -1344
    prednisone | -1344
    sodium diclofenac | -1344
    ill-looking cushingoid | 0
    pale | 0
    cyanotic extremities | 0
    decreased tissue perfusion | 0
    marked lower limbs edema | 0
    slightly disoriented | 0
    blood pressure 50/30 mmHg | 0
    pulse 110 beats/minute | 0
    respiratory rate 24 respiratory movements/minute | 0
    axillary temperature 37 °C | 0
    distended abdomen | 0
    diffusely tender abdomen | 0
    decreased bowel sounds | 0
    negative rebound tenderness test | 0
    liver palpable up to 1 cm below the right costal margin | 0
    unremarkable heart examination | 0
    unremarkable lungs examination | 0
    extracellular volume repletion with saline | 0
    ceftriaxone | 0
    metronidazole | 0
    hydrocortisone | 0
    noradrenaline | 0
    referred to ICU | 0
    hemoglobin 12.6 g/dL | 0
    creatinine 2.9 mg/dL | 0
    hematocrit 37.4% | 0
    potassium 4.7 mEq/L | 0
    leucocytes 19100 103/mm3 | 0
    sodium 110 mEq/L | 0
    bands 17% | 0
    ALT 28 U/L | 0
    segmented 72% | 0
    AST 44 U/L | 0
    eosinophils 1% | 0
    LDH 336 U/L | 0
    basophils 0% | 0
    CK 933 U/L | 0
    lymphocytes 8% | 0
    amylase 11 U/L | 0
    monocytes 2% | 0
    lipase 15 U/L | 0
    platelets 382.103/mm3 | 0
    total protein 4.9 g/dL | 0
    CRP 142 mg/L | 0
    albumin 2.3 g/dL | 0
    BUN 62 mg/dL | 0
    PT (INR) 1.21 | 0
    minimal free fluid in abdominal cavity | 0
    diffuse decrease of small bowel peristaltic movements | 0
    liquid distention | 0
    negative anti-HIV serology | 0
    hemodynamically unstable | 0
    continuous administration of norepinephrine | 0
    continuous administration of vasopressin | 0
    no initial clinical improvement | 0
    petechiae | 72
    ecchymoses | 72
    abdomen lesions | 72
    upper limbs lesions | 72
    worsened mental status | 96
    orotracheal intubation | 96
    mechanical ventilation | 96
    multi sensitive E. coli in blood culture | 96
    no clinical improvement | 96
    death | 96
    multiple petechial skin lesions | 96
    generalized edema of limbs | 96
    mild ascites | 96
    S. stercoralis larvae in dermis | 96
    foci of hemorrhage in skin | 96
    no inflammatory cells in skin | 96
    boggy and heavy lungs | 96
    diffuse alveolar damage | 96
    areas of alveolar hemorrhage | 96
    hemosiderin-laden macrophages | 96
    S. stercoralis larvae in lungs | 96
    giant cell granulomatous reaction | 96
    flat lesions in small bowel | 96
    petechial foci of hemorrhage in small bowel mucosa | 96
    hemorrhage on abdominal serous surfaces | 96
    S. stercoralis larvae in duodenal mucosa | 96
    S. stercoralis larvae in omentum | 96
    acute hematogenous pyelonephritis | 96
    subcapsular abscesses in left kidney | 96
    acute inflammation in spleen | 96
    septic emboli in spleen | 96
    acute infarction in spleen | 96
    adrenal gland lipid depletion | 96
    adrenal gland hemorrhagic foci | 96
    liver necrosis on zone 3 | 96
    acute tubular necrosis | 96
    ischemic pancreatitis | 96
    diffuse dilatation of heart chambers | 96
    myocardial softening | 96
    focal hyaline thrombi in lungs | 96
    focal hyaline thrombi in glomeruli | 96
    S. stercoralis hyperinfection syndrome | 96
    Gram-negative bacterial septicemia | 96
    septic shock | 96
    
