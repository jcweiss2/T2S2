69 years old | 0 | 0 
female | 0 | 0 
admitted to the hospital | 0 | 0 
stabbed herself in the abdomen | -1 | -1 
self-inflicted stab wound | -1 | -1 
kitchen knife | -1 | -1 
suicidal intent | -1 | -1 
blood pressure could not be measured | 0 | 0 
pulseless electrical activity | 0 | 0 
body temperature was 35.0 °C | 0 | 0 
oxygen saturation was 99 % | 0 | 0 
Glasgow Coma Scale score of 3 | 0 | 0 
agonal respiration | 0 | 0 
wound measuring 5 cm | 0 | 0 
intra-abdominal fluid collection | 0 | 0 
emergency thoracotomy | 0 | 1 
aortic cross-clamping | 0 | 15 
open cardiac massage | 0 | 15 
epinephrine administration | 0 | 15 
temporary return of spontaneous circulation | 15 | 15 
hemodynamically unstable | 15 | 15 
laparotomy | 15 | 30 
injuries to the common hepatic and splenic arteries | 15 | 30 
injuries to the pancreas | 15 | 30 
injuries to the spleen | 15 | 30 
injuries to the liver | 15 | 30 
ligation of the injured arteries | 15 | 30 
distal pancreatectomy | 30 | 45 
splenectomy | 30 | 45 
liver sutured | 30 | 45 
norepinephrine administration | 30 | 48 
second-look surgery | 24 | 24 
no signs of active bleeding | 24 | 24 
no ischemic change | 24 | 24 
abdominal wall closure | 72 | 72 
regular examinations | 72 | 168 
enhanced computed tomography scan | 96 | 96 
disruption of the celiac artery | 96 | 96 
gastroduodenal artery arising from the superior mesenteric artery | 96 | 96 
gastroscopy | 216 | 216 
patchy mucosal necrosis | 216 | 216 
conservative treatment | 216 | 336 
fever | 552 | 552 
pain in the stomach | 552 | 552 
white blood cell count of 34,000/mm3 | 552 | 552 
C reactive protein of 13.4 mg/dL | 552 | 552 
CT scan | 552 | 552 
air in the gastric wall | 552 | 552 
intra-abdominal free air | 552 | 552 
gastric necrosis | 552 | 552 
emergency surgery | 552 | 576 
total gastrectomy | 552 | 576 
Roux-en-Y reconstruction | 552 | 576 
histological findings of the stomach | 576 | 576 
diffuse necrotic changes | 576 | 576 
inflammatory cell infiltrations | 576 | 576 
no evidence of invasive fungal infection | 576 | 576 
leakage on the duodenal stump | 696 | 696 
continuous tube drainage | 696 | 696 
sepsis | 1680 | 1680 
multidrug-resistant Pseudomonas aeruginosa infection | 1680 | 1680 
disseminated intravascular coagulation | 1680 | 1680 
death | 1680 | 1680