18 years old | 0
male | 0
pregnant | 0
primigravida | 0
34-week pregnancy | 0
spontaneous pregnancy | 0
admitted to hospital | 0
recurrent vomiting | -24
epigastric pain | -24
diagnosed with uterine fibroid | -24
history of weight loss | -24
no change in bowel habits | -24
no hematemesis or rectal bleeding | -24
no history of hematuria or passing stones | -24
using iron tablets | -24
ill | -24
markedly dehydrated | -24
drowsy | -24
blood pressure 126/76 mmHg | -24
pulse rate 94 min–1 | -24
respiratory rate 30 min–1 | -24
temperature 36.6°C | -24
no lymphadenopathy | -24
no thyromegaly | -24
no edema | -24
uterus size of 40 weeks | -24
tender epigastric area | -24
drowsy and hypotonic | -24
brisk deep tendon reflexes | -24
no obvious focal neurological sign | -24
down-going planter reflexes | -24
chest and cardiovascular systems unremarkable | -24
hemoglobin (Hb) 8.7 g/dl | -24
WBCs 7000 μl–1 | -24
platelets 445 000 μl–1 | -24
ESR 109 mm/h | -24
toxic granulation of WBCs | -24
BUN 4.4 mmol/l | -24
creatinine 59 μmol/l | -24
HCO3 22 mmol/l | -24
Na 138 mmol/l | -24
Ca 4.8 mmol/l | -24
uric acid 508 μmol/l | -24
lactic acid 1.2 mmol/l | -24
phosphorous 0.8 mmol/l | -24
HIV serology negative | -24
calcium at 14 weeks’ gestation 2.43 mmol/l | -672
ALT 4 u/l | -24
AST 11 u/l | -24
ALP 150 u/l | -24
total protein 72 g/l | -24
albumen 30 g/l | -24
cholesterol 4.05 mmol/l | -24
triglyceride 3.59 mmol/l | -24
PTH 3 pg/ml | -24
TSH 0.68 mIU/l | -24
free thyroxin 16.6 pmol/l | -24
cortisol 1849 nmol/l | -24
vitamin D 15 ng/ml | -24
serum protein electrophoresis normal | -24
serum level of angiotensin-converting enzyme normal | -24
normal saline infusion | 0
calcitonin | 0
hemodialysis | 0
rupture membrane | 12
urgent cesarean section | 12
bleeding | 12
hypotension | 12
blood transfusion | 12
delivery of a baby girl | 12
removal of uterine masses | 12
histopathological examination | 12
leiomyoma with calcifications | 12
septicemia | 12
septic shock | 12
vasopressors | 12
broad-spectrum antibiotics | 12
serum calcium 2.34 mmol/l | 24
phosphorus 1.1 mmol/l | 24
BUN 6.2 mmol/l | 24
Cr 75 mmol/l | 24
Na 143 mmol/l | 24
K 4.2 mmol/l | 24
HCO3 16 mEq/l | 24
chloride 113 mEq/l | 24
albumin 21 g/l | 24
serum lactate 5.19 | 24
serum PTH 155 pg/ml | 24
serum amylase 88 u/l | 24
serum lipase 73 u/l | 24
Hb 5.8 g/dl | 24
platelets 125 000 μl1 | 24
CT scan of the chest and pelvis | 24
MRI of the brain | 24
vasospasm of the internal carotid, the middle and the anterior carotid arteries | 24
diffuse ischemic changes | 24
generalized muscle weakness and stiffness | 24
discharged home | 168
final diagnosis of humoral hypercalcemia associated with a uterine fibroid | 168
serum calcium remained within the normal range | 504