15 years old | 0
male | 0
admitted to the hospital | 0
short stature | 0
hydrocephalus | 0
blurring of vision | -360
drowsy | 0
Glasgow coma scale 12/15 | 0
tubercular meningitis | -720
hypertelorism | 0
downslanting prominent eyes | 0
thick lips | 0
high palatal arch | 0
Mallampati score 3 | 0
limited neck extension | 0
mouth opening 4 cm | 0
scoliosis of dorsal spine | 0
reduced volume of thorax | 0
systolic murmur at left sternal edge | 0
sinus tachycardia | 0
systemic hypertension | 0
high BP detected | -720
no antihypertensives | -720
mild motor delay | -13140
growth retardation | -13140
physical deformities | -13140
no symptoms of cardiac or respiratory decompensation | 0
haemoglobin level 12.8 g/dl | 0
normal serum electrolytes | 0
normal glucose | 0
normal liver function tests | 0
normal renal function tests | 0
normal coagulation profile | 0
normal platelet counts | 0
chest X-ray | 0
X-ray neck anterior-posterior and lateral view | 0
non-contrast computed tomography head | 0
magnetic resonance imaging of the brain | 0
basilar invagination | 0
atlantoaxial dislocation | 0
sinus tachycardia | 0
left ventricular hypertrophy | 0
Q-waves in lead II, III, aVF, V5 and V6 | 0
hypertrophic cardiomyopathy | 0
no left ventricular outflow tract obstruction | 0
no systolic anterior motion of the mitral valve | 0
standard monitors attached | 0
HR 130 beats per min | 0
BP 180/100 mm Hg | 0
SPO2 100% | 0
antibiotic prophylaxis | 0
cefuroxime 50 mg/kg | 0
resuscitation and difficult airway cart ready | 0
premedicated with midazolam | 0
right radial artery cannulated | 0
esmolol administered | 0
induction of anaesthesia | 0
preoxygenation for 5 min | 0
morphine administered | 0
thiopentone administered | 0
bag mask ventilation | 0
check laryngoscopy | 0
Cormack Lehane Grade 2b | 0
vecuronium bromide administered | 0
fentanyl administered | 0
lignocaine administered | 0
trachea intubated | 0
left internal jugular vein cannulated | 0
anaesthesia maintained | 0
O2/N2O and sevoflurane | 0
small tidal volumes | 0
high respiratory rates | 0
end tidal CO2 concentration monitored | 0
estimated blood loss 50 ml | 120
duration of surgery 120 min | 120
intraoperative blood gas analysis | 120
pH 7.5 | 120
PaO2 97 mm Hg | 120
PaCO2 29 mm Hg | 120
HCO3 22 mmol/L | 120
urine output monitored | 0
temperature monitored | 0
reversal of residual paralysis | 120
glycopyrrolate administered | 120
neostigmine administered | 120
trachea extubated | 120
GCS 12 | 120
transferred to ICU | 120
shunt obstruction | 24
GCS deteriorated | 24
re-intubated | 24
septic shock | 360
multi organ dysfunction syndrome | 360
died | 360