69 years old | 0
male | 0
admitted to the hospital | 0
paraumbilical hernia | -672
abdominal distension | -672
diarrhoea | -672
weight loss | -672
lung fibrosis | 0
obstructive airway disease | 0
atrial fibrillation | 0
cardiomyopathy | 0
heart failure | 0
biventricular pacemaker | 0
systemic sclerosis | 0
steroids | 0
methotrexate | 0
CT scan | 0
free fluid | 0
air in the abdomen | 0
perforation | 0
ischaemic bowel necrosis | 0
emergency laparotomy | 24
small bowel ischaemia | 24
pockets of subserosal gas | 24
PI | 24
probable self-sealed perforations | 24
abdominal cavity irrigated | 24
drained | 24
hernia repaired | 24
intensive care | 24
nutritional support | 48
ileus | 48
discharged | 168
oral antibiotics | 168
outpatient review | 168
Rheumatology team | 168
severe epigastric pain | 744
metabolic acidosis | 744
tachycardic | 744
tachypneic | 744
normotensive | 744
white cell count | 744
haemoglobin | 744
creatinine | 744
INR | 744
urgent CT | 744
conservative approach | 744
p-possum score | 744
morbidity | 744
mortality | 744
deteriorated | 768
acidotic | 768
lactate | 768
re-operate | 768
died | 768
post mortem | 768
small bowel perforation | 768
PI | 768