64 years old | 0  
    male | 0  
    end-stage liver disease | 0  
    secondary biliary cirrhosis | 0  
    non-alcoholic steatohepatitis | 0  
    robotic cholecystectomy | -6720  
    hepatic duct leak | -6720  
    open choledochojejunostomy | -6720  
    elevated liver function tests | -6720  
    magnetic resonance cholangiopancreatography | -6720  
    choledochojejunostomy stricture | -6720  
    intrahepatic biliary tree dilation | -6720  
    liver biopsy | -6720  
    cirrhosis | -6720  
    chronic biliary obstruction | -6720  
    non-alcoholic steatohepatitis | -6720  
    liver transplantation | 0  
    extensive adhesions | 0  
    extended two-hepatic vein piggy-back technique | 0  
    portal vein anastomosis | 0  
    common hepatic artery anastomosis | 0  
    reconstruction of accessory right hepatic artery | 0  
    biliary reconstruction | 0  
    steroid taper | 0  
    Myfortic | 0  
    Tacrolimus | 0  
    Micafungin | 0  
    Valcyte | 0  
    Bactrim | 0  
    thrombus of the accessory right hepatic artery | 24  
    computed tomography angiography | 24  
    common hepatic artery patent | 24  
    therapeutic low molecular weight heparin | 24  
    perihepatic hematoma | 24  
    percutaneous drain | 24  
    drain fluid cultures negative | 24  
    nonbilious drain output | 24  
    therapeutic anticoagulation | 24  
    transition to Apixaban | 192  
    discharge | 192  
    perihepatic drain removed | 240  
    sudden onset severe right upper quadrant abdominal pain | 528  
    lightheadedness | 528  
    hemodynamically unstable | 528  
    tachycardic | 528  
    hypotensive | 528  
    abdominal distension | 528  
    massive transfusion protocol | 528  
    resuscitation initiated | 528  
    sepsis protocol | 528  
    severe lactic acidosis | 528  
    bicarbonate 8 mmol/L | 528  
    lactate 9.8 mmol/L | 528  
    acute blood loss anemia | 528  
    hemoglobin 6.5 g/dl | 528  
    acute kidney injury | 528  
    creatinine 3.1 mg/dl | 528  
    worsening liver function tests | 528  
    blood product resuscitation | 528  
    computed tomography | 528  
    main hepatic artery pseudoaneurysm | 528  
    active extravasation | 528  
    hemoperitoneum | 528  
    endovascular therapy | 528  
    acute decompensation | 528  
    mean arterial pressure 30-40 mmHg | 528  
    pulseless electrical activity | 528  
    advanced cardiac life support | 528  
    intubation | 528  
    right femoral arterial line | 528  
    REBOA sheath | 528  
    REBOA inflated | 528  
    spontaneous cardiac activity recovery | 528  
    emergency transport to operating room | 528  
    rapid laparotomy | 528  
    fresh blood clot | 528  
    hematoma | 528  
    no biloma | 528  
    no bile leak | 528  
    no enteric leak | 528  
    no abscess formation | 528  
    hepatic allograft ischemic | 528  
    REBOA occlusion | 528  
    identification and control of recipient hepatic artery | 528  
    REBOA deflation | 528  
    reperfusion injury | 528  
    recurrent pulseless electrical activity | 528  
    REBOA re-inflation | 528  
    ACLS resumed | 528  
    pulse resumption | 528  
    additional aortic occlusion | 528  
    donor proper hepatic artery thrombosed | 528  
    donor proper hepatic artery damaged | 528  
    donor hepatic artery ruptured | 528  
    mycotic change | 528  
    recipient hepatic artery ligation | 528  
    open abdomen negative pressure therapy | 528  
    transfer to surgical intensive care unit | 528  
    continuous renal replacement therapy | 528  
    goal-directed resuscitation | 528  
    refractory septic shock | 528  
    severe acidosis | 528  
    electrolyte abnormalities | 528  
    coagulopathy | 528  
    hepatic ischemic insult | 528  
    hemorrhagic insult | 528  
    stabilization for re-transplant | 528  
    condition decline | 528  
    multiorgan failure | 528  
    allograft non-function | 528  
    bradycardic | 542  
    pulseless | 542  
    resuscitation discontinued | 542  
    deceased | 542  
    Streptococcus Constellatus bacteremia | 528  
    Klebsiella Pneumoniae colonization | 528  
    postmortem microbiology results | 542  

