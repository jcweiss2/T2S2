55 years old | 0
male | 0
morbidly obese | 0
diabetes mellitus | 0
end-stage renal disease | 0
hemodialysis | 0
peripheral vascular disease | 0
left below knee amputation | 0
right above knee amputation | 0
right extra anatomical axillobifemoral bypass graft | 0
admitted to emergency department | 0
right-sided abdominal pain | -48
vomiting | -48
fever | -48
conscious | 0
alert | 0
oriented | 0
pale | 0
sick | 0
temperature 37.8°C | 0
blood pressure 150/90 mmHg | 0
oxygen saturation 95% | 0
abdomen distended | 0
tympanic | 0
right upper quadrant tenderness | 0
right flank tenderness | 0
total leukocyte count 20 × 10^3 | 0
hemoglobin 10.7 gm% | 0
acidotic pH 7.33 | 0
end-stage renal disease | 0
chest X-ray | 0
air under the right hemi-diaphragm | 0
evaluated by general surgeon | 0
impression of perforated viscous | 0
computed tomography scan | 0
right perinephric collection | 0
extension into the right sub-phrenic region | 0
gas in the right collecting system | 0
gas in the urinary bladder | 0
no gas in the renal parenchyma | 0
right atrial thrombus | 0
started on parenteral antibiotics | 0
admitted to intensive care unit | 0
trial of percutaneous drainage | 12
percutaneous drainage failed | 12
evaluated by anesthetist | 12
not fit for general anesthesia | 12
open drainage | 24
epidural anesthesia | 24
sedation | 24
loculated perinephric and sub-phrenic collection | 24
cystoscopy | 24
abnormal bladder mucosa | 24
multiple cystic lesions | 24
air “bubbles” in bladder | 24
ureteric Double J stent | 24
urethral catheter | 24
reasonably well during procedure | 24
condition deteriorated | 48
culture of collection | 48
Klebsiella pneumonia extended-spectrum β-lactamase | 48
severe sepsis | 72
multiple organ failure | 72
died | 72