55 years old | 0
male | 0
no significant past medical history | 0
dyspnea | -744
dry cough | -744
joint pain | -744
diffuse joint pain | -744
bilateral distribution | -744
fingers | -744
hands | -744
wrists | -744
elbows | -744
shoulders | -744
hips | -744
knees | -744
ankles | -744
shoveling snow | -744
persistent symptoms | -336
ibuprofen | -336
oxycodone-acetaminophen | -336
methylprednisolone | -336
worsened joint pain | -336
dyspnea with dry cough | -336
multiple home tests for SARS-CoV-2 | -336
negative SARS-CoV-2 tests | -336
shortness of breath with exertion | 0
joint pain | 0
dry cough | 0
unintentional weight loss | 0
15 lb weight loss | 0
no fever | 0
no headache | 0
no sore throat | 0
no chest pain | 0
no hemoptysis | 0
no gastrointestinal symptoms | 0
no calf swelling | 0
no calf pain | 0
former smoker | 0
20-year pack history | 0
quit smoking 10 years prior | 0
no recent travel | 0
no sick contacts | 0
no occupational or environmental toxic fume exposure | 0
Moderna SARS-CoV-2 vaccine | -744
third dose | -744
blood pressure 98/63 mm Hg | 0
heart rate 93 beats/min | 0
respirations 18/min | 0
temperature 36.8 °C | 0
oxygen saturation 93% | 0
oxygen saturation 98% | 0
bibasilar rales | 0
tenderness | 0
swelling | 0
erythematous papules | 0
erythematous macules | 0
no muscle tenderness | 0
D-dimer 1,702 | 0
aspartate aminotransferase 86 | 0
alanine aminotransferase 65 | 0
C-reactive protein 3.70 | 0
erythrocyte sedimentation rate 52 | 0
admitted to hospital | 0
rheumatology consult | 0
pulmonology consult | 0
complete infectious workup | 0
complete rheumatologic workup | 0
azithromycin | 0
ceftriaxone | 0
fluticasone-vilanterol | 0
tiotropium bromide | 0
prednisone | 0
discharged | 72
oral cefuroxime | 72
follow-up appointment with rheumatology | 168
diagnosed with CADM | 168
elevated anti-MDA5 antibody | 168
mycophenolate mofetil | 168
prednisone | 168
follow-up appointment with pulmonology | 168
6-min walk test | 168
pulmonary function testing | 168
diagnosed with asthma | 168
mild ILD | 168
fluticasone-salmeterol | 168
tiotropium bromide | 168
new cough | 504
foamy sputum production | 504
outpatient bronchoscopy | 504
bronchoalveolar lavage | 504
transbronchial biopsy | 504
fever | 504
readmitted | 504
vancomycin | 504
piperacillin-tazobactam | 504
sulfamethoxazole/trimethoprim | 504
methylprednisone | 504
high resolution CT scan | 504
traction bronchiectasis | 504
interval worsening of bilateral mixed interstitial alveolar infiltrates | 504
ground glass opacities | 504
septal thickening | 504
clinical status deterioration | 510
increasing supplemental oxygen requirements | 510
persistent hypoxia | 510
transbronchial biopsy results | 510
normal lung tissue | 510
BAL results | 510
Pneumocystis jirovecii | 510
Pneumocystis pneumonia | 510
immunosuppressive therapy | 510
trimethoprim-sulfamethoxazole | 510
plasma exchange therapy | 510
intubated | 516
pneumothorax | 516
pneumomediastinum | 516
cardiothoracic surgery consult | 516
no chest tube placement | 516
full ventilator support | 516
norepinephrine | 516
pulseless electrical activity arrest | 522
death | 522