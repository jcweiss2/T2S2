85 years old | 0 | 0 
male | 0 | 0 
admitted to the hospital | 0 | 0 
farmer | 0 | 0 
active lifestyle | 0 | 0 
atrial fibrillation | -720 | 0 
benign prostatic hypertrophy | -720 | 0 
trismus | -144 | -144 
hypertonia | -144 | -144 
C. tetani infection | -144 | 0 
injured his leg | -144 | -144 
immunoglobulins | -144 | -120 
tetanus vaccination | -144 | -120 
metronidazole | -144 | -134 
transferred to ICU | -120 | -120 
tracheostomy | -120 | -120 
mechanical ventilation | -120 | -120 
vasoactive support | -120 | -120 
respiratory failure | -120 | -120 
seizures | -120 | -120 
baclofen | -120 | -120 
midazolam | -120 | -120 
diazepam | -120 | -120 
electroencephalography | -120 | -120 
severely slow cerebral activity | -120 | -120 
opacity on chest radiography | -120 | -120 
peripheral leukocytosis | -120 | -120 
ventilator-associated pneumonia | -120 | -120 
blood cultures | -120 | -120 
tracheal secretion samples | -120 | -120 
Klebsiella pneumoniae | -120 | -120 
methicillin-sensitive Staphylococcus aureus | -120 | -120 
piperacillin-tazobactam | -120 | -110 
transferred to geriatric unit | -110 | -110 
coma | -110 | -90 
breathed spontaneously | -90 | -90 
supplemental oxygen | -90 | 0 
linezolid | -90 | -76 
VAP exacerbation | -90 | -90 
meropenem | -76 | -59 
septic shock | -76 | -76 
awoke | -59 | -59 
feeding tube removed | -59 | -59 
cholestasis | -59 | -59 
acute edematous pancreatitis | -59 | -59 
endoscopic treatment postponed | -59 | -59 
urinary tract infection | -59 | -52 
multidrug-resistant organisms | -59 | -52 
K. pneumoniae | -59 | -52 
Acinetobacter baumannii | -59 | -52 
Enterococcus faecalis | -59 | -52 
colistin | -59 | -52 
amoxicillin-clavulanate | -59 | -52 
clinical condition improved | -52 | -52 
transferred to rehabilitation unit | -52 | -52 
MDRO isolation | -52 | 0 
tracheal supplemental oxygen | -52 | 0 
bladder catheter | -52 | 0 
pressure ulcers | -52 | 0 
sarcopenic | -52 | 0 
low handgrip strength | -52 | 0 
appendicular skeletal mass | -52 | 0 
rehabilitation | -52 | 0 
Clostridioides difficile infection | -24 | -14 
oral vancomycin | -24 | -14 
atrial fibrillation | -14 | -14 
third-degree atrioventricular block | -14 | -14 
heart rate 30 beats/min | -14 | -14 
transferred to cardiac ICU | -14 | -14 
single-chamber pacemaker implantation | -14 | -14 
hyperkinetic delirium | -14 | -14 
Pseudomonas aeruginosa bloodstream infection | -10 | -3 
ceftazidime-avibactam | -10 | -3 
amikacin | -10 | -3 
SARS-CoV-2 | -7 | -7 
remdesivir | -7 | -4 
droplet isolation | -7 | 0 
second recurrence of C. difficile | -4 | -4 
fidaxomicin | -4 | 6 
bloodstream infection | 6 | 6 
Candida parapsilosis | 6 | 6 
MSSA | 6 | 6 
Candida tropicalis | 6 | 6 
caspofungin | 6 | 23 
cefazolin | 6 | 23 
intravenous catheter replaced | 6 | 6 
P. aeruginosa | 23 | 23 
piperacillin-tazobactam | 23 | 30 
aztreonam | 30 | 30 
ceftazidime-avibactam | 30 | 30 
cefepime | 30 | 40 
tracheostomy closure | 40 | 40 
nutritional supplementation | -52 | 0 
malnutrition | -52 | 0 
sarcopenia | -52 | 0 
postural transition | 0 | 0 
aided transfers | 0 | 0 
axial stability | 0 | 0 
balance improvement | 0 | 0 
breath-movement coordination | 0 | 0 
thoracic expansion | 0 | 0 
girdle opening | 0 | 0 
inhalation-exhalation | 0 | 0 
wheelchairs | 0 | 0 
walkers | 0 | 0 
rehabilitation follow-up | 0 | 0 
ENT follow-up | 0 | 0 
geriatric follow-up | 0 | 0 
discharged | 0 | 0