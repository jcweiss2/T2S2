45 years old | 0
right-handed | 0
man | 0
HIV | -672
CD4+ T-cell count 556 | -672
not on anti-retroviral medications | -672
presented to hospital | -24
acute onset of horizontal diplopia | -24
weakness of left face | -24
weakness of right arm | -24
weakness of right leg | -24
hemiparesis alternans | -24
history unremarkable | 0
vital signs unremarkable | 0
physical exam unremarkable | 0
routine laboratory tests normal | 0
initial MRI | 0
FLAIR signal hyperintensity left pons | 0
DWI restriction left pons | 0
acute ischemic stroke | 0
Millard-Gubler syndrome | 0
extra-axial curvilinear FLAIR hyperintensity | 0
T1 high signal | 0
DWI high signal subarachnoid space | 0
ADC low signal subarachnoid space | 0
unclear etiology extra-axial entity | 0
MRA unremarkable | 0
admitted to neuroscience ICU | 0
cardiac telemetry sinus tachycardia | 0
transthoracic echocardiography normal | 0
transesophageal echocardiography normal | 0
normal ejection fraction | 0
normal valves | 0
normal chambers | 0
no clot | 0
no vegetation | 0
no patent foramen ovale | 0
no septal defect | 0
young age (>55) | 0
lack of traditional stroke risk factors | 0
hypercoagulable serum panel ordered | 0
anticardiolipin antibodies negative | 0
lupus anticoagulant negative | 0
protein C normal | 0
protein S normal | 0
anti-thrombin III normal | 0
fibrinogen normal | 0
factor VIII normal | 0
prothrombin 20210 normal | 0
homocystine normal | 0
lipoprotein (a) normal | 0
sickle cell screen negative | 0
developed severe headache | 24
headache progression over few days | 24
meningismus | 24
stupor | 24
lumbar puncture | 24
opening pressure 230 mm H2O | 24
250 red blood cells CSF | 24
75 white blood cells CSF | 24
neutrophils 79% CSF | 24
glucose 80 CSF | 24
protein 54 CSF | 24
ruled out Cryptococcus | 24
ruled out tuberculosis | 24
ruled out syphilis | 24
low suspicion due to CD4 556 | 24
acid-fast bacilli test negative | 24
PPD negative | 24
chest X-rays no lesions | 24
RPR non-reactive | 24
VDRL non-reactive | 24
FTA-ABS non-reactive | 24
HSV PCR negative | 24
CMV PCR negative | 24
VZV PCR negative | 24
no dermatomal vesicles | 24
seeping pustular furuncles knees | 24
cultured MRSA | 24
blood cultures positive MRSA | 24
intravenous vancomycin started | 24
second MRI | 72
intra-axial FLAIR hyperintensities bilateral pons | 72
DWI restriction bilateral pons | 72
intra-axial FLAIR hyperintensities left cerebellum | 72
DWI restriction left cerebellum | 72
new cerebral infarctions | 72
exacerbating cerebral infarctions | 72
subarachnoid DWI restriction increased | 72
subarachnoid DWI restriction expanded | 72
communicating hydrocephalus | 72
effacement fourth ventricle | 72
dilation lateral ventricles | 72
dilation third ventricle | 72
CSF trans-exudation | 72
another lumbar puncture | 72
4 red blood cells CSF | 72
112 white blood cells CSF | 72
neutrophils 74% CSF | 72
glucose 130 CSF | 72
protein 2126 CSF | 72
high-dose antibiotics | 72
vancomycin | 72
ceftriaxone | 72
ampicillin | 72
aggressive intravenous fluids | 72
pressor agents | 72
ventriculostomy | 72
supportive care | 72
continued deterioration | 72
comatose | 72
third MRI | 96
diffusion restriction spread | 96
FLAIR hyperintensity spread | 96
brainstem parenchyma involvement | 96
pons involvement | 96
medulla involvement | 96
left cerebellum involvement | 96
MRA irregularity vertebro-basilar circulation | 96
MRA narrowing vertebro-basilar circulation | 96
lack of flow-related enhancement left vertebral artery | 96
lack of flow-related enhancement posterior cerebral arteries | 96
expired | 96
autopsy | 96
brain weight 1212 g | 96
basilar artery patent | 96
posterior cerebral arteries patent | 96
cerebellar arteries patent | 96
arteritis | 96
lymphoplasmocytic infiltration | 96
partial large-vessel occlusion | 96
partial small-vessel occlusion | 96
fibrointimal proliferation | 96
basilar meninges thickened | 96
white purulent material | 96
inferior brainstem infarcts | 96
left cerebellum infarcts | 96
inflammation cervical spinal cord leptomeninges | 96
vasculitis cervical spinal cord leptomeninges | 96
dilatation lateral ventricles | 96
dilatation third ventricle | 96
aqueduct dilatation | 96
compression fourth ventricle | 96
Gram stain GPC chains | 96
GMS stain GPC chains | 96
MRSA in blood | 96
MRSA in furuncles | 96
GPC in brain insufficient DNA | 96
broad-spectrum antibiotic use | 96
paraffin block PCR beta-globin genes | 96
