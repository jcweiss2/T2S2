69 years old | 0 | 0 
female | 0 | 0 
admitted to the hospital | 0 | 0 
high-grade fever | -72 | 0 
pleuritic right lower chest pain | -72 | 0 
cough | -72 | 0 
elevated temperature | 0 | 0 
bibasilar crackles | 0 | 0 
lower extremity edema | 0 | 0 
grade 3 holosystolic apical murmur | 0 | 0 
mitral valve regurgitation | 0 | 0 
long-term venous access port | -672 | 0 
anemia | -672 | 0 
transfusion-dependent anemia | -672 | 0 
hemoglobin 12.1 g/dL | 0 | 0 
white blood cell count 15.1×10^3/µL | 0 | 0 
absolute neutrophil count 13.2×10^3/µL | 0 | 0 
b-type natriuretic peptide 788 pg/mL | 0 | 0 
congestive heart failure | 0 | 0 
left bundle branch pattern | 0 | 0 
Corynebacterium CDC group G bacteremia | 0 | 0 
gram positive rods | 0 | 0 
moderate mitral valve regurgitation | 0 | 0 
thickened anterior mitral leaflet | 0 | 0 
vegetations | 0 | 0 
severely elevated pulmonary artery systolic pressure | 0 | 0 
bacterial IE | 0 | 0 
vancomycin | 0 | 168 
clindamycin | 0 | 168 
discharged | 120 | 120 
readmitted | 168 | 168 
shortness of breath | 168 | 168 
hypoxic | 168 | 168 
elevated white blood cell count | 168 | 168 
severe mitral valve regurgitation | 168 | 168 
large and mobile vegetation | 168 | 168 
mitral valve replacement | 168 | 168 
coronary artery bypass grafting | 168 | 168 
oliguric acute renal failure | 168 | 168 
respiratory failure | 168 | 168 
mechanical ventilation | 168 | 168 
vancomycin resistant enterococcus | 168 | 168 
urinary tract infection | 168 | 168 
daptomycin | 168 | 504 
worsening congestive heart failure | 360 | 360 
transesophageal echocardiogram | 408 | 408 
severe mitral valve regurgitation | 408 | 408 
recurrent endocarditis | 408 | 408 
doxycycline | 504 | 504 
aztreonam | 504 | 504 
anidulafungin | 504 | 504 
bioprosthetic mitral valve replaced | 504 | 504 
St. Jude’s mechanical mitral valve | 504 | 504 
limb ischemia | 552 | 552 
disseminated intravascular coagulation | 552 | 552 
multi-organ failure | 552 | 552 
expired | 552 | 552 
diphtheroids | -672 | 0 
native valve endocarditis | 0 | 552 
prosthetic valve endocarditis | 168 | 552 
Corynebacterium CDC group G | -672 | 552 
line-associated bacteremia | -672 | 0 
pneumonia | -672 | -672 
levofloxacin | -672 | -656 
chronic implanted venous access device | -672 | 0 
infective endocarditis | 0 | 552 
mitral valve | 0 | 552 
aortic valve | 0 | 0 
porcine valves | 0 | 0 
Bjork-Shiley prosthetic valves | 0 | 0 
rheumatic fever | 0 | 0 
degenerative valve disease | 0 | 0 
mitral valve prolapse | 0 | 0 
intravenous drug misuse | 0 | 0 
vascular instrumentation | 0 | 0 
health-care associated infections | 0 | 552 
nosocomial bloodstream infections | 0 | 552 
polymicrobial infections | 0 | 552 
contaminants | 0 | 552 
colonizers | 0 | 552 
clinician communication | 0 | 552 
microbiology laboratory | 0 | 552 
adequate identification | 0 | 552 
adequate therapy | 0 | 552 
fatal illness | 552 | 552 
high rate of mortality | 552 | 552 
native valve | 0 | 168 
prosthetic valve | 168 | 552 
bioprosthetic valve | 168 | 504 
mechanical valve | 504 | 552 
Edwards-Carpentier pericardial valve | 168 | 504 
St. Jude’s prosthesis | 504 | 552 
reverse saphenous vein graft | 168 | 168 
distal right coronary artery | 168 | 168 
fibrinopurulent exudate | 168 | 168 
granulation tissue | 168 | 168 
endocarditis | 0 | 552 
diphtheroids | -672 | 552 
Corynebacterium CDC group G-1 | 0 | 0 
Corynebacterium CDC group G-2 | 0 | 0 
Corynebacterium CDC group G | 0 | 552 
vancomycin resistant enterococcus | 168 | 168 
VRE | 168 | 168 
daptomycin | 168 | 504 
doxycycline | 504 | 504 
aztreonam | 504 | 504 
anidulafungin | 504 | 504 
mechanical ventilation | 168 | 504 
acute kidney injury | 168 | 504 
respiratory failure | 168 | 504 
sepsis | 504 | 552 
fever | 0 | 552 
hypotension | 504 | 552 
transesophageal echocardiography | 408 | 408 
mitral regurgitation | 408 | 552 
recurrent vegetations | 408 | 552 
bioprosthetic mitral valve | 168 | 504 
St. Jude’s mechanical mitral valve | 504 | 552 
limb ischemia | 552 | 552 
disseminated intravascular coagulation | 552 | 552 
multi-organ failure | 552 | 552 
expired | 552 | 552 
native mitral valve | 0 | 168 
mitral valve leaflet | 168 | 168 
endocarditis | 0 | 552 
fibrinopurulent exudate | 168 | 168 
granulation tissue | 168 | 168 
diphtheroids | -672 | 552 
Corynebacterium CDC group G | -672 | 552 
line-associated bacteremia | -672 | 0 
pneumonia | -672 | -672 
levofloxacin | -672 | -656 
chronic implanted venous access device | -672 | 0 
infective endocarditis | 0 | 552 
mitral valve | 0 | 552 
aortic valve | 0 | 0 
porcine valves | 0 | 0 
Bjork-Shiley prosthetic valves | 0 | 0 
rheumatic fever | 0 | 0 
degenerative valve disease | 0 | 0 
mitral valve prolapse | 0 | 0 
intravenous drug misuse | 0 | 0 
vascular instrumentation | 0 | 0 
health-care associated infections | 0 | 552 
nosocomial bloodstream infections | 0 | 552 
polymicrobial infections | 0 | 552 
contaminants | 0 | 552 
colonizers | 0 | 552 
clinician communication | 0 | 552 
microbiology laboratory | 0 | 552 
adequate identification | 0 | 552 
adequate therapy | 0 | 552 
fatal illness | 552 | 552 
high rate of mortality | 552 | 552 
native valve | 0 | 168 
prosthetic valve | 168 | 552 
bioprosthetic valve | 168 | 504 
mechanical valve | 504 | 552 
Edwards-Carpentier pericardial valve | 168 | 504 
St. Jude’s prosthesis | 504 | 552 
reverse saphenous vein graft | 168 | 168 
distal right coronary artery | 168 | 168 
fibrinopurulent exudate | 168 | 168 
granulation tissue | 168 | 168 
endocarditis | 0 | 552 
diphtheroids | -672 | 552 
Corynebacterium CDC group G-1 | 0 | 0 
Corynebacterium CDC group G-2 | 0 | 0 
Corynebacterium CDC group G | 0 | 552 
vancomycin resistant enterococcus | 168 | 168 
VRE | 168 | 168 
daptomycin | 168 | 504 
doxycycline | 504 | 504 
aztreonam | 504 | 504 
anidulafungin | 504 | 504 
mechanical ventilation | 168 | 504 
acute kidney injury | 168 | 504 
respiratory failure | 168 | 504 
sepsis | 504 | 552 
fever | 0 | 552 
hypotension | 504 | 552 
transesophageal echocardiography | 408 | 408 
mitral regurgitation | 408 | 552 
recurrent vegetations | 408 | 552 
bioprosthetic mitral valve | 168 | 504 
St. Jude’s mechanical mitral valve | 504 | 552 
limb ischemia | 552 | 552 
disseminated intravascular coagulation | 552 | 552 
multi-organ failure | 552 | 552 
expired | 552 | 552 
native mitral valve | 0 | 168 
mitral valve leaflet | 168 | 168 
endocarditis | 0 | 552 
fibrinopurulent exudate | 168 | 168 
granulation tissue | 168 | 168 
diphtheroids | -672 | 552 
Corynebacterium CDC group G | -672 | 552 
line-associated bacteremia | -672 | 0 
pneumonia | -672 | -672 
levofloxacin | -672 | -656 
chronic implanted venous access device | -672 | 0 
infective endocarditis | 0 | 552 
mitral valve | 0 | 552 
aortic valve | 0 | 0 
porcine valves | 0 | 0 
Bjork-Shiley prosthetic valves | 0 | 0 
rheumatic fever | 0 | 0 
degenerative valve disease | 0 | 0 
mitral valve prolapse | 0 | 0 
intravenous drug misuse | 0 | 0 
vascular instrumentation | 0 | 0 
health-care associated infections | 0 | 552 
nosocomial bloodstream infections | 0 | 552 
polymicrobial infections | 0 | 552 
contaminants | 0 | 552 
colonizers | 0 | 552 
clinician communication | 0 | 552 
microbiology laboratory | 0 | 552 
adequate identification | 0 | 552 
adequate therapy | 0 | 552 
fatal illness | 552 | 552 
high rate of mortality | 552 | 552 
native valve | 0 | 168 
prosthetic valve | 168 | 552 
bioprosthetic valve | 168 | 504 
mechanical valve | 504 | 552 
Edwards-Carpentier pericardial valve | 168 | 504 
St. Jude’s prosthesis | 504 | 552 
reverse saphenous vein graft | 168 | 168 
distal right coronary artery | 168 | 168 
fibrinopurulent exudate | 168 | 168 
granulation tissue | 168 | 168 
endocarditis | 0 | 552 
diphtheroids | -672 | 552 
Corynebacterium CDC group G-1 | 0 | 0 
Corynebacterium CDC group G-2 | 0 | 0 
Corynebacterium CDC group G | 0 | 552 
vancomycin resistant enterococcus | 168 | 168 
VRE | 168 | 168 
daptomycin | 168 | 504 
doxycycline | 504 | 504 
aztreonam | 504 | 504 
anidulafungin | 504 | 504 
mechanical ventilation | 168 | 504 
acute kidney injury | 168 | 504 
respiratory failure | 168 | 504 
sepsis | 504 | 552 
fever | 0 | 552 
hypotension | 504 | 552 
transesophageal echocardiography | 408 | 408 
mitral regurgitation | 408 | 552 
recurrent vegetations | 408 | 552 
bioprosthetic mitral valve | 168 | 504 
St. Jude’s mechanical mitral valve | 504 | 552 
limb ischemia | 552 | 552 
disseminated intravascular coagulation | 552 | 552 
multi-organ failure | 552 | 552 
expired | 552 | 552 
native mitral valve | 0 | 168 
mitral valve leaflet | 168 | 168 
endocarditis | 0 | 552 
fibrinopurulent exudate | 168 | 168 
granulation tissue | 168 | 168 
diphtheroids | -672 | 552 
Corynebacterium CDC group G | -672 | 552 
line-associated bacteremia | -672 | 0 
pneumonia | -672 | -672 
levofloxacin | -672 | -656 
chronic implanted venous access device | -672 | 0 
infective endocarditis | 0 | 552 
mitral valve | 0 | 552 
aortic valve | 0 | 0 
porcine valves | 0 | 0 
Bjork-Shiley prosthetic valves | 0 | 0 
rheumatic fever | 0 | 0 
degenerative valve disease | 0 | 0 
mitral valve prolapse | 0 | 0 
intravenous drug misuse | 0 | 0 
vascular instrumentation | 0 | 0 
health-care associated infections | 0 | 552 
nosocomial bloodstream infections | 0 | 552 
polymicrobial infections | 0 | 552 
contaminants | 0 | 552 
colonizers | 0 | 552 
clinician communication | 0 | 552 
microbiology laboratory | 0 | 552 
adequate identification | 0 | 552 
adequate therapy | 0 | 552 
fatal illness | 552 | 552 
high rate of mortality | 552 | 552 
native valve | 0 | 168 
prosthetic valve | 168 | 552 
bioprosthetic valve | 168 | 504 
mechanical valve | 504 | 552 
Edwards-Carpentier pericardial valve | 168 | 504 
St. Jude’s prosthesis | 504 | 552 
reverse saphenous vein graft | 168 | 168 
distal right coronary artery | 168 | 168 
fibrinopurulent exudate | 168 | 168 
granulation tissue | 168 | 168 
endocarditis | 0 | 552 
diphtheroids | -672 | 552 
Corynebacterium CDC group G-1 | 0 | 0 
Corynebacterium CDC group G-2 | 0 | 0 
Corynebacterium CDC group G | 0 | 552 
vancomycin resistant enterococcus | 168 | 168 
VRE | 168 | 168 
daptomycin | 168 | 504 
doxycycline | 504 | 504 
aztreonam | 504 | 504 
anidulafungin | 504 | 504 
mechanical ventilation | 168 | 504 
acute kidney injury | 168 | 504 
respiratory failure | 168 | 504 
sepsis | 504 | 552 
fever | 0 | 552 
hypotension | 504 | 552 
transesophageal echocardiography | 408 | 408 
mitral regurgitation | 408 | 552 
recurrent vegetations | 408 | 552 
bioprosthetic mitral valve | 168 | 504 
St. Jude’s mechanical mitral valve | 504 | 552 
limb ischemia | 552 | 552 
disseminated intravascular coagulation | 552 | 552 
multi-organ failure | 552 | 552 
expired | 552 | 552 
native mitral valve | 0 | 168 
mitral valve leaflet | 168 | 168 
endocarditis | 0 | 552 
fibrinopurulent exudate | 168 | 168 
granulation tissue | 168 | 168 
diphtheroids | -672 | 552 
Corynebacterium CDC group G | -672 | 552 
line-associated bacteremia | -672 | 0 
pneumonia | -672 | -672 
levofloxacin | -672 | -656 
chronic implanted venous access device | -672 | 0 
infective endocarditis | 0 | 552 
mitral valve | 0 | 552 
aortic valve | 0 | 0 
porcine valves | 0 | 0 
Bjork-Shiley prosthetic valves | 0 | 0 
rheumatic fever | 0 | 0 
degenerative valve disease | 0 | 0 
mitral valve prolapse | 0 | 0 
intravenous drug misuse | 0 | 0 
vascular instrumentation | 0 | 0 
health-care associated infections | 0 | 552 
nosocomial bloodstream infections | 0 | 552 
polymicrobial infections | 0 | 552 
contaminants | 0 | 552 
colonizers | 0 | 552 
clinician communication | 0 | 552 
microbiology laboratory | 0 | 552 
adequate identification | 0 | 552 
adequate therapy | 0 | 552 
fatal illness | 552 | 552 
high rate of mortality | 552 | 552 
native valve | 0 | 168 
prosthetic valve | 168 | 552 
bioprosthetic valve | 168 | 504 
mechanical valve | 504 | 552 
Edwards-Carpentier pericardial valve | 168 | 504 
St. Jude’s prosthesis | 504 | 552 
reverse saphenous vein graft | 168 | 168 
distal right coronary artery | 168 | 168 
fibrinopurulent exudate | 168 | 168 
granulation tissue | 168 | 168 
endocarditis | 0 | 552 
diphtheroids | -672 | 552 
Corynebacterium CDC group G-1 | 0 | 0 
Corynebacterium CDC group G-2 | 0 | 0 
Corynebacterium CDC group G | 0 | 552 
vancomycin resistant enterococcus | 168 | 168 
VRE | 168 | 168 
daptomycin | 168 | 504 
doxycycline | 504 | 504 
aztreonam | 504 | 504 
anidulafungin | 504 | 504 
mechanical ventilation | 168 | 504 
acute kidney injury | 168 | 504 
respiratory failure | 168 | 504 
sepsis | 504 | 552 
fever | 0 | 552 
hypotension | 504 | 552 
transesophageal echocardiography | 408 | 408 
mitral regurgitation | 408 | 552 
recurrent vegetations | 408 | 552 
bioprosthetic mitral valve | 168 | 504 
St. Jude’s mechanical mitral valve | 504 | 552 
limb ischemia | 552 | 552 
disseminated intravascular coagulation | 552 | 552 
multi-organ failure | 552 | 552 
expired | 552 | 552 
native mitral valve | 0 | 168 
mitral valve leaflet | 168 | 168 
endocarditis | 0 | 552 
fibrinopurulent exudate | 168 | 168 
granulation tissue | 168 | 168 
diphtheroids | -672 | 552 
Corynebacterium CDC group G | -672 | 552 
line-associated bacteremia | -672 | 0 
pneumonia | -672 | -672 
levofloxacin | -672 | -656 
chronic implanted venous access device | -672 | 0 
infective endocarditis | 0 | 552 
mitral valve | 0 | 552 
aortic valve | 0 | 0 
porcine valves | 0 | 0 
Bjork-Shiley prosthetic valves | 0 | 0 
rheumatic fever | 0 | 0 
degenerative valve disease | 0 | 0 
mitral valve prolapse | 0 | 0 
intravenous drug misuse | 0 | 0 
vascular instrumentation | 0 | 0 
health-care associated infections | 0 | 552 
nosocomial bloodstream infections | 0 | 552 
polymicrobial infections | 0 | 552 
contaminants | 0 | 552 
colonizers | 0 | 552 
clinician communication | 0 | 552 
microbiology laboratory | 0 | 552 
adequate identification | 0 | 552 
adequate therapy | 0 | 552 
fatal illness | 552 | 552 
high rate of mortality | 552 | 552 
native valve | 0 | 168 
prosthetic valve | 168 | 552 
bioprosthetic valve | 168 | 504 
mechanical valve | 504 | 552 
Edwards-Carpentier pericardial valve | 168 | 504 
St. Jude’s prosthesis | 504 | 552 
reverse saphenous vein graft | 168 | 168 
distal right coronary artery | 168 | 168 
fibrinopurulent exudate | 168 | 168 
granulation tissue | 168 | 168 
endocarditis | 0 | 552 
diphtheroids | -672 | 552 
Corynebacterium CDC group G-1 | 0 | 0 
Corynebacterium CDC group G-2 | 0 | 0 
Corynebacterium CDC group G | 0 | 552 
vancomycin resistant enterococcus | 168 | 168 
VRE | 168 | 168 
daptomycin | 168 | 504 
doxycycline | 504 | 504 
aztreonam | 504 | 504 
anidulafungin | 504 | 504 
mechanical ventilation | 168 | 504 
acute kidney injury | 168 | 504 
respiratory failure | 168 | 504 
sepsis | 504 | 552 
fever | 0 | 552 
hypotension | 504 | 552 
transesophageal echocardiography | 408 | 408 
mitral regurgitation | 408 | 552 
recurrent vegetations | 408 | 552 
bioprosthetic mitral valve | 168 | 504 
St. Jude’s mechanical mitral valve | 504 | 552 
limb ischemia | 552 | 552 
disseminated intravascular coagulation | 552 | 552 
multi-organ failure | 552 | 552 
expired | 552 | 552 
native mitral valve | 0 | 168 
mitral valve leaflet | 168 | 168 
endocarditis | 0 | 552 
fibrinopurulent exudate | 168 | 168 
granulation tissue | 168 | 168 
diphtheroids | -672 | 552 
Corynebacterium CDC group G | -672 | 552 
line-associated bacteremia | -672 | 0 
pneumonia | -672 | -672 
levofloxacin | -672 | -656 
chronic implanted venous access device | -672 | 0 
infective endocarditis | 0 | 552 
mitral valve | 0 | 552 
aortic valve | 0 | 0 
porcine valves | 0 | 0 
Bjork-Shiley prosthetic valves | 0 | 0 
rheumatic fever | 0 | 0 
degenerative valve disease | 0 | 0 
mitral valve prolapse | 0 | 0 
intravenous drug misuse | 0 | 0 
vascular instrumentation | 0 | 0 
health-care associated infections | 0 | 552 
nosocomial bloodstream infections | 0 | 552 
polymicrobial infections | 0 | 552 
contaminants | 0 | 552 
colonizers | 0 | 552 
clinician communication | 0 | 552 
microbiology laboratory | 0 | 552 
adequate identification | 0 | 552 
adequate therapy | 0 | 552 
fatal illness | 552 | 552 
high rate of mortality | 552 | 552 
native valve | 0 | 168 
prosthetic valve | 168 | 552 
bioprosthetic valve | 168 | 504 
mechanical valve | 504 | 552 
Edwards-Carpentier pericardial valve | 168 | 504 
St. Jude’s prosthesis | 504 | 552 
reverse saphenous vein graft | 168 | 168 
distal right coronary artery | 168 | 168 
fibrinopurulent exudate | 168 | 168 
granulation tissue | 168 | 168 
endocarditis | 0 | 552 
diphtheroids | -672 | 552 
Corynebacterium CDC group G-1 | 0 | 0 
Corynebacterium CDC group G-2 | 0 | 0 
Corynebacterium CDC group G | 0 | 552 
vancomycin resistant enterococcus | 168 | 168 
VRE | 168 | 168 
daptomycin | 168 | 504 
doxycycline | 504 | 504 
aztreonam | 504 | 504 
anidulafungin | 504 | 504 
mechanical ventilation | 168 | 504 
acute kidney injury | 168 | 504 
respiratory failure | 168 | 504 
sepsis | 504 | 552 
fever | 0 | 552 
hypotension | 504 | 552 
transesophageal echocardiography | 408 | 408 
mitral regurgitation | 408 | 552 
recurrent vegetations | 408 | 552 
bioprosthetic mitral valve | 168 | 504 
St. Jude’s mechanical mitral valve | 504 | 552 
limb ischemia | 552 | 552 
disseminated intravascular coagulation | 552 | 552 
multi-organ failure | 552 | 552 
expired | 552 | 552 
native mitral valve | 0 | 168 
mitral valve leaflet | 168 | 168 
endocarditis | 0 | 552 
fibrinopurulent exudate | 168 | 168 
granulation tissue | 168 | 168 
diphtheroids | -672 | 552 
Corynebacterium CDC group G | -672 | 552 
line-associated bacteremia | -672 | 0 
pneumonia | -672 | -672 
levofloxacin | -672 | -656 
chronic implanted venous access device | -672 | 0 
infective endocarditis | 0 | 552 
mitral valve | 0 | 552 
aortic valve | 0 | 0 
porcine valves | 0 | 0 
Bjork-Shiley prosthetic valves | 0 | 0 
rheumatic fever | 0 | 0 
degenerative valve disease | 0 | 0 
mitral valve prolapse | 0 | 0 
intravenous drug misuse | 0 | 0 
vascular instrumentation | 0 | 0 
health-care associated infections | 0 | 552 
nosocomial bloodstream infections | 0 | 552 
polymicrobial infections | 0 | 552 
contaminants | 0 | 552 
colonizers | 0 | 552 
clinician communication | 0 | 552 
microbiology laboratory | 0 | 552 
adequate identification | 0 | 552 
adequate therapy | 0 | 552 
fatal illness | 552 | 552 
high rate of mortality | 552 | 552 
native valve | 0 | 168 
prosthetic valve | 168 | 552 
bioprosthetic valve | 168 | 504 
mechanical valve | 504 | 552 
Edwards-Carpentier pericardial valve | 168 | 504 
St. Jude’s prosthesis | 504 | 552 
reverse saphenous vein graft | 168 | 168 
distal right coronary artery | 168 | 168 
fibrinopurulent exudate | 168 | 168 
granulation tissue | 168 | 168 
endocarditis | 0 | 552 
diphtheroids | -672 | 552 
Corynebacterium CDC group G-1 | 0 | 0 
Corynebacterium CDC group G-2 | 0 | 0 
Corynebacterium CDC group G | 0 | 552 
vancomycin resistant enterococcus | 168 | 168 
VRE | 168 | 168 
daptomycin | 168 | 504 
doxycycline | 504 | 504 
aztreonam | 504 | 504 
anidulafungin | 504 | 504 
mechanical ventilation | 168 | 504 
acute kidney injury | 168 | 504 
respiratory failure | 168 | 504 
sepsis | 504 | 552 
fever | 0 | 552 
hypotension | 504 | 552 
transesophageal echocardiography | 408 | 408 
mitral regurgitation | 408 | 552 
recurrent vegetations | 408 | 552 
bioprosthetic mitral valve | 168 | 504 
St. Jude’s mechanical mitral valve | 504 | 552 
limb ischemia | 552 | 552 
disseminated intravascular coagulation | 552 | 552 
multi-organ failure | 552 | 552 
expired | 552 | 552 
native mitral valve | 0 | 168 
mitral valve leaflet | 168 | 168 
endocarditis | 0 | 552 
fibrinopurulent exudate | 168 | 168 
granulation tissue | 168 | 168 
diphtheroids | -672 | 552 
Corynebacterium CDC group G | -672 | 552 
line-associated bacteremia | -672 | 0 
pneumonia | -672 | -672 
levofloxacin | -672 | -656 
chronic implanted venous access device | -672 | 0 
infective endocarditis | 0 | 552 
mitral valve | 0 | 552 
aortic valve | 0 | 0 
porcine valves | 0 | 0 
Bjork-Shiley prosthetic valves | 0 | 0 
rheumatic fever | 0 | 0 
degenerative valve disease | 0 | 0 
mitral valve prolapse | 0 | 0 
intravenous drug misuse | 0 | 0 
vascular instrumentation | 0 | 0 
health-care associated infections | 0 | 552 
nosocomial bloodstream infections | 0 | 552 
polymicrobial infections | 0 | 552 
contaminants | 0 | 552 
colonizers | 0 | 552 
clinician communication | 0 | 552 
microbiology laboratory | 0 | 552 
adequate identification | 0 | 552 
adequate therapy | 0 | 552 
fatal illness | 552 | 552 
high rate of mortality | 552 | 552 
native valve | 0 | 168 
prosthetic valve | 168 | 552 
bioprosthetic valve | 168 | 504 
mechanical valve | 504 | 552 
Edwards-Carpentier pericardial valve | 168 | 504 
St. Jude’s prosthesis | 504 | 552 
reverse saphenous vein graft | 168 | 168 
distal right coronary artery | 168 | 168 
fibrinopurulent exudate | 168 | 168 
granulation tissue | 168 | 168 
endocarditis | 0 | 552 
diphtheroids | -672 | 552 
Corynebacterium CDC group G-1 | 0 | 0 
Corynebacterium CDC group G-2 | 0 | 0 
Corynebacterium CDC group G | 0 | 552 
vancomycin resistant enterococcus | 168 | 168 
VRE | 168 | 168 
daptomycin | 168 | 504 
doxycycline | 504 | 504 
aztreonam | 504 | 504 
anidulafungin | 504 | 504 
mechanical ventilation | 168 | 504 
acute kidney injury | 168 | 504 
respiratory failure | 168 | 504 
sepsis | 504 | 552 
fever | 0 | 552 
hypotension | 504 | 552 
transesophageal echocardiography | 408 | 408 
mitral regurgitation | 408 | 552 
recurrent vegetations | 408 | 552 
bioprosthetic mitral valve | 168 | 504 
St. Jude’s mechanical mitral valve | 504 | 552 
limb ischemia | 552 | 552 
disseminated intravascular coagulation | 552 | 552 
multi-organ failure | 552 | 552 
expired | 552 | 552 
native mitral valve | 0 | 168 
mitral valve leaflet | 168 | 168 
endocarditis | 0 | 552 
fibrinopurulent exudate | 168 | 168 
granulation tissue | 168 | 168 
diphtheroids | -672 | 552 
Corynebacterium CDC group G | -672 | 552 
line-associated bacteremia | -672 | 0 
pneumonia | -672 | -672 
levofloxacin | -672 | -656 
chronic implanted venous access device | -672 | 0 
infective endocarditis | 0 | 552 
mitral valve | 0 | 552 
aortic valve | 0 | 0 
porcine valves | 0 | 0 
