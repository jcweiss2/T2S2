55 years old | 0
male | 0
admitted to the hospital | 0
right femoropopliteal bypass | -1296
intermittent claudication | -1296
arterial insufficiency | -1296
stenosis of graft | -624
recurrence of symptoms | -624
right iliac artery - right popliteal artery bypass | -624
polytetrafluoroethylene (PTFE) graft | -624
gross hematuria | -48
sepsis | -48
insertion of three-way Foley catheter | -48
irrigation | -48
computed tomography (CT) scan | 0
angiography | 0
fistulous communication between right iliac artery and right ureter | 0
surrounding inflammatory changes | 0
covered stenting with PTFE graft | 0
antibiotic coverage | 0
monitored in intensive care unit | 0
Foley catheter removed | 120
afebrile | 120
discharged | 168
follow-up | 336
watery discharge from scar of previous surgery | 336
fistulous communication between the right ureter and overlying skin | 336
no communication with iliac artery | 336
cystoscopy | 336
retrograde pyelography | 336
JJ stent placed | 336
discharged | 448
no discharge | 504
no signs of arterial insufficiency | 504
no lower urinary tract symptoms | 504
JJ stent removed | 1008
stable on subsequent follow-ups | 1008