52 years old | 0
female | 0
admitted to the emergency department | 0
generalized abdominal discomfort | -96
altered mental status | -96
diarrhea | -96
fevers | -96
chills | -96
alcohol abuse | -96
alcohol-related liver cirrhosis | -96
blood pressure of 74/42 mmHg | 0
heart rate of 112 beats/min | 0
respiratory rate of 20 breaths/min | 0
temperature of 98.6 F | 0
jaundice | 0
abdominal distention | 0
tenderness to palpation | 0
right upper quadrant tenderness | 0
no rash | 0
no ulcers | 0
no recent travels | 0
no exposure to sick people | 0
no domestic animals at home | 0
no contact with pets | 0
mechanical ventilation | 0
admitted to the medical intensive care unit | 0
systemic inflammatory response syndrome | 0
sepsis | 0
septic shock | 0
multi-organic dysfunction syndrome | 0
community-acquired pneumonia | 0
possible biliary tract infection | 0
ascending cholangitis | 0
probable spontaneous bacterial peritonitis | 0
alcoholic hepatitis | 0
aggressive intravenous fluids resuscitation | 0
crystalloids | 0
vasopressors | 0
blood cultures | 0
urine cultures | 0
respiratory cultures | 0
legionella urine antigen | 0
empiric intravenous antimicrobial therapy | 0
piperacillin/tazobactam | 0
azithromycin | 0
complete blood cell count of 21,000/mm3 | 0
90% neutrophils | 0
platelet count of 51,000/mm3 | 0
sodium level of 127 mEq/L | 0
potassium level of 5.3 mEq/L | 0
bicarbonate level of 15 mEq/L | 0
creatinine level of 6.3 mg/dl | 0
aspartate aminotransferase level of 121 IU/L | 0
alanine aminotransferase level of 65 IU/L | 0
alkaline phosphatase level of 290 IU/L | 0
gamma-glutamyl transpeptidase level of 290 U/L | 0
lactate dehydrogenase level of 482 U/L | 0
total bilirubin level of 14.5 mg/dl | 0
direct bilirubin level of 10.1 mg/dl | 0
lactic acid level of 6.4 mg/dl | 0
prothrombin time of 25.2 s | 0
INR of 2.29 | 0
serum alcohol level within normal limits | 0
arterial blood gases pH of 7.15 | 0
pCO2 of 23 | 0
pO2 of 132 | 0
FIO2 of 60% | 0
chest X-ray left lung infiltrate | 0
pleural effusion | 0
blood cultures grew P. multocida | 24
isolate sensitive to piperacillin/tazobactam | 24
isolate sensitive to azithromycin | 24
medical condition deteriorated | 24
patient expired | 72
