41 years old | 0
male | 0
no significant past medical history | 0
lower extremity edema | -504
fatigue | -504
shortness of breath | -504
pale | 0
melenic stool | 0
admitted to the medical intensive care unit | 0
resuscitation | 0
urgent endoscopy | 0
multiple gastric ulcers | 0
diffuse lymphadenopathy | 0
metastatic lymphoma | 0
excisional biopsy | 0
Hodgkin lymphoma | 0
acute renal failure | 0
temporary hemodialysis | 0
acute respiratory failure | 0
intubation | 0
septic shock | 0
vasopressor support | 0
norepinephrine | 0
sedated | 0
propofol | 0
fentanyl | 0
ventilator | 0
telemetry displayed a sudden onset of ST-segment elevations | 0
abdominal distention | 0
no murmurs | 0
blood pressure of 101/57 mm Hg | 0
heart rate of 112 beats/min | 0
respiratory rate of 23 breaths/min | 0
oxygen saturation of 99% | 0
sinus tachycardia | 0
ST-segment elevations in the precordial leads | 0
deep T-wave inversions | 0
J-point depression in the inferior leads | 0
marked QT prolongation | 0
STEMI | 0
emergency cardiology consultation | 0
troponin-T level of <0.01 ng/ml | 0
potassium of 4.3 mEq/l | 0
calcium of 7.6 mg/dl | 0
anion gap of 12 mEq/l | 0
hemoglobin of 10.1 g/dl | 0
hematocrit of 29.4% | 0
arterial blood gas showed a pH of 7.40 | 0
bicarbonate of 21 mmol/l | 0
lactate of 3.1 mmol/l | 0
left ventricular ejection fraction to be 60% to 65% | 0
no regional wall motion abnormalities | 0
no pericardial effusion | 0
abrupt resolution of ST-segment elevations on telemetry | 0
gentle palpation of the abdomen | 0
resolution of ST-segment elevations | 0
gastric distention | 0
ileus | 0
gastric decompression with nasogastric tube placement | 24
resolution of ST-segment elevations | 24
coronary angiography was deferred | 24
new-onset seizures | 48
focal neurological deficits | 48
magnetic resonance imaging of the brain | 48
leptomeningeal enhancement | 48
metastatic spread | 48
comfort care | 72
died | 72