39 years old | 0
male | 0
admitted to the hospital | 0
fever | -168
diffuse myalgia | -168
pleuritic type precordial chest pain | -72
dyspnea | -72
diabetes mellitus type 1 | -6720
insulin treatment | -6720
apyrexial | 0
dyspneic at rest | 0
blood pressure of 160/90 mmHg | 0
pulse rate of 130 beats per minute | 0
distended jugular veins | 0
pericardial friction rub | 0
heart sounds were not muffled | 0
diminished sounds in bases | 0
electrocardiogram (ECG) showed sinus tachycardia | 0
normal amplitude QRS complexes | 0
concaved ST elevation | 0
concordant T waves | 0
reciprocal ST depression | 0
PR elevation | 0
PR depression | 0
chest radiography revealed a massively enlarged globular cardiac shadow | 0
left pleural effusion | 0
white-blood-cell count of 10 800/μl | 0
83% segmented cells | 0
9% lymphocytes | 0
hemoglobin of 10.5 g/dl | 0
platelet count of 182 000/μl | 0
CRP was 192 U/l | 0
renal and liver function tests were normal | 0
NT-proBNP levels was 1155 pg/ml | 0
admitted to the intensive care unit | 0
arterial line was placed | 0
pulsus paradoxus was observed | 0
echocardiogram performed | 24
good left ventricular function | 24
ejection fraction of 78% | 24
no signals of valve dysfunctions | 24
massive pericardial effusion | 24
right ventricular systolic collapse | 24
cardiac tamponade | 24
pericardiocentesis was performed | 24
hemodynamic stability was achieved | 24
direct aspiration of 160 ml purulent fluid | 24
laboratory analysis of the pericardial fluid showed 500 000 nucleated cells/μl | 24
80% segmented cells | 24
8% lymphocytes | 24
2% eosinophils | 24
1000 red blood cells/μl | 24
lactate dehydrogenase of 19 523 U/l | 24
triglycerides of 90 mg/dl | 24
glucose of 36 mg/dl | 24
protein of 5.9 g/dl | 24
pH of 6.0 | 24
gram-positive cocci | 24
no acid-fast bacilli were present | 24
vancomycin (1 g IV every 12 hours) was started | 24
rapid HIV test was performed | 24
positive result | 24
follow-up echocardiogram performed | 48
substantial reaccumulation of fluid in the pericardial sac | 48
right ventricular collapse | 48
urgent surgical approach was indicated | 48
drain was placed in the pericardial sac | 48
bacterial, fungal and tuberculous culture from pericardial fluid were set up | 48
Methicilin-sensitive S. aureus | 72
high levels of adenosine deaminase (ADA) | 72
>200 U/l | 72
episodes of fever | 120
continuous drainage of purulent fluid | 120
tuberculostatic drugs were initiated | 120
testing for human immunodeficiency virus was positive | 120
CD4 count was 28 cells/μl | 120
HIV viral load 347 609 copies/mm3 | 120
pericardial biopsy revealed non-specific inflammation pattern | 120
culture negative | 120
thoracic drain was placed | 120
large pleural effusion | 120
no evidence of empyema | 120
chest computed tomography (CT) did not reveal any pulmonary parenchymal lesion | 120
lymphadenopathy | 120
abdominal CT scan was normal | 120
fluid aspect reduced | 168
pericardial drain was removed | 168
pending pericardial fluid cultures persisted negatives | 168
fungal and tuberculous etiologies | 168
cytology for malignant cells of pericardial fluid was negative | 168
corticosteroids were not prescribed | 168
another echocardiogram was performed | 168
no fluid reaccumulation | 168
constrictive pericarditis patterns | 168
rifampin, isoniazid, pyrazinamide and ethambutol were prescribed | 168
elective pericardiectomy | 240