87 years old | 0
male | 0
presented to the emergency department | 0
right hand cellulitis | 0
bitten by pet dog | 0
coronary artery disease | 0
TIA | 0
hypertension | 0
hyperlipidemia | 0
osteoporosis | 0
glaucoma | 0
previously smoked a few cigarettes per day | -525600
quit smoking | -525600
denied illicit drug use | 0
intravenous ampicillin/sulbactam | 0
wound washed | 0
discharged | 0
oral amoxicillin/clavulanate | 0
orthopedic clinic follow up | 72
continued significant erythema | 72
edema | 72
warmth of the wound and hand | 72
hospitalized | 72
intravenous ampicillin/sulbactam | 72
vancomycin | 72
improvement | 72
discharged | 168
oral amoxicillin/clavulanate | 168
minocycline | 168
presented to emergency room | 336
ankle pain | 336
loose non-bloody bowel movements | 336
fever 102.7 F | 336
hypotension 90/62 | 336
tachycardia 108 bpm | 336
tachypnea 22 bpm | 336
oxygen saturation 87% | 336
breathing comfortably | 336
speaking comfortably | 336
faint crackles | 336
3/6 systolic murmur | 336
flat JVP | 336
mild erythema | 336
eschar on dorsal hand | 336
mild left ankle warmth | 336
mild left ankle edema | 336
leukocytosis 20.8 k/uL | 336
74% neutrophils | 336
20% lymphocytes | 336
2.8% eosinophils | 336
creatinine 1.38 mg/dL | 336
normal liver enzymes | 336
chest radiograph bilateral effusions | 336
bilateral upper lobe lung infiltrates | 336
diagnosed with ankle sprain | 336
hospitalized for severe sepsis | 336
pneumonia | 336
acute kidney injury | 336
intravenous ertapenem | 336
vancomycin | 336
azithromycin | 336
oral metronidazole | 336
worsening tachypnea | 480
hypoxia | 480
ongoing fevers | 480
supplemental oxygen 4 L/min | 480
leukocytosis 17.3 k/uL | 480
eosinophilia 22.8% | 480
chest film diffuse alveolar filling | 480
bilateral pleural effusions persisted | 480
CT chest diffuse bilateral airspace disease | 480
ground glass attenuation | 480
moderate bilateral pleural effusions | 480
trachea intubated | 480
flexible fiberoptic bronchoscopy | 480
BAL | 480
transbronchial biopsies | 480
liberation from mechanical ventilation failed | 480
reintubated | 480
mechanical ventilatory support | 480
FiO2 0.80 | 528
pneumothorax | 528
chest tube placed | 528
streptococcus parasanguinus | 528
urine culture Klebsiella | 528
C. difficile toxin negative | 528
urine legionella antigen negative | 528
coccidiodes IgG negative | 528
coccidiodes IgM negative | 528
antimicrobials tailored | 528
ampicillin/sulbactam | 528
ciprofloxacin | 528
BAL nucleated cells 515/uL | 528
6% neutrophils | 528
5% lymphocytes | 528
15% eosinophils | 528
transbronchial biopsies eosinophilia | 528
bacterial stains negative | 528
fungal stains negative | 528
mycobacterial stains negative | 528
viral stains negative | 528
methylprednisolone started | 528
leukocytosis 13.5 k/uL | 624
eosinophilia 8.3% | 624
defervesced | 720
marked gas exchange improvement | 720
liberated from mechanical ventilation | 720
supplemental oxygen 3 L/min | 720
eosinophilia 0.1% | 720
improvement in air space disease | 720
solumedrol transitioned to prednisone | 720
ciprofloxacin discontinued | 720
chest tube removed | 1008
transthoracic echocardiogram no endocarditis | 1008
repeat blood cultures sterile | 1008
vancomycin completed | 1008
discharged | 720
pulmonary clinic follow up | 1080
denied respiratory symptoms | 1080
prednisone taper | 1080
inhaled mometasone | 1080
denied illicit drug use |+0
