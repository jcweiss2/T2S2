29 years old | 0
    male | 0
    muscle pain | -144
    joint pain | -144
    general weakness | -144
    fever up to 39°C | -144
    pronounced liver dysfunction | -144
    total bilirubin 5.7 mg/dl | -144
    serum glutamic oxaloacetic transaminase 633 U/L | -144
    serum glutamic pyruvate transaminase 412 U/L | -144
    gamma-glutamyl transferase 161 U/L | -144
    lactate dehydrogenase 1668 U/L | -144
    C-reactive protein 519 mg/l | -144
    procalcitonin 1.28 ng/ml | -144
    increased leukocyte levels 14.8 × 10³/μl | -144
    acute respiratory failure | 0
    altered state of consciousness | 0
    continuous sedation | 0
    muscle relaxation | 0
    intubation | 0
    mechanical ventilation | 0
    FiO2 of 100% | 0
    SpO2 of 88.7% | 0
    hemodynamic instability | 0
    norepinephrine 0.6 μg/kg/min | 0
    broad-spectrum empirical antimicrobial therapy | 0
    meropenem 1 g every 8 h IV | 0
    azithromycin 500 mg once daily IV | 0
    oseltamivir 75 mg every 12 h | 0
    methylprednisolone 80 mg every 12 h IV | 0
    stress ulcer prophylaxis | 0
    thromboprophylaxis (UFH) | 0
    drug doses adjusted for renal function | 0
    continuous sedation | 168
    paralyzed | 168
    intubated | 168
    controlled mechanical ventilation (lung-protective ventilation) | 168
    continuous respiratory monitoring | 168
    hemodynamic monitoring | 168
    regular monitoring of arterial blood gases | 168
    prone positioning | 0
    chest CT showing massive bilateral pneumonia | 0
    minimal pleural effusions | 0
    bedside focus ultrasound | 0
    acute renal failure | 144
    CRRT started | 144
    progressing hemodynamic instability | 144
    uncontrolled inflammatory response | 144
    CytoSorb® adsorber installed into CRRT circuit | 144
    recurring septic episode | 240
    second CytoSorb® therapy session | 240
    norepinephrine requirements lowered to 0.15 μg/kg/min | 144
    norepinephrine discontinued 2 days later | 192
    deterioration of clinical condition | 240
    increase in norepinephrine demand | 240
    second CytoSorb® application | 240
    norepinephrine cessation 1 day later | 264
    CRP decreased to 330 mg/L | 144
    further decrease in CRP levels | 240
    leukocyte levels normalized | 240
    ventilation parameters improved | 144
    lung function improved | 144
    ICU delirium | 264
    treated with antipsychotics | 264
    prolonged intubation | 264
    inadequate state of consciousness | 264
    percutaneous tracheostomy | 264
    hemodynamic status stable | 264
    gradual recovery | 264
    satisfactory state of consciousness | 264
    successfully weaned off ventilator | 264
    transferred to general ward | 1152
    sent to rehabilitation clinic | 1200
    influenza A (H1N1) | -144
    multiorgan failure | 144
    CVVHDF mode | 144
    hemodynamic stabilization | 144
    decrease in circulating pro-inflammatory cytokines | 144
    rapid fall in white blood cells | 144
    removal of antibiotics monitored | 144
    inability to measure cytokine levels | 0
    therapeutic drug monitoring | 144
    bilateral pneumonia | -144
    control of inflammatory response | 144
    significant decrease in inflammation markers | 144
    gradual improvement in ventilation parameters | 144
    improved lung function | 144
    vasopressors discontinued | 192
