64 years old | 0
    male | 0
    diabetes | -24
    insulin | -24
    hypertension | -24
    amlodipine | -24
    admitted to intensive care unit | 0
    septic shock | 0
    undetermined cause of infection | 0
    leukocyturia | -24
    no individualized germs | -24
    normal chest X-ray | -24
    normal lumbar puncture | -24
    somnolent | 0
    febrile 38.5°C | 0
    desaturated 90% | 0
    hypotensive 80/40 mmHg | 0
    tachycardic 110 bpm | 0
    blood sugar level 3 g/l | 0
    sugar in urine | 0
    no acetone | 0
    positive inflammatory syndrome | 0
    white blood cells 20,000/µl | 0
    C-reactive protein 270 mg/l | 0
    platelets 100,000/µl | 0
    normal renal function | 0
    creatinine 9.97 mg/l | 0
    urea 0.15 g/l | 0
    painful infiltration left iliac fossa | 0
    crepitus left iliac fossa | 0
    abdomino-pelvic CT scan | 24
    destroyed left kidney | 24
    oval cavity hydrous content | 24
    aerial collection left iliac fossa 75x26 mm | 24
    fluid resuscitation ringer lactate 30 ml/kg | 24
    vasoactive drugs noradrenaline | 24
    initial dose noradrenaline 1 mg/h | 24
    noradrenaline gradually decreased | 24
    noradrenaline weaned at day 3 | 72
    glycemic control insulin infusion | 24
    empirical antibiotic therapy 10 days | 24
    imipenem 1 g/8h | 24
    ciprofloxacin 200 mg/12h | 24
    clinical improvement | 168
    medical treatment continued | 168
    no percutaneous drainage | 168
    transferred to urology department | 240
    C-reactive protein 60 mg/l | 240
    discharged | 312
    no impairment of renal function | 312
    <|eot_id|>