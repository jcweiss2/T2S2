27 years old | 0
female | 0
admitted to the hospital | 0
fever | -48
abdomen pain | -48
vomiting | -48
severe dehydration | -48
altered sensorium | 0
high plasma blood sugar | 0
severe metabolic acidosis | 0
severe hypokalemia | 0
urine ketone bodies were large | 0
acute onset flaccid paralysis | 24
paradoxical breathing | 28
intubated | 28
mechanical ventilation | 28
failure to wean off from mechanical ventilation | 48
neurophysician opinion | 48
nerve conduction velocity studies | 48
electromyography studies | 48
primary muscle disease with axonal polyneuropathy | 48
HBA1C | 72
GAD antibodies were positive | 72
CPK total increased | 72
blood cultures isolated coagulase-negative Staphylococcus | 72
urine culture isolates budding yeast cells | 72
cerebrospinal fluid examination was within normal limit | 72
magnetic resonance imaging brain revealed diffuse cerebral edema | 72
tracheostomy | 432
ventilator-associated pneumonia | 432
chest roentgenogram showed nonhomogeneous patches | 432
high-resolution computed tomography of chest suggested bilateral infiltration | 432
sputum culture was positive for Klebsiella pneumoniae | 432
diagnosis of type 1 diabetes mellitus | 120
diabetic ketoacidosis | 120
sepsis | 120
severe hypokalemia | 120
CIPNM | 120
hyperglycemia was controlled | 120
diabetic ketoacidosis was corrected | 120
pneumonia and sepsis were treated with antibiotics | 120
large potassium deficits were corrected | 120
intravenous immunoglobulins | 120
parenteral nutritional support | 120
antioxidant therapy | 120
physiotherapy | 120
clinically improved | 720
power was regained | 720
reflexes were present | 720
weaned off mechanical ventilation | 720
repeat electrophysiological studies suggested recovery | 720
discharged | 1080
grade 4/5 power in all the limbs | 1080
regular physiotherapy | 1080
insulin analogs | 1080