71 years old | 0
female | 0
admitted to the hospital | 0
unconscious state | 0
hypertension | -672
ischaemic heart disease | -672
peripheral vascular disease | -672
stroke | 0
head computed tomographic scan | 0
inotropic support | 24
septic shock | 24
elevated levels of inflammatory markers | 24
erythrocyte sedimentation rate | 24
C-reactive protein | 24
blood obtained | 24
yeast in both aerobic and anaerobic BacT/ALERT culture bottles | 24
caspofungin administered | 24
died | 72
yeast isolate identified as C. parapsilosis | 24
VITEK 2 yeast identification system | 24
referred to the Mycology Reference Laboratory | 24
CHROMagar Candida | 48
turquoise blue colonies | 48
acetate ascospore agar | 168
long ellipsoidal-shaped ascospores | 168
internally transcribed spacer region of ribosomal DNA amplified and sequenced | 168
DNA sequence data comparisons | 168
Lodderomyces elongisporus | 168
antifungal susceptibility determined | 168
Etest | 168
RPMI 1640 medium | 168
glucose | 168
amphotericin B | 168
fluconazole | 168
voriconazole | 168
posaconazole | 168
itraconazole | 168
flucytosine | 168
caspofungin | 168
micafungin | 168
lower limb ischaemia | -336
hospitalized | -336
discharged | -336
inoculation of the yeast from the skin | -672
translocation from the gastrointestinal tract | -672
endocarditis | -672
global prevalence | -672
Mexico | -672
Malaysia | -672
China | -672
Australia | -672
Middle East | -672
Japan | -672
Spain | -672
Korea | -672