22 years old | 0
female | 0
Rett syndrome | -6840
seizure disorders | -6840
constipation | -6840
air swallowing | -6840
difficulty in evacuation of stool | -6840
rectal enema | -672
rectal digitation for defecation | -672
abdominal distention | -168
vomiting | -168
hyperventilation episodes | -168
no stool discharge | -96
abdominal distension | 0
abdominal tenderness | 0
rebound | 0
septic appearance | 0
bloody discharge | 0
increased sphincter tonus | 0
decreased Turgol-tonus | 0
dilated bowel segments with air-fluid levels | 0
coffee-bean sign | 0
sigmoid volvulus | 0
acute abdomen | 0
increased Blood Urea Nitrogen | 0
increased creatinine | 0
increased white blood cell count | 0
increased serum sodium | 0
increased blood glucose | 0
increased plasma CRP levels | 0
acute metabolic acidosis | 0
sinus tachycardia | 0
QT interval 500 ms | 0
urgent laparotomy | 0
sigmoid volvulus | 0
colon tumor | 0
liver mass | 0
Hartman procedure | 0
liver biopsy | 0
septic shock | 24
pulmonary and cardiac functions deteriorated | 48
death | 48
musinous adenocarcinoma | 48
adenocarcinoma metastasis | 48