57 years old | 0
male | 0
admitted to the emergency department | 0
right flank pain | 0
high fever | 0
poor health | 0
urosepsis | 0
right nephrolithotomy | -672
stenting during angiography | -672
coronary heart disease | -672
kidney stones | -672
multiple kidney stones | 0
pyonephrosis | 0
renal cyst | 0
nephrostomy catheter inserted | -24
intravenous antibiotic therapy | -24
nephrectomy | 0
cyst excision | 0
preoxygenation with 100% oxygen | 0
anesthesia induced with thiopental | 0
anesthesia induced with rocuronium | 0
anesthesia maintained with sevoflurane | 0
endotracheal intubation | 0
nephrectomy operation started under laparoscopy | 0
operation converted to open surgery | 0
cyst ruptured | 50
content of the cyst diffused to the retroperitoneal area | 50
surgeon aspirated and irrigated the area | 50
operation continued | 50
anaesthesia ended | 100
patient extubated | 100
patient had difficulty in breathing | 115
patient agitated | 115
blood gas analysis | 118
hypoxaemia | 118
pH: 7.49 | 118
pO2: 54 mmHg | 118
pCO2: 30 mmHg | 118
HCO3: 23 | 118
SpO2: 88 | 118
patient taken to the intensive care unit | 120
respiratory distress | 120
decreased right lung sounds | 120
pleural effusion | 120
thoracentesis | 120
chest tube insertion | 120
cultures of the pleural effusion | 120
cultures of cyst fluid | 120
Klebsiella pneumoniae | 120
imipenem administered | 120
linezolid administered | 120
metronidazole administered | 120
diaphragm intact during surgery | 120
no defect on CT | 120
retroperitoneal fluid transition through the diaphragmatic pores | 120
patient's general condition improved | 192
antibiotic therapy | 192
drainage of the pleural fluid | 192
pathology report indicated chronic pyelonephritis | 192
patient referred to the urology department | 96
improvement in blood gas values | 96
pH: 7.35 | 96
pO2: 88 mmHg | 96
pCO2: 36 mmHg | 96
HCO3: 24 | 96
SpO2: 96 | 96
respiratory parameters improved | 96
chest radiography improved | 96
chest tube removed | 288
patient discharged | 288