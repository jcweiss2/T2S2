pre-term birth | -2600
developmental delays in growth and motor function | -2600
short stature | -2080
Russell–Silver syndrome | -2080
proteinuria | -2080
hypoalbuminemia | -2080
nephrotic syndrome | -2080
high-dose steroid treatment | -2080
calcineurin inhibitor treatment | -2080
renal function deterioration | -2080
right renal vein thrombosis | -1040
pulmonary embolism | -1040
anticoagulant treatment | -1040
persistent pulmonary hypertension | -1040
sildenafil treatment | -1040
living donor kidney transplantation | 0
immunosuppression with prednisolone, mycophenolate mofetil (MMF), and tacrolimus | 0
discontinuation of MMF | 70
tapering of steroid | 70
pneumocystis pneumonia | 90
mechanical ventilation | 90
intravenous sulfamethoxazole/trimethoprim treatment | 90
increase in steroid dose | 90
discharge | 104
dysuria | 135
gross hematuria | 135
elevated blood urea nitrogen (BUN) | 135
elevated creatinine (Cr) | 135
elevated C-reactive protein (CRP) | 135
urinalysis with red blood cell (RBC) count > 100/high power fields (HPF) | 135
urinalysis with white blood cell (WBC) count > 100/HPF | 135
negative urine culture for bacteria and BK virus | 135
positive urine John Cunningham (JC) virus polymerase chain reaction (PCR) | 135
positive urine adenovirus culture | 135
diagnosis of hemorrhagic cystitis | 135
hydration and pain control treatment | 135
persistent dysuria and hematuria | 142
elevated RBC count | 142
elevated WBC count | 142
fever | 159
general weakness | 159
chest tightness | 159
mild cough | 159
persistent dysuria | 159
persistent hematuria | 159
elevated BUN | 159
elevated Cr | 159
elevated CRP | 159
emergent hemodialysis | 159
empirical treatment with piperacillin/tazobactam | 159
negative sputum, blood, and urine culture results | 159
positive adenovirus real-time PCR of sputum | 159
positive blood cytomegalovirus (CMV) antigen | 159
presumed diagnosis of disseminated adenovirus infection | 159
reduction of immunosuppression | 159
ganciclovir treatment | 159
renal allograft biopsy | 159
diffuse necrotizing granulomatous tubulointerstitial nephritis | 159
negative staining for CD3 and C4d | 159
positive JC virus PCR | 159
positive serum CMV PCR | 159
coinfection | 159
treatment with ganciclovir, antibiotic therapy, granulocyte colony-stimulating factor, immunoglobulin, transfusion, and hemodialysis | 159
persistent high inflammatory marker and fever | 167
initiation of cidofovir treatment | 167
nephrotoxicity | 167
administration of 4 doses of cidofovir | 170
change in cidofovir regimen to 2 mg/kg every 2 weeks | 170
positive serum adenovirus PCR | 174
positive cerebrospinal fluid adenovirus PCR | 174
unrecovered renal function | 174
generalized tonic-clonic seizure | 174
treatment with vancomycin, meropenem, and acyclovir | 174
deterioration of general condition | 174
anemia | 180
leukopenia | 180
thrombocytopenia | 180
bone marrow suppression | 180
intensive care, including mechanical ventilation and continuous renal replacement therapy | 180
death | 215