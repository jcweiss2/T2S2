83 years old | 0
female | 0
weight loss | -72
dyspepsia | -72
abdominal pain | -72
fever | -48
admitted to the emergency department | 0
hypertension | 0
diabetes mellitus | 0
no history of trauma | 0
no history of surgery | 0
no history of alcoholism | 0
no history of smoking | 0
blood pressure 110/70 mmHg | 0
no history of coronary artery disease | 0
normal heart sounds | 0
diminished bowel sounds | 0
abdomen distended | 0
diffuse defense | 0
rebound | 0
sensitivity | 0
white blood cell 10.8 10^3/ml | 0
hemoglobin 8.1 g/dl | 0
urea 38 mg/dL | 0
creatinin 1.6 mg/dL | 0
potassium 5.7 mmol/L | 0
normal blood amylase level | 0
normal electrocardiogram | 0
free air under the right diaphragm | 0
widespread free abdominal fluid | 0
admitted to the intensive care unit | 0
supportive therapy | 0
operating room | 0
midline laparotomy | 0
giant perforation | 0
purulent material aspirated | 0
peritoneal cavity washed | 0
biopsies from the edges of the perforation | 0
gastric resection not suitable | 0
purse-string sutures | 0
omental flap prepared | 0
omental flap transfixed | 0
leaking areas checked | 0
methylene blue test | 0
drains placed | 0
operation time 40 min | 0
intubated | 0
Meropenem 3*1 gr/iv | 0
infection diseases department consultation | 0
white blood cell count reduced | 24
pre-renal failure improved | 24
inotropic agents decreased | 24
inotropic agents stopped | 48
abdomen smooth | 120
abdomen free from distension | 120
abdomen free from rigidity | 120
methylene blue test | 120
no leakage | 120
abdominal drains withdrawn | 120
pulmonary problems not recovered | 120
acquired pneumonia | 120
sedation given up | 120
mechanical ventilator weaning | 120
pulmonary failure | 360
died | 360
histopathology examination | 360
moderately differentiated adenocarcinoma | 360