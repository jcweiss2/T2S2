sports-related injury to her left shoulder | -1080
surgical revisions | -1080
recurrent and prolonged shoulder infections | -1080
Pseudomonas aeruginosa infection | -1080
Sphingomonas paucimobilis infection | -1080
Candida colliculosa infection | -1080
Staphylococcus aureus infection | -1080
left shoulder tendon release and revision | -240
development of CRPS | -240
severe pain | 0
allodynia | 0
edema | 0
muscle spasms | 0
temperature changes of her LUE | 0
electromyography evaluation | 0
brachial plexus injury | 0
asthma | 0
selective IgG3 deficiency | 0
oral medical management | 0
opioids | 0
antidepressants | 0
antispasmodics | 0
left stellate ganglion blockade | 0
continuous cervical epidural infusions | 0
placement of a left C6–C7 interlaminar epidural catheter | 0
transfer to the postanesthesia care unit | 0
preprocedure labs | 0
antibiotic prophylaxis with vancomycin | -1
epidural infusion of 0.25% bupivacaine with hydromorphone and clonidine | 0
oral home medications | 0
methadone | 0
hydromorphone | 0
diazepam | 0
baclofen | 0
amitriptyline | 0
decrease in pain | 24
less muscle spasms | 24
improved sleep | 48
increased infusion to 6 mL per hour | 48
demand dose of 2 mL every 15 minutes | 48
febrile to 38.1°C | 120
wean the infusion | 120
remove the epidural catheter | 126
progressive headache | 130
neck pain | 130
increase in temperature to 40.0°C | 130
neurological examination | 130
blood and urine cultures | 130
chest x-ray | 130
laboratory workup | 130
increase in white count | 130
cephalosporin | 130
abatement of fever | 130
decrease in white count | 130
MRI of the cervical spine | 132
epidural collection | 132
interstitial edema in the left paraspinal muscles | 132
transfer to the neurosciences intensive care unit | 132
hourly neurological examination | 132
intractable nausea and vomiting | 156
left arm weakness | 156
emergent decompression and evacuation | 156
intraoperative cultures | 156
P aeruginosa infection | 156
vancomycin stopped | 156
cefepime continued | 156
resolution of arm weakness | 180
uneventful postoperative course | 180
discharged home | 180
intravenous cefepime | 180