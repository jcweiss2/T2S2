8 years old | 0
male | 0
admitted to hospital | 0
flame burn injury | -72
intubated and ventilated | -72
debridement of burns | -72
Total Body Surface Area affected by burns 61% | -72
retrieved to tertiary Paediatric Intensive Care Unit | -72
donor sites harvested | -48
burns debrided | -48
significant blood loss | -48
no grafting completed | -48
Split Skin Graft | -42
posterior torso | -42
buttocks | -42
posterior upper thighs | -42
right lower leg | -42
bilateral upper arms | -42
prone position | -42
minimal movement and repositioning | -42
septic | -30
systemic inflammatory response | -30
respiratory deterioration | -30
difficult to ventilate | -30
multifocal regions of atelectasis change | -30
no spontaneous cough | -30
increasing ventilator requirements | -30
raised peak inspiratory pressures | -30
retained secretions | -30
hemodynamic instability | -30
episodes of hypotension | -30
fluid resuscitation | -30
inotropes | -30
repositioning using bed tilt | -24
manual hyperinflation | -24
saline lavage | -24
suction | -24
passive mobility of unaffected joints | -24
limited effectiveness | -24
secretions remained difficult to access | -24
palpable secretions persisting | -24
MetaNeb treatment implemented | 0
consultation with LCCH PICU Medical Consultants | 0
consultation with USA centres | 0
MetaNeb attached to oxygen source | 0
open-ended bagging circuit | 0
Continuous High Frequency Oscillation mode | 0
occlusion ring placed in circuit | 0
inline nebuliser | 0
pressure maintained | 0
variable volume breaths delivered | 0
secretion mobilization evaluated | 0
manual Hyperinflation with expiratory flow bias | 0
suction via ETT | 0
cycle of treatment repeated | 0
sputum volume and quality measured | 0
CXR measured | 0
PIP values measured | 0
vital signs monitored | 0
blood pressure monitored | 0
transient decrease in MAP | 12
recovery without intervention | 12
resolution of focal changes on CXR | 96
reduction in secretions load | 96
reduction in PIP | 96
extubated without incident | 96
trial of MetaNeb via mouthpiece | 120
poorly tolerated | 120
discontinued due to behavioural issues | 120
lip pain and swelling | 120
inhibited lip seal | 120
skin grafting | 192
required intubation | 192
ventilation and immobility | 192
MetaNeb utilized | 192
optimization of secretion clearance | 192
decrease risk of retained secretions | 192
decrease risk of lung infection | 192
no respiratory deterioration | 240
successful extubation | 240