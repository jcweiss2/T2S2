62 years old | 0
male | 0
admitted to the intensive care unit | 0
septic shock | -24
transrectal ultrasound-guided prostate biopsy | -24
elevated prostate-specific antigen | -24
urosepsis | -24
extended spectrum beta lactamase Escherichia coli | -24
pyelonephritis | -24
phenylephrine | -24
vasopressin | -24
norepinephrine | -24
hypoxemic respiratory failure | -24
shock liver | -24
acute renal failure | -24
acalculous cholecystitis | -24
transferred to the medicine ward | 288
bilateral upper extremities distal pressor-induced ischemia | -288
bilateral lower extremities distal pressor-induced ischemia | -288
gangrene | -288
topical nitroglycerin | -216
hyperbaric oxygen therapy | 24
bilateral amputations of all fingers | -240
bilateral below the knee amputations consideration | -240
bilateral transmetatarsal amputations | -192
necrotic calcanei removal | -192
soft tissues removal | -192
Integra Bilayer Matrix Wound Dressing | -192
debridement | -192
intravenous antibiotics | -192
bilayered bovine collagen | -192
porcine xenografts | -192
bilateral free flap planning | 1092
anterior tibial arteries patent | 1092
peroneal arteries patent | 1092
sensate anterolateral thigh flap left foot | 1092
end-to-side anastomosis posterior tibial artery | 1092
end-to-end venous anastomosis saphenous vein | 1092
deep vena comitantes | 1092
neurotization lateral femoral cutaneous nerve | 1092
split-thickness skin graft left thigh | 1092
neurotized ALT flap right foot | 1320
end-to-side anastomosis posterior tibial artery | 1320
2-vein anastomosis | 1320
coaptation lateral circumflex femoral nerve | 1320
non-weight-bearing | 1344
ankle foot orthoses | 1344
custom braces | 1344
intensive physical therapy | 1680
protective sensation bilateral heels | 1680
ambulatory | 2208
ExoSym prosthesis | 2208
retained sensation bilateral free flaps | 2208
functionally ambulatory | 2208
