62 years old | 0
    woman | 0
    presented | 0
    sudden onset shortness of breath at rest | -168
    hemoptysis | -168
    intermittent yellow sclera | -720
    heavy alcohol consumption | 0
    migrated from Mexico more than 30 years ago | 0
    no contact with known tuberculosis case | 0
    illegal alien immigrant status | 0
    limited access to health care | 0
    no regular follow-ups with primary care physicians | 0
    tachypneic | 0
    tachycardiac | 0
    significant respiratory distress | 0
    nonrebreather mask | 0
    broad-spectrum antibiotic therapy | 0
    transferred to progressive care unit | 0
    bilevel positive airway pressure | 0
    scleral icterus | 0
    dried blood on lips and chin | 0
    diffuse crackles over bilateral lower lung fields | 0
    bilateral lower extremity pitting edema | 0
    white blood cell count 25.7 k/mm3 | 0
    hemoglobin 10.1 g/dL | 0
    platelet count 71,000 k/mm3 | 0
    albumin 2.9 g/dL | 0
    alkaline phosphatase 172 IU/L | 0
    aspartate aminotransferase 133 IU/L | 0
    alanine aminotransferase 32 IU/L | 0
    bilirubin 12.4 mg/dL |$|0
    lactate 2.2 mmol/L | 0
    BNP 886 pg/mL | 0
    high-sensitivity troponin 449 pg/mL | 0
    D-Dimer 29,578 ng/mL | 0
    fibrinogen 183 mg/dL | 0
    INR 1.8 | 0
    PT 20.9 sec | 0
    chest x-ray bilateral multifocal patchy opacities | 0
    CT chest extensive patchy parenchymal airspace opacities | 0
    CT abdomen diffusely heterogeneous enhancement and nodularity of liver | 0
    liver cirrhosis | 0
    severe respiratory acidosis | 0
    pH 7.24 | 0
    pCO2 68.9 | 0
    intubation | 0
    transferred to ICU | 0
    IV steroids | 0
    bronchoalveolar lavage | 0
    erythematous airways | 0
    bloody lavage return | 0
    alveolar hemorrhage | 0
    benign respiratory epithelium | 0
    reactive changes | 0
    acute inflammation | 0
    macrophages | 0
    red blood cells | 0
    negative acid-fast stain | 0
    negative cultures | 0
    negative Pneumocystis jiroveci smear | 0
    negative autoimmune disease testing | 0
    normal IgG and IgM cardiolipin antibodies | 0
    normal Beta-2-Glycoprotein IgG and IgM antibodies | 0
    negative ANA | 0
    negative P$ANCA and C$ANCA | 0
    negative rheumatoid factor | 0
    negative anti-glomerular basement membrane antibody | 0
    negative HIV-1/2 antibodies | 0
    negative HIV-1 antigen | 0
    negative Histoplasma galactomannan urine antigen | 0
    negative Legionella urinary antigen | 0
    negative pneumococcal urinary antigen | 0
    negative Epstein-Barr DNA PCR | 0
    negative hepatitis viral panel | 0
    negative Blastomyces dermatitidis antibodies | 0
    negative Aspergillus galactomannan antigen | 0
    negative Mycoplasma | 0
    negative West Nile virus | 0
    negative cytomegalovirus | 0
    negative dengue virus serum IgM and IgG antibodies | 0
    negative blood cultures | 0
    negative urine cultures | 0
    negative bronchial brushing cultures | 0
    negative fungal cultures | 0
    respiratory viral panel positive for human metapneumovirus | 0
    COVID-19 testing denied | 0
    no recent travels | 0
    no sick contacts | 0
    no community transmission suspected | 0
    started on vasopressors | 96
    prone position | 192
    worsening hypoxia | 192
    hemodialysis | 216
    severe acute kidney injury | 216
    creatinine 4.83 mg/dL | 216
    acidosis pH 7.21 | 216
    disseminated intravascular coagulation | 264
    platelet count 19 k/mm3 | 264
    D-Dimer 36,469 ng/mL | 264
    fibrinogen 91 mg/dL | 264
    CT head scattered small bilateral subarachnoid hemorrhages | 264
    multi-organ failure | 264
    cardiac arrest | 264
    death | 264
    