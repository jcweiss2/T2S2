57 years old | 0
male | 0
industrial accident | -15840
C2 vertebral body fracture | -15840
high cervical SCI at C3 level | -15840
no key muscle activity in all extremities | -15840
last intact sensory level C3 dermatome | -15840
deep anal pressure | -15840
no voluntary anal contraction | -15840
classified as C3 AIS B | -15840
pulmonary function tested | -15840
tidal volume 220 mL | -15840
vital capacity 800 mL | -15840
peak cough flow 130 L/min | -15840
continuous hypercapnia | -15840
PaCO2 over 45 mmHg | -15840
diaphragm fluoroscopy | -15840
decreased diaphragm apex length | -15840
portable ventilator applied | -15840
volume controlled assisted ventilation mode | -15840
respiratory function improved | -15840
pulmonary rehabilitation techniques | -15840
air stacking exercise | -15840
sputum expectoration | -15840
mechanical insufflation-exsufflation | -15840
accessory respiratory muscle training | -15840
readmitted to intensive care unit | 0
septic shock | 0
urinary tract infection | 0
tracheostomy performed | 0
pulmonary rehabilitation program | 0
tracheostomy tube removed | 0
total weaning not achieved | 0
respiratory insufficiency | 0
concomitant sleep apnea | 0
aging | 0
intermittent NIV applied | 0
pressure support ventilation mode | 0
nasal mask used | 0
mouth opening during sleep | 0
full face mask applied | 0
oral air leak reduced | 0
inability to take off mask | 0
communication limitation | 0
anxiety | 0
novel alarm system designed | 0
microcontroller board used | 0
sound generator | 0
pressure transducer | 0
endotracheal tube | 0
programmed with open-source software | 0
neck rotation motion | 0
pressure transducer sensor | 0
pressure exceeded 10 cm H2O | 0
single beep sound | 0
loud alarm sound | 0
adapted to full face mask | 0
discharged home | 24
no complications | 24
