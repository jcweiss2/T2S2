33 years old | 0
male | 0
abdominal pain | -672
abdominal distension | -672
bowel obstruction | -672
enterolysis | -672
omentum majus biopsy | -672
relapse of abdominal pain | -336
exploratory laparotomy | -336
bypass operation | -336
intermittent fever | -168
cachexia | -168
severe intra-abdominal infection | -168
hypoalbuminemia | -168
hydrothorax | -168
poor incisions healing | -168
suspected fistula | -168
intestinal juice flowing from the incision | -168
admitted to the hospital | 0
intermittent high fever | 0
cachexia | 0
anti-infection therapy | 0
acid suppression therapy | 0
digestive juices secretion suppression therapy | 0
total parenteral nutrition | 0
double-pipe drainage | 0
open abdomen | 0
enteroatmospheric fistula | 0
high-resolution computed tomography | 0
contrast-mediated fistula angiography | 0
fistula stent implantation | 216
implantation of fistula stent | 216
contrast-mediated fistula angiography after implantation | 216
restored enteral nutrition | 220
nasal feeding | 220
skin grafting | 504
follow-up | 720
definitive intestinal anastomosis | 720
abdominal closure | 720
fistula stent removal | 720