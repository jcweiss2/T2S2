50 years old | 0
male | 0
admitted to the hospital | 0
perianal swelling | -144
anal pain | -144
discomfort | -144
perianal abscess | -48
incision and drainage | -48
high fever | -24
scrotal swelling | -24
purulence | -24
wound discharge | -24
flatulence | -24
body temperature 38.2 °C | 0
respiratory rate 21 breaths/min | 0
heart rate 81 beats/min | 0
blood pressure 105/69 mmHg | 0
dysuresia | 0
perianal necrotizing fasciitis | 0
perineal necrotizing fasciitis | 0
cryptoglandular infection | 0
inadequate drainage | 0
multiple incisions | 0
thread-dragging therapy | 0
urethra catheter surgery | 0
spinal anesthesia | 0
lithotomy position | 0
anal gland defect | 0
internal opening | 0
necrotic tissue removal | 0
rubber catheters | 0
loose setons | 0
fourth-generation cephalosporin | 0
metronidazole | 0
human blood albumin | 0
vitamins | 0
lipids | 0
nutrition support | 0
daily laboratory examination | 0
wound cleaning | 0
wound dressing | 0
necrotic tissue trimming | 0
hydrogen peroxide | 0
oxygenate | 0
CT scan | 0
urine retention | 0
lymph nodes | 0
Proteus mirabilis | 0
surgical area rinsing | 24
necrotic perineal skin removal | 72
final drainage incision | 72
local anesthesia | 72
perianal magnetic resonance imaging | 168
laboratory examinations | 168
antibiotic treatment stopped | 168
nutrition support continued | 168
daily dressing changes | 168
discharged | 336
follow-up | 504
anorectal manometry | 1008
perianal morphology retained | 1008
function recovered | 1008
satisfied with treatment | 1008