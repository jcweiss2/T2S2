backache | 0
calculi in both kidneys associated with ureteral calculi | 0
admitted | 0
HLL combined with double J catheterization | 0
purulent urine | 0.5
severe fever | 0.5
chill | 0.5
low blood pressure | 0.5
empiric anti-infection drugs | 0.5
fluid resuscitation | 0.5
vasoactive agent | 0.5
Hydrocortisone sodium succinate hormone | 0.5
anuric | 48
ARDS | 48
invasive ventilatory support with endotracheal intubation | 48
CRRT | 48
transferred to ICU | 48
sedated state | 48
cold, clammy extremities | 48
loud bubbling sound in the lung | 48
arterial blood gas analysis | 48
cardiac function detected through the chest wall | 48
diffuse dysfunction | 48
severe functional damage in the left ventricle | 48
LVEF 20.3% | 48
normal function in the right ventricle | 48
sinus tachycardia | 48
broad ST depression | 48
elevated troponin I | 48
elevated amino-terminal brain natriuretic peptide precursor | 48
elevated creatinine | 48
anuria | 48
multiple organ function failure | 48
VA-ECMO treatment | 48
ECMO venous leading-out end used a 20F catheter | 48
arterial leading-in end used a 17F catheter | 48
No. 6 arterial catheter | 48
ECMO ran normally | 48
Norepinephrine stopped | 48.5
Epinephrine stopped | 48.5
CRRT performed | 49
Imipenem and Cilastatin sodium combined with Vancomycin | 49
lactic acid level declined | 51
vasoactive drugs completely stopped | 58
arterial blood lactate level normal | 60
extended-spectrum β-lactamase-positive Escherichia coli | 72
inflammatory indices diminished | 72
anti-infection regimen continued | 72
minimum serum trough concentration of Vancomycin monitored | 72
LVEF 35% | 120
black and necrotic skin | 120
weaned from ECMO therapy | 144
renal function scaled as acute kidney injury grade 3 | 144
CRRT discontinued | 144
urinating | 144
vascular ultrasonography | 168
computed tomography angiography | 168
vascular surgery consultation | 168
necrotic tissues amputated | 168
spontaneous breathing | 120
trachea opened | 240
anti-infection combination replaced | 240
bedside physical rehabilitation | 240
weaned from ventilator | 480
tracheotomy tube sealed | 600
discharged | 768
intermittent hemodialysis | 768
follow-up | 1056