62 years old | 0
female | 0
aortobifemoral bypass | -6720
abdominal aortic aneurysm | -6720
coronary artery stenting | -240
unstable angina | -240
fatigue | -72
myalgia | -72
left flank pain | -72
left flank pain irradiating to the left thigh | -72
fever | 0
urinary symptoms | 0
severe leukocytosis | 0
elevated CRP | 0
altered liver function test | 0
positive urinalysis | 0
leukocyturia | 0
microscopic hematuria | 0
bacteriuria | 0
CT-urography | 0
left retroperitoneal hemato-urinoma | 0
ureteral rupture | 0
urinary extravasation | 0
renal pelvis and calyceal blood clots | 0
medical and supportive treatment | 0
intravenous hydration | 0
antibiotics | 0
analgesics | 0
endoscopic drainage | 0
JJ stent insertion | 0
Foley urinary catheter | 0
urine culture | 0
multi-sensitive Escherichia Coli | 0
discharged home | 240
Foley catheter removal | 240
septic shock | 336
intensive care unit admission | 336
CT-guided left 8F nephrostomy | 336
left 10F percutaneous drain | 336
fungal infection | 336
Candida Kefyr | 336
persistent ureteral fistula | 504
laparoscopic nephrectomy | 1440
subtotal ureterectomy | 1440
necrotic and inflamed ureter | 1440
stone extraction | 1440