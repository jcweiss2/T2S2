45 years old | 0
    male | 0
    presented to the Emergency Department | 0
    epigastric pain | -72
    no diarrhea | 0
    no fever | 0
    no history of travel | 0
    no sick contact | 0
    unremarkable systemic history | 0
    temperature of 36.2°C | 0
    respiratory rate of 16 per minute | 0
    blood pressure of 167/90 mm Hg | 0
    heart rate of 62 beats per minute | 0
    normal oxygen saturation | 0
    abdominal tenderness in the epigastric area | 0
    no guarding | 0
    no rebound tenderness | 0
    normal per rectal examination | 0
    no melena | 0
    normal chest exam | 0
    normal heart exam | 0
    elevated serum creatinine | 0
    elevated blood urea | 0
    urine output 600 mL per day | 0
    no urgent dialysis indication | 0
    unremarkable abdominal CT scan | 0
    unremarkable chest X-ray | 0
    severe abdominal pain | 0
    fentanyl | 0
    paracetamol | 0
    abdominal pain persisted during days 1–3 | 0
    high serum creatinine | 0
    fever of 38.5°C | 72
    non-productive cough | 72
    dyspnea with minimal exertion | 72
    lymphopenia | 72
    COVID-19 suspected | 72
    airborne isolation | 72
    nasopharyngeal swab RT-PCR positive | 72
    oropharyngeal swab RT-PCR positive | 72
    respiratory status worsened | 168
    wheezes | 168
    temperature of 39.3°C | 168
    respiratory rate of 33 per minute | 168
    heart rate of 115 beats per minute | 168
    required 5L oxygen | 168
    oxygen saturation 94% | 168
    chest X-ray bilateral infiltrates | 168
    lymphopenia | 168
    elevated CRP | 168
    elevated liver enzymes | 168
    elevated urea | 168
    elevated creatinine | 168
    desaturated on 15L oxygen | 168
    shifted to ICU | 168
    intubated | 168
    hydroxychloroquine | 168
    azithromycin | 168
    tocilizumab | 168
    methylprednisolone | 168
    respiratory symptoms improved | 216
    abdominal pain improved | 216
    extubated | 216
    discharged | 840
    hypertension diagnosed | 0
    chronic kidney disease | 0
    acute kidney injury | 0
    bilateral increased renal parenchymal echotexture | 0
    normal size kidneys | 0
    dehydration | 0
    improvement with hydration | 0
    acute respiratory distress syndrome | 168
    COVID-19 diagnosis | 72
    ARDS precipitated by COVID-19 | 168
    surgical abdomen excluded | 0
    acute pancreatitis excluded | 0
    normal serum lipase | 0
    normal serum amylase | 0
    negative CT for pancreatitis | 0
    normal chest X-ray on day 1 | 0
    bilateral lung infiltrates on day 8 | 168
    elevated D-dimer | 168
    elevated ferritin | 168
    no further complications | 840
    hospital stay 35 days | 840

    45 years old | 0
    male | 0
    presented to the Emergency Department | 0
    epigastric pain | -72
    no diarrhea | 0
    no fever | 0
    no history of travel | 0
    no sick contact | 0
    unremarkable systemic history | 0
    temperature of 36.2°C | 0
    respiratory rate of 16 per minute | 0
    blood pressure of 167/90 mm Hg | 0
    heart rate of 62 beats per minute | 0
    normal oxygen saturation | 0
    abdominal tenderness in the epigastric area | 0
    no guarding | 0
    no rebound tenderness | 0
    normal per rectal examination | 0
    no melena | 0
    normal chest exam | 0
    normal heart exam | 0
    elevated serum creatinine | 0
    elevated blood urea | 0
    urine output 600 mL per day | 0
    no urgent dialysis indication | 0
    unremarkable abdominal CT scan | 0
    unremarkable chest X-ray | 0
    severe abdominal pain | 0
    fentanyl | 0
    paracetamol | 0
    abdominal pain persisted during days 1–3 | 0
    high serum creatinine | 0
    fever of 38.5°C | 72
    non-productive cough | 72
    dyspnea with minimal exertion | 72
    lymphopenia | 72
    COVID-19 suspected | 72
    airborne isolation | 72
    nasopharyngeal swab RT-PCR positive | 72
    oropharyngeal swab RT-PCR positive | 72
    respiratory status worsened | 168
    wheezes | 168
    temperature of 39.3°C | 168
    respiratory rate of 33 per minute | 168
    heart rate of 115 beats per minute | 168
    required 5L oxygen | 168
    oxygen saturation 94% | 168
    chest X-ray bilateral infiltrates | 168
    lymphopenia | 168
    elevated CRP | 168
    elevated liver enzymes | 168
    elevated urea | 168
    elevated creatinine | 168
    desaturated on 15L oxygen | 168
    shifted to ICU | 168
    intubated | 168
    hydroxychloroquine | 168
    azithromycin | 168
    tocilizumab | 168
    methylprednisolone | 168
    respiratory symptoms improved | 216
    abdominal pain improved | 216
    extubated | 216
    discharged | 840
    hypertension diagnosed | 0
    chronic kidney disease | 0
    acute kidney injury | 0
    bilateral increased renal parenchymal echotexture | 0
    normal size kidneys | 0
    dehydration | 0
    improvement with hydration | 0
    acute respiratory distress syndrome | 168
    COVID-19 diagnosis | 72
    ARDS precipitated by COVID-19 | 168
    surgical abdomen excluded | 0
    acute pancreatitis excluded | 0
    normal serum lipase | 0
    normal serum amylase | 0
    negative CT for pancreatitis | 0
    normal chest X-ray on day 1 | 0
    bilateral lung infiltrates on day 8 | 168
    elevated D-dimer | 168
    elevated ferritin | 168
    no further complications | 840
    hospital stay 35 days | 840