53 years old | 0
male | 0
admitted to the emergency department | 0
mild COVID-19 | -240
severe and sharp abdominal pain | -48
abdominal pain located in the epigastrium | -48
fever | -48
arterial hypertension | 0
dyslipidemia | 0
previous myocardial infarction | -0 
coronary bypass surgery | -0 
febrile | 0
stable patient | 0
blood pressure 125/82 mmHg | 0
hazard ratio 89 bpm | 0
cardiopulmonary auscultation was normal | 0
abdomen was non-distended | 0
tender mass in the epigastrium | 0
localized guarding | 0
hypoactive bowel sounds | 0
no abdominal hernias | 0
normal white blood cell count | 0
hemoglobin level of 13.80 g/dl | 0
C-reactive protein level of 22.10 mg/dl | 0
d-dimer level of 0.94 μg/ml | 0
normal hepatobiliopancreatic, cardiac and renal biochemical parameters | 0
normal urinalysis | 0
normal arterial-blood gas test | 0
ultrasonography was not performed | 0
computed tomography scan with intravenous contrast of the abdomen | 0
inflammatory signs and localized free peritoneal fluid | 0
residual ground-glass opacities related to COVID-19 | 0
cholecystitis was ruled out | 0
pancreatitis was ruled out | 0
perforation of hollow viscus was ruled out | 0
diagnostic and potentially therapeutic exploratory laparotomy | 0
suppurative Meckel’s diverticulitis | 0
local abscess | 0
drainage | 0
segmental ileal resection with primary anastomosis | 0
inflammatory markers were responding positively to intravenous antibiotics | 24
no further rises in temperature | 24
no complications | 24
discharged on postoperative Day 6 | 144
anatomopathological examination | 144
small bowel with active inflammation | 144
gangrenous Meckel’s diverticulum | 144