75 years old | 0
male | 0
diabetes mellitus | 0
hypertension | 0
admitted to the Department of Urology | 0
left flank pain | 0
dysuria | 0
high fever | 0
increased BUN | 0
increased creatinine | 0
glycosuria | 0
albuminuria | 0
leukocyturia | 0
Candida albicans infection | 0
fluconazole treatment | 0
meropenem treatment | 0
multiple bilateral kidney stones | 0
left early hydronephrosis | 0
persistent oliguria | 0
left pyelostomy | 72
transferred to ICU | 72
septic shock | 72
improved renal function | 168
readmitted to urology department | 168
double J ureteral stent placed | 168
stent removed | 1344
discharged home | 1344
sensory obtundation | -72
blurred speech | -72
weakness in the right arm and leg | -72
stuporous | 0
right hemiparesis | 0
sensory-motor aphasia | 0
increased ESR | 0
monocytosis | 0
left parietal epidural mass | 0
midline shift | 0
leptomeningeal enhancement | 0
diagnosis of epidural abscess | 0
progression of hemiparesis to hemiplegia | 0
coma | 0
left anisocoria | 0
emergency surgery | 0
fronto-temporal-parietal craniotomy | 0
mass involving dura mater | 0
durotomy | 0
en bloc removal | 0
bone unaffected | 0
duroplasty | 0
bone repositioned | 0
postoperative course uneventful | 120
ICU stay | 120
conscious | 120
aphasic | 120
right hemiparesis | 120
improved symptoms | 120
Candida albicans hyphae | 0
amphotericin B treatment | 120
meropenem treatment | 120
midline re-alignment | 336
subdural hygroma | 336
discharged to rehabilitation | 336
high fever | 3360
impaired consciousness | 3360
aphasia | 3360
subcutaneous collection | 3360
skin reddening | 3360
tenderness | 3360
subcutaneous empyema | 3360
epidural empyema | 3360
purulent collection | 3360
eroded bone | 3360
scar tissue removal | 3360
ceftriaxone treatment | 3360
teicoplanin treatment | 3360
no bacterial or fungal growth | 6720
therapy interrupted | 6720
discharged to rehabilitation | 6720
contrast enhanced MRI negative | 8064
titanium cranioplasty | 8064
discharged home | 8064
no residual deficits | 8064
no complications | 8064
