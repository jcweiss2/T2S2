17 years old | 0
    female | 0
    fever | -264
    altered behavior | -264
    abnormal body movement | -264
    altered sensorium | -264
    agitation | -264
    suspiciousness | -264
    aggression | -264
    restlessness | -264
    disturbed sleep | -264
    violence with family members | -264
    focal abnormal movement | -264
    generalized abnormal movement | -264
    up rolling of eyes | -264
    clenching of teeth | -264
    clenching of the fist | -264
    tongue biting | -264
    altered level of consciousness | -264
    olanzapine 5 mg | -264
    phenytoin 900 mg | -264
    temperature of 101°F | 0
    blood pressure of 130/70 mmHg | 0
    tachycardia | 0
    heart rate 117 beats/min | 0
    tachypnea | 0
    respiratory rate 20 breaths/min | 0
    oxygen saturation 92% | 0
    Glasgow Coma Scale score 8 | 0
    Antibody Prevalence in Epilepsy and Encephalopathy score 7 | 0
    absence of nuchal rigidity | 0
    bilaterally mute plantar reflex | 0
    cognitive function not assessed | 0
    lumbar puncture | 0
    intravenous fluids | 0
    anticonvulsants | 0
    antibiotics | 0
    transfer to ICU | 0
    CT scan head | 0
    MRI brain | 0
    CT scan abdomen and pelvis | 0
    CSF lymphocytic pleocytosis | 0
    normal CSF protein | 0
    normal CSF glucose | 0
    RT-PCR HSV-1 negative | 0
    RT-PCR HSV-2 negative | 0
    RT-PCR Mycobacterium tuberculosis negative | 0
    autoimmune encephalitis panel | 0
    anti-NMDA receptor antibodies positive | 0
    intravenous methylprednisolone 1 g per day | 0
    intravenous immunoglobulins 16 g per day | 0
    ventilator-associated pneumonia | 0
    septic shock | 0
    unresponsive to vasopressor therapy | 0
    intractable cardiac failure | 0
    death | 0
    