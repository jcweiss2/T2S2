24 years old| 0
male | 0
admitted to the hospital | 0
fever | -72
cough | -72
fatigue | -72
blood in nasopharynx | 0
no oral injury | 0
no urinary incontinence | 0
no bowel incontinence | 0
no neck stiffness | 0
vomiting 500 mL coffee ground emesis | 0
hematemesis | 0
oxygen saturation 99% | 0
blood pressure 126/84 mmHg | 0
temperature 39.4°C | 0
deteriorated consciousness | 0
intubation | 0
normal lung parenchyma | 0
severe deranged liver function | 0
SARS-CoV-2 positive | 0
severe disease | 0
chloroquine | 0
azithromycin | 0
oseltamivir | 0
tocilizumab | 0
acetylcysteine infusion | 0
lactulose | 0
vitamin K | 0
rifaximin | 0
intravenous pantoprazole | 0
4-factor prothrombin complex concentrate | 0
fresh frozen plasma | 0
fibrinogen | 0
sustained low-efficiency dialysis | 0
no intracranial hemorrhage | 0
normal brain parenchyma | 0
no hydrocephalus | 0
no midline shift | 0
no mass effect | 0
normal liver size | 0
coarse parenchymal echotexture | 0
no liver foci | 0
patent common bile duct | 0
normal spleen size | 0
homogeneous spleen echotexture |-
no spleen focal lesions | 0
normal kidney size | 0
no kidney calculus | 0
no hydronephrosis | 0
fluctuating temperature | 0
ventilatory settings CMV | 0
PEEP 5 cm H2O | 0
FiO2 25% | 0
oxygen saturation 99-100% | 0
disseminated intravascular coagulation | 168
bleeding from IV site | 168
bleeding from endotracheal tube | 168
ICU admission | 0
multiorgan failure | 240
acute liver failure | 240
acute renal failure | 240
death | 240
hepatitis B infection | 0
coagulopathy | 0
high INR | 0
low platelets | 0
low fibrinogen | 0
high d-dimer | 0
elevated liver enzymes | 0
H score 172 | 0
hemophagocytic syndrome risk | 0
cytokine storm | 0
immunosuppression | 0
hepatitis B viral replication | 0
hypothermia | 0
poor neurological outcome | 0
inverse neutrophil to lymphocyte ratio | 240
