Here is the table of events and timestamps:

31 years old | 0
female | 0
non-smoking | 0
Caucasian | 0
no past medical history | 0
sudden-onset severe headache | -5
left arm numbness | -5
cranial computed tomography (CT) scan | -5
grade 2 (Hunt and Hess scale) SAH | -5
admitted to the neurosurgical ward | -5
digital subtraction angiography (DSA) | -5
ruptured right middle cerebral artery aneurysm | -5
percutaneous endovascular coil embolization | -5
fever | -61
chills | -61
constant abdominal pain | -61
purulent uterine discharge | -61
denies urinary or respiratory symptoms | -61
sepsis | -57
septic shock | -57
transferred to the intensive care unit | -57
body temperature 38.3°C | -57
invasive blood pressure 90/65 mmHg | -57
heart rate 135/min | -57
arterial oxygen saturation 82% | -57
mild disorientation | -57
slower capillary refill | -57
coarse rales | -57
sequential organ failure assessment (SOFA) score 4 | -57
hemoglobin 6.8 g/dL | -57
d-dimers 4.58 μg/mL | -57
C-reactive protein 322 mg/L | -57
fibrinogen concentration 6.4 mL | -57
blood culture E. coli | -57
chest radiography pulmonary nodules | -57
CT of the thorax pulmonary nodules | -57
transvaginal ultrasound enlarged uterus | -57
abdominal magnetic resonance imaging (MRI) enlarged heterogenous myometrial mass | -57
splenic metastatic lesion | -57
serum β-human chorionic gonadotrophin (β-hCG) 232,085 mUI/mL | -57
suction evacuation and curettage | -57
choriocarcinoma diagnosis | -57
International Federation of Gynecology and Obstetrics (FIGO) modified WHO prognostic scoring system for gestational trophoblastic disease (GTN) | -57
total score 12 | -57
diagnosed with metastatic choriocarcinoma at high risk | -57
low-dose etoposide (100 mg/m2) in combination with cisplatin (20 mg/m2) | -57
EMA/CO regimen | -50
etoposide, methotrexate, and actinomycin D, alternating on a weekly basis with cyclophosphamide and vincristine | -50
completed six cycles | -50
β-hCG levels plateaued above normal | -50
MRI of the brain and 18F-fluorodeoxyglucose (FDG) positron emission tomography (PET)/CT scan | -50
decreased pulmonary nodules and a uterine mass | -50
revised FIGO score 7 | -50
therapeutic regimen changed to EP/EMA | -43
etoposide plus cisplatin on day 1, followed by etoposide, methotrexate, and actinomycin D on day 8 | -43
β-hCG normalization | -43
grade 3 neutropenia | -43
grade 2 fatigue | -43
grade 2 nausea | -43
grade 2 hair loss | -43
discharged | 24