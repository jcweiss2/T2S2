6 years old | 0
female | 0
102 cm tall | 0
17 kg | 0
admitted to the hospital | 0
chronic intestinal pseudo-obstruction | 0
gastric volvulus | -8760
congenital megacolon | -8760
gastropexy | -8760
segmental resection of the transverse colon | -8760
transverse colostomy | -365
mechanical ileus | -365
malnutrition | -365
electrolyte imbalance | -365
total parenteral nutrition | -365
abdominal distension | -120
malfunctioning colostomy | -120
colostomy function normalized | -118
conservative medical care | -118
scheduled for multivisceral organ transplantation | 0
multivisceral organ transplantation | 0
liver transplantation | 0
spleen transplantation | 0
stomach transplantation | 0
duodenum transplantation | 0
small bowel transplantation | 0
colon transplantation | 0
pancreas transplantation | 0
cadaveric donor | 0
brain death | -672
medulloblastoma | -672
increased intracranial pressure | -672
histidine-tryptophan-ketoglutarate solution | 0
ischemic time | 0
intraoperative gross finding | 0
no significant abnormality | 0
premedication | 0
blood pressure 120/64 mmHg | 0
heart rate 120 beats/min | 0
oxygen saturation 100% | 0
hemoglobin 9.4 g/dl | 0
Na+ 142 mmol/L | 0
K+ 3.7 mmol/L | 0
creatinine 0.34 mg/dl | 0
AST 43 IU/L | 0
ALT 35 IU/L | 0
total bilirubin 0.5 mg/dl | 0
albumin 4.4 g/dl | 0
prothrombin time 1.00 INR | 0
anesthesia induced | 0
pentothal sodium | 0
rocuronium | 0
fentanyl | 0
tracheal intubation | 0
sevoflurane | 0
continuous infusion of fentanyl | 0
continuous infusion of vecuronium | 0
brachial artery cannulation | 0
central venous catheter | 0
femoral venous pressure monitoring | 0
MAP 86 mmHg | -10
heart rate 90 bpm | -10
central venous pressure 4 mmHg | -10
femoral venous pressure 16 mmHg | -10
body temperature 36.7℃ | -10
pH 7.32 | -10
base excess -9.5 mEq/L | -10
arterial lactate concentration 5.6 mmol/L | -10
Na+ 142 mmol/L | -10
K+ 2.5 mmol/L | -10
Ca2+ 0.83 mmol/L | -10
hemoglobin 10.8 g/dl | -10
blood glucose 98 mg/dl | -10
NaHCO3 injection | 0
graft reperfusion | 0
MAP 39 mmHg | 0
femoral venous pressure 4 mmHg | 0
central venous pressure 4 mmHg | 0
epinephrine injection | 0
MAP 44 mmHg | 0
hypotension | 0
volume replacement | 0
MAP 38 mmHg | 5
arterial blood gas analysis | 5
severe metabolic acidosis | 5
pH 7.09 | 5
base excess -17.9 mEq/L | 5
arterial lactate concentration 8.5 mmol/L | 5
K+ 4.8 mmol/L | 5
Ca2+ 0.84 mmol/L | 5
glucose 114 mg/dl | 5
hemoglobin 8.5 g/dl | 5
NaHCO3 injection | 5
epinephrine injection | 5
hypothermia | 5
body temperature 33.4℃ | 5
norepinephrine infusion | 10
MAP within acceptable range | 10
body temperature 35.7℃ | 540
metabolic acidosis | 540
arterial pH 7.23 | 540
base excess -10.0 mEq/L | 540
fluid infusion | 540
balanced crystalloid solution | 540
half-normal saline | 540
5% dextrose water | 540
5% albumin | 540
packed red blood cells | 540
transferred to intensive care unit | 540
AST 2108 IU/L | 540
ALT 2351 IU/L | 540
prothrombin time 3.07-5.69 INR | 540
total bilirubin 3.4 mg/dl | 540
primary hepatic graft failure | 540
re-transplantation of the liver | 72
adult to child living donor liver transplantation | 72
vital signs stable | 72
MAP 70-80 mmHg | 72
arterial blood pH 7.49 | 72
base excess -0.1 mEq/L | 72
arterial lactate concentration 3.8 mmol/L | 72
Na+ 137 mmol/L | 72
K+ 3.3 mmol/L | 72
Ca2+ 0.97 mmol/L | 72
hemoglobin 8.2 g/dl | 72
blood glucose 170 mg/dl | 72
PRS | 72
epinephrine injection | 72
phenylephrine injection | 72
arterial lactate concentration 3.1 mmol/L | 72
pH 7.44 | 72
base excess -2.2 mEq/L | 72
Na+ 138 mmol/L | 72
K+ 2.9 mmol/L | 72
Ca2+ 1.00 mmol/L | 72
hemoglobin 6.8 g/dl | 72
packed red blood cells transfusion | 72
vital signs stable | 72
MAP 70-76 mmHg | 72
plasma hemoglobin concentration 11.9 g/dl | 168
AST 453 IU/L | 168
ALT 695 IU/L | 168
total bilirubin 3.6 mg/dl | 168
creatinine 0.6 mg/dl | 168
albumin 2.9 g/dl | 168
prothrombin time 1.74 INR | 168
AST 69 IU/L | 168
ALT 150 IU/L | 168
total bilirubin 1.4 mg/dl | 168
prothrombin time 1.07 INR | 168
feeding through gastrostomy tube | 168
discharged | 139 × 24