17 years old|0  
    male|0  
    admitted to the intensive care unit|0  
    shortness of breath|0  
    pleuritic chest pain|0  
    dry cough|-720  
    fatigue|-720  
    weight loss of 2 kg|-720  
    fever|-24  
    chills|-24  
    pleuritic chest pain (rated 3 points)|-24  
    shortness of breath development|-2  
    pleuritic chest pain aggravated|-2  
    pain radiation to shoulder and jaw|-2  
    fever (39.0℃)|0  
    blood pressure 107/70 mmHg|0  
    heart rate 110 beats/min|0  
    respiratory rate 30/min|0  
    oxygen saturation 98%|0  
    white blood cell count 20,100/mm3|0  
    neutrophils 88.4%|0  
    hemoglobin 12.6 g/dL|0  
    hematocrit 37.3%|0  
    platelet count 394,000/mm3|0  
    C-reactive protein 21.7 mg/dL|0  
    aspartate aminotransferase 84 U/L|0  
    alanine aminotransferase 177 U/L|0  
    D-dimer 2.97 mg/L|0  
    B-type natriuretic peptide 97 pg/mL|0  
    troponin I 0.04 ng/mL|0  
    HIV antibody test negative|0  
    sinus tachycardia|0  
    PR segment elevation in aVR|0  
    PR depression in other leads|0  
    cardiac silhouette enlargement|0  
    left lower lobar consolidation|0  
    pericardial effusion|0  
    pericardial enhancement|0  
    multiple necrotic lymph nodes|0  
    air in mediastinal area|0  
    broncho-lymph nodal fistula suspected|0  
    TB pericarditis presumed|0  
    lymphadenitis presumed|0  
    intravenous ceftriaxone administration|0  
    increased respiratory rate (40 breaths/min)|6  
    blood pressure drop to 90/50 mmHg|6  
    jugular venous distention|6  
    cardiac tamponade presumed|6  
    emergency pericardiocentesis|6  
    pericardial fluid drained (200 mL)|6  
    pericardial catheter placement|6  
    white blood cell count 197,840/mm3|6  
    neutrophils 98%|6  
    red blood cell count 70,000/mm3|6  
    lactate dehydrogenase 1,894 U/L|6  
    triglycerides 31 mg/dL|6  
    glucose 3 mg/dL|6  
    adenosine deaminase 91.8 U/L|6  
    TB PCR positive|24  
    AFB staining negative|24  
    Gram staining negative|24  
    isoniazid administration|24  
    rifampin administration|24  
    ethambutol administration|24  
    pyrazinamide administration|24  
    pyridoxine administration|24  
    yeast growth in culture|72  
    fluconazole administration|72  
    Candida parapsilosis identified|96  
    pericardial fluid decreased to 70 mL/day|96  
    fever persisted|96  
    gram-positive bacterium growth|96  
    vancomycin administration|96  
    ciprofloxacin administration|96  
    fever (38.1℃)|168  
    blood pressure 110/75 mmHg|168  
    heart rate 98 beats/min|168  
    respiratory rate 18/min|168  
    cardiac silhouette decreased|168  
    pneumopericardium development|168  
    pericardial wall thickening|168  
    septated pericardium|168  
    vancomycin and ciprofloxacin switched to ertapenem|168  
    Peptostreptococcus asaccharolyticus identified|216  
    Streptococcus anginosus identified|216  
    Methicillin-sensitive S. aureus identified|216  
    Prevotella oralis identified|216  
    multiple organisms from oral cavity suspected|216  
    pericardiectomy performed|240  
    pericardial irrigation|240  
    septation removal|240  
    thickened pericardium removal|240  
    acute and chronic inflammation|240  
    liquefactive necrosis|240  
    patient improvement postoperatively|240  
    TB cultures negative|720  
    discharge|720  
    oral antifungal medication|720  
    oral antibiotic medication|720  
    oral anti-TB medication|720  
    amoxicillin/clavulanic acid stopped|2160  
    fluconazole stopped|4320  
    anti-TB medication continued|4320  
    return to normal activity|4320  
    ejection fraction minimally decreased|4320  
    no cardiac relaxation abnormality|4320  
