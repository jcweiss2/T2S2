58 years old | 0
diabetic | 0
female | 0
transferred to intensive care unit | 0
emergency coronary angiogram | -48
normal coronaries | -48
treated for urinary tract infection | -72
treated for diabetic ketoacidosis | -72
pulseless ventricular tachycardia | -48
advanced cardiac life support protocol | -48
transferred for coronary angiogram | -48
raised troponin levels | -48
2D echocardiography showing left ventricular hypokinesia | -48
mechanically ventilated | 0
receiving vasopressors (norepinephrine 0.18 μg/kg/minute) | 0
easily arousable to call | 0
no neurological deficit | 0
episodes of ill-sustained ventricular tachycardia | 0
optimal oxygenation | 0
high anion gap acidosis | 0
neutrophilic leukocytosis | 0
intravenous amiodarone infusion | 0
correction of hypokalemia (2.9 mEq/dL) | 0
correction of hypomagnesemia (1.2 mEq/dL) | 0
intravenous meropenem | 0
human insulin infusion | 0
blood sugar levels between 140 mg/dL and 180 mg/dL | 0
general condition improved over the next 12 hours | 12
resolution of shock | 12
correction of acidosis | 12
restoration of normal sinus rhythm | 12
extubated | 12
computed tomography urography confirmed pyelonephritis | 12
bedside 2D echocardiography suggestive of Takotsubo cardiomyopathy | 12
apical ballooning of the left ventricle | 12
speckle tracking echocardiography suggested apical hypokinesia | 12
electrophysiologist opinion sought | 12
oral bisoprolol added | 12
oral amiodarone added | 12
shifted to step-down unit | 12
cardiac magnetic resonance imaging done | 12
ruled out structural abnormality | 12
Takotsubo cardiomyopathy appearance in mid and apical cavity | 12
shifted back to intensive care unit | 24
episodes of ill-sustained ventricular tachycardia with pulse | 24
managed with advanced cardiac life support guidelines | 24
synchronized cardioversion | 24
intravenous antiarrhythmic bolus doses of amiodarone | 24
intravenous antiarrhythmic bolus doses of lignocaine | 24
episodes of ill-sustained ventricular tachycardia continued | 24
thoracic epidural catheter inserted | 24
sympathetic blockade administered | 24
hypokalemia (3.2 mEq/dL) | 24
no further episodes of ventricular tachycardia | 72
stabilized | 72
epidural catheter removed | 72
discharged from the hospital | 216
oral propefenone | 216
oral amiodarone | 216
oral bisoprolol | 216
2D echocardiography at discharge | 216
mild apical hypokinesia | 216
mild distal interventricular septal hypokinesia | 216
ejection fraction 45% | 216
