61 years old|0
    male|0
    presented to emergency room|0
    flank pain on right side|0
    dysuria|0
    urgency|0
    frequency|0
    occasional hematuria|-72
    fever|-72
    chills|-72
    rigors|-72
    admitted for renal colic|-504
    new staghorn calculus in the kidney|-504
    managed conservatively with 7 days of oral antibiotics|-504
    40 pounds weight loss over 3 months|-2160
    drenching night sweats|-2160
    occasional low grade fevers|-2160
    multiple episodes of renal colic secondary to nephrolithiasis treated with lithotripsy|-several years ago
    30 pack year history of smoking|0
    occasional alcohol consumption|0
    no substance abuse|0
    no high risk behavior|0
    hypotension|0
    blood pressure 78/49 mmHg|0
    MAP 59 mmHg|0
    hypotension did not correct with bolus of 3 liters of 0.9% normal saline|0
    diagnosed with urinary tract infection leading to urosepsis and septic shock|0
    admitted to medical intensive care unit|0
    pressor support with norepinephrine|0
    broad spectrum antibiotic coverage with vancomycin|0
    piperacillin-tazobactam|0
    temperature 97.3°F|0
    heart rate 80/min|0
    respiratory rate 18/min|0
    SpO2 98-99% on room air|0
    averaged sized man in mild distress|0
    mild pallor|0
    no icterus|0
    no cyanosis|0
    no edema|0
    mild right costovertebral angle tenderness|0
    hemoglobin 9.2 g/dL|0
    MCV 77.6 fL|0
    leukocyte count 5.1 k/µL|0
    77% neutrophils|0
    alkaline phosphatase 212 U/L|0
    ALT 80 U/L|0
    AST 96 U/L|0
    total protein 3.6 g/dL|0
    albumin 1.5 g/dL|0
    urine dipstick positive for blood (1+)|0
    proteins (30)|0
    glucose (50)|0
    urine microscopy 109 RBC|0
    urine microscopy 12 WBC|0
    cortisol level 182.6 mg/dL|0
    two sets of blood culture done|0
    urine culture done|0
    CT scan abdomen showed numerous ill defined lesions in the liver|0
    staghorn calculus|0
    no evidence of obstruction|0
    no radiographic evidence of pyelonephritis|0
    no renal abscess|0
    received 2 days of pressor support with norepinephrine|24
    blood pressure improved to MAP over 70 mmHg|24
    intermittent episodes of hypotension|24
    frequent boluses of 1000 to 500 mL of 0.9% NS|24
    day 5 of admission|120
    increased shortness of breath|120
    hypoxic|120
    trans-thoracic echocardiogram showed normal ejection fraction|120
    normal inferior vena cava|120
    diagnosed with fluid overload secondary to frequent fluid boluses|120
    given 20 mg i.v. lasix|120
    resolution of shortness of breath|120
    intermittent episodes of hypotension|0
    colonoscopy done|0
    EGD done|0
    2 polyps|0
    tubular adenoma|0
    thick gastric folds with chronic gastritis|0
    liver biopsy planned|0
    day 9 of hospitalization|216
    declined liver biopsy|216
    deferred liver biopsy|216
    discharged|216
    4 blood cultures|0
    3 urine cultures|0
    discharged with oral levofloxacin|216
    14 days of antibiotics for complicated UTI|216
    returned to emergency room|264
    acute onset weakness|264
    fatigue|264
    single episode of fever|264
    received ibuprofen at home|264
    rectal temperature 94.1°F|264
    BP 84/49 mmHg|264
    MAP 60 mmHg|264
    breathing rate 18/min|264
    heart rate 59/min|264
    saturating 97% on room air|264
    unremarkable examination|264
    readmitted to MICU|264
    provisional diagnosis of urosepsis|264
    given vancomycin|264
    piperacillin-tazobactam|264
    blood culture done|264
    urine culture done|264
    biopsy of liver lesions showed extensive lymphocytic and histiocytic infiltrates|264
    abnormal large cells|264
    positive stains for CD15|264
    positive stains for CD30|264
    bone marrow biopsy showed residual trilineage hematopoesis|264
    40% cellularity|264
    para-trabecular infiltrates composed of large atypical cells|264
    Reed-Sternberg cells|264
    mixed inflammatory background|264
    immunohistochemical stains positive for CD15|264
    CD30|264
    negative for CD45|264
    CD3|264
    CD20|264
    bone marrow aspirate showed trilineage hematopoesis|264
    orderly maturation|264
    100 cell count granulocytes 56%|264
    monocytes 1%|264
    eosinophils 6%|264
    erythroid precursors 34%|264
    lymphocytes 2%|264
    plasma cells 1%|264
    presence of Reed-Sternberg cells|264
    diagnosis of Hodgkin lymphoma|264
    confirmed by IHC stain for CD15|264
    CD30|264
    negative IHC for CD45|264
    CD3|264
    CD20|264
    CT chest for staging|264
    no hilar lymphadenopathy|264
    started on chemotherapy|264
    doxorubicin|264
    dacarbazine|264
    vinblastine|264
    bleomycin withheld|264
    added later after pulmonary function test normal|264
    blood pressure improved to MAP over 80 mmHg after 1st cycle of chemotherapy|264
    6 month follow up|12960
    free of hypotension|12960
    free of hypothermia|12960
