24 years old | 0
male | 0
admitted to the hospital | 0
sore throat | -240
difficulty in swallowing | -240
pain and swelling on the left side of the neck | -96
severe throbbing headache | -48
vomiting | -48
restlessness | -48
bulge in the posterior pharyngeal wall | 0
uvula deviated to the right | 0
febrile | 0
tachycardic | 0
tender swelling on the left side of the neck | 0
Hb 13.3 gm% | 0
total count of 9800 cells/cumm | 0
platelet count 282,210 cells/cumm | 0
ESR 37 mm/h | 0
HIV negative | 0
left parapharyngeal abscess | 0
thrombosis of the left IJV | 0
reduced flow or stasis in left transverse and sigmoid sinuses | 0
diagnosis of Lemierre's syndrome | 0
parapharyngeal abscess drained | 0
imipenem started | 0
fondaparinux started | 0
persistent hypotension | 48
systolic pressures between 70 and 90 mmHg | 48
total count decreased to 3720 cell/cu mm | 48
platelet count dropped to 35,000/cu mm | 48
Activated partial thromboplastin time prolonged | 48
serum procalcitonin 1.4 ng/mL | 48
diagnosis of septic shock | 48
imipenem stopped | 48
vancomycin started | 48
clindamycin started | 48
metronidazole started | 48
single donor platelet units transfused | 48
central venous access obtained via the right femoral vein | 48
fondaparinux stopped | 48
noradrenaline infusion started | 48
cultures of pus and devitalized tissue grew S. aureus | 48
blood culture was negative | 48
no anaerobes isolated | 48
progressively tachypneic | 72
hypoxemic | 72
bilateral lower zone opacities on chest X-ray | 72
intubated and ventilated | 72
weaned off the inotrope | 120
weaned off the ventilator support | 120
platelet count improved to 379,000/cu mm | 120
coagulation normalized | 120
chest X-ray normalized | 120
discharged to ward | 168
oral linezolid continued for 3 weeks | 168
discharged from the hospital | 504