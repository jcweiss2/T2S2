10 years old | 0
male | 0
born by caesarean section | -720
birth weight 2100 g | -720
birth length 48 cm | -720
prominent forehead | -720
relative macrocephaly | -720
limb asymmetry | -720
5th finger clinodactyly of both hands | -720
2/3 toe syndactyly of both legs feet | -720
hypomethylation of the 11p15 region of the paternal chromosome | -504
delayed motor development | -336
walked independently in 16th month of life | -336
hepatic dysfunction | -336
increased concentration of alanine aminotransferase | -336
increased concentration of aspartate aminotransferase | -336
increased creatine kinase level | -336
diagnosis of Duchenne muscular dystrophy | -336
mutation of the maternal DMD gene located on the X chromosome | -336
exon deletion 49–50 | -336
often falling | -240
tiptoed | -240
Achilles tendon contractures | -240
Gover’s syndrome | -240
enlarged calves | -240
corticosteroids treatment | -240
prednisone | -240
deflazacort | -192
qualified for G-CSF treatment | -192
G-CSF treatment | -192
sepsis | -144
hypoglycaemia | -144
neurological symptoms | -144
glucose level of 14 mg/dl | -144
hypospadias | -144
episodes of sinus tachycardia | -72
heart murmur | -72
cardiological diagnostics | -72
propranolol | -72
growth hormone deficiency | -72
rhGH treatment | -72
dysmorphic features | -72
slightly limb asymmetry | -72
hypotonia | -72
malocclusion | -72
hypospadias | -72
pubertal status | -72
auxological examination | -72
height 115.9 cm | -72
weight 19.9 kg | -72
body mass index 14.8 kg/m2 | -72
target height 182.5 cm | -72
height velocity 4.3 cm/year | -72
glucose and insulin levels in oral glucose tolerance test | -72
IGF-1 and IGFBP-3 concentrations | -72
MRI of the hypothalamic-pituitary region | -72
transparent septum cyst | -72
rhGH treatment started | 0
improvement of auxological parameters | 12
height velocity increased | 12
level of IGF-1 increased | 12
BMI increased | 12
worsening of glucose metabolism | 12
increasing insulin resistance | 12
HbA1c elevated | 12
distance covered in 6MWT decreased | 12
abnormal, weakened gait | 12
behavioural treatment with lifestyle modification | 12
rhGH dose reduced | 12
growth 2.8 cm | 6
rhGH therapy discontinued | 18
auxological and hormonal evaluation | 18
change of height during life and rhGH treatment | 18
change of BMI during life and rhGH treatment | 18
body mass composition | 12
densitometry | 12
bone density test of the lumbar spine | 12
Z-score –2.2 | 12