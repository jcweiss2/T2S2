65 years old | 0
male | 0
diet-controlled type 2 diabetes mellitus | -8760
hyperlipidemia | -8760
stage 3 chronic kidney disease | -8760
cardiac arrest | -720
chills | -48
body aches | -48
shortness of breath | -48
cough productive of yellow sputum tinged with blood | -48
denies sick contacts | -48
denies travel | -48
heavy alcohol use | -8760
smoking | -8760
admitted to the hospital | 0
confused | 0
hypoxemic | 0
chest radiograph | 0
moderately dense consolidation in the right mid-lung | 0
treatment with azithromycin | 0
treatment with ceftriaxone | 0
intubated | 24
blood and respiratory cultures grew non-lactose fermenting Gram-negative rods | 24
meropenem | 24
levofloxacin | 24
amikacin | 24
lymphopenia | 24
persistent elevation in blood lactate | 24
worsening thrombocytopenia | 24
acute kidney injury (AKI) | 24
high oxygen requirements | 24
mechanical ventilation | 24
repeat chest radiograph | 24
progression of disease | 24
transferred to the intensive care unit (ICU) | 72
septic shock | 72
unresponsive to 3 vasopressors | 72
coarse breath sounds | 72
lower extremities and digits were cool and mottled | 72
administration of 100% oxygen | 72
saturations above 88% | 72
Acinetobacter baumannii | 72
sensitive to all antimicrobials tested | 72
therapy narrowed to cefepime | 72
repeat cultures remained negative | 72
inexorable decline | 72
persistent lactic acidosis | 72
disseminated intravascular coagulopathy (DIC) | 72
AKI necessitating hemodialysis | 72
bullae on his legs | 240
dry gangrene on his digits | 240
life support withdrawn | 264
expired | 264