54 years old | 0  
    male | 0  
    autism | 0  
    bipolar disorder | 0  
    intellectual disability | 0  
    urinary incontinence | 0  
    presented to the emergency department | 0  
    scrotal swelling | -24  
    blood pressure 131/83 | 0  
    febrile | 0  
    temperature 101.2F | 0  
    maximum temperature 103F | 0  
    tachycardic | 0  
    heart rate 111 beats/min | 0  
    respiratory rate 16 breaths/min | 0  
    saturation 100% on room air | 0  
    awake | 0  
    disheveled | 0  
    disoriented | 0  
    not following commands | 0  
    unremarkable cardiac exam | 0  
    unremarkable respiratory exam |)