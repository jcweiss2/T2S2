27 years old | 0
male | 0
admitted to the hospital | 0
car accident | -5760
neck fracture | -5760
quadriplegic | -5760
tracheostomy intubation | -5760
nasogastric tube inserted | -5760
discharge of food from the foramen of tracheostomy tube | -672
massive bleeding from the tracheostomy tube | 0
unstable vital signs | 0
blood pressure below 80/60 | 0
peripheral pulse not palpable | 0
urgent surgery | 0
general anesthesia | 0
rigid bronchoscopy | 0
tracheal stenosis | 0
tracheoesophageal fistula (TEF) | 0
bleeding stopped | 0
division and ligature of the innominate artery | 0
separation of the trachea from the divided artery | 0
repair of trachea | 0
reinforcement with strap muscle | 0
tracheostomy tube reinserted | 0
jejunostomy tube inserted | 0
vital signs stabilized | 0
neurologic examination not changed | 0
right radial pulse weaker than left radial pulse | 0
discharged from hospital | 312
admitted to the hospital again | 744
endoscopy | 744
large foramen in anterior wall of esophagus | 744
deep vein thrombosis in the left leg | 744
heparin administered | 744
colored Doppler sonography | 751
deep vein thrombosis resolved | 751
purulent discharge from the tracheostomy tube | 758
bronchiectasis and pneumonia | 758
septic shock | 772
expired | 1104