14 years old | 0
female | 0
obesity | 0
admitted to the hospital | 0
confluent and reticulated papillomatosis (CARP) | -672
minocycline 100 mg daily | -672
acute multiorgan dysfunction | 0
acute kidney injury | 0
hepatic dysfunction | 0
pneumonia | 0
shock | 0
fever | -336
lymphadenopathy | -336
facial edema | -336
diffuse exanthematous eruption | 0
pseudovesicular erythematous papules | 0
significant facial edema | 0
hyperpigmented, reticulated plaques | 0
white blood cell 65.0 | 0
eosinophil differential of 17% | 0
creatinine 1.85 | 0
aspartate aminotransferase 2650 | 0
alanine transaminase 767 | 0
alkaline Phosphatase 181 | 0
prothrombin time 25.1 | 0
partial thromboplastin time 62.1 | 0
ferritin 9259.2 | 0
lactate dehydrogenase 7326 | 0
procalcitonin 82.18 | 0
fibrin 90 | 0
erythrocyte sedimentation rate 26 | 0
elevated human herpesvirus 6 polymerase chain reaction | 0
minocycline discontinued | -336
broad-spectrum antibiotics administered | -336
broad-spectrum antibiotics discontinued | 48
high dose steroids | 48
IL-1 blockade (anakinra) | 48
IL-6 blockade (siltuximab) | 48
Janus kinase-signal transducer and activator of transcription (JAK-STAT) blockade (ruxolitinib) | 96
total plasma exchange | 72
total plasma exchange | 96
DRESS syndrome diagnosed | 0
HLH diagnosed | 0
Registry of Severe Cutaneous Adverse Reaction (RegiSCAR) score calculated | 0
patient passed away | 168
recalcitrant hypotension | 168
asystole | 168