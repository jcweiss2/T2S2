52 years old | 0
female | 0
high risk AML | -720
recurrent Clostridioides difficile infection | -720
admitted to the hospital | 0
match-unrelated donor hematopoietic stem cell transplant | 0
reduced intensity fludarabine-melphalan | 0
tacrolimus | 0
methotrexate | 0
graft-versus-host prophylaxis | 0
sepsis | 0
metabolic encephalopathy | 0
chronic diarrhea | 0
transaminitis | 0
acute kidney injury | 0
bone graft failure | 0
febrile neutropenia | 0
encephalopathy | 0
Klebsiella bacteremia | 0
J. hoylei bacteremia | -720
afebrile | 0
normotensive | 0
blood pressure 143/104 | 0
pulse 104 beats per minute | 0
respiratory rate 22 breaths per minute | 0
oxygen saturation 97% | 0
diffuse anasarca | 0
bruising throughout her extremities | 0
bleeding gums | 0
oral ulcers | 0
mucositis | 0
course bilateral breath sounds | 0
hypoactive bowel sounds | 0
no thrush | 0
PICC site clean, dry and intact | 0
peripheral line | 0
decompensation | 0
oral mucositis hemorrhage | 0
transferred to the intensive care unit | 0
airway management | 0
aerobic blood culture | -720
sheep blood agar | -720
Gram-positive | -720
coryneform | -720
MALDI-TOF MS | -720
16S ribosomal RNA gene PCR/sequencing | -720
cefepime | -192
vancomycin | -264
imipenem | 0
linezolid | 0
susceptibility results | 0
MICs | 0
follow-up blood cultures | 168
negative | 168
pancytopenia worsened | 168
repeat bone marrow biopsy | 168
severely aplastic bone marrow | 168
no signs of leukemia | 168
poor prognosis | 168
deterioration in functional status | 168
elected for comfort and hospice care | 168
died | 192
acyclovir | -720
inhaled pentamidine | -720
levofloxacin | -720
oral vancomycin | -720
fluconazole | -720
voriconazole | -720
parenteral vancomycin | -720
piperacillin-tazobactam | -720
aztreonam | -720
febrile neutropenia | -720