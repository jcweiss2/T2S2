40 years old | 0
female | 0
admitted to the hospital | 0
acute severe epigastric pain | 0
leukocytosis | 0
neutrophils 91% | 0
serum amylase 1,309 U/l | 0
total bilirubin 1.9 mg/dl | 0
direct bilirubin 0.5 mg/dl | 0
AST 126 U/l | 0
ALT 343 U/l | 0
alkaline phosphatase 104 U/l | 0
endoscopic retrograde cholangiopancreatography | 0
common bile duct sludge | 0
high-grade fever | -336
abdominal pain | -336
CT scan showed pancreatic necrosis | -336
fluid collection at the pancreatic body | -336
intravenous antibiotics | -336
EUS-guided drainage | -336
10 Fr × 7 cm double pigtail stent | -336
prophylactic antibiotics | -336
re-admitted | -168
severe abdominal pain | -168
sepsis | -168
CT scan of the upper abdomen | -168
enlargement of the pancreatic collection | -168
increased enhancement of the rim | -168
septation | -168
air inside | -168
repeat EUS-guided drainage | -168
partially clogged stent | -168
large collection with turbid content | -168
air inside | -168
punctured the abscess | -168
19-gauge needle | -168
aspirated fluid purulent | -168
culture | -168
contrast injection | -168
8.5 and 10 Fr tapered tip Teflon catheters | -168
dilatation | -168
10 Fr × 7 cm double pigtail stent | -168
two additional stents | -168
better drainage | -168
extended course of intravenous antibiotics | -168
discharged | 792
follow-up MRI | 1008
small pancreatic fluid collection | 1008