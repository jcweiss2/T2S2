45 years old | 0
male | 0
admitted to the hospital | 0
severe COVID-19 symptoms | 0
ground-glass pattern on thoracic computed tomography | 0
history of hypertension | -672
nasopharyngeal swab test concluded positive for ribonucleic acid | 0
oseltamivir | 0
hydroxychloroquine | 0
broad-spectrum antibiotics | 0
mechanical ventilation | 48
transferred to intensive care unit | 48
endotracheal intubation | 48
favipiravir | 48
rehabilitation program planned | 48
passive range of motion exercises | 48
bed positioning | 48
prone position | 48
sepsis | 72
broad-spectrum antibiotherapy continued | 72
tracheostomy | 720
mechanical ventilator | 0-1320
oxygen support | 0-1440
discharged from ICU | 1440
discharged from hospital | 1504
rehabilitation program planned | 1512
physical medicine and rehabilitation outpatient clinic | 1512
complaints of walking disability | 1512
stiffness in both hips, elbows, and shoulders | 1512
unable to stand up and move comfortably | 1512
dependent on daily living activities | 1512
physical examination | 1512
no red, warm and swollen joint | 1512
pain in elbows and hips | 1512
hard and fixed growth masses in hips | 1512
total ankylosis of both elbows | 1512
decreased range of motion in shoulders | 1512
flexion deformity in hips | 1512
difficulty in lying in prone position | 1512
normal range of motion in other joints | 1512
muscle strength could not be evaluated | 1512
X-rays revealed heterotopic ossification | 1512
increased alkaline phosphatase | 1512
normal serum calcium | 1512
chronic sensory-motor polyneuropathy | 1512
cranial magnetic resonance imaging | 1512
mild cerebral atrophy | 1512
home-based rehabilitation program | 1512
slight stretching exercises | 1512
submaximal muscle strengthening exercises | 1512
pulmonary exercises | 1512
physiotherapist supervised | 1512
written informed consent | 1512