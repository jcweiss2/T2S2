69 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
high-grade fever | -72 | 0 | Factual
pleuritic right lower chest pain | -72 | 0 | Factual
cough | -72 | 0 | Factual
elevated temperature | 0 | 0 | Factual
bibasilar crackles | 0 | 0 | Factual
lower extremity edema | 0 | 0 | Factual
grade 3 holosystolic apical murmur | 0 | 0 | Factual
mitral valve regurgitation | 0 | 0 | Factual
long-term venous access port | -672 | 0 | Factual
anemia | -672 | 0 | Factual
hemoglobin 12.1 g/dL | 0 | 0 | Factual
white blood cell count 15.1×10^3/µL | 0 | 0 | Factual
absolute neutrophil count 13.2×10^3/µL | 0 | 0 | Factual
b-type natriuretic peptide 788 pg/mL | 0 | 0 | Factual
congestive heart failure | 0 | 0 | Factual
left bundle branch pattern | 0 | 0 | Factual
Corynebacterium CDC group G bacteremia | -672 | 0 | Factual
blood cultures positive for Corynebacterium CDC group G | 0 | 0 | Factual
gram stain positive for gram positive rods | 0 | 0 | Factual
Corynebacterium CDC group G identified | 0 | 0 | Factual
moderate mitral valve regurgitation | 0 | 0 | Factual
thickened anterior mitral leaflet | 0 | 0 | Factual
vegetations | 0 | 0 | Factual
severely elevated pulmonary artery systolic pressure | 0 | 0 | Factual
bacterial IE | 0 | 0 | Factual
vancomycin treatment | 0 | 168 | Factual
clindamycin treatment | 0 | 168 | Factual
discharged | 120 | 120 | Factual
readmitted | 168 | 168 | Factual
shortness of breath | 168 | 168 | Factual
hypoxic | 168 | 168 | Factual
elevated white blood cell count | 168 | 168 | Factual
severe mitral valve regurgitation | 168 | 168 | Factual
large and mobile vegetation | 168 | 168 | Factual
mitral valve replacement | 216 | 216 | Factual
coronary artery bypass grafting | 216 | 216 | Factual
oliguric acute renal failure | 216 | 216 | Factual
respiratory failure | 216 | 216 | Factual
mechanical ventilation | 216 | 216 | Factual
vancomycin resistant enterococcus | 240 | 240 | Factual
urinary tract infection | 240 | 240 | Factual
daptomycin treatment | 240 | 504 | Factual
worsening congestive heart failure | 360 | 360 | Factual
transesophageal echocardiogram | 408 | 408 | Factual
severe mitral valve regurgitation | 408 | 408 | Factual
recurrent endocarditis | 408 | 408 | Factual
doxycycline treatment | 600 | 504 | Factual
aztreonam treatment | 600 | 504 | Factual
anidulafungin treatment | 600 | 504 | Factual
bioprosthetic mitral valve replacement | 624 | 624 | Factual
mechanical St. Jude’s prosthesis | 624 | 624 | Factual
limb ischemia | 696 | 696 | Factual
disseminated intravascular coagulation | 696 | 696 | Factual
multi-organ failure | 696 | 696 | Factual
expired | 696 | 696 | Factual