9 years old | 0
    girl | 0
    referred to the Almokala University Hospital | -48
    low-grade fever | -72
    sore throat | -72
    swelling of the neck | -24
    dysphagia | -24
    born at a rural hospital in Yemen | -262080
    received Bacillus Calmette-Guérin vaccination | 0
    received hepatitis B vaccination | 0
    no other additional vaccinations | 0
    no known previous medical problems | 0
    lived with mother | 0
    lived with father | 0
    lived with aunt | 0
    lived with cousin | 0
    history of close contact with sick patients | -48
    brother died | -48
    acute febrile illness (brother) | -48
    ill-looking | 0
    not in respiratory distress | 0
    normal color appearance | 0
    febrile (38.5°C) | 0
    tachycardia (130 bpm) | 0
    average respiratory rate (20 breaths/min) | 0
    normal blood pressure (110/70 mm Hg) | 0
    weight 22 kg (10th centile) | 0
    swelling of the right side of the neck tissue | 0
    soft | 0
    tender | 0
    without fluctuation | 0
    healthy skin overlying | 0
    inflamed pharyngotonsillar area | 0
    white patches | 0
    enlarged tonsils | 0
    lungs bilaterally clear to auscultation | 0
    hemoglobin 13.5 g/dL | 0
    white blood cell count 11,700 cells/mm3 | 0
    neutrophils 88% | 0
    lymphocytes 3% | 0
    platelet count 95,000/mm3 | 0
    blood urea nitrogen elevated (51 mg/dL) | 0
    creatinine elevated (1.0 mg/dL) | 0
    throat swab Gram stain showed gram-positive bacilli | 0
    throat swab culture showed Corynebacterium diphtheriae | 0
    troponin T level 74 ng/mL | 0
    creatine kinase-MB level 7.6 ng/mL | 0
    pro-brain natriuretic peptide 1236 ng/L | 0
    started on DAT (20,000 units intravenously) | 0
    penicillin G (200,000 U/kg/day intravenously) | 0
    ceftriaxone (100 mg/kg/day intravenously) | 0
    abdominal pain | 48
    vomiting | 48
    ultrasound showed mild ascetic fluid collection | 48
    blood urea nitrogen increased (67 mg/dL) | 48
    creatinine increased (2.2 mg/dL) | 48
    creatine kinase-MB level 66 IU/L | 48
    improper initial dose of DAT | 0
    contacted CDC | 72
    recommended redosing DAT at 80,000 units | 72
    clinical deterioration | 72
    generalized edema | 192
    hypotension | 192
    diminished urine output | 192
    declared dead | 216
    acute myocarditis | 216
    cardiogenic shock | 216
    no DAT remaining dose | 216
    
    
    