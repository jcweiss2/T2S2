74 years old | 0 | 0 
female | 0 | 0 
admitted to the hospital | 0 | 0 
low-grade fever | -48 | 0 
dry cough | -48 | 0 
shortness of breath | -48 | 0 
elective right total knee replacement | -168 | -168 
post-operative course | -168 | -168 
pain | -168 | 0 
redness | -168 | 0 
swelling | -168 | 0 
essential hypertension | 0 | 0 
obesity | 0 | 0 
myasthenia gravis | 0 | 0 
osteoarthritis | 0 | 0 
body temperature | 0 | 0 
blood pressure | 0 | 0 
pulse | 0 | 0 
respiratory rate | 0 | 0 
oxygen saturation | 0 | 0 
lung auscultation | 0 | 0 
bilateral rhonchi | 0 | 0 
rales | 0 | 0 
chest radiography | 0 | 0 
patchy air space opacity | 0 | 0 
pneumonia | 0 | 0 
rapid nucleic acid amplification test | 0 | 0 
nasopharyngeal swab | 0 | 0 
broad-spectrum antibiotics | 0 | 96 
cefepime | 0 | 96 
levofloxacin | 0 | 96 
supportive care | 0 | 0 
supplemental oxygen | 0 | 0 
mild diarrhea | 72 | 72 
generalized weakness | 72 | 72 
fatigue | 72 | 72 
intravenous immunoglobulin | 72 | 120 
mild MG exacerbation | 72 | 120 
MG crises | 72 | 120 
arterial blood gases | 0 | 0 
complete blood count | 0 | 0 
basic metabolic profile | 0 | 0 
mild absolute lymphopenia | 0 | 0 
anemia | 0 | 0 
pH | 0 | 0 
pCO2 | 0 | 0 
pO2 | 0 | 0 
bicarbonate | 0 | 0 
increasing SOB | 0 | 96 
oxygen requirements | 0 | 96 
high-flow nasal cannula | 0 | 96 
nasopharyngeal swab results | 96 | 96 
SARS-CoV-2 | 96 | 96 
hydroxychloroquine | 96 | 240 
azithromycin | 96 | 240 
zinc sulfate | 96 | 240 
oral vitamin C | 96 | 240 
blood cultures | 0 | 96 
sputum cultures | 0 | 96 
septic shock | 144 | 144 
ARDS | 144 | 144 
mechanical ventilation | 144 | 240 
norepinephrine | 144 | 192 
colchicine | 144 | 192 
cytokine storm | 144 | 192 
elevated interleukin-6 | 144 | 192 
intubation | 144 | 144 
emergent basis | 144 | 144 
pressure-regulated volume-controlled mechanical ventilation | 144 | 240 
high-dose vitamin C | 168 | 240 
clinical condition improvement | 168 | 240 
norepinephrine support | 192 | 192 
CXR improvement | 240 | 240 
spontaneous breathing trial | 240 | 240 
CPAP/PS | 240 | 240 
PEEP | 240 | 240 
PS above PEEP | 240 | 240 
fraction of inspired oxygen | 240 | 240 
ABGs | 240 | 240 
pH | 240 | 240 
pCO2 | 240 | 240 
pO2 | 240 | 240 
bicarbonate | 240 | 240 
extubation | 240 | 240 
oxygen saturation | 384 | 384 
CXR | 384 | 384 
inpatient physical rehabilitation | 240 | 384 
occupational rehabilitation | 240 | 384 
isolation room | 240 | 384 
discharge | 384 | 384 
quarantine | 384 | 398