23 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
history of methicillin-resistant Staphylococcus aureus (MRSA) impetigo | -8760 | -8760 | Factual
right tibia fracture | -8760 | -8760 | Factual
intramedullary fixation (IMN) | -8760 | -8760 | Factual
interlocking screws removed | -720 | -720 | Factual
skin irritation | -720 | -720 | Factual
pain | -720 | -720 | Factual
referred to the emergency room (ER) | -720 | -720 | Factual
redness and swelling at the surgical site | -720 | -720 | Factual
diagnosed with stitch abscess | -720 | -720 | Factual
cultures from the surgical site were positive for MRSA | -720 | -720 | Factual
prescribed an oral antibiotic treatment | -720 | -720 | Factual
discharged home | -720 | -720 | Factual
returned to the ER with a fever | -504 | -504 | Factual
right groin pain | -504 | -504 | Factual
discharged home with the diagnosis of viral infection | -504 | -504 | Factual
returned to the ER with a systemic fever | -504 | -504 | Factual
myalgia | -504 | -504 | Factual
difficult and painful ambulation | -504 | -504 | Factual
right forearm cellulitis | -504 | -504 | Factual
right sudden onset uveitis | -504 | -504 | Factual
systemic rash | -504 | -504 | Factual
right hip lymphadenopathy | -504 | -504 | Factual
increased CRP level | -504 | -504 | Factual
elevated WBC count | -504 | -504 | Factual
hepatic enzymes elevated | -504 | -504 | Factual
lactic dehydrogenase (LDH) elevated | -504 | -504 | Factual
creatine phosphokinase (CPK) elevated | -504 | -504 | Factual
radiograph of both hips in anterior-posterior view was unremarkable | -504 | -504 | Factual
advised to start the treatment with intravenous (IV) antibiotics | -504 | -504 | Factual
medical condition continued to deteriorate | -504 | 0 | Factual
positron emission tomography-computed tomography (PET-CT) scan | 0 | 0 | Factual
OIM abscess with systemic manifestations | 0 | 0 | Factual
blood cultures were positive for MRSA bacteria | 0 | 0 | Factual
hemodynamic deterioration | 0 | 0 | Factual
fulminant MRSA sepsis | 0 | 0 | Factual
admitted to the intensive care unit (ICU) | 0 | 0 | Factual
underwent ultrasound-guided drainage | 0 | 48 | Factual
no improvement | 48 | 48 | Factual
underwent a full-body CT scan | 72 | 72 | Factual
enlargement of the abscesses diameter | 72 | 72 | Factual
persistent fever | 72 | 72 | Factual
CRP level of 36 mg/dL | 72 | 72 | Factual
WBC count of 20,000 | 72 | 72 | Factual
consulting the orthopaedic team | 72 | 72 | Factual
surgical intervention was considered | 72 | 72 | Factual
combined approach of Smith-Peterson and modified Stoppa | 72 | 72 | Factual
surgery | 96 | 96 | Factual
general condition was improving | 96 | 120 | Factual
less frequent fever spikes | 96 | 120 | Factual
decrease in CRP and WBC levels | 96 | 120 | Factual
additional antibiotic treatment support for 6 weeks | 120 | 360 | Factual
almost complete recovery | 720 | 720 | Factual
able to ambulate normally without any pain or functional limitations | 720 | 720 | Factual
returned to his daily activities | 720 | 720 | Factual