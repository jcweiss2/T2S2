46 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
obesity | 0 | 0 | Factual
psoriatic arthritis | 0 | 0 | Factual
hypoparathyroidism | -7200 | 0 | Factual
hypothyroidism | -7200 | 0 | Factual
total thyroidectomy | -7200 | -7200 | Factual
multinodular goitre | -7200 | -7200 | Factual
elective sleeve gastrectomy | 0 | 0 | Factual
gastric perforations | 0 | 0 | Factual
friable mucosa | 0 | 0 | Factual
abdominal sepsis | 0 | 0 | Factual
transfer to intensive care | 96 | 96 | Factual
critically low calcium level | 96 | 96 | Factual
ionised calcium 0.78 mmol/L | 96 | 96 | Factual
continuous intravenous calcium gluconate infusion | 96 | 0 | Factual
maintenance intermittent IV calcium boluses | 96 | 0 | Factual
prolonged ICU admission | 96 | 6048 | Factual
multiple abdominal operations | 96 | 6048 | Factual
weight loss 14 kg | 96 | 6048 | Factual
endocrinology advice | 96 | 6048 | Factual
intravenous triiodothyronine | 336 | 0 | Factual
euthyroidism | 336 | 0 | Factual
high dose intravenous calcium | 336 | 0 | Factual
ionised calcium measured daily | 336 | 0 | Factual
serum phosphate level 1.07 mmol/L | 336 | 0 | Factual
intravenous calcitriol | 1008 | 1012 | Factual
limited stock and high cost | 1012 | 1012 | Factual
intramuscular cholecalciferol | 1344 | 1344 | Factual
low 1,25(OH)vitamin D3 level | 1344 | 1344 | Factual
normal renal function | 1344 | 1344 | Factual
additional intravenous calcitriol | 1824 | 0 | Factual
reduced calcium gluconate requirements | 1824 | 0 | Factual
intramuscular thyroxine | 1904 | 1904 | Factual
intravenous thyroxine | 1908 | 0 | Factual
maintenance schedule established | 1908 | 0 | Factual
discharge | 6048 | 6048 | Factual
normocalcaemia on review | 6480 | 6480 | Factual
weight 71.8 kg | 6480 | 6480 | Factual
BMI 29 kg/m2 | 6480 | 6480 | Factual