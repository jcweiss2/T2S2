66 years old | 0
female | 0
admitted to the hospital | 0
fever | 0
hypotension | 0
tachycardia | 0
elevated inflammation values | 0
leukocytes 18.8 Gpt/L | 0
CRP 405 mg/L | 0
acute renal failure | 0
creatinine 212 μmol/L | 0
glomerular filtration rate (GFR) 20 mL/min/1.73 qm | 0
leukocyturia | 0
proteinuria | 0
bacteria in urine | 0
horseshoe kidney | 0
second-degree urinary retention | 0
urosepsis | 0
stent insertion | 0
renal function restricted | 0
GFR 60 mL/min/1.73 qm | 0
inhomogeneous mass | 0
cystic parts adjacent to the right ovary | 0
contact to the right ureter | 0
contact to iliac vessels | 0
contact to bladder | 0
suspicion of infiltration of the sacrum | 0
diverticulosis | 0
no metastases on 18F-FDG-PET | 0
sarcoma suspected | 0
neoadjuvant radiotherapy | 0
tumor operation | 0
iliac vascular resection | 0
partial ureteral resection | 0
NET G2 (Ki67 10%) | 0
liver metastases | 128
refused further treatment | 128
multiple liver lesions | 160
NET G2 (Ki67 15%) | 160
somatostatin receptor expression | 160
pathologic lymph node adjacent to the head of the pancreas | 160
no tumor of the pancreas | 160
dose-reduced 177Lu–DOTATATE | 192
lanreotide | 192
disease stabilization | 192
progression | 240
everolimus | 240
NET G3 (Ki67 34%) | 240
capecitabine plus temozolomide | 272
PRRT | 304
oxaliplatin and capecitabine | 336
dose reduction | 336
discontinuation of chemotherapy | 360
molecular testing | 360
BRCA1 Mutation R691fs*10 | 360
tumor mutational burden zero | 360
microsatellite stability | 360
germline analysis | 360
Olaparib | 432
stable liver metastases | 432
upper abdominal pain | 432
PRRT with 225Ac-DOTATATE | 464
abdominal complaints disappeared | 464
Olaparib restarted | 496
restaging with 68Ga-Dotatate PET/MRI | 496
decrease in liver metastases | 496
stable large liver metastasis | 624
progression of smaller hepatic metastases | 624
TAT planned | -672 
acne | -672 
minocycline | -672 
increased WBC count | 0
eosinophilia | 0
systemic involvement | 0
diffuse erythematous or maculopapular eruption | 0
pruritis | 0
DRESS syndrome | 0
fever persisted | 0
rash persisted | 0
discharged | 24