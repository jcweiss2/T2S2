10 years old | 0
male | 0
admitted to the hospital | 0
born | -8760
birth weight 2100 g | -8760
birth length 48 cm | -8760
prominent forehead | -8760
relative macrocephaly | -8760
limb asymmetry | -8760
5th finger clinodactyly | -8760
2/3 toe syndactyly | -8760
hypomethylation of the 11p15 region | -504
genetic examination | -504
diagnosis of SRS | -504
delayed motor development | -384
walked independently | -384
hepatic dysfunction | -420
increased concentration of alanine aminotransferase | -420
increased concentration of aspartate aminotransferase | -420
increased creatine kinase level | -420
diagnosis of Duchenne muscular dystrophy | -420
genetic test | -396
mutation of the maternal DMD gene | -396
corticosteroids treatment | -288
prednisone treatment | -288
deflazacort treatment | -192
G-CSF treatment | -144
sepsis | -144
hypoglycaemia | -144
neurological symptoms | -144
glucose level 14 mg/dl | -144
urological care | -144
hypospadias | -144
cardiological diagnostics | -12
episodes of sinus tachycardia | -12
heart murmur | -12
propranolol treatment | -12
growth hormone deficiency | -12
rhGH treatment | 0
growth hormone therapy | 0
impaired glucose tolerance | 12
insulin resistance | 12
weight gain | 12
discontinuation of rhGH therapy | 18
muscle weakness | 18
paediatric neurologist | 18
hypoglycaemia | -144
fasting hypoglycaemia | -144
glucocorticoid therapy | -288
disturbances of carbohydrate metabolism | -288
growth hormone therapy | 0
hepatic gluconeogenesis | 0
insulin resistance | 12
hyperinsulinaemia | 12
diabetes | 12
scoliosis | 0
bone mineral density | 12
dual-energy X-ray absorptiometry | 12
BMD assessment | 12
lumbar spine | 12
Z-score -2.2 | 12