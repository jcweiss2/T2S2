20 years old | 0
male | 0
relapsed acute myeloid leukemia | -1680
myelodysplasia-related features | -1680
chemotherapy administered | -1680
recto-cecal abscess | -1176
appendectomy | -1176
admitted to the hospital | -1176
febrile neutropenia | -1176
septic shock | -1176
thrombocytopenia | -1176
broad spectrum antibiotics | -1176
meropenem | -1176
vancomycin | -1176
micafungin | -1176
amikacin started | -1176
amikacin discontinued | -1176
right arm cellulitis | -1176
abscess | -1176
ESBL | -1176
CRE Escherichia coli | -1176
colistin started | -1176
loading dose colistin | -1176
maintenance dose colistin | -1176
amphotericin B | -1176
ICU admission | 0
colistin continued | 0
meropenem continued | 0
tigecycline added | 0
micafungin switched to amphotericin B | 0
blood pressure improved | 24
norepinephrine discontinued | 24
febrile | 0
colistin administration day 28 | 672
hypotension | 672
norepinephrine re-initiated | 672
shortness of breath | 672
hypoxia | 672
tachycardia | 672
tachypnea | 672
flushed face | 672
colistin held | 672
adrenaline administered | 672
chlorpheniramine administered | 672
hydrocortisone administered | 672
leukocytosis | 672
acute kidney injury | 672
colistin treatment continued | 672
leukocytosis resolved | 96
renal function baseline | 96
norepinephrine discontinued | 96
colistin resumed | 96
day 5 ICU admission | 120
day 31 colistin treatment | 744
hypotension | 744
norepinephrine re-initiated | 744
shortness of breath | 744
hypoxia | 744
flushed face | 744
generalized erythema | 744
adrenaline administered | 744
hydrocortisone administered | 744
chlorpheniramine administered | 744
leukocytosis | 744
acute kidney injury | 744
increased total bilirubin | 744
colistin discontinued | 744
meropenem continued | 744
tigecycline continued | 744
amikacin started | 744
norepinephrine discontinued | 168
laboratory results resolved | 168
condition stabilized | 216
transferred to floor | 216
piperacillin/tazobactam | 216
tigecycline | 216
amikacin | 216
ventricular fibrillation | 240
death | 240
