27 years old | 0
G2P1 | 0
healthy female | 0
40 weeks of pregnancy | 0
emergency cesarean section | 0
arrest of labor | 0
uncomplicated pregnancy | 0
no gestational hypertension | 0
no diabetes | 0
episode of bradycardia | 0
hypotension | 0
postpartum hemorrhage | 0
estimated blood loss of 2 L | 0
progressive hypoxemia | 0
refractory hypotension | 0
urgent surgical exploration | 0
no significant ongoing bleeding | 0
hemodynamic instability | 0
heart rate 150 bpm | 0
blood pressure 70/50 mm Hg | 0
oxygen saturation 90% | 0
on 100% nonrebreather | 0
oliguric | 0
resuscitation | 0
transferred to intensive care unit | 0
evidence of DIC | 0
hemoglobin 115 g/L | 0
platelet count 81 x 10E9/L | 0
fibrinogen 0.4 g/L | 0
international normalized ratio 1.8 | 0
acute kidney injury | 0
creatinine 130 μmol/L | 0
arterial blood gas | 0
pH 7.38 | 0
pCO2 26 mm Hg | 0
pO2 91 mm Hg | 0
HCO3 15 mmol/L | 0
lactate 1.7 mmol/L | 0
baseline electrocardiogram | 0
sinus tachycardia | 0
nonspecific T-wave changes | 0
elevated troponin level | 0
492 ng/L | 0
differential diagnosis | 0
AFE | 0
pulmonary embolism | 0
peripartum cardiomyopathy | 0
acute respiratory distress syndrome | 0
anaphylaxis | 0
septic shock | 0
obstetrical causes excluded | 0
transthoracic echocardiogram | 0
left ventricle normal | 0
preserved systolic function | 0
RV dilation | 0
severely reduced systolic function | 0
McConnell’s sign | 0
akinesis of mid RV wall | 0
hypercontractility of RV apex | 0
moderate tricuspid regurgitation | 0
TR max velocity 310.8 cm/sec | 0
linear structure in IVC | 0
consistent with thrombus | 0
computed tomographic pulmonary angiography | 0
low-burden pulmonary embolism | 0
lateral basal segmental pulmonary artery | 0
right lower lobe | 0
abdominal and pelvic computed tomography | 0
thrombosis in right gonadal vein | 0
thrombus extending into IVC | 0
bilateral renal cortical necrosis | 0
norepinephrine | 0
mean arterial pressure | 0
at least 60 mm Hg | 0
acute right heart failure | 0
epinephrine | 0
dobutamine | 0
RV dysfunction | 0
invasive pulmonary artery pressure monitoring | 0
therapeutic anticoagulation | 0
unfractionated heparin | 0
hemodynamics improved | 24
weaning off pressor support | 24
continuous renal replacement therapy | 24
anuric renal failure | 24
refractory volume overload | 24
intermittent hemodialysis | 48
discharge | 168
follow-up | 2160
doing well clinically | 2160
no longer dialysis dependent | 2160
repeat echocardiogram | 2160
normal biventricular function | 2160
repeat computed tomography imaging | 2160
not performed | 2160