37 years old | 0
female | 0
type 2 diabetes mellitus | -672
peripheral neuropathy | -672
morbid obesity | -672
obstructive sleep apnea | -672
gastroesophageal reflux disease | -672
depression | -672
intellectual disability | -672
metformin | -672
hemoglobin A1c 9.8% | -672
sitagliptin | -30
canagliflozin | -30
pain in the left gluteal region | -30
dysuria | -30
trimethoprim/sulfamethoxazole | -25
urinary tract infection | -25
admitted to the hospital | 0
afebrile | 0
tachycardic | 0
blood pressure 144/79 mmHg | 0
respiratory rate 19 breaths/minute | 0
lethargic | 0
in distress | 0
suprapubic tenderness | 0
induration to the left gluteal region | 0
blood glucose 402 mg/dL | 0
serum bicarbonate 12 mmol/L | 0
elevated anion gap 24 mmol/L | 0
lactate 1.8 mmol/L | 0
glycosuria | 0
ketonuria | 0
b-hydroxybutyrate 2.49 mmol/L | 0
arterial blood gas analysis | 0
pH 7.23 | 0
PCO2 34 mmHg | 0
computed tomography of the abdomen and pelvis | 0
Fournier’s gangrene | 0
IV normal saline | 0
IV ceftazidime | 0
IV clindamycin | 0
vancomycin | 0
debridement | 0
incision and drainage | 0
hypotensive | 24
tachycardic | 24
sepsis | 24
surgical exploration | 24
vasopressors | 24
antibiotics switched | 24
surgical re-explorations | 48
laparoscopic transverse loop colostomy | 168
DKA management | 72
subcutaneous insulin | 72
insulin infusion | 72
aggressive fluid resuscitation | 72
anion gap closed | 96
acidosis resolved | 96
transferred to the general medical floor | 408
discharged | 672
canagliflozin discontinued | 672
sitagliptin-metformin discontinued | 672
insulin glargine | 672
urinary catheter | 672
vacuum dressing | 672
colostomy | 672