17 years old | 0
female | 0
school-going | 0
admitted to the hospital | 0
acute onset of behavioral change | -72
extreme politeness | -72
obedience | -72
excessive and irrelevant talks | -72
disinhibition | -72
verbal and physical aggression | -240
muttering to herself | -240
marked delusional thoughts | -240
tendency to run amok | -240
diagnosis of acute functional psychosis | -240
oleanzapine started | -240
stiffness of whole body | -168
akinesia | -168
mutism | -168
MRI Brain | -168
non-diffusion restricted, non-contrast-enhancing T2 and FLAIR hyper intensities | -168
CSF examination | -168
no cells | -168
normal protein | -168
normal glucose levels | -168
CSF viral markers negative | -168
Venereal Diseases Research Laboratory test negative | -168
gram stain negative | -168
acid fast bacillus stain negative | -168
India ink negative | -168
cryptococcal antigen negative | -168
bacterial, mycobacterial and fungal cultures negative | -168
Electroencephalogram | -168
non-specific diffuse theta delta slowing | -168
low grade fever | -168
serum Creatinine Phosphokinase raised | -168
diagnosis of NMS | -168
dantrolene and hydration started | -168
clinical worsening | -168
frequent bouts of tachypnea | -48
tachycardia | -48
hypotension | -48
sweating | -48
gasping for breath | -24
oxygen desaturation | -24
endotracheal intubation | -24
mechanical ventilation | -24
widely fluctuating heart rate | 0
blood pressure fluctuations | 0
stimulus-induced sinus tachycardia | 0
tachypnea | 0
diaphoresis | 0
sedative infusion | 0
provisional diagnosis of sepsis syndrome | 0
bilateral aspiration pneumonia | 0
critical care and medical support | 0
re-evaluation by neurology team | 0
possibility of immune encephalitis | 0
MRI Brain repeated | 0
similar changes as noted before | 0
work up for infectious meningoencephalitis | 0
CSF samples sent for anti-NMDA receptor antibody | 0
anti-Voltage gated potassium channel VGKC | 0
anti-α-amino-3-hydroxy-5-methyl-4-isoxazolepropionic acid receptor antibody levels | 0
vasculitic work up | 0
anti nuclear antibody negative | 0
anti-double stranded DNA negative | 0
anti phospholipid antibody negative | 0
lupus anti-coagulant negative | 0
cytoplasmic and perinuclear anti neutrophilic cytoplasmic antibody negative | 0
anti-thyroid peroxidase antibody negative | 0
anti-thyroglobulin antibody negative | 0
CT scan of chest, abdomen, and pelvis | 0
no ovarian teratoma | 0
no other malignancy | 0
tonic-clonic seizures | 0
intravenous immunoglobulin | 0
20 g/day | 0
5 days | 0
improvement of sensorium | 24
ability to spontaneously open eyes | 24
fixate gaze | 24
ventilator-associated bilateral pneumothorax | 48
bilateral intercostal tube drainage | 48
oro-lingual dyskinesias | 48
subsided over next 10 days | 120
weaned off the ventilator | 168
anti-NMDA antibody in CSF positive | 168
anti-VGKC and anti-AMPA antibodies negative | 168
diagnosis of anti-NMDARE confirmed | 168
remarkable and quick neurological recovery | 336
full recovery of sensorium | 336
normal higher mental functions | 336
distal acral lower motor neuron deficit | 336
critical illness polyneuropathy | 336
follow-up and periodic screening for teratoma | 336