57 years old | 0
male | 0
admitted to the hospital | 0
fever | -168
cough | -168
ischaemic stroke | -17520
patent foramen ovale | -17520
percutaneous closure | -17520
temperature 38°C | 0
dyspnoea | 0
bilateral lung crackles | 0
no murmur | 0
no sign of heart failure | 0
SARS-CoV-2 infection | 0
bilateral ground-glass and crazy paving pulmonary involvement | 0
hydroxychloroquine | 0
antiviral agents | 0
lopinavir/ritonavir | 0
hypoxaemia | 72
non-responsive to ventilation with continuous positive air pressure (CPAP) | 72
PaO2/FiO2 ratio <100 | 72
acute respiratory distress syndrome | 72
ICU admission | 72
mechanical ventilation | 72
paroxysmal atrial fibrillation | 72
low molecular weight heparin | 72
fever | 336
haemoculture positive for MRSA | 336
transthoracic echocardiography | 336
poor ultrasound window | 336
mild mitral regurgitation | 336
mild impairment of left ventricular systolic function | 336
ejection fraction 45% | 336
sepsis-related myocardial dysfunction | 336
ARDS-related myocardial dysfunction | 336
high clinical suspicion for IE | 336
transoesophageal echocardiography | 480
endocarditis vegetation | 480
no paravalvular abscess | 480
no abnormalities on PFO closure device | 480
no significant dysfunction in other cardiac valves | 480
tiny perforation | 480
mild eccentric aortic valve regurgitation | 480
ventilator-associated pneumonia | 480
Klebsiella pneumoniae infection | 480
bilateral areas of increased density | 480
teicoplanin | 504
ceftazidime/avibactam | 504
linezolid | 504
fosfomycin | 528
reduction of inflammatory markers | 528
improvement of clinical status | 528
SARS-CoV-2 infection | 504
no severe aortic valve dysfunction | 504
no endocarditis-related complications | 504
ICU discharge | 720
rehabilitation hospital transfer | 888
transthoracic echocardiography | 1200
residual vegetation of smaller dimension | 1200
no significant regurgitation | 1200
