48 years old | 0
male | 0
chronic pancreatitis | 0
alcohol dependency | 0
presented with septic shock | 0
cellulitic genitalia | 0
oedematous genitalia | 0
mottled discoloration of genitalia | 0
cellulitic perineum | 0
oedematous perineum | 0
mottled discoloration of perineum | 0
transferred to tertiary centre | 0
radical debridement by urology | 0
radical debridement by plastic surgery | 0
radical debridement by general surgery | 0
copious pus from left inguinal canal | 0
large left-sided retroperitoneal collection | 0
placement of two large drains | 0
no intra-peritoneal collection | 0
computed tomography scan | 0
acute-on-chronic pancreatitis | 0
focal necrosis at head of pancreas | 0
fluid tracking to retroperitoneum | 0
fluid tracking to perineum | 0
subcutaneous emphysema in left flank | 0
stabilized in ICU | 0
inotropic support | 0
intravenous antibiotic therapy | 0
further debridement of non-viable soft tissues | 0
medial thigh pouches for testes | 0
VAC dressing | 0
polymicrobial growth isolated | 0
sensitive to piperacillin/tazobactam | 0
histology confirmed necrotizing fasciitis | 0
3-week intravenous therapy | 0
switched to oral antibiotics for 3 weeks | 168
acute pancreatitis | 0
Imrie Score 4 | 0
managed conservatively | 0
nasogastric feeding | 0
diabetes mellitus type 2 | 0
commenced oral treatment | 0
multiple debridements | 0
VAC changes | 0
abdomino/perineal skin defect ready for resurfacing | 504
split-skin grafting | 504
100% graft uptake by Day-7 | 504
discharged | 504
follow-up at 2 months | 1344
excellent recovery | 1344
