42 years old | 0
male | 0
Caucasian | 0
bilateral lung transplant | -12000
cystic fibrosis | -12000
admitted to the ICU | 0
fever | -24
flu-like symptoms | -24
acute hypoxemic respiratory failure | -24
PaO2/FiO2 ratio = 81 | -24
computed tomogram of the chest | 0
diffuse bilateral ground-glass nodular opacities | 0
areas of mosaic attenuation | 0
mechanical ventilation | 24
low tidal volume | 24
positive end-expiratory pressure | 24
septic shock | 24
refractory hypoxemia | 24
neuromuscular blockade | 24
cisatracurium | 24
pulmonary vasodilator therapy | 24
inhaled epoprostenol | 24
vasopressor support | 24
immunosuppression curtailed | 24
broad-spectrum antimicrobial therapy | 24
vancomycin | 24
piperacillin-tazobactum | 24
azithromycin | 24
voriconazole | 24
PPV initiated | 24
manual proning | 24
improvement in hypoxemia | 48
PaO2 of 81 mmHg to 168 mmHg | 48
bronchoscopic sampling deferred | 24
patient's daughter tested positive for Bordetella pertussis | 192
patient tested positive for Bordetella pertussis | 216
levofloxacin added | 216
mechanically rotating bed | 216
PPV for approximately 16 hours a day | 216
ventilator dyssynchrony | 432
deep sedation | 432
intermittent neuromuscular blockade | 432
tracheostomy | 648
liberated from mechanical ventilation | 1536
severe neuromuscular weakness | 648
critical illness neuropathy/myopathy | 648
ICU delirium | 648
non-reactive pupils | 744
cessation of neuromuscular blockade | 744
neurological work-up | 744
magnetic resonance imaging of the brain | 744
multifocal lesions | 744
left occipital lobe | 744
central and peripheral enhancement | 744
septic emboli | 744
lumbar puncture | 744
MR angiography | 744
trans-esophageal echocardiogram | 744
serial blood cultures | 744
fundoscopic examination | 744
bilateral visual loss | 744
optic nerve pallor | 744
hypoxia-induced cerebral infarction | 744
increased intraocular pressure | 744
decrease in ocular perfusion pressure | 744
optic nerve injury | 744
A2B0 rejection | -12000
peak FEV1 post-transplant = 3.32 liters | -12000
pre-ICU FEV1 = 3.17 liters | 0
FEV1 = 1.74 liters | 4320
legally blind | 4320
bilateral optic atrophy | 4320
retinal vascular attenuation | 4320