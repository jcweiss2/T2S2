59 years old | 0
male | 0
resident of Riyadh | 0
visited Karachi | -672
arrival back to Saudi Arabia | -48
persistent fever | -48
seen in clinic in King Faisal Specialized Hospital | -24
prescribed antipyretics | -24
failed to improve fever | -24
symptoms progressed | -24
continuous vomiting | -24
nonprojectile vomiting | -24
headaches | -24
no contact with sick individuals | -672
no URTI symptoms | 0
no ear problems | 0
no animal contact | 0
no swimming | 0
no bathing ponds | 0
CSF sample taken | 0
assessed by neurology team | 0
awake | 0
confused | 0
agitated | 0
became drowsy | 1
barely responsive to painful stimuli | 1
no longer protecting airway | 1
intubated | 1
admitted to ICU | 1
septic shock | 1
primary central nervous system infection | 1
laboratory investigations | 0
CT brain angiogram | 0
no acute intracranial insult | 0
CTA | 0
no significant stenosis | 0
no focal occlusion | 0
CT brain without contrast | 24
new onset diffuse brain edema | 24
moderate diffuse narrowing of CSF spaces | 24
scattered hyperattenuating foci | 24
leptomeningeal process | 24
physical examination | 24
coma | 24
fixed dilated pupils | 24
vital signs stable | 24
inotropic support | 24
other examinations within normal limits | 24
started on broad antimicrobial coverage | 24
lumbar puncture | 24
cultures negative | 24
CSF preserved for metagenomics | 24
clinical condition worsened | 72
antimicrobial regimen modified | 72
technetium-99m HMPO brain perfusion scan | 72
confirmed brain death | 72
clinical situation persisted | 72
biochemical situation deteriorated | 72
passed away | 216
metagenomic sequencing | 216
identified PAM | 216
Naegleria fowleri | 216
developed symptoms after return from Karachi | -48
acquired infection in Karachi | -48
draft assembly of Karachi-NF001 genome | 216
unique genetic features | 216
rare disease | 0
no high index of suspicion | 0
trophozoites detection | 0
culture-based detection | 0
PCR methods | 0
immunohistochemistry methods | 0
signs similar to bacterial meningitis | 0
signs similar to viral meningitis | 0
metagenomics protocol | 216
PAM detection within 24 hours | 216
mNGS-based diagnosis | 216
access to NGS facilities limitation | 216
efforts for mNGS facilities | 216
study reveals mNGS valuable | 216
no acute intracranial insult |= 0
