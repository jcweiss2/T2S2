44 years old | 0
male | 0
admitted to the hospital | 0
shortness of breath | -48
nonproductive cough | -48
obesity | 0
type 2 diabetes | 0
bacterial pneumonia | 0
viral upper or lower respiratory tract infection | 0
pulmonary embolism | 0
COVID-19 illness | 0
temperature 99.3°F | 0
heart rate 152 beats/min | 0
blood pressure 102/84 mm Hg | 0
respiratory rate 44 breaths/min | 0
hypoxic | 0
peripheral oxygenation saturation 86% | 0
supplemental oxygen via nasal cannula | 0
non-rebreather mask | 0
diffuse bilateral hazy opacities | 0
SARS-CoV-2 nasopharyngeal swab polymerase chain reaction test positive | 0
venous blood gas analyses | 0
pH 7.09 | 0
partial arterial pressure of carbon dioxide 41 mm Hg | 0
partial arterial pressure of oxygen 33 mm Hg | 0
lactate level 12 mmol/l | 0
intubation | 0
arterial blood gas analysis | 0
pH 7.14 | 0
partial arterial pressure of carbon dioxide 53 mm Hg | 0
partial arterial pressure of oxygen 193 mm Hg | 0
fraction of inspired oxygen 100% | 0
Pao2:fraction of inspired oxygen ratio 193 | 0
acute respiratory distress syndrome | 0
white blood cell count 27.8 × 10^3/μl | 0
serum creatinine 1.88 mg/dl | 0
high-sensitivity troponin-T level 46 ng/l | 0
N-terminal B-type natriuretic peptide 14,535 pg/ml | 0
ferritin 3,495 ng/l | 0
D-dimer >20 μg/ml | 0
transthoracic echocardiography | 0
left ventricular ejection fraction 45% | 0
global hypokinesis | 0
right ventricle moderate to severely dilated | 0
right ventricular systolic function moderate to severely reduced | 0
flattening of the interventricular septum | 0
clot in transit | 0
norepinephrine 40 μg/min | 6
vasopressin 2.4 U/h | 6
methylprednisolone 1 mg/kg | 6
tissue plasminogen activator 100 mg | 6
unfractionated heparin | 8
dobutamine infusion | 8
venoarterial extracorporeal membrane oxygenation | 8
weaned off pressors | 24
weaned off inotropic support | 72
repeat transthoracic echocardiography | 72
normal left ventricular systolic function | 72
mild dilation of the right ventricle | 72
preserved right ventricular systolic function | 72
clot in transit no longer visualized | 72
right ventricular function improving | 72
bilateral lower extremity venous Doppler ultrasounds | 72
deep vein thrombosis negative | 72
bleeding within the oropharynx | 120
compression packing | 120
continued systemic anticoagulation | 120
plan for oral anticoagulation | 120