34 years old | 0
female | 0
admitted to the hospital | 0
complaints of epigastric pain | -48
dyspnoea | -48
diaphoresis | -48
nausea | -48
vomiting | -48
weight loss | -4320
left flank pain | 0
mild abdominal tenderness | 0
ascites | 0
palpable painful mass | 0
hypotension | 0
ventricular fibrillation | 0
cardiac arrest | 0
defibrillation | 0
cardiopulmonary resuscitation | 0
adrenaline administration | 0
sinus rhythm | 0
coronary angiogram | 0
high thrombus burden | 0
no reflow | 0
tirofiban infusion | 0
stent deployment | 0
echocardiogram | 24
regional wall motion abnormalities | 24
hypokinesia | 24
ejection fraction | 24
right atrial mass | 24
inferior vena cava mass | 24
anticoagulation | 48
rivaroxaban | 48
dual antiplatelet therapy | 48
acetylsalicylic acid | 48
clopidogrel | 48
investigation of diseases | 48
haematological parameters | 48
biochemical parameters | 48
lipid profile | 48
tumour markers | 48
connective tissue markers | 48
thrombophilia panel | 48
cancer antigen 125 | 48
abdominal CT scan | 168
necrotic mass | 168
left adrenal gland bed | 168
tumour thrombus | 168
hepatic veins | 168
right atrium | 168
iliac vein bifurcation | 168
venous Doppler | 168
24-hour urine analyses | 216
vanillylmandelic acid | 216
5 hydroxy indole acetic acid | 216
homovanillic acid | 216
image-guided tissue sampling | 312
histopathological analysis | 312
PHEOs diagnosis | 312
surgical procedure | 408
metastatic foci | 408
intensive anticoagulant therapy | 408
177Lu-DOTATATE-based PRRT | 480
treatment initiation | 480
septic shock | 720
nosocomial infections | 720
vancomycin-resistant enterococci | 720
discharge | 720
readmission | 2160
death | 2160