34 years old | 0
male | 0
alcohol dependence | 0
left-sided, cramping abdominal pain | -24
abdominal pain radiating to the back | -24
denied prior episodes | 0
denied any inciting incidents | 0
denied any known history of diabetes mellitus | 0
denied medication use | 0
denied pancreatitis | 0
denied family history of genetic dyslipidemias | 0
not obese | 0
body mass index (BMI) 24.4 | 0
tachycardia | 0
tachycardia at 112/min | 0
moderate tenderness to palpation in the right upper quadrant | 0
moderate tenderness to palpation in the left upper quadrant | 0
moderate tenderness to palpation in the left lower quadrant | 0
leukocytes 12 k/µL | 0
neutrophils 81.8% | 0
potassium 3.2 mEq/L | 0
random glucose 136 mg/dL | 0
calcium 6.8 mg/dL | 0
alanine aminotransferase 73 U/L | 0
aspartate aminotransferase 80 U/L | 0
alkaline phosphatase 135 IU/L | 0
TGs 9708 mg/dL | -24
low-density lipoprotein 373 mg/dL | 0
lipase 245 U/L | 0
acute interstitial pancreatitis | 0
peripancreatic fluid surrounding the pancreatic tail | 0
fatty infiltration of the terminal ileum submucosa | 0
admitted to the medical ICU | 0
nil per os | 0
insulin drip | 0
dextrose 10% in water drip | 0
high-volume intravenous fluids | 0
electrolyte replenishment | 0
analgesia | 0
serum TG level 4025 mg/dL | 0
plasmapheresis | 24
volume replacement of 1250 cm3 of fresh frozen plasma | 24
volume replacement of 1250 cm3 of 5% albumin | 24
TG level 603 mg/dL | 24
insulin drip continued | 24
TG level 304 mg/dL | 48
transferred to the medical floors | 48
discharged | 72