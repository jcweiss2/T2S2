36 years old | 0
male | 0
black | 0
admitted to the hospital | 0
low back pain | -96
bruised hips | -96
macroscopic hematuria | -96
gingival bleeding | -96
conscious | 0
oriented | 0
pale | 0
tachycardic | 0
blood pressure 120/90 mmHg | 0
mild edema | 0
varicose veins of the lower limbs | 0
chronic malleolar ulcers | 0
bleeding and bruising in the pelvic region | 0
denies personal or family history of bleeding diathesis | 0
renal and urological diseases ruled out | 0
hemoglobin level 4.8 g/dL | 0
platelet count 270 × 10^9/L | 0
incoagulable blood | 0
prothrombin time (PT) | 0
activated partial thromboplastin time (APTT) | 0
transfusion of red blood cells | 0
transfusion of cryoprecipitate | 0
transfusion of fresh frozen plasma | 0
transferred to the intensive care unit | 0
hematuria | 48
ecchymosis | 48
incoagulable blood | 48
patient-to-control APTT ratio 1.79 | 48
transfusion support continued | 48
positive results for lupus anticoagulant antibodies | 48
negative results for anticardiolipin immunoglobulin (Ig)M | 48
negative results for anticardiolipin immunoglobulin (Ig)G | 48
negative results for anticardiolipin immunoglobulin (Ig)A | 48
negative results for antinuclear antibodies | 48
negative results for rheumatoid factors | 48
activity levels of coagulation factors | 48
factor VII 3% | 48
factor II 130% | 48
factor V 150% | 48
factor VIII >200% | 48
factor IX 47% | 48
factor X 75.8% | 48
intravenous pulse therapy with methylprednisolone | 48
prothrombin complex concentrate | 48
recovered well | 72
no bleeding | 72
corticotherapy maintained with oral administration of 1 mg/kg/day prednisone | 72
discharged | 408
follow-up in an outpatient clinic | 408
corticoid dose reduced | 504
consecutive PT test results showed a progressive tendency toward normality | 504
condition stabilized | 504
no new hemorrhagic episodes | 504
corticoid treatment suspended | 816
PT 83.2% | 816
patient-to-control APTT ratio 1.05 | 816
fibrinogen level 248.7 mg/dL | 816
factor VII activity level 60.6% | 816
factor II 130% | 816
factor V 180% | 816
factor VIII >200% | 816
factor IX 47% | 816
factor X 75.8% | 816
lupus anticoagulant negative | 816