44 years old | 0
African-American | 0
female | 0
admitted to the Hematology/Oncology clinic | 0
complaints of weakness | 0
complaints of fatigue | 0
past medical history of HTLV associated T-cell lymphoma/leukemia | -672
underwent allogenic bone marrow transplant | -672
disease relapse | -168
graft failure | -168
blood transfusion dependence | -168
recently admitted due to disseminated aspergillosis | -24
involving the skin | -24
involving the lungs | -24
on treatment with oral posaconazole | -24
on treatment with high dose micafungin | -24
via left tunneled internal jugular catheter | -24
prophylaxis regimen included oral acyclovir | -24
prophylaxis regimen included oral levofloxacin | -24
prophylaxis regimen included monthly inhaled pentamidine | -24
hypotensive | 0
tachycardic | 0
afebrile | 0
non-tender ulceration of 2 cm in diameter in right distal leg | 0
without erythema | 0
without discharge | 0
without induration | 0
left internal jugular tunneled catheter | -120
catheter exit site without erythema | 0
catheter exit site without drainage | 0
admitted to the intensive care unit | 0
presumptive diagnosis of sepsis | 0
blood cultures obtained from the central line | 0
blood cultures obtained from periphery | 0
empirically treated with cefepime | 0
empirically treated with vancomycin | 0
leukopenia | 0
absolute neutrophil count of 0.04 K/uL | 0
low hemoglobin | 0
thrombocytopenia | 0
high creatinine | 0
marked elevation of transaminases | 0
AST 505 U/L | 0
ALT 477 U/L | 0
bilateral perihilar and pulmonary nodules | 0
hypotension worsened | 24
norepinephrine infusion | 24
antibiotic therapy escalated from cefepime to meropenem | 24
vancomycin continued | 24
intravenous isavuconazole substituted for posaconazole | 24
intravenous micafungin continued | 24
four sets of blood cultures grew gram-positive rods | 48
identified as Cellulosimicrobium sp. | 48
in vitro susceptibility testing performed by E-test | 48
Benzyl penicillin minimum inhibitory concentration (MIC) = 0.012 ug/mL | 48
levofloxacin MIC >32 ug/mL | 48
vancomycin MIC = 0.38 ug/mL | 48
tunneled catheter removed | 48
catheter tip grew Cellulosimicrobium sp. | 48
clinically improved | 72
resolution of hypotension | 72
resolution of acute renal failure | 72
resolution of transaminitis | 72
meropenem discontinued | 72
oral levofloxacin resumed for neutropenic prophylaxis | 72
repeat blood cultures became negative | 96
intravenous vancomycin therapy | 0
discharged | 168
readmitted | 216
pneumonia | 216
death | 216