71 years old | 0
female | 0
admitted to the hospital | 0
unconscious state | 0
history of hypertension | 0
history of ischaemic heart disease | 0
history of peripheral vascular disease | 0
stroke | 0
head computed tomographic scan | 0
inotropic support | 24
septic shock | 24
elevated levels of inflammatory markers | 24
erythrocyte sedimentation rate | 24
C-reactive protein | 24
blood culture | 24
yeast in both aerobic and anaerobic BacT/ALERT culture bottles | 24
caspofungin | 24
died | 72
identification of yeast | 24
VITEK 2 yeast identification system | 24
CHROMagar Candida | 24
acetate ascospore agar | 168
internally transcribed spacer region of ribosomal DNA | 168
sequencing | 168
Lodderomyces elongisporus | 168
Candida parapsilosis | 168
antifungal susceptibility | 168
Etest | 168
amphotericin B | 168
fluconazole | 168
voriconazole | 168
posaconazole | 168
itraconazole | 168
flucytosine | 168
caspofungin | 168
micafungin | 168