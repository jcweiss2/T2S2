25 years old | 0
African American | 0
female | 0
presenting to the emergency department | 0
found on the floor at home | 0
verbally incomprehensible | 0
complete bilateral vision loss | 0
altered mental status | 0
systemic hypertension of unknown cause | -672
stage 4 chronic kidney disease | -672
idiopathic intracranial hypertension | -672
ventriculoperitoneal shunt | -672
hypertensive retinopathy | -672
optic neuropathy | -672
loss of peripheral vision in right eye | -672
loss of central vision in left eye | -672
third admission for acute kidney injury on chronic kidney disease | 0
blood pressure of 168/98 mmHg | 0
pulse of 100 beats per minute | 0
minimally verbal | 0
obtunded | 0
total bilateral vision loss | 0
left sided rib pain | 0
coughing | 0
hypodensities in the cerebellum | 0
hyperdensities extending to the cortex in the posterior occipital lobe | 0
vasogenic edema in the cerebellum | 0
posterior parietal and occipital lobes bilaterally | 0
blood urea nitrogen of 92.0 mg/dL | 0
creatinine of 17.56 mg/dL | 0
right-sided atrial septum vegetation | 0
culture-negative endocarditis | 0
PRES diagnosis | 0
controlled blood pressure with labetalol and hydralazine | 0
clevidipine initiation | 0
carvedilol regimen | 24
lisinopril regimen | 24
nifedipine regimen | 24
tunneled catheter placement | 24
dialysis treatment | 24
sevelamer carbonate initiation | 24
vancomycin initiation | 24
ceftazidime initiation | 24
regained baseline cognition | 168
regained baseline vision | 168
cerebral metamorphopsia | 168
metamorphopsia resolution | 168
outpatient follow-up MRI | 336
vasogenic edema resolution | 336
