75 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
fever | -168 | 0 | Factual
chills | -168 | 0 | Factual
dizziness | -168 | 0 | Factual
remission after fever | -168 | 0 | Factual
no headache | 0 | 0 | Negated
no abdominal pain | 0 | 0 | Negated
no diarrhea | 0 | 0 | Negated
no sputum | 0 | 0 | Negated
no nasal congestion | 0 | 0 | Negated
no runny nose | 0 | 0 | Negated
hypertension | -672 | 0 | Factual
body temperature 39.0 °C | -168 | 0 | Factual
levofloxacin | 0 | 72 | Factual
body temperature above 39.0 °C | 0 | 72 | Factual
blood culture indicated penicillin-resistant Staphylococcus | 72 | 72 | Factual
Vancomycin | 72 | 168 | Factual
body temperature returned to normal | 168 | 168 | Factual
discharged | 168 | 168 | Factual
high fever again | 168 | 168 | Factual
chills | 168 | 168 | Factual
cough | 168 | 168 | Factual
sputum | 168 | 168 | Factual
no chest pain | 168 | 168 | Negated
no limb twitching | 168 | 168 | Negated
pupils sluggish in light reflection | 168 | 168 | Factual
confused | 168 | 168 | Factual
mentally soft | 168 | 168 | Factual
diarrhea | 168 | 168 | Factual
hospitalized in ICU | 168 | 168 | Factual
high-frequency oxygen inhalation | 168 | 168 | Factual
piperacillin and tazobactam | 168 | 240 | Factual
methylprednisolone | 168 | 240 | Factual
body temperature above 38.3 °C | 168 | 240 | Factual
levofloxacin | 240 | 240 | Factual
body temperature returned to normal | 240 | 240 | Factual
CRP dropped to 76.4 mmol/L | 240 | 240 | Factual
transferred to general ward | 240 | 240 | Factual
atrial fibrillation | 240 | 240 | Factual
unresponsiveness | 240 | 240 | Factual
slurred speech | 240 | 240 | Factual
shortness of breath | 240 | 240 | Factual
slow light reflexes | 240 | 240 | Factual
stiff neck | 240 | 240 | Factual
increased muscle tone | 240 | 240 | Factual
wet rales in both lungs | 240 | 240 | Factual
septic shock | 240 | 240 | Factual
norepinephrine micropump | 240 | 288 | Factual
vancomycin and meropenem | 240 | 288 | Factual
methylprednisolone stopped | 240 | 288 | Factual
unconscious | 288 | 288 | Factual
base of tongue fell back | 288 | 288 | Factual
shortness of breath | 288 | 288 | Factual
stiff neck | 288 | 288 | Factual
tremor of limbs | 288 | 288 | Factual
heart rate dropped to 40 beats per minute | 288 | 288 | Factual
trachea intubated | 288 | 288 | Factual
breathing assisted by ventilator | 288 | 288 | Factual
condition deteriorated rapidly | 288 | 288 | Factual
multiple organ failure | 288 | 288 | Factual
discontinuation of treatment | 288 | 288 | Factual
death | 288 | 288 | Factual
L. monocytogenes | -168 | 288 | Factual
meningoencephalitis | 0 | 288 | Factual
sepsis | 0 | 288 | Factual
lung infection | 0 | 288 | Factual
respiratory failure | 0 | 288 | Factual
electrolyte imbalance | 0 | 288 | Factual
hyponatremia | 0 | 288 | Factual
hypokalemia | 0 | 288 | Factual
autoimmune disease | 0 | 288 | Factual
cerebrospinal fluid metagenomic test | 0 | 0 | Factual
bilateral blood culture test | 0 | 0 | Factual
cerebrospinal fluid examination | 0 | 0 | Factual
metagenomic detection technology | 0 | 0 | Factual
sensitive antibiotics | 0 | 288 | Factual
early identification | 0 | 0 | Factual
timely application of antibiotics | 0 | 288 | Factual