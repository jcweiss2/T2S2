15 years old | 0
male | 0
admitted to the hospital | 0
fever | -24
confusion | -24
sweating | -24
vomiting | -24
myalgias | -24
cutaneous rash | -24
mildly confused | -24
body temperature 38.6 °C | 0
blood pressure 60/30 mmHg | 0
heart rate 170 bpm | 0
oxygen saturation 98% | 0
diffuse cutaneous exanthema | 0
moderate abdominal tenderness | 0
elevated inflammatory markers | 0
WBC 21 000/mm³ | 0
CRP 250 mg/L | 0
coagulopathy | 0
acute renal failure | 0
transferred to the Intensive Care Unit | 0
intravenous fluids | 0
vasopressors | 0
empirical amoxicillin-clavulanate | 0
blood cultures positive for staphylococci | 24
Staphylococcus aureus identified | 29
PBP2a test negative | 29
antibiogram confirmed multi-sensitive bacterial strain | 29
treatment with intravenous antibiotics | 0
treatment with oral antibiotics | 168
hand and feet desquamation | 336
molecular analysis confirmed tsst-1 gene | 168
typing of the strain showed t2509 Staphylococcus aureus | 168
discharged | 168
ate meat in a fast food restaurant | -28
food intoxication syndrome | -24
emesis | -24
diarrhea | -24