31 years old | 0
G1P0 | 0
primary infertility | 0
cystic fibrosis | 0
preconception counseling | -52
trying to conceive | -52
infertility work-up | -52
ovulation predictor kits | -52
timed intercourse | -52
hysterosalpingogram | -52
semen analysis | -52
mild teratospermia | -52
pelvic ultrasound | -52
antral follicle count | -52
arcuate uterus | -52
polycystic ovarian syndrome work-up | -52
serum hormone levels | -52
ovulation induction protocol | -36
letrozole | -36
cycle day 12 ultrasound | -36
luteinizing hormone | -36
progesterone levels | -36
combined oral contraceptive pills | -24
increase in breast size | -24
in vitro fertilization | -17
follicle stimulating hormone | -17
gonadotropin-releasing hormone antagonist | -17
estradiol | -14
progesterone supplementation | -7
embryo transfer | -1
pregnancy | 0
breast pain | 4
breast ultrasound | 4
Endocrinology referral | 5
bromocriptine | 5
cabergoline | 8
surgical oncology consultation | 10
plastic surgery consultation | 13
physical therapy | 13
manual lymphatic drainage | 13
superficial skin breakdown | 15
oxycodone | 17
tylenol | 17
admitted to antepartum unit | 17
methadone | 17
deep venous thrombosis prophylaxis | 17
enoxaparin | 17
breast ulceration | 20
hemorrhage from exposed venous sinuses | 20
suture ligation | 20
betamethasone | 24
bilateral IV access | 24
crossmatched for packed red blood cells | 24
intravenous iron infusions | 24
visual hallucinations | 24
psychiatry consultation | 24
venlafaxine | 24
citalopram | 24
induction of labor | 31
primary C-section | 31
neonatal intensive care unit | 31
respiratory distress syndrome | 31
necrotizing enterocolitis | 31
Zosyn | 31
postoperative day 5 | 36
breast size decrease | 36
methadone weaning | 36
narcotic withdrawal | 36
postpartum hospitalization | 36
wound care | 36
plastic surgery follow-up | 36
breast surgery follow-up | 36
MFM follow-up | 36
3-week postpartum visit | 42
narcotic-free | 42
breast reduction | 69
free nipple grafts | 69
surgery | 69
postoperative day 1 | 70
Jackson-Pratt drains | 70