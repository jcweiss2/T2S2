female | 0
infant | 0
born at 36+6 weeks gestation | 0
birth weight of 3776 g | 0
conceived via in-vitro fertilization | -672
Apgar scores were 8 and 9 at 1 and 5 min of life | 0
high vaginal swab tested negative for group B streptococcal colonization | -672
no history of prolonged rupture of membranes | -672
no maternal pyrexia | -672
mother is a hepatitis B carrier | -672
Hepatitis B immunoglobulin and vaccine soon after birth | 0
grunting with nasal flaring and subcostal retractions | 0
borderline saturations in room air at 5 min of life | 0
required continuous positive airway pressure (CPAP) support | 0
transferred to the Neonatal Intensive Care Unit (NICU) | 0
intubated at 13 h of life | 13
respiratory support was graded up to High Frequency Oscillatory Ventilation and nitric oxide | 13
Chest X-ray suggested hyaline membrane disease | 13
required two doses of surfactant | 13
Umbilical venous (UVC) and arterial catheters were inserted | 13
malpositioning of the UVC into the right portal vein | 13
septic work up was performed | 24
treated for presumed sepsis with intravenous Penicillin and Gentamicin | 24
Gentamicin was discontinued after the first dose | 24
intravenous Cefotaxime was added | 24
full blood count (FBC) and C-reactive protein (CRP, 0.2 mg l−1) were unremarkable | 0
infective markers showed an upward trend by 12 h (CRP, 24 mg l−1) | 12
infective markers showed an upward trend by day 2 of life (CRP, 170 mg l−1) | 48
blood culture at birth grew SGp | 0
SGp was sensitive to Penicillin and Clindamycin | 0
ear swab cultures showed light mixed growth of SGp | 0
ear swab cultures showed light mixed growth of Escherichia coli | 0
lumbar puncture was deferred due to increasing lability | 24
lumbar puncture was performed | 96
cerebrospinal fluid (CSF) studies returned negative for meningitis | 96
CRP showed a downward trend (48 mg l−1) | 96
developed fever (38.6 °C) | 120
Infectious Disease (ID) team was involved in the care | 120
liver function test revealed conjugated hyperbilirubinemia | 120
renal function normalized | 120
CRP showed a second spike again to 165 mg l−1 | 120
blood culture was repeated | 120
amikacin was added | 120
umbilical lines were removed | 120
urine analysis was unremarkable | 120
echocardiogram was negative for structural heart disease and infective endocarditis | 120
imaging of the abdomen using ultrasound (US) scan showed the presence of a multi-loculated cystic structure | 120
liver abscess | 120
became afebrile | 144
successfully extubated | 144
Penicillin and Amikacin were stopped | 240
continued on Cefotaxime | 240
serial follow-up US scan of the liver showed slow regression of the abscess | 240
needle aspiration and biopsy of the lesion was performed under US guidance | 840
aspirate yield was scanty | 840
biopsy was obtained from the solid hypo-to-isoechoic component of the solid-cystic nodule | 840
histopathological findings are compatible with an abscess cavity | 840
Gram-stain, acid-fast stain and special stains for fungi were negative | 840
bacterial and fungal cultures were sterile | 840
follow-up US on day 37 of life showed further resolution of the abscess cavity | 888
parenteral antibiotics were discontinued | 1080
continued with oral Co-amoxiclav | 1080
imaging at 3 months of age revealed significant resolution of the liver abscess | 2160
sequential liver US scans were done | 4896
abscess cavity to be 0.9×0.3×0.4 cm with dystrophic calcification | 4896
growth and neurodevelopmental assessments were appropriate for age | 4896
Hepatitis B surface antibody was 947 miu l−1 at 9 months of age | 6480