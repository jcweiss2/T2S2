63 years old | 0
    man | 0
    right median nerve epithelioid hemangioendothelioma | -3504
    wide local excision | -3504
    pain along right arm below shoulder | -96
    radiograph of right elbow | -96
    radiograph of chest | -96
    benign muscular pathology | -96
    rotator cuff tendons | -96
    conservative treatments | -96
    pain persisted | -96
    pain worsened | -96
    tumor recurrence concern | -96
    CT scan of right upper extremity | -672
    post-surgical changes | -672
    pain intensified | -672
    PET-CT | -1056
    abnormal uptake in right forearm | -1056
    biopsy of FDG avid area of right forearm | -1056
    traumatic neuroma | -1056
    advised to continue conservative treatments | -1056
    intensifying pain | -2616
    radiograph of right upper extremity | -2616
    abnormality over cortical surface of distal aspect of humeral shaft | -2616
    new lytic lesion | -2616
    repeat PET-CT | -3168
    FDG avidity of mid to distal right humeral shaft | -3168
    associated periosteal changes | -3168
    medial soft tissue mass | -3168
    two satellite nodules in humeral neck area | -3168
    CT-guided biopsy of right humeral mass | -3168
    recurrence of high-grade epithelioid hemangioendothelioma | -3168
    soft tissue recurrence | 0
    local bone metastasis | 0
    discussed with multidisciplinary team | 0
    surgical resection | 0
    progressive dyspnea on exertion | -96
    lower extremity swelling | -96
    difficult to take deep breath | -96
    CT imaging of chest with angiography | -96
    new interstitial-nodular opacities | -96
    negative for acute pulmonary embolism | -96
    cardiac work-up unremarkable | -96
    no symptoms at rest | -96
    discharged home | -96
    symptoms improved | -96
    no longer huffing | -96
    dyspnea when climbing stairs | -96
    pre-anesthesia medical evaluation | 0
    lungs clear to auscultation | 0
    able to lay flat without dyspnea | 0
    resting oxygen saturation 96% on room air | 0
    pre-procedure chest radiograph | 0
    bilateral pulmonary opacities | 0
    predominantly interstitial/septal thickening | 0
    upper lung predominant fine reticulation/micronodularity | 0
    surgical removal of tumor | 0
    pathology revealed high-grade epithelioid hemangioendothelioma | 0
    nodal involvement | 0
    clear margins | 0
    post-operative period | 0
    successfully extubated | 0
    required supplemental oxygen | 0
    chest CT angiogram with PE protocol | 0
    segmental pulmonary embolism | 0
    right diaphragm paralysis | 0
    worsening interstitial-nodular opacities | 0
    progression of prior pulmonary edema | 0
    carcinomatosis could not be ruled out | 0
    transthoracic echocardiogram | 0
    new severe right heart failure | 0
    fully anticoagulated with heparin | 0
    received diuretics | 0
    clinical status continued to decline | 0
    respiratory failure | 0
    septic shock | 0
    transfer to intensive care unit | 0
    intubated | 0
    treated with broad spectrum antibiotics | 0
    bronchoscopy | 0
    bloody secretions | 0
    mildly edematous airway | 0
    no focal endobronchial abnormality | 0
    no area of bleeding | 0
    bronchoalveolar lavage negative for malignancy | 0
    chest imaging | 0
    diffuse alveolar filling process | 0
    treated empirically with high-dose steroids | 0
    no response | 0
    succumbed to hypoxia | 0
    autopsy | 0
    acute bronchopneumonia | 0
    organizing fibrinous pneumonia | 0
    right pulmonary artery thromboembolism | 0
    epithelioid hemangioendothelioma in lymphangitic and intraparenchymal distribution | 0
    death | 0
    