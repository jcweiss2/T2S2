73 years old | 0
    woman | 0
    hypertension | 0
    admitted to emergency department | 0
    melena | -24
    blood pressure 110/70 mmHg | 0
    heart rate 108 beats/min | 0
    body temperature 36.8 °C | 0
    respiratory rate 18 breaths/min | 0
    no pain complaint | 0
    no abdominal mass | 0
    red blood cell 2.51 × 1012/L | 0
    hemoglobin 8 g/dL | 0
    white blood cell count 21.75 G/L | 0
    89% neutrophils | 0
    prothrombin 80% | 0
    urea 14 mmol/L | 0
    creatinine 127 µmol/L | 0
    abdominal ultrasound | 0
    infrarenal AAA 33 × 46 mm | 0
    partially thrombosed 60 × 16 mm | 0
    esophagogastroduodenoscopy | 24
    small curvilinear ulcer | 24
    red scars | 24
    atrophic gastritis | 24
    colonoscopy | 24
    no bleeding point | 24
    diagnosed with moderate upper GI bleeding | 24
    gastric ulcer | 24
    resuscitated | 24
    intravenous fluid administration | 24
    350 mL red blood cells transfusion | 24
    350 mL platelets transfusion | 24
    proton pump inhibitor infusion | 24
    fasting | 24
    hemodynamic stability | 36
    no hematochezia | 36
    upper abdominal pain | 72
    dizziness | 72
    hypotension | 72
    systolic pressure 60 mmHg | 72
    heart rate 120 beats/min | 72
    SpO2 90% | 72
    gastric drainage with bright red blood | 72
    transferred to ICU | 72
    coma | 72
    second endoscopy | 72
    aggressive resuscitation | 72
    normal saline | 72
    700 mL packed red blood cells | 72
    500 mL fresh plasma | 72
    vasopressor | 72
    tracheal intubation | 72
    endoscopy with blood clots | 72
    inadequate gastric visualization | 72
    abdominal CT scan | 72
    infrarenal fusiform AAA 75 × 53 mm | 72
    25 mm thick anterior wall thrombus | 72
    ruptured into second part of duodenum | 72
    hemorrhage | 72
    aortoduodenal fistula | 72
    EVAR | 72
    3 stent graft components | 72
    plugging ruptured aneurysm with histoacryl | 72
    successful intervention | 72
    no contrast leak | 72
    died | 82
    multiple organ failure | 82
    reversible hypovolemic shock | 82
    