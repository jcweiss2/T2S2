73 years old | 0
male | 0
admitted to the hospital | 0
altered mental status | -72
feeling weak | -720
feeling lethargic | -720
agitated | 0
confused | 0
not oriented to person, place, or time | 0
febrile | 0
tachycardic | 0
hypotensive | 0
respiratory rate of 20/min | 0
oxygen saturation of 99% on room air | 0
multiple stage 3 to 4 draining ulcers | 0
bilateral lower-extremity +2 pitting edema | 0
leukocytosis | 0
bandemia | 0
dehydration | 0
elevated lactate | 0
urinary tract infection | 0
received a 4-liter bolus of normal saline | 0
maintenance at a rate of 250 ml/h | 0
broad-spectrum IV antibiotics | 0
vasopressors | 0
cardiac markers normal | 0
EKG revealed normal sinus rhythm with tachycardia | 0
echocardiography showed an ejection fraction of 55% | 0
mild diastolic dysfunction | 0
central venous pressure of 8 cmH2O | 0
transferred to the intensive care unit | 0
surgical debridement of the infected decubitus ulcer | 0
initial blood and wound cultures grew Streptococcus agalactiae | 0
urine culture grew Citrobacter amalonaticus | 0
WBC count slightly trended down | 0
lactic acid normalized | 0
Doppler studies showed an extensive right lower-extremity occluding thrombus | 0
started on a weight-based therapeutic dose of unfractionated heparin | 0
cell counts, PT, INR, aPTT and anti-Factor Xa activity were measured daily | 0
normal lab values for fibrinogen | 0
normal lab values for fibrinogen degradation product | 0
normal lab values for D-dimer | 0
continued to have altered consciousness | 0
remained hypotensive | 0
lab values remained stable | 0
significant drop in hemoglobin value | 72
heparin discontinued | 72
coagulopathy reversed with 2 units of fresh frozen plasma | 72
4 units of packed red blood cells were transfused | 72
hemoglobin remained steady at about 10 g/dL | 72
CT of the abdomen and pelvis showed a retroperitoneal hematoma | 72
expansion of the left iliopsoas musculature | 72
inferior vena cava filter placed | 96
no increase in size of the iliopsoas hematoma | 96
died on day 7 of hospitalization | 168
multi-organ failure | 168