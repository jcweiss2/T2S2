51 years old | 0
male | 0
motorcycle accident | 0
hemodynamic instability | 0
pelvic fracture | 0
catastrophic soft tissue injury | 0
scrotum injury | 0
perineum injury | 0
anus injury | 0
absent anal reflex | 0
extended EcoFast | 0
no fluid collection in abdomen | 0
no pneumothorax | 0
pelvis X-ray | 0
ischiopubic fracture | 0
ileopubic fracture | 0
symphyseal disruption | 0
anterior posterior fracture APII | 0
resuscitation | 0
full-body computed tomography | 0
pelvis fixed with external screws | 0
exploratory laparotomy | 0
exclude abdominal organ damage | 0
loop colostomy | 0
anal incompetence | 0
admitted to ICU | 0
no bowel function | -144
post-operative day 7 | 168
abdominal distension | 168
elevated inflammatory indices | 168
fever | 168
abdominal CT with oral and intravenous contrast | 168
intestinal obstruction | 168
dilated small bowel loops | 168
air/fluid levels | 168
ileum segment trapped in sacral fracture | 168
exploratory laparotomy | 168
small bowel resection | 168
end-to-end manual anastomosis | 168
second post-operative period uneventful | 168
discharged from ICU | 168
evaluation of rectal sphincter | 168
normal rectal sphincter function | 168
peroneal wound healed | 168
colostomy closed | 168
