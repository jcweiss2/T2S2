75 years old | 0
Hispanic | 0
male | 0
hypertension | -672
hyperlipidaemia | -672
nephrolithiasis | -672
right flank pain | -48
dysuria | -168
frequency | -168
admitted to the hospital | 0
antibiotics | 0
fluids | 0
emergency ureteral stent placement | 12
acute respiratory distress syndrome | 12
severe hypoxaemia | 12
intubated | 12
intravenous fluids | 12
vasopressors | 12
dopamine | 12
norepinephrine | 12
lactate | 12
vasopressin | 24
bluish discolouration | 48
capillary refill | 48
radial and dorsalis pedis pulses | 48
skin intact and cool to touch | 48
gangrenous changes | 72
intravenous argatroban | 72
dialysed | 72
fluid-filled bullae | 216
gangrenous changes | 216
discharged to a nursing home | 216
local wound care | 216
monitoring for gangrene demarcation | 216
necrosis of both feet | 720
left heel cellulitis | 720
intravenous antibiotics | 720
discharged | 726
left hand digits 1, 4 and 5 amputated | 1440
transmetatarsal amputations | 2160
Veraflow wound vacuum-assisted closure | 2170
split-thickness skin graft | 2880
recovery as an outpatient | 2880
full ambulation | 2880