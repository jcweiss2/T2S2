history of mucosal resection for early gastric cancer | -1000
history of partial resection for left lung cancer | -1000
collected knee-high wild grass from a riverbed for 10 days | -240
developed systemic pain and fatigue | -168
developed fever, chills, watery diarrhea, loss of appetite, and mildly disturbed consciousness | -168
visited the department of internal medicine at a nearby hospital | -14
hospitalized | 0
decreased white blood cells and platelet counts | 0
elevated hepatic enzyme levels | 0
referred to our department for further examination | 0
Glasgow Coma Scale of 14: E3, V5, M6 | 0
blood pressure of 130/79 mmHg | 0
heart rate of 96/min | 0
respiratory rate of 20/min | 0
O2 saturation of 94% | 0
temperature of 38.9°C | 0
crusted skin lesions on the medial surface of the left thigh | 0
freely movable adenopathy | 0
aggregated papules in the right inguinal region | 0
no remarkable head-and-neck or chest abnormalities | 0
no remarkable neurological abnormalities | 0
administered antibiotics | 24
elevated ferritin levels | 48
performed bone marrow biopsy | 48
diagnosed with HLH | 48
administered prednisolone | 48
developed chest pain, shivering, and fever | 72
elevated CK levels | 72
elevated LDH levels | 72
elevated high-sensitivity troponin I | 72
severe left ventricular dysfunction | 72
ST elevation in the V1-2 leads | 72
suspected acute myocarditis | 72
moved to negative-pressure room | 72
submitted serum and urine samples and throat swabs to a responsible public health center | 72
RT-PCR analysis detected SFTSV RNA | 96
infected cells stained positively by an anti-SFTSV-nucleoprotein antibody | 96
withdrew from circulatory agonist and ventilator management | 336
ECG showed improvement of ST elevation | 336
re-submitted serum and confirmed negativity for viremia | 408
released from quarantine | 408
performed CAG and EMB | 576
pathological evaluation of the EMB specimen revealed myocardial inflammation | 576
discharged | 696
follow-up visit | 744
transthoracic echocardiography showed a slight improvement | 744
no heart failure | 744