73 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
hypertension | 0 | 0 | Factual
syphilis | 0 | 0 | Factual
type 2 diabetes mellitus | 0 | 0 | Factual
mechanical fall | -720 | -720 | Factual
pruritic scalp | -720 | 0 | Factual
purulent drainage from sinuses on the scalp | -720 | 0 | Factual
altered mental status | 0 | 0 | Factual
temperature of 97.9°F | 0 | 0 | Factual
heart rate of 127 bpm | 0 | 0 | Factual
respiratory rate of 22 breaths/min | 0 | 0 | Factual
blood pressure of 144/80 mmHg | 0 | 0 | Factual
oxygen saturation of 98% on room air | 0 | 0 | Factual
oriented to person and place, but not to time | 0 | 0 | Factual
face, scalp and right ear were erythematous and edematous | 0 | 0 | Factual
large fluctuant mass with purulent drainage over the occipital and parietal portions of the scalp | 0 | 0 | Factual
posterior auricular mass without signs of active drainage | 0 | 0 | Factual
hyperglycemia to 700 | 0 | 0 | Factual
anion gap metabolic acidosis with serum bicarbonate of 20 | 0 | 0 | Factual
ketonuria | 0 | 0 | Factual
non-contrast head computed tomography (CT) showed extensive multifocal scalp swelling | 0 | 0 | Factual
admitted to the intensive care unit | 0 | 0 | Factual
diabetic ketoacidosis | 0 | 0 | Factual
cellulitis of the scalp | 0 | 0 | Factual
concern for underlying abscesses | 0 | 0 | Possible
continuous infusion of insulin | 0 | 720 | Factual
intravenous Vancomycin | 0 | 720 | Factual
intravenous Cefepime | 0 | 720 | Factual
incision and drainage of scalp lesion | 48 | 48 | Factual
10-cm subgaleal abscess with large amounts of purulence evacuated | 48 | 48 | Factual
initial admission blood cultures grew MRSA | 72 | 72 | Factual
paranasal sinus CT with intravenous contrast did not show involvement | 72 | 72 | Factual
transesophageal echocardiogram without evidence for endocarditis | 72 | 72 | Factual
pulse irrigation of the wounds | 96 | 120 | Factual
sharp debridement | 96 | 120 | Factual
serial bedside debridements | 96 | 720 | Factual
scalp wound ultimately measured 20 cm in length, 10 cm in width and 2 cm depth | 120 | 720 | Factual
right posterior auricular wound measured 7 × 7 × 2 cm | 120 | 720 | Factual
split-thickness skin grafts harvested from the right thigh | 120 | 120 | Factual
100% take of the grafts on postoperative day 7 | 168 | 168 | Factual
discharged on hospital day 32 | 768 | 768 | Factual
intravenous Vancomycin to complete a full 7-week course | 768 | 1008 | Factual