78 years old | 0
woman | 0
requested re-fabrication of upper and lower partial dentures | 0
hypertension | -4320
hyperlipidemia | -4320
renal calculi | -4320
trichlormethiazide | -4320
warfarin potassium | -4320
fluvastatin sodium | -4320
blood pressure within normal ranges | 0
lipid levels within normal ranges | 0
renal calculi within normal ranges | 0
re-fabrication of lower partial dentures | -4320
re-fabrication of upper partial dentures planned | -4320
intense instability (tooth mobility level 3) in upper left molar region | -4320
marked alveolar bone resorption | -4320
spontaneous pain in upper left molar region | -144
swelling in upper left molar region | -144
pus discharge from periodontal pocket | -144
cleaned and sterilized with normal saline solution | -144
iodo-glycol paste | -144
loxoprofen sodium prescribed | -144
swelling spread to left buccal region | -144
spontaneous pain became more intense | -144
difficulty while eating for 2–3 days | -144
referred to visit hospital | -72
Glasgow Coma Scale score 11 | 0
facial pallor | 0
cold hands and fingers | 0
shivering | 0
weak radial artery pulse | 0
axillary temperature 41°C | 0
systolic blood pressure 80–90 mmHg | 0
diastolic blood pressure 40–50 mmHg | 0
pulse rate 130–160 bpm | 0
SpO2 75%–85% | 0
dehydration suspected | 0
septic shock suspected | 0
oxygen administration at 10 L/min initiated | 0
venous line secured to cubital fossa | 0
blood drawn for rapid blood examination | 0
drip infusion of acetate linger solution 500 mL | 0
normal saline solution 100 mL | 0
ampicillin sodium 2 g | 0
albumin 2.3 g/dL | 0
sodium 127 mEq/L | 0
white blood cell count 29,830/µL | 0
C-reactive protein levels 22.86 mg/dL | 0
improvement after venous infusion of antibacterial drugs | 0
Glasgow Coma Scale score 14 | 0
axillary temperature 38.5°C | 0
systolic blood pressure 120–130 mmHg | 0
diastolic blood pressure 80–90 mmHg | 0
pulse rate 120–140 bpm | 0
SpO2 100% | 0
transferred to nearby general hospital | 24
D-dimer 23.98 µg/mL | 24
fibrin degradation products 38.6 µg/mL | 24
disseminated intravascular coagulation (DIC) suspected | 24
systemic management in intensive care unit | 24
condition worsened | 48
death confirmed | 72
pleural effusion | 72
pulmonary infiltration | 72
pulmonary shadows | 72
possible lung cancer | 72
no histopathological testing | 72
no pathological autopsy | 72
informed consent obtained | 72
septic shock symptoms caused by infectious dental disease | 0
emergency treatment | 0
death the following day | 24
periodontal abscess | -144
gram-negative anaerobic bacteria spread | -144
alveolar abscess requiring prompt medical intervention | -144
rapid progression from dental infection to dehydration and septicemia | -144
decreased immune function related to age | -4320
accompanying malnutrition | -4320
high mortality rate associated with infection | -4320
oral cavity as source of infection | -144
complications of diabetes or malignant neoplasms | -4320
chronic lymphocytic leukemia | -4320
malignant neoplasm possibility | -4320
early intensive treatment | 0
no improvement of symptoms | 0
asymmetric dimethylarginine (ADMA) association | -4320
soluble urokinase-type plasminogen activator receptor (suPAR) association | -4320
Aggregatibacter actinomycetemcomitans (AA) association | -4320
infection worsens prognosis in HIV-positive patients | -4320
follow-up of patients with oral implants | -4320
biomaterial to cover wound surface | -4320
implant placement techniques | -4320
life-threatening periodontal abscess | 0
decreased immune function | -4320
suboptimal nutritional state | -4320
various systemic complications | -4320
oral infections prone to develop into septicemia or DIC | -144
administration of antibacterial drugs | 0
local and systemic states confirmation | 0
daily sterilization | 0
co-operation of medical department sought | 0
