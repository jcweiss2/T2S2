Here is the extracted table of events and timestamps:

63 years old | 0
female | 0
168 cm height | 0
53 kg weight | 0
papillary thyroid carcinoma | -9720
resection | -9720
radiotherapy | -9720
stenosis of the esophagus | -7200
repeated aspiration | -7200
respiratory insufficiency | -7200
pneumonia | -7200
purulent pleurisy | -7200
pleurectomy | -7200
restrictive ventilation pattern | -7200
recurrent nerve palsy | -7200
percutaneous endoscopic gastrostomy | -7200
tracheostoma | -7200
home ventilation | -7200
mobility decreased | -4320
secondary depression | -4320
mandible nearly fixed | -4320
cannot open mouth over 20 degrees | -4320
left axis vertebralis stented | -2190
stenosis of the internal axis carotis | -2190
arterial hypertension | -2190
secondary lactase deficiency | -2190
esophageal stenosis dilated | -720
fistula between esophagus and tracheal membrane | -720
decreasing general condition | -720
referred to University of Erlangen | -720
examined by several chiefs and consultants | -720
deemed too unstable for open surgery | -720
inability to open mouth | -720
recurrent nerve palsy | -720
minimal invasive orthograde approach impossible | -720
referred to hospital on surgical intensive care unit | -720
pneumonia by 4-multiresistente gramnegative Pseudomonas aeruginosa | -720
veno-venous extracorporeal membrane oxygenation (vv-ECMO) | -720
partial thromboplastin time of 60 seconds | -720
preseptic status | -720
ventilated through tracheostoma with low ventilation forces | -720
thoracic computed tomography | -720
big fistula of the tracheal membrane | -720
tracheal cannula ended shortly beneath lower limit of mediastinal fistula | -720
decision to try endobronchial stenting | -720
plan to close fistula with pedicled omentum majus replacement | -720
surgical plastic needed abutment and secured continuous airway replacement | -720
procedure performed | -24
vv-ECMO began to be partly ineffective | -24
high volume input of physiological saline needed | -24
oral approach only allowed small flexible bronchoscope | -24
approach for upper part of trachea had to be performed through percutaneous tracheostoma | -24
trying different Dumon and one-hybrid self expandable metalic y-stent | -24
plan to changeover to more floppy Freitag stent (FS) | -24
successful retrograde stenting performed in four steps | -24
Step I | -24
manually compressed “y” of FS pushed downward on main carina | -24
Step II | -24
frontal surface of stent cut with at least 1 cm opening in longitudinal axis | -24
stent surface reduced ~40% in sagittal axis | -24
new stoma for regular tracheal cannula created | -24
lower new edge of stoma fixed subcutaneously | -24
Step III | -24
jagwire introduced through mouth into trachea | -24
jagwire running out of new FS stoma | -24
soft-tip stiff DLET introduced for more stability | -24
DLET dragged out of new stoma of cut FS | -24
distal jagwire introduced into oral orifice of FS | -24
FS flipped with upper part over soft-tip stiff DLET into upper third of trachea | -24
whole fistula bridged by FS up to level of vocal cords | -24
upper edge of new FS stoma fixed subcutaneously | -24
Step IV | -24
regular tracheal cannula introduced for ventilation | -24
lungs not aerated at that point of time | -24
spontaneous breathing work increased | 24
vv-ECMO support reduced | 24
lungs became re-aerated again | 24
patient woke up again | 24
patient could communicate with family by writing and eyes | 24
infections continued to be very severe | 24
spontaneous work of breathing never exceeded tidal ventilation of 170 mL per breath | 24
reduction of intravenous saline injection limited | 24
vv-ECMO support mandatory but reduced | 24
patient and family decided to actively reduce vv-ECMO support | 48
patient died | 72