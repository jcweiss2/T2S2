65 years old | 0
male | 0
admitted to hospital | 0
chest pain | 0
shortness of breath | 0
history of smoking | -8760
history of hypertension | -8760
on antihypertensive medication | -8760
mild chest discomfort | -48
ECG showed ST-segment elevation | 0
elevated troponin levels | 0
diagnosed with AMI | 0
underwent PCI with stent placement | 24
started on dual antiplatelet therapy | 24
developed fever | 72
diagnosed with sternal wound infection | 72
treated with intravenous antibiotics | 72
condition stabilized | 240
discharged | 240
advised to quit smoking | 240
advised to manage hypertension | 240