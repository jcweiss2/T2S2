2 years old | 0
female | 0
born full term | 0
spontaneous vaginal delivery | 0
prolonged obstructive jaundice | 0
steatorrhea | 0
generalized itchiness | 0
ultrasound abdomen | 0
contrast-enhanced computed tomography scan | 0
choledochol cyst | 0
scheduled for portoenterostomy | 0
liver biopsy | 0
on-table cholangiogram | 0
caudal epidural catheter insertion | 0
Perifix ONE Paed | 0
skin to space distance 1.5 cm | 0
left lateral position | 0
catheter advanced 10 cm | 0
minimal twisting | 0
T7 dermatome | 0
ultrasound guidance used | 0
confirm cephalad movement of catheter tip | 0
surgery | 0
extubated | 24
discharged to ward | 24
epidural infusion functioning well | 24
continuous infusion 2-4 ml/h | 24
pain well-controlled | 24
epidural catheter removal planned | 48
resistance encountered during removal | 48
full flexion of trunk | 48
repositioned to extension | 48
epidural catheter fell off | 48
end segment sheared off | 48
6 cm left inside space | 48
segment twisted | 48
segment crimped | 48
segment fractured | 48
no remnant around skin area | 48
informed surgeon | 48
informed parents | 48
urgent MRI thoracolumbar | 48
non-contrast CT scan spine | 48
CT scan showed retained catheter tip | 48
retained from upper border of L4 | 48
posterior part of thecal sac at S4 | 48
retained segment approximately 6 cm | 48
no other remnant in thoracic region | 48
no other remnant in lumbar region | 48
persistent vomiting | 72
fever | 72
total white count increased from 17.15 to 23x10^9/L | 72
no neurological deficit | 72
differential diagnosis includes laparotomy pathology | 72
differential diagnosis includes sepsis | 72
differential diagnosis includes retained catheter tip | 72
CT brain urgent | 72
normal finding | 72
no mass effect | 72
no hydrocephalus | 72
repeated CT scan spine | 72
no catheter migration | 72
no abnormal findings | 72
no focal swelling | 72
no collection | 72
fever subsided | 72
vomiting persists | 72
relaparotomy on postoperative day 18 | 432
adhesions found | 432
adhesiolysis | 432
small bowel resection | 432
side-to-side anastomosis | 432
extubated on second postoperative day | 456
discharged home 9 days after re-laparotomy | 576
asymptomatic | 576
risk of surgery high | 576
decided to leave fragment in situ | 576
follow-up | 576
advised parents to report symptoms | 576
clinic review over past year | 8784
no symptoms of complication | 8784
generalized itchiness |>
