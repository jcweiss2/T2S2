40 years old | 0
female | 0
161 cm | 0
67 kg | 0
36 and 6/7 weeks gestation | 0
placenta previa totalis | 0
Cesarean section | 0
myomectomy | -7560
myoma in the low portion of uterus | -7560
preoperative laboratory tests were normal | 0
invasive arterial blood pressure monitoring | 0
anesthesia induced with thiopental sodium | 0
anesthesia induced with succinylcholine | 0
intubation | 0
anesthesia maintained with sevoflurane | 0
anesthesia maintained with nitrous oxide | 0
volume-controlled mode with 50% oxygen | 0
electrocardiogram monitoring | 0
BIS monitoring | 0
pulse oximetry | 0
ventilator set to end-tidal carbon dioxide partial pressure 30-35 mmHg | 0
atracurium injected intravenously | 0
baby delivered | 9
Apgar scores at 1 and 5 min were 8 and 9 points | 9
no complications with the fetus | 9
bleeding observed in the uterus at placental attachment sites | 109
methyl ergonovine injected intravenously | 109
central venous catheter inserted | 109
packed RBCs administered | 109
vital sign remained stable | 109
surgeon finished the uterine suture | 100
EtCO2 partial pressure dropped | 100
blood pressure dropped | 100
ventricular fibrillation appeared | 100
chest compression started | 100
defibrillation attempted | 100
epinephrine injected | 100
atropine injected | 100
bicarbonate injected | 100
cardiac compression continued | 100
BIS values maintained above 40 | 100
systolic blood pressure maintained at approximately 60-100 mmHg | 100
arterial oxygen saturation was 86% | 100
blood-like secretion exited the endotracheal tube | 100
EtCO2 partial pressure checked as apnea | 100
cardiac compression attempted for 40 min | 100
defibrillation performed three times | 140
epinephrine 60 mg injected | 140
atropine 5 mg injected | 140
bicarbonate 120 mEq injected | 140
calcium chloride 1,200 mg injected | 140
corrugating tube exchanged five times | 140
EtCO2 partial pressure monitoring stopped | 140
manual ventilation maintained with 100% oxygen | 140
return of a normal sinus rhythm | 150
blood pressure was 90/50 mmHg | 150
heart rate was 110 beats/min | 150
mannitol 100 ml injected | 150
lasix 20 mg injected | 150
methylprednisolone 500 mg injected | 150
obstetricians completed the operation | 150
no urine output during CPR | 150
urine excreted at a rate higher than 200 ml/hour | 150
vaginal bleeding developed | 170
heart rate increased to 120-130 beats/min | 170
hysterectomy performed | 170
transesophageal echocardiography probe inserted | 170
thrombus in the heart not found | 170
global hypokinesia in the left ventricle | 170
platelet count of 39,000 | 170
prothrombin time of 28.6 sec | 170
activated partial thrombin time of 129.1 sec | 170
fibrinogen at 60 mg/dl | 170
d-dimer > 20 µg/ml | 170
disseminated intravascular coagulation suspected | 170
3 units of whole blood transfused | 170
10 units of pack cells transfused | 170
20 units of platelets transfused | 170
10 units of fresh frozen plasma transfused | 170
total anesthesia time was 8 hours and 40 minutes | 520
patient transferred to the intensive care unit | 520
chest radiography showed pulmonary edema | 520
treated with transfusion and fluid therapy | 520
recovered to a drowsy state | 580
responded to pain stimulation | 580
pulmonary edema showed a slight improvement | 620
transthoracic echocardiography revealed no obvious regional wall motion abnormality | 620
returned to an alert mental state | 700
cooperative | 700
extubation performed | 700
vital signs were stable | 700
pH 7.605 | 700
PaCO2 25.3 mmHg | 700
PaO2 98.5 mmHg | 700
HCO3- 24.6 mmol/L | 700
SaO2 98.4% | 700
hemoglobin 9.9 g/dl | 700
platelet 108,000 | 700
PT/aPTT, 16.6/48.5 sec | 700
fibrinogen 263 mg/dl | 700
d-dimer 4.51 µg/ml | 700
experienced a sudden loss of consciousness | 730
cardiac arrest developed | 730
defibrillation performed | 730
mental state and heart rhythm recovered | 730
tachyarrhythmia and cardiac arrest | 790
multi-organ failure | 1180
extracorporeal membrane oxygenation | 1180
continuous renal replacement therapy | 1180
died | 1440