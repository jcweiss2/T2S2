58 years old | 0
male | 0
admitted to the hospital | 0
sore throat | 0
COVID-19 | 0
moderate pneumonia | 0
oxygen therapy | 0
glucocorticoids | 0
increased oxygen requirements | -17
worsened pneumonia | -17
severe respiratory fatigue | -17
acute respiratory distress syndrome (ARDS) | -17
hypertension | -672
intubation | -17
mechanical ventilation | -17
tocilizumab | -17
venovenous ECMO | -17
prone position | -17
computed tomography (CT) | -17
bilateral and peripheral ground-glass and consolidative pulmonary opacities | -17
intra-abdominal bleed | -9
hypotension | -9
right hemicolectomy | -9
ileostoma creation | -9
ischemic changes | -18
stomal reconstruction | -18
necrotic changes | -18
repeated debridement | -18
Mucorales infection | -18
thrombi | -18
vessel thrombosis | -18
tissue necrosis | -18
multi-organ failure | -46
death | -46
autopsy | -46
necrosis of reconstructed stoma | -46
necrosis of skin | -46
necrosis of abdominal wall muscles | -46
thrombus in common iliac vein | -46
necrosis of multiple abdominal organs | -46
Rhizopus oryzae infection | -46
histopathological examination | -46
immunohistochemical analysis | -46
cytomegalovirus infection | -46
sepsis | -46
disseminated mucormycosis | -46
COVID-19-associated mucormycosis | -46
early suspicion and diagnosis | 0
treatment | 0
better outcomes | 0
increased risk of mucormycosis | 0
uncontrolled diabetes mellitus | 0
steroids | 0
numerous cytokines during ARDS | 0
drugs such as lopinavir, ritonavir, and remdesivir | 0
glucocorticoid use | 0
surgical stress | 0
ARDS | 0
mucormycosis | 0
systemic dissemination | 0
routine serological tests | 0
histopathological examination | 0
antigen-antibody reactions | 0
beta-D-glucan test | 0
cell-free DNA next-generation sequencing | 0
posaconazole | 0
liposomal amphotericin B | 0
quantitative polymerase chain reaction examination | 0
novel serum-based techniques | 0
better outcomes in patients with systemic mucormycosis | 0
initiation of treatment | 0
tissue necrosis | 0
disseminated mucormycosis | 0
rare report | 0
autopsy for disseminated COVID-19-associated mucormycosis | 0
flowchart of autopsy diagnosis | 0
opportunistic infections triggered by COVID-19 | 0
critical problem | 0
delayed diagnosis | 0
mucormycosis | 0
increased risk | 0
COVID-19 patients | 0
early suspicion | 0
timely diagnosis | 0
treatment | 0
better outcomes | 0
affected individuals | 0