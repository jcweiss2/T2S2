80 years old | 0
male | 0
admitted to the hospital | 0
septic shock | 0
P. aeruginosa necrotizing CAP | 0
bacteremia | 0
three day history of severe right sided chest pain | -72
dyspnea | -72
fever | -72
denies any use of alcohol | 0
denies any use of tobacco | 0
hypertension | -504
hypothyroidism | -504
calcified pleural plaques | -504
autoimmune hemolytic anemia (AIHA) | -504
treated with oral prednisone 70 mg daily | -504
negative HIV | -504
negative hepatitis B | -504
negative hepatitis C | -504
antinuclear antibodies were positive | -504
anti double-stranded DNA titer 1:360 | -504
plasma protein electrophoresis was normal | -504
Positron emission tomography (PET) scan was normal | -504
chest-abdomen-pelvis computed tomography (CT) was normal | -504
dyspneic | 0
respiratory rate of 27 breaths/min | 0
heart rate of 93 beats/ min | 0
fever of 39 °C | 0
lung auscultation was negative for crackles | 0
hypotensive | 0
blood pressure of 80/60 mmHg | 0
required vasopressor support with norepinephrine | 0
leukocytosis | 0
white blood cell count of 27,100/mm3 | 0
hemoglobin level of 14.5 g/dL | 0
platelet count of 187,000/mm3 | 0
arterial blood gas showed pH of 7.48 | 0
PaO2 of 62 mmHg | 0
PaCO2 of 35 mmHg | 0
C-reactive protein (CRP) was elevated at 130 mg/L | 0
acute kidney injury | 0
creatinine at 1.386 mg/dL | 0
lactic acid was elevated to 31.53 mg/dL | 0
procalcitonin (PCT) was increased to 14.6 ng/mL | 0
blood cultures were obtained | 0
pneumococcal and Legionella urine antigens were negative | 0
pulmonary consolidation in the right upper lobe (RUL) with a cavity | 0
RUL consolidation associated with septated cavitation | 0
empiric antimicrobial therapy was started with intravenous (IV) cefotaxime 2 g x 3 daily | 0
IV levofloxacin 500 mg twice daily | 0
blood cultures became positive for pan-sensitive P. aeruginosa | 24
antimicrobials were changed to IV cefepime 2 g over eight hours twice daily | 24
bronchoscopy with bronchoalveolar lavage (BAL) | 48
positive culture of P. aeruginosa at the concentration of 105/mL | 48
respiratory strain susceptibility pattern was identical to the blood culture | 48
acid-fast bacilli stain was negative | 48
clinical condition improved on IV cefepime | 48
vasopressor was rapidly weaned | 48
oxygen therapy was stopped | 96
transferred out of the ICU to the pulmonology floor | 120
discharged from the hospital | 504
repeat chest x-ray at 2 weeks showed dramatic decrease of the pulmonary consolidation | 336
residual 10 cm cavity | 336