24 years old | 0
    female | 0
    primigravida | 0
    gestational age 26 weeks | 0
    referred | -720
    persistent abdominal pain | -720
    recurrent vaginal bleeding | -720
    admitted repeatedly | -720
    abdominal pain | -720
    denied previous pelvic inflammatory disease | 0
    denied intrauterine contraceptive device use | 0
    denied pelvic surgery | 0
    abruptio placenta suspected | -720
    induced with oxytocin | -720
    transferred | -24
    arrival | 0
    conscious | 0
    severe pain | 0
    pale | 0
    afebrile | 0
    distended abdomen | 0
    uterine fundus 30 cm | 0
    generalized tenderness | 0
    fetal heartbeats not detected | 0
    closed cervix | 0
    uneffaced cervix | 0
    firm cervix | 0
    posterior cervix | 0
    presenting part not found | 0
    transabdominal ultrasound | 0
    live intrauterine diamniotic-dichorionic twins | 0
    estimated gestational age 26 weeks | 0
    enlarged cystic placentas | 0
    retro-placental clots | 0
    hemoglobin 7.0g/dl | 0
    blood group A | 0
    Rhesus positive | 0
    concealed abruptio placenta | 0
    live twin pregnancy | 0
    emergency abdominal delivery | 0
    laparotomy | 0
    thickened peritoneum | 0
    hematoma | 0
    cystic mass | 0
    normal-sized intact uterus | 0
    pregnant sac engulfed by thickened omentum | 0
    normal fallopian tubes | 0
    normal ovaries | 0
    live female twins extracted | 0
    placenta attached to ceacum | 0
    placenta attached to ascending colon | 0
    placenta adhered to posterior aspect of omentum | 0
    placenta adhered to transverse colon | 0
    placenta adhered to sigmoid colon | 0
    profuse bleeding | 0
    ligation of placental blood vessels | 0
    placentas left in situ | 0
    umbilical cords cut | 0
    estimated blood loss 2000ml | 0
    transfused 4 units of whole blood | 0
    first twin weight 700g | 0
    second twin weight 800g | 0
    Apgar score 5 at first minute | 0
    Apgar score 6 at fifth minute | 0
    no congenital abnormalities | 0
    admitted to neonatal intensive care unit | 0
    babies died | 168
    covered with broad spectrum antibiotics | 0
    admitted to intensive care unit | 0
    septicemia | 72
    treated with meropenem | 72
    improved | 72
    discharged | 336
    readmitted | 504
    peritonitis | 504
    repeat laparotomy | 504
    attempt to remove placentas | 504
    massive hemorrhage | 504
    controlled by intra-abdominal packing | 504
    transfused 3 units of blood | 504
    abdominal packs removed | 552
    no active bleeding | 552
    fascial dehiscence | 624
    taken to operating room | 624
    placentas detached without bleeding | 624
    postoperative recovery | 624
    discharged | 744
    outpatient follow-up | 744
    three visits | 2448
    discharged from clinic | 2448
    good condition | 2448
    