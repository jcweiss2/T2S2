multiple blisters and erosions all over body | -156
superadded maggot infection | -156
previous episodes of lesions | -312
lesions subsided after treatment with steroids | -156
lesions developed all over body | -156
febrile | 0
numerous flaccid blisters and erosions | 0
Nikolsky sign strongly positive | 0
diagnosis of PV confirmed by skin biopsy | 0
tzanck smear | 0
IV dexamethasone pulse | 0
supportive care | 0
IV antibiotics | 0
adjuvant immunosuppressors held back | 0
oozing from skin ulcerations | 24
hemorrhagic excoriation | 24
peeling of skin | 24
oral methyl prednisolone | 72
hypoproteinemia | 168
pleural effusion | 168
blood culture showed enterobacter | 168
pus culture from erosions showed Staphylococcus aureus and Proteus mirabilis | 168
intravenous Tigecycline and vancomycin | 168
sepsis | 168
high grade fever | 168
albumin levels fell | 168
TPE planned | 216
TPE performed | 216
Nikolsky sign became negative | 240
no new lesions appeared | 240
exudation from lesions reduced | 240
dressings started to remain dry | 240
lesions showed re-epithelization | 240
lesions showed healing | 288
oral lesions healed completely | 288
little erosions on back, anterior aspect of thigh and buttocks persisted | 288
IV methyl prednisolone pulse | 288
cyclophosphamide | 288
patient clinically stable | 312
plan for one more TPE cycles | 312
patient discharged | 336
monthly IV dexamethasone pulse | 336
daily oral prednisolone | 336