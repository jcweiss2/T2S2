38 years old | 0
male | 0
admitted to the hospital | 0
long-term problems with food intake | -5040
previous surgery for congenital pylorostenosis | -52560
native X-ray | -672
ultrasound examination | -672
computed tomography (CT) scan | -672
suspicion of gastrostasis | -672
suspicion of recurrent pylorostenosis | -672
contrast-enhanced examination of upper gastrointestinal tract | -672
barium sulphate as contrast agent | -672
stenosis of the pylorus | -672
gastrostasis | -672
stasis of all contrast agent in the stomach | -672
benign stenosis of the pylorus | -672
scheduled for planned surgical intervention | -672
unplanned return to surgeon’s office | -120
substantial and increasing pain in left epigastrium | -120
left epigastric region tender | -120
pain on palpation | -120
X-ray examination | -120
stasis of large amount of contrast agent in the stomach | -120
inflammation parameters not elevated | 0
CRP 0.3 mg/L | 0
procalcitonine 0.086 µg/L | 0
admitted to surgery ward | 0
nasogastric tube inserted | 0
unsuccessful attempt to evacuate contrast agent | 0
condition deteriorated | 24
immediate laparotomy indicated | 24
tumorous lesion on pylorus | 24
diameter 5 cm | 24
dilated stomach | 24
adhesions | 24
precipitated and sedimented barium sulphate | 24
BII partial stomach resection | 24
histological examination | 24
Roux-en-Y gastrojejunal anastomosis | 24
repeated lavage of peritoneal cavity | 24
Tygon tube 27 drainage inserted | 24
moved to central intensive care unit | 24
intense antibiotics therapy | 24
infusions | 24
nutritional support | 24
condition worsened | 48
elevation of inflammation markers | 48
CRP 78.9 mg/L | 48
procalcitonine 4.45 µg/L | 48
suspected leak of anastomosis | 48
suspected contrast agent spillage | 48
suspected peritonitis | 48
CT scan | 48
no contrast agent spillage intraperitoneally | 48
no anastomosis failure | 48
methylene blue administered | 48
no methylene blue in drained exudate | 48
drainage bags contained sanguinolent fluid | 48
CT exam on third day | 72
small amount of contrast agent in paragastric intraperitoneal region | 72
same amount of contrast agent next to stomach | 72
active leak not suspected | 72
worsening laboratory results | 72
CRP 267.60 mg/L | 72
procalcitonine 25.90 µg/L | 72
sepsis suspected | 72
patient remained afebrile | 72
anastomosis dehiscence unconfirmed | 72
antibiotic therapy revised | 72
vasopressor support introduced | 72
condition improved | 96
amount of exudate drained significantly lower | 96
surgical wound dehiscent and phlegmonous | 96
local therapy applied | 96
condition improving further | 168
stools being passed | 168
vasopressors discontinued | 168
inflammation parameters improved | 168
CRP 78.60 mg/L | 168
procalcitonine 2.85 µg/L | 168
two weeks after surgery | 336
CRP 13.80 mg/L | 336
discharged | 336
histological exam confirmed malignant stenosis of pylorus | 336
moderately differentiated adenocarcinoma | 336
resection margin positive for carcinoma | 336
repeated resection indicated | 336
revision of anastomosis | 336
surgical wound healed per secundam | 336
referred to department of clinical oncology | 336
chemotherapy initiated | 336
PET/CT exam on July 9, 2018 | 336
no metastatic lesions | 336
