42 years old | 0
male | 0
extensive alcohol abuse | 0
fatty liver disease | 0
admitted to the hospital | 0
acute necrotizing pancreatitis | 0
catheter-guided implantation of a self-expanding nitinol stent | -336
sigmoid colon perforation | -336
resection of sigmoid colon | -320
transversostoma application | -320
extubated | -304
white blood cell count increased | -288
C-reactive protein levels increased | -288
new onset of fever | -288
computed tomography (CT) performed | -240
peripancreatic abscess | -240
CT scan | -216
CT-guided percutaneous catheter | -168
drained brownish, partly solid pus | -168
Candida albicans detected | -144
Bordetella hinzii detected | -144
deep skin swab sample taken | -144
B. hinzii detected in skin swab | -144
Staphylococcus epidermidis detected | -120
B. hinzii detected again | -120
16S ribosomal RNA gene sequencing | -120
antimicrobial susceptibility testing | -120
cefotaxime resistant | -120
levofloxacin resistant | -120
trimethoprim/sulfamethoxazole resistant | -120
piperacillin/tazobactam susceptible | -120
ceftazidime susceptible | -120
meropenem susceptible | -120
tigecycline susceptible | -120
empirical therapy initiated | -168
piperacillin/tazobactam administered | -168
allergic skin reactions | -168
therapy switched to meropenem | -160
allergic skin reactions | -160
levofloxacin administered | -144
anaphylactic reaction | -144
tigecycline initiated | -136
defervescence | -120
reduction of drained secretion | -120
intravenous tigecycline stopped | -96
whole genome sequencing | -96
genetic relation elucidated | -96
core genome multilocus sequence typing | -96
genetic distance compared | -96
no acquired antimicrobial resistance genes | -96
discharged | 0