58 years old | 0
male | 0
pancreatogenic diabetes | 0
cholecystectomy | 0
admitted to the emergency room | 0
severe episodes of bright red blood stool | -48
abdominal pain | -48
difficulty breathing | -48
dehydrated | 0
tachycardic | 0
hypotensive | 0
confused | 0
severe anemia | 0
lactate 5 mmol/L | 0
bicarbonate 12 meq/L | 0
creatinine level 3.5 mg/dl | 0
mildly elevated liver chemistries | 0
normal coagulation profile | 0
admitted to the intensive care unit | 0
treated with vigorous volume resuscitation | 0
transfused 4 units of blood | 0
vasopressors | 0
colonoscopy | 0
inconclusive colonoscopy | 0
enhanced abdominal computed tomography | 0
10 × 11 mm aneurysm of the left colic artery | 0
angiography | 0
transcatheter arterial embolization | 0
bleeding controlled | 0
improved | 0
vasopressors phased out | 0
discharged | 48
high fever | 336
acute abdominal pain | 336
diffuse abdominal tenderness | 336
leukocytosis | 336
neutrophilia | 336
elevated C-reactive protein | 336
increased levels of serum procalcitonin | 336
contrast-enhanced abdominal CT | 336
enlarged spleen | 336
hypodense low-density lesion filled with gas | 336
free liquid in the abdomen | 336
surgery | 336
laparotomy | 336
1000 cc of purulent fluid | 336
necrosis and purulent discharge | 336
extensive lavage of the peritoneal cavity | 336
splenectomy | 336
drain left in place | 336
readmitted to the ICU | 336
Escherichia coli identified | 336
10-day scheme of carbapenems | 336
recovered | 360
pathology reported extensive necrosis of the splenic tissue | 360
spleen abscess | 360
postoperative course uneventful | 360
discharged | 432
full diet initiated | 432
drain removed | 432
low and serous output | 432
doing well on follow-ups | 720