68 years old | 0
female | 0
admitted to the hospital | 0
metastatic adenocarcinoma of the ampulla of Vater | 0
pancreaticoduodenectomy and lymphadenectomy | 0
central venous catheter placement | 0
drains placement | 0
bile culture positive for Enterococcus faecalis | 24
bile culture positive for Klebsiella pneumoniae | 24
bi-antibiotherapy with meropenem and vancomycine | 24
fever | 528
shivering | 528
blood cultures drawn | 528
blood cultures negative | 592
blood cultures drawn from central venous catheter | 552
blood cultures positive | 624
microscopic examination of blood cultures | 624
unusual fungal elements | 624
treatment with intravenous fluconazole | 624
treatment switched to liposomal amphotericin B | 648
central venous catheter withdrawn | 552
control blood cultures negative | 576
septic shock | 648
blood cultures positive to Candida albicans | 648
blood cultures positive to Candida glabrata | 648
transferred to intensive care unit | 648
evolution favorable | 720
admitted back to digestive surgery unit | 720
liposomal amphotericin B continued | 720
identification of Pseudozyma aphidis | 720
sequencing of ITS region | 720
susceptibility testing | 720
MIC values | 720
treatment with liposomal amphotericin B successful | 1008
discharged | 1008