44 years old | 0
male | 0
hypothyroidism | 0
bronchial asthma | 0
low mood | -2160
anxiety | -2160
increasing social withdrawal | -2160
difficulty sleeping | -2160
change in employment status | -2160
brain biopsy left frontal lesion | -2160
craniotomy | -2160
discharged home | -2160
dexamethasone | -2160
weaker right side | -960
weakness worse in right leg | -960
behavioral changes initial | -2880
readmitted | -480
denied fever | 0
denied weight loss | 0
denied night sweats | 0
denied nausea | 0
denied vomiting | 0
denied raw milk ingestion | 0
denied smoking | 0
denied drug use | 0
denied alcohol use | 0
contact with sick cats | 0
normal higher mental functions | 0
normal language | 0
normal speech | 0
normal cranial nerve function | 0
minimally spastic muscle tone right-sided limbs | 0
weak elbow flexion right side | 0
weak wrist flexion right side | 0
0/5 power right lower limb | 0
normal power left side | 0
normal reflexes | 0
stand with support | 0
sit with support | 0
normal complete blood count | 0
normal differential | 0
brain MRI multiple intracranial focal mass lesions | 0
rim enhancement | 0
restricted diffusion periphery | 0
perilesional vasogenic edema | 0
spine MRI no intramedullary lesions | 0
spine MRI no leptomeningeal enhancement | 0
dexamethasone initiated | 0
levetiracetam initiated | 0
escitalopram | 0
quetiapine | 0
infectious diseases team consulted | 0
unrevealing autoimmune antibodies | 0
unrevealing paraneoplastic auto-antibodies | 0
unrevealing lymphoma | 0
unrevealing zoonoses | 0
unrevealing Brucella | 0
unrevealing Bartonella | 0
unrevealing Q-fever | 0
unrevealing Treponema | 0
unrevealing Histoplasma | 0
unrevealing HIV | 0
no systemic malignancy | 0
lumbar puncture opening pressure 14 cmH2O | 0
normal lumbar puncture results | 0
malignant cells negative | 0
lymphoma panel flow cytometry negative | 0
first brain biopsy necroinflammatory process | 0
no acid-fast bacilli | 0
no fungi | 0
no toxoplasma | 0
CD3-positive T-lymphocytes | 0
second brain biopsy performed | 720
occult malignancy workup negative | 0
negative tumor markers | 0
CT chest normal | 0
CT abdomen normal | 0
CT pelvis normal | 0
enlarged mesenteric lymph nodes | 0
central necrosis mesenteric lymph nodes | 0
thyroid ultrasound no malignancy | 0
scrotum ultrasound no malignancy | 0
whole-body FDG-PET scan postoperative changes left frontal | 0
right frontal hypometabolic lesion | 0
no abnormal FDG uptake rest of body | 0
follow-up MRI brain minimal regression lesions | 0
microhemorrhages | 0
MRI with perfusion reduced rCBV | 0
reduced rCBF | 0
high rMTT | 0
reduced NAA peak | 0
high Ch peak | 0
high glutamate peak | 0
variable lipid lactate peaks | 0
changes fraction anisotropy | 0
changes tractography | 0
cerebral angiogram beading anterior cerebral artery | 0
pulse steroids methylprednisolone | 0
improvement mood | 0
improvement right side power | 0
walking with cane | 0
foot orthosis | 0
over anxiety | 0
hyper-alertness | 0
low mood | 0
right distal leg weakness | 0
foot drop | 0
polyuria | 0
rituximab 1000 mg | 0
chest infection | 0
neurological deterioration | 0
focal seizures | 0
encephalopathic | 0
follow-up MRI increased enhancing lesions | 0
increased vasogenic edema | 0
necrotic brain tissue | 0
angiocentric lymphoproliferative process | 0
CD2 expression | 0
CD3 expression | 0
CD7 expression | 0
granzyme B expression | 0
TIA 1 expression | 0
negative CD4 | 0
negative CD5 | 0
negative CD8 | 0
negative CD56 | 0
negative TCR beta F1 | 0
negative TCR delta | 0
EBER negative | 0
peripheral T-cell lymphoma diagnosis | 0
pulmonary embolism | 0
sepsis | 0
disseminated intravascular coagulation | 0
multiorgan failure | 0
brain CT large left frontoparietal hematoma | 0
significant vasogenic edema | 0
midline shift | 0
diffuse loss gray-white differentiation | 0
effacement sulci | 0
cardiopulmonary arrest | 2160
deceased | 2160
