18 years old | 0
male | 0
autoimmune cirrhosis | -1560
ostium secundum | -730
percutaneous Amplatzer | -730
propranolol | -672
azathioprine | -672
vitamin E | -672
multivitamin supply | -672
leukopenia | 0
lymphocytes | 0
anemia | 0
thrombocytopenia | 0
alkaline phosphatase | 0
total serum bilirubin | 0
direct bilirubin | 0
indirect bilirubin | 0
severity score of CHILD A | 0
MELD 11 | 0
variceal banding | 0
desaturation | 0
right superior and inferior lobar atelectasis | 0
purulent tracheal secretions | 0
clinical sepsis | 120
intensive care unit | 120
increased cholestasis | 120
endoscopic retrograde cholangiopancreatography | 120
biliary stenting | 120
cardiothoracic focus search | 120
transesophageal echocardiography | 120
persistent tracheal secretions | 720
sputum cultures | 720
Aspergillus spp | 720
thoracic CT scan | 720
multiple nodes in both lungs | 720
tree-in-bud opacities | 720
posaconazole | 720
caspofungin | 720
amphotericin B | 720
aciclovir | 720
neurological symptoms | 840
left hemiplegia | 840
severe headache | 840
mental status changes | 840
magnetic resonance imaging of the brain | 840
multiple right frontal and right parietal lesions | 840
perilesional edema | 840
biopsy of brain lesions | 840
stereotactic guidance | 840
multiple organ failure | 1152
death | 1152
abundant copper deposits | 1152
aldehyde fuchsin | 1152
periodic acid-Schiff | 1152
hepatic parenchyma | 1152
copper | 1152
binding protein | 1152
periseptal location | 1152
focal intracanalicular cholestasis | 1152
Mallory bodies | 1152
nuclear pseudoinclusions | 1152
Trucut liver biopsy | 96
hepatocanalicular cholestasis | 96
apoptotic hepatocytes | 96
Kupffer cells | 96
sinusoidal congestion | 96
trichrome staining | 96
fibrosis | 96
PAS-D-positive material | 96
intracytoplasmic iron deposits | 96
cytomegalovirus | 96
mild acute cellular rejection | 96
Banff score 4/9 | 96
portal swelling | 96
ductulitis | 96
endotheliitis | 96
cerebral collection | 840
frontal right abscesses | 840
H&E | 840
PAS-D | 840
Ziehl-Neelsen | 840
Gram | 840
Gomori | 840
edema | 840
extensive necrosis | 840
neutrophil infiltration | 840
apoptotic cells | 840
septate hyphae | 840
necrotizing encephalitis | 840
Aspergillus structures | 840