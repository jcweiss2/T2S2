26 years old | 0
twin pregnancy | 0
36 weeks and one day gestation | 0
gravida 1 | 0
0 abortions | 0
malaise | -144
fever | -144
non-productive cough | -144
febrile | 0
tachycardic | 0
hypoxic | 0
O2 saturation of 92% | 0
diffuse rhonchi | 0
increased erythrocyte sedimentation rate | 0
non-stress-test reactive for both fetuses | 0
biophysical profiles 6/8 | 0
decreased fetal movement | 0
chest computed tomography scan | 0
multifocal sub-pleural patchy consolidative opacities | 0
COVID-19 pneumonia | 0
cesarean section | 0
good condition of infants | 0
first minute APGAR score of 9/10 | 0
infants isolated from mother | 0
infants transferred to Neonatal Intensive Care Unit | 0
COVID-19 infection confirmed in mother | 0
RT-PCR negative in infants | 0
infants asymptomatic at two-week follow-up | 0
meropenem | 0
azithromycin | 0
hydroxychloroquine | 0
supplemental oxygen | 0
lack of favorable response to treatment | 6
plasma transfusion from cured COVID-19 patients | 144
Favipiravir added | 144
clinical course improved | 168
second chest CT scan | 288
very faint residual ground-glass opacities | 288
dramatic response to treatment | 288
COVID-19 with pulmonary involvement | 0
discharged after 2 weeks | 336
newborns no COVID-19 symptoms | 336
negative PCR results in newborns | 336
