40 years old | 0
male | 0
presented to the hospital | 0
new-onset uncontrolled seizures | 0
unresponsive | 0
intubated | 0
sedated | 0
admitted to the neurological critical care unit | 0
no significant past medical history | 0
lived in Hardin County, Texas | 0
worked in swimming pool maintenance | 0
had not traveled outside of the state | 0
progressively worsening migraines | -3360
pharmacologic therapy | -3360
nausea | -3360
vomiting | -3360
intermittent neck stiffness | -3360
decreased appetite | -3360
30-pound unintentional weight loss | -3360
severe headaches | -192
photophobia | -192
neck pain | -192
back pain | -192
slurred speech | -192
tremors | -192
drooling | -192
left facial droop | -192
discharged home | -192
noncontrast computed tomography imaging of head and spine | 0
elevated white blood cell count | 0
electroencephalogram showed diffuse slowing | 0
lumbar puncture | 0
elevated opening pressure | 0
low glucose | 0
elevated protein | 0
elevated WBCs in CSF | 0
vancomycin administered | 0
piperacillin-tazobactam administered | 0
Gram stain of CSF | 0
India Ink stain of CSF | 0
BioFire FilmArray Meningitis/Encephalitis Panel positive | 0
CrAg LFA cryptococcal antigen positive in CSF | 0
CrAg LFA cryptococcal antigen positive in serum | 0
intravenous amphotericin B administered | 24
flucytosine administered | 24
CSF cultures grew C gattii | 24
l-canavanine, glycine, 2-bromothymol blue agar test | 24
multilocus sequence typing | 24
worsening fevers | 24
shivering | 24
neck stiffness | 24
thoracic CT identified left lung consolidation | 24
bronchoalveolar lavage performed | 24
continuation of antifungal therapy | 24
serial lumbar punctures | 24
evaluation of immune status | 24
repeated lumbar punctures | 24
elevated opening pressures | 24
persistently elevated protein | 24
decreased glucose | 24
elevated leukocyte counts | 24
no evidence of immunocompromised state | 24
negative HIV 1/2 Ag-Ab | 24
negative hepatitis A/B/C panel | 24
negative QuantiFERON-TB Gold | 24
normal alpha-1-antitrypsin | 24
negative antimitochondrial Ab | 24
negative antinuclear Ab | 24
normal IgA | 24
mildly decreased IgG | 24
mildly decreased IgM | 24
normal CD4/CD8 ratio | 24
mildly decreased absolute lymphocyte count | 24
absence of lymphoproliferation | 24
absence of leukemia | 24
normal CSF angiotensin-converting enzyme | 24
reduced absolute CD4 | 48
reduced absolute CD8 | 48
reduced IgG | 72
reduced IgM | 72
normal chromosomal analysis | 24
serial MRI revealed cerebral diffusion restriction | 24
leptomeningeal enhancement | 24
hemorrhagic transformation of left posterior parietal lobe | 24
restricted diffusion in right upper cervical spinal cord | 24
unable to follow commands | 24
neurological decompensation to eye-opening | 24
purposeful withdrawal from pain | 24
abnormal decerebrate posturing | 24
compromise of brainstem reflexes | 24
discharged to inpatient hospice | 336
died | 336
granulomatous meningitis | 336
cryptococcal organisms in brain | 336
cryptococcal organisms in spinal cord | 336
cryptococcal organisms in posterior pituitary | 336
diffuse bilateral cerebral cortical infarcts | 336
hemorrhage in left posterior parieto>occipital region | 336
small infarct in cervical spinal cord | 336
large cryptococcoma in left lung | 336
cryptococcal organisms in bilateral lungs | 336
disseminated cryptococcosis | 336
cryptococcal meningitis | 336
cause of death complications | 336
