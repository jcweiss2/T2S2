22 years old | 0  
male | 0  
admitted to the hospital | 0  
late-onset multiple acyl-CoA dehydrogenase deficiency (MADD) | 0  
homozygous c.1074G > C variant in the ETFDH gene | 0  
arginine substitution with serine | 0  
reduction of myristate oxidation | 0  
standard treatment of diet | 0  
supplementation of riboflavin | 0  
supplementation of L-carnitine | 0  
numerous crises of hypoglycemia | -...  
numerous crises of metabolic decompensation | -...  
acute kidney failure | -...  
acute respiratory distress syndrome | -...  
hemodialysis | -...  
assisted ventilation | -...  
moderate liver steatosis | 0  
lipid storage myopathy | 0  
mild exercise intolerance | 0  
muscle weakness | 0  
muscle pain | 0  
elevations of plasma-creatine kinase | 0  
normal concentration of free carnitine | 0  
increased concentrations of acyl-carnitines | 0  
hospitalized with acute hypoglycemia | -...  
metabolic acidosis | -...  
intestinal Clostridium difficile infection (CDI) | -...  
recovered on intravenous glucose | -...  
recovered on antibiotics | -...  
hospitalized for acute hypoglycemia | -...  
hospitalized for metabolic acidosis | -...  
recurrent CDI | -...  
abdominal pain | -...  
CT scan of the abdomen | -...  
significantly enlarged spleen | -...  
fecal microbiota transplantation | -...  
admitted to the hospital in a state of hypoglycemia | -...  
admitted to the hospital in a state of metabolic decompensation | -...  
septicemia caused by staphylococcal bacteria | -...  
treated with glucose | -...  
treated with antibiotics | -...  
hospitalized due to progressive abdominal pain | -...  
bloating | -...  
mushy stools | 0  
jaundiced | 0  
febrile | 0  
abdomen distended | 0  
prolonged coagulation | 0  
elevated transaminases | 0  
elevated bilirubin | 0  
impaired synthesis function | 0  
acute necrosis of liver cells | 0  
CT scan of the abdomen | 0  
cirrhotic-looking liver | 0  
multiple small hypodense lesions | 0  
large-volume ascites | 0  
rectal portosystemic shunt | 0  
collaterals to the inferior mesenteric vein | 0  
consistent splenomegaly | 0  
severe colitis | 0  
no stigmata of chronic liver disease | 0  
routine hepatitis tests were negative | 0  
profiles of amino acids remained unchanged | 0  
profiles of acylcarnitines remained unchanged | 0  
ultrasound images of the liver | 0  
CT angiography of the liver | 0  
patent vessels | 0  
no biliary dilatation | 0  
severe degree of portal hypertension | 0  
hepato-fugal portal venous flow | 0  
liver biopsy | 0  
severe macro-vesicular steatosis | 0  
severe micro-vesicular steatosis | 0  
accumulation of glycogen | 0  
accumulation of copper | 0  
accumulation of Mallory bodies | 0  
cirrhotic liver | 0  
no signs of malignancy | 0  
no signs of infection | 0  
liver function rapidly deteriorated | 0  
died from acute liver failure (ALF) | 0  
not a candidate for liver transplant surgery | 0  
not a candidate for trans-jugular intrahepatic portosystemic shunt insertion | 0  
family declined autopsy | 0  
sudden and rapid progression of hepatopathy | 0  
severe steatosis | 0  
beginning cirrhosis of the liver | 0  
overall immunocompromised state | 0  
advanced liver disease | 0  
cholestasis | 0  
hyperbilirubinemia | 0  
no sign of Kayser-Fleischer ring | 0  
recurring hypoglycemic events | -...  
decline in liver function | 0  
impairment of glycogenolysis | 0  
impairment of gluconeogenesis | 0  
habitually elevated transaminases | 0  
increase in transaminases | 0  
increase ascribed to lipid storage myopathy | 0  
liver biopsy not performed | 0  
early stage in development of cirrhosis | 0  
distinguish isoenzymes of transaminases | 0  
initiate appropriate treatment | 0  
decompensated cirrhosis | 0  
portal hypertension | 0  
acute liver failure (ALF) | 0  
death | 0  
