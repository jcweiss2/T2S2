48 years old | 0
    man | 0
    admitted to the emergency department | 0
    cough | -96
    dyspnea | -96
    fever | -48
    highest temperature of 39.3°C | -48
    yellowish sputum | -48
    chills | -48
    sweats | -48
    denied hemoptysis | 0
    took oral cefixime | -96
    took diclofenac sodium | -96
    prior to admission | -96
    in good health | 0
    no history of hypertension | 0
    no history of diabetes | 0
    no history of stroke | 0
    no history of myocardial infarction | 0
    no prior illnesses | 0
    no hospitalizations before present illness | 0
    no known drug allergies | 0
    living in Chengdu | 0
    denied tobacco abuse | 0
    denied alcohol abuse | 0
    denied drug abuse | 0
    married | 0
    three healthy daughters | 0
    family history negative for genetic disease | 0
    body temperature 40.0°C | 0
    heart rate 130 beats/min | 0
    breathing rate 41 breaths/min | 0
    blood pressure 111/59 mmHg | 0
    oxygen saturation 93% | 0
    chest CT revealed diffuse bilateral interstitial infiltrates | 0
    WBC count 6.88×109/L | 0
    neutrophil percentage 85.4% | 0
    lymphocyte percentage 11.0% | 0
    ESR 23 mm/h | 0
    PCT 0.12 ng/mL | 0
    PT 12.5 s | 0
    INR 1.16 | 0
    Fbg 7.01 g/L | 0
    TT 148 s | 0
    D2 1.66 µg/mL | 0
    FDP 6.80 µg/mL | 0
    blood gas analysis pH 7.492 | 0
    PCO2 36 mmHg | 0
    PO2 60.4 mmHg | 0
    oxygenation index 234 mmHg | 0
    electrolytes not significantly abnormal | 0
    renal function not significantly abnormal | 0
    myocardial injury markers not significantly abnormal | 0
    tumor markers not significantly abnormal | 0
    infection markers not significantly abnormal | 0
    Chlamydia pneumoniae not significantly abnormal | 0
    Mycoplasma pneumoniae not significantly abnormal | 0
    developed respiratory failure | 24
    transferred to intensive care unit | 24
    received mechanical ventilation | 24
    received supportive care | 24
    no pleural effusion | 0
    no subsegmental pulmonary embolisms | 0
    no history of cardiac vegetation | 0
    urine tests indicated glucose | 0
    re-examination showed no pathogenic bacteria | 0
    treated with moxifloxacin | 0
    treated with piperacillin tazobactam | 0
    treated with oseltamivir | 0
    body temperature reached 40.0°C | 0
    fever continued | 0
    pulmonary infection progression on repeat CT | 0
    moxifloxacin replaced with linezolid | 72
    moxifloxacin replaced with meropenem | 72
    fever subsided | 96
    symptoms and signs persisted | 96
    WBC count indicated inflammatory activity | 96
    PCT indicated inflammatory activity | 96
    inspiratory crackles in both lungs | 96
    WBC total count 10.11×109/L | 144
    neutrophil count 6.38×109/L | 144
    neutrophils 81.8% | 144
    lymphocytes 32.5% | 144
    lymphocytes 1.51×109/L | 144
    CRP 20 mg/L | 144
    ESR 51 mm/h | 144
    PCT 15.4 ng/mL | 144
    tests for influenza A virus negative | 144
    tests for influenza B virus negative | 144
    tests for cytomegalovirus negative | 144
    tests for Toxoplasma negative | 144
    tests for Epstein–Barr virus negative | 144
    tests for rubella virus negative | 144
    tests for herpes simplex virus negative | 144
    cryptococcal antigen negative | 144
    galactomannan test negative | 144
    β-D-glucan test negative | 144
    anti-nuclear antibody negative | 144
    anti-extractable nuclear antigen antibody negative | 144
    anti-neutrophilic cytoplasmic antibody negative | 144
    peripheral blood cultures showed no abnormalities | 144
    contact with domestic pigeons | 0
    mNGS of BALF identified C. psittaci | 0
    antibacterial agents switched to doxycycline | 168
    moxifloxacin continued | 168
    meropenem continued | 168
    empirical antiviral agents ceased | 168
    PCT decline | 168
    WBC count decline | 168
    fever returned to normal | 360
    no abnormalities in lower limb vascular ultrasonography | 24
    acrocyanosis of both lower extremities | 72
    palpable purpura progressively worsened | 72
    left dorsalis pedis artery occlusion | 144
    right peroneal vein thrombosis | 144
    pulse of left dorsal pedal artery not palpable | 144
    no pathogens detected in sputum | 0
    no pathogens detected in BALF | 0
    no pathogens detected in blood culture | 0
    survived multiple organ failure | 0
    amputation of both legs | 0
    repatriated for further rehabilitation | 0
    doing well at one-year follow-up | 0
    no further symptoms | 0
    C. psittaci pneumonia | 0
    atherosclerotic occlusive disease | 144
    severe infection | 0
    destruction of endothelial cell layer | 0
    serious hemodynamic disorder | 0
    arterioocclusive sclerosis | 0
    sepsis | 0
    multiple organ failure | 0
    confirmed presence of C. psittaci | 96
    tetracycline antibiotics | 168
    macrolides | 168
    quinolones | 168
    combined anti-infective therapy | 168
    lower limb arterial occlusion | 72
    disease progression leading to amputation | 168
    endothelial cell layer destruction | 0
    hemodynamic disorder | 0
    arterioocclusive sclerosis | 0
    first case of C. psittaci pneumonia with lower extremity atherosclerotic occlusive disease | 0
    contact with birds | 0
    mNGS confirmed C. psittaci infection | 96
    treatment with doxycycline | 168
    treatment with moxifloxacin | 168
    treatment with meropenem | 168
    cessation of antiviral agents | 168
    patient recovery | 360
    one-year follow-up | 8784
