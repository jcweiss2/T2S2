36 years old | 0
female | 0
admitted to the hospital | 0
dry cough | -96
shortness of breath | -96
dyspnea | -2
heart palpitations | -2
myalgia | -96
arthralgia | -96
orthopnea | -48
tobacco consumption | -13000
type 2 diabetes in mother | -0
arterial hypertension in mother | -0
no allergies | 0
no controlled substances | 0
no past blood transfusions | 0
no traveling to endemic regions | 0
no tattoos | 0
no body piercings | 0
no history of lung disease | 0
no asthma | 0
no chronic or degenerative diseases | 0
four pregnancies | -0
one delivery | -0
two cesarean surgeries | -0
normal evolution of 33-week pregnancy | 0
recumbent patient | 0
Glasgow coma score of 15 | 0
no focal neurologic deficits | 0
no meningeal signs | 0
diaphoretic | 0
skin and mucosae dehydrated | 0
tachypnea | 0
thoracic and abdominal dissociation | 0
decreased expansion | 0
no vibrations or fremitus | 0
no asymmetries | 0
disseminated bilateral crepitant crackles | 0
bilateral decreased inspiratory breath sounds | 0
tachycardia | 0
heart sounds of good intensity | 0
no extra heart sounds | 0
globous abdomen | 0
live single product | 0
fetal heart rate of 158 bpm | 0
no visceromegaly | 0
no abnormalities upon palpation | 0
filiform pulse | 0
augmented in frequency | 0
decreased in amplitude | 0
no trophic changes | 0
BP of 130/90 mm Hg | 0
HR of 100 bpm | 0
RR of 21 rpm | 0
SO2 with noninvasive ventilation at a rate of 10 L/min of 74% | 0
temperature of 36°C | 0
body-weight of 70 kg | 0
height of 165 cm | 0
BMI of 25.7 | 0
type one respiratory insufficiency | 2
invasive artificial airway with an endotracheal tube | 2
thoracic and abdominal dissociation | 2
intercostal retractions | 2
diaphoresis | 2
cesarean emergency procedure | 4
live newborn male of 1940gr | 4
no malformations | 4
400 cc hemorrhage | 4
admitted to the Intensive Care Unit | 4
bilateral opacities with predominance in the lower lobes | 4
bilateral alveolar infiltrates | 4
areas of consolidation | 4
right predominance at the bases | 4
antimicrobial treatment | 4
one gram of intravenous ceftriaxone | 4
clarithromycin 500 mg orally | 4
consecutive blood cultures | 8
culture of bronchial secretions | 8
IgG antibodies against Mycoplasma pneumonie | 8
galactomannan assay | 8
serum procalcitonin levels | 8
urinalysis | 8
abundant bacteria | 8
erythrocytes 118 per field | 8
leukocytes of 163 per high power field | 8
immunoassays | 8
negative | 8
extubated | 48
adequate respiratory mechanics | 48
discharged to Internal Medicine Department | 48
echocardiogram | 48
left ventricular ejection fraction of 66% | 48
normal systolic function | 48
mild diastolic dysfunction | 48
global pericardial effusion | 48
CT-guided percutaneous lung biopsy | 168
moderately differentiated malignant neoplasia | 168
invasive pulmonary adenocarcinoma | 168
lepidic growth pattern | 168
immunohistochemistry studies | 168
pneumothorax | 168
tube thoracostomy | 168
endopleural tube | 168
pleural effusion | 168
exudate | 168
evaluated by the Oncology Department | 168
completely disabled | 168
ECOG 4 | 168
chemotherapy administration contraindicated | 168
sepsis of unknown origin | 168
palliative care protocol | 168
morphine | 168
dyspnea | 168
pain control | 168
torpid clinical evolution | 240
orthopnea | 240
temperature of 39°C | 240
leukocytosis | 240
extreme bradycardia | 720
asystole | 720
death | 720