56 years old | 0  
    male | 0  
    diagnosed with pancreatic cancer | -5760  
    multiple liver metastases | -5760  
    chemotherapy | -5760  
    stent insertion | -408  
    biliary tract obstruction | -408  
    febrile sense | -336  
    chills | -336  
    antipyretics | -336  
    analgesics | -336  
    admitted to nursing care hospital | -240  
    emergency room visit | -240  
    unresolved fever | -240  
    chill | -240  
    abdominal pain | -240  
    diabetes mellitus | 0  
    vidagliptin/metformin | 0  
    acutely ill | 0  
    blood pressure 100/60 mmHg | 0  
    blood pressure 90/60 mmHg | 1  
    respiratory rate 20 breaths per minute | 0  
    pulse rate 90 beats per minute | 0  
    body temperature 38.8°C | 0  
    WBC count 1,250/mm3 | 0  
    hemoglobin 5.9 g/dL | 0  
    platelet count 14,000/mm3 |%0  
    C-reactive protein 19.75 mg/dL | 0  
    aspartate aminotransferase 274 UI/L | 0  
    alanine aminotransferase 143 IU/L | 0  
    total/direct bilirubin 4.11/2.71 mg/dL | 0  
    total protein 4.4 g/dL | 0  
    albumin 2.0 g/dL | 0  
    prothrombin time (international normalized ratio) 25.3 second (2.21) | 0  
    active partial thromboplastin time 60.7 second | 0  
    blood urea nitrogen 34.5 mg/dL | 0  
    creatinine 1.9 mg/dL | 0  
    arterial blood gas analysis pH 7.515 | 0  
    pCO2 31.6 mmHg | 0  
    pO2 78.8 mmHg | 0  
    HCO3 25.5 mmol/L | 0  
    O2 saturation 96.9% | 0  
    abdomen CT showed pancreatic cancer | 0  
    metallic stent inserted | 0  
    no evidence of bleeding | 0  
    acute cholangitis | 0  
    septic shock | 0  
    intravenous piperacillin/tazobactam | 0  
    teicoplanin | 0  
    norepinephrine | 0  
    packed red cells transfusion | 0  
    platelets transfusion | 0  
    admitted to ICU | 8  
    APACHE II score 19 | 8  
    WBC count deteriorated to 250/mm3 | 48  
    platelet count deteriorated to 8,000/mm3 | 48  
    died | 120  
    carbapenem-resistant K. pneumoniae blood culture | 0  
    antimicrobial resistance | 0  
    KPC2 producing Klebsiella pneumoniae | 0  
    MCR1 possessing ST307/Tn4401a[blaKPC2] K. pneumoniae | 120  
    no hospital outbreak | 120  
    IRB approval | 120  
    community-onset bacteremia | 0  
    fatal outcome | 120  
    inter-regional spread | 120  
    inter-facility spread | 120  
    community-onset infections | 120  

