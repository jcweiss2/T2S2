63 years old | 0
woman | 0
psychiatric disorders | 0
coma | 0
septic shock | 0
mild traumatic brain injury | -432
fall | -432
aspiration pneumonia | -432
no loss of consciousness | -432
computed tomography (CT) performed | -432
normal CT | -432
no bleeding | -432
thin ventricles | -432
median structure in place | -432
pneumonia evolved to ARDS | -72
prone positioning sessions | -72
deep sedation with midazolam | -72
deep sedation with sufentanil | -72
bispectral index (BIS) monitoring | -72
low BIS values (25–34) | -72
low sedative doses | -72
discontinuation of sedative drugs | 0
spontaneous ventilation recovery | 72
no signs of waking up | 72
low BIS (20–30) | 72
no acute kidney injury | 72
no liver failure | 72
sluggish reaction to pain on left arm | 72
intermediate pupils | 72
reactive pupils | 72
ultrasonography for brain perfusion | 72
TCD on left MCA | 72
pulsatility index = 1.09 | 72
end diastolic velocity = 52.11 cm/s | 72
right MCA not identifiable | 72
ONSD measurements: right eye 7.4 mm, left eye 7.05 mm | 72
elevated ICP suspected | 72
new brain CT performed | 72
osmotherapy initiated | 72
blood pressure elevation | 72
head elevation | 72
temperature control | 72
carbon dioxide control | 72
glycemia control | 72
multiple deep parenchymal hematomas | 72
bilateral cerebellar ischemia | 72
diffuse cerebral edema | 72
brain coning | 72
optimal brain perfusion treatment | 72
unfavorable evolution | 168
brain death | 192
backflow in MCA | 192
two electroencephalograms confirming brain death | 192
