84 years old | 0
female | 0
Alzheimer's dementia | -936
admitted to the hospital | 0
fever | 0
pulmonary thromboembolism | -936
deep vein thrombosis | -936
blood pressure 87/44 mm Hg | 0
heart rate 105 bpm | 0
body temperature 38.2° | 0
leukocytosis | 0
elevated levels of C-reactive protein | 0
serum lactate level 3.57 mmoL/L | 0
septic shock | 0
methicillin-resistant Staphylococcus aureus bacteremia | 0
contrast-enhanced chest and abdominal CT | 4
multiple peripheral nodules in both lungs | 4
septic embolism | 4
mild swelling and heterogeneous enhancement of the thyroid gland | 4
perithyroidal fluid collection | 4
admitted to the intensive care unit | 4
glycopeptide antibiotic | 4
fluid resuscitation | 4
diluted norepinephrine | 4
central venous catheter | 4
hemodynamically stable | 4
follow-up neck CT | 22
thyroid function tests | 22
normal concentrations of serum free thyroxine | 22
normal concentrations of serum thyroid-stimulating hormone | 22
low concentration of serum triiodothyronine | 22
moved to the general ward | 96
discharged | 120