27 years old | 0
female | 0
admitted to the hospital | 0
seizure | -24
loss of consciousness | -24
acute psychosis | -72
cold-like symptoms | -168
runny nose | -168
low-grade fever | -168
stable vital signs | 0
Glasgow coma scale 6 | 0
mild signal changes in the bilateral hippocampus and left temporal cortex | 0
local meningeal congestion | 0
anti-NMDA receptor antibodies detected | 0
abdominal ultrasound screening | 0
weak liquid echo of the right ovary | 0
teratoma suspected | 0
tumor removal | 24
pathology report confirmed teratoma containing nerve tissues | 24
comatose | 24
facial involuntary movement | 24
lip peristalsis | 24
uncontrolled eye blinking | 24
first-line therapy initiated | 24
IVMP | 24
IVIG | 48
plasmapheresis | 72
immunoadsorption | 120
second-line therapy initiated | 168
rituximab | 168
cyclophosphamide | 192
septicemia with Staphylococcus caprae | 240
septicemia with klebsiella pneumoniae | 360
bilateral salpingo-oophorectomy | 336
inflammation found | 336
no teratoma found | 336
immunosuppressant therapy initiated | 336
mycophenolate mofetil | 336
intrathecal MTX and DXM | 432
antibody titer decreased | 432
recovered consciousness | 1020
GCS score 9T | 1020
physical therapy | 1020
good prognosis | 1104
mRS score 1 | 1104
diffuse muscular ossification | 1104
X-ray examination | 1104