3 years old | 0
male | 0
admitted to the hospital | 0
cough | -168
nasal congestion | -168
sore throat | -24
no fever | 0
no dyspnea | 0
no trauma | 0
no recent travel | 0
tolerating solids | 0
tolerating liquids | 0
cough suppressant | -168
ibuprofen | -168
symptomatic relief | -168
well appearing | 0
afebrile | 0
hemodynamically stable | 0
temperature 36.7°C | 0
pulse 113 | 0
respiratory rate 23 | 0
pulse oximetry 98% | 0
nasal congestion | 0
erythematous pharynx | 0
drink fluids | 0
discharged home | 0
viral syndrome | 0
congestion | 72
sore throat | 72
torticollis | 72
limited range of motion of the neck | 72
drooling | 72
tactile fever | 48
self-resolved fever | 48
no vomiting | 72
temperature 37.5°C | 72
pulse 121 | 72
blood pressure 102/60 | 72
respiratory rate 24 | 72
pulse oximetry 100% | 72
well appearing | 72
well-hydrated | 72
diffuse neck tenderness | 72
no lymphadenopathy | 72
left-sided torticollis | 72
no significant trismus | 72
no evidence of meningismus | 72
elevated WBC (24.1 K/µL) | 72
elevated CRP (2.07 mg/dL) | 72
mild hypoglycemia (65 mg/dL) | 72
slightly low serum bicarbonate level (18 mmol/L) | 72
retropharyngeal abscess concern | 72
soft tissue neck plain film | 72
diffuse paravertebral swelling | 72
2.2 cm linear radiopaque density | 72
foreign body concern | 72
eating fish earlier in the week | -168
antibiotics | 72
transferred to another pediatric facility | 72
ENT consultation | 72
repeat soft tissue neck plain film | 72
rigid esophagoscopy | 72
purulent fluid in the cervical esophagus | 72
drainage of purulent fluid | 72
2 cm fish bone | 72
fish bone removed | 72
Penrose drain placed | 72
esophageal perforation | 72
abscess | 72
postoperative CT scan of the neck | 72
no residual foreign body | 72
no residual abscess | 72
admitted to pediatric intensive care unit | 72
broad-spectrum antibiotics | 72
clindamycin | 72
ampicillin/sulbactam | 72
positive wound cultures | 72
gram-positive cocci in pairs | 72
Penrose drain removed | 72
discharged home | 72
tolerating feeds | 72
oral clindamycin | 72
no evidence of persistent abscess | 72
no esophageal perforation | 72
ENT follow up | 72
