52 years old| 0
male | 0
admitted to the hospital | 0
right upper quadrant pain | -168
discomfort | -168
abdominal fullness | -168
distention | -168
worsened after meals | -168
denied nausea | -168
denied vomiting | -168
denied stiffness | -168
denied fever | -168
hepatic puncture | -24
drainage | -24
afebrile | 0
pulse rate 80 beats/minute | 0
blood pressure 118/73 mmHg | 0
respiratory rate 26 breaths/minute | 0
leukocyte count 16.4×109/L | 0
neutrophil 94.5% | 0
haemoglobin 85 g/L | 0
platelet count 240×109/L | 0
procalcitonin 2.3 ng/mL | 0
plasma fibrinogen 7.48 g/L | 0
serum glutamic oxalacetic transaminase 67 U/L | 0
glutamic-pyruvic transaminase 83 U/L | 0
cholinesterase 1360 U/L | 0
total protein 50.8 g/L | 0
albumin 21.5 g/L | 0
blood urea nitrogen 10.8 mmol/L | 0
creatinine 51.3 umol/L | 0
HIV negative | 0
syphilis negative | 0
abdominal distension | 48
mild bellyache | 48
extreme thirst | 48
right abdominal tenderness | 48
no rebound | 48
no guarding | 48
temperature 36.8°C | 48
drainage catheter yield 150 mL fulvous fluid | 48
abdominal CT scan | 48
pelvic CT scan | 48
irregular low-density lesion in right posterior hepatic lobe | 48
gas density shadow inside liver lesion | 48
liquid density shadow around lower margin of liver | 48
high-density drainage tube shadow | 48
round-like low-density lesion in right lobe of liver | 48
appendix thickened 20 mm diameter | 48
ascending colon disorganised structure | 48
multiple gas accumulation in bowel | 48
dilation in bowel | 48
air-fluid levels inside abdomen | 48
blood pressure 93/59 mmHg | 48
exploratory laparotomy | 48
fulvous purulent exudate | 48
necrotic tissue in extraperitoneal space | 48
necrotic tissue in abdominal cavity | 48
partial postnecrotic defect in peritoneum | 48
massive epiploon adhesion | 48
perforation under right side of liver | 48
perforation in right ascending colon | 48
ileocecal resection | 48
partial resection of ascending colon | 48
ileostomy | 48
drainage of hepatic abscess | 48
drainage of abdominal abscess | 48
drainage of extraperitoneal abscess | 48
orotracheal intubation | 48
hypotension | 48
anemia | 48
fever | 48
transferred to ICU | 48
noradrenaline pumped | 48
ventilator used | 48
intravenous hydration | 48
nutritional support therapy | 48
blood transfusion | 48
blood cultures sent | 48
drainage fluids sent | 48
intravenous tigecycline | 48
intravenous piperacillin/tazobactam | 48
temperature monitoring | 48
routine blood count monitoring | 48
procalcitonin monitoring | 48
CRP monitoring | 48
temperature 39.3°C | 72
pulse rate 130 beats/minute | 72
leukocyte count 35.9×109 cells/L | 72
neutrophil 92.4% | 72
PCT 8.15 ng/mL | 72
CRP 174 mg/L | 72
blood cultures for aerobic culture | 72
blood cultures for anaerobic culture | 72
continued tigecycline | 72
continued piperacillin/tazobactam | 72
anaerobic blood culture positive | 120
Gram-positive bacillus | 120
blood agar base medium culture | 120
anaerobic incubation | 120
E. lenta identified | 120
plasma fibrinogen 1.0 g/L | 120
tigecycline replaced by teicoplanin | 120
piperacillin/tazobactam discontinued | 120
ertapenem added | 120
drainage fluid cultures | 120
Escherichia coli isolated | 120
treated with ertapenem | 120
treated with teicoplanin | 120
fever improved | 120
leukocytosis improved | 120
PCT improved | 120
CRP improved | 120
transferred to general ward | 168
ertapenem continued | 168
teicoplanin continued | 168
debridement | 168
dressing change | 168
symptomatic supportive treatment | 168
negative blood cultures | 168
CT showed decreased hepatic abscess | 168
CT showed decreased ascites | 168
intravenous ertapenem continued | 168
intravenous teicoplanin continued | 168
symptoms alleviated | 168
discharged | 240
oral clindamycin | 240
no recurrence of fever | 240
complete resolution of abscess | 240
six-week course of ertapenem | 240
