33 years old | 0
male | 0
good general health | 0
good nutritional status | 0
185 cm | 0
80 kg | 0
minor superficial injury on lower left leg | -240
acquired during ski vacation | -240
no pre-existing diseases | 0
no significant medical history | 0
local self-treatment | -240
deterioration of wound conditions | -240
visited centre for general medicine | -192
initiation of antibiotic therapy with oral Cefuroxime | -192
progressive clinical deterioration of wound conditions | -192
aching hematoma | -192
admitted to hospital | 0
surgical treatment of hematoma | 0
two further wound debridements | 24
application of vacuum-assisted closure | 24
antibiotic therapy escalated to Clindamycin | 0
antibiotic therapy escalated to Tazobactam | 0
transferred to university hospital | 216
awake | 0
oriented | 0
stable respiratory condition | 0
stable circulatory condition | 0
temperature 37.2 °C | 0
blood pressure 171/85 mmHg | 0
pulse 140 beats per minute | 0
oxygen saturation 95% | 0
somnolent | 0
easily aroused | 0
severe pain | 0
swellings in both axillae | 0
swellings in both groins | 0
increased white blood cell count | 0
C-reactive protein 298.8 mg/dL | 0
surgical wound excisions | 0
large debridement | 0
empirical antibiotic therapy changed to Meropenem | 0
empirical antibiotic therapy changed to Penicillin G | 0
empirical antibiotic therapy changed to Clindamycin | 0
tissue samples taken | 0
swabs taken | 0
blood cultures taken | 0
no causative pathogen identified | 0
anti-infective therapy supplemented by Levofloxacin | 48
anti-infective therapy supplemented by Daptomycin | 48
Caspofungin added | 48
hole-body computed tomography scan | 72
fasciitis of left upper and lower leg | 72
bilateral pulmonary oedema | 72
bilateral pleural effusions | 72
basal atelectasis | 72
generalized barrier disruption | 72
mechanical ventilation | 96
operational inspection | 96
large debridement of both axillae | 96
fasciotomy of left thigh | 96
necrotic area increased | 96
microbiological analyses negative | 96
positive serological evidence of Herpes simplex virus-I | 96
therapy with Acyclovir | 96
Corynebacterium tuberculostearicum detected | 120
Acinetobacter baumanii detected | 120
cortisone therapy initiated | 120
intravenous immunoglobulin therapy initiated | 120
hyperinflammation diminished | 144
general condition improved | 144
weaning from respirator | 144
CRP dropped | 144
WBC dropped | 144
pro-calcitonin dropped | 144
need for hemodynamic support reduced | 144
vacuum assisted wound closure | 240
wound conditions improved | 240
wounds closed | 312
split-skin graft from right thigh | 312
discharged from hospital | 432
follow-up examination | 4320
healthy | 4320
sufficient wound conditions | 4320