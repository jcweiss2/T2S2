60 years old | 0
male | 0
admitted to the hospital | 0
recurrent episodes of fever | -1728
recurrent episodes of cough | -1728
most recent episode of fever | -144
most recent episode of cough | -144
most recent episode of chills | -144
treatment with clarithromycin (first episode) | -1728
cruise trip to the Baltic Sea | -1728
febrile (temperature 40.1°C) | 0
tachycardic (109 beats/min) | 0
normotensive (138/81 mmHg) | 0
tachypneic (28 breaths/min) | 0
basal rales over the left lung | 0
perioral grouped blisters | 0
leukocytosis (13×109/L) | 0
elevated C-reactive protein (303 mg/mL) | 0
elevated total protein (97 g/L) | 0
low albumin (26 g/L) | 0
moderate hyponatremia (sodium 127 mmol/L) |B0
chest X-ray showing retrocardiac consolidation of the left lower lobe | 0
community-acquired pneumonia | 0
empirical antimicrobial therapy with piperacillin/tazobactam | 0
empirical antimicrobial therapy with clarithromycin | 0
blood cultures positive for S. pneumoniae | 24
sputum cultures positive for S. pneumoniae | 24
de-escalated to intravenous benzylpenicillin | 24
de-escalated to oral amoxicillin | 24
treated for a total duration of 14 days | 336
presumed cutaneous herpes simplex type 1 (HSV-1) infection | 0
treatment with valaciclovir | 0
confirmed HSV-1 infection (positive PCR) | 24
detailed history revealed night sweats | 0
detailed history revealed weight loss of 4 kg | 0
HIV test negative | 0
suspected multiple myeloma (MM) | 0
serum electrophoresis identified IgG kappa monoclonal gammopathy | 24
immunofixation identified IgG kappa monoclonal gammopathy | 24
bone marrow biopsy showing plasma cell infiltration >60% | 24
whole-body computed tomography showing lytic lesions | 24
diagnosis of MM IgG kappa | 24
recovery from bacteremic pneumonia | 336
induction treatment with bortezomib | 336
induction treatment with lenalidomide | 336
induction treatment with dexamethasone | 336
scheduled for autologous hematopoietic stem cell transplantation | 336
treatment with intravenous immunoglobulin discussed | 336
received 13-valent pneumococcal vaccination | 720
discharged | 336
