diagnosed with Hodgkin lymphoma | -192
treated with chemotherapy | -192
treated with mantle field radiation | -192
diagnosed with inflammatory colitis | -192
treated with mesalazine | -192
last flare of inflammatory colitis | -12
diagnosed with breast cancer | 0
palpable mass on right breast | 0
radiological examination of breast | 0
pathological examination confirmed invasive ductal carcinoma | 0
staging CT scan of thorax and abdomen | 0
started neoadjuvant chemotherapy | 14
completed first cycle of chemotherapy | 24
underwent port-à-cath insertion | 27
presented to emergency room with fever | 38
started broad-spectrum i.v. antibiotic therapy | 38
underwent PORT rimotion and necrosectomy | 38
defervescence and improvement in subcutaneous cellulitis | 41
new febrile seizure | 44
underwent second necrosectomy | 44
modified antibiotic therapy | 44
transferred to Thoracic Surgery Unit | 44
underwent left thoracoscopy with pleural and mediastinal drainage | 44
admitted to Intensive Care Unit | 44
started systemic methylprednisolone | 50
started topical cyclosporine | 50
showed progressive resolution of mediastinitis and pleural effusion | 50
showed wound improvement with scar | 50
underwent breast ultrasound | 65
underwent right mastectomy and axillary dissection | 65
breast surgical wound healing was regular | 70
pathology assessment revealed fibroelastosis and chronic inflammation | 70
restaging brain/chest/abdomen CT was negative for distant metastasis | 70
released from hospital | 83
underwent autologous skin graft | 83
resumed chemotherapy with carboplatin and paclitaxel | 90
completed fourth and last cycle of chemotherapy | 200
started follow-up | 200