61 years old | 0
male | 0
admitted to the hospital | 0
pleuritic chest pain | 0
paroxysmal AF | -720
pulmonary vein isolation | -240
cryothermal ablation | -240
diabetes mellitus | 0
hypertension | 0
empagliflozin | 0
dabigatran | 0
bisoprolol | 0
pericardial friction rub | 0
diffuse ST-elevation | 0
PR depression | 0
normal troponin levels | 0
preserved ventricular function | 0
small to medium circumferential pericardial effusion | 0
0.5 mg/kg/day of prednisone | 0
0.5 mg colchicine twice daily | 0
discharged | 96
severe weakness | 144
fatigue | 144
single syncopal episode | 144
blood-tinted vomitus | 144
pleuritic chest pain | 144
low blood pressure | 144
high temperature | 144
high oxygen saturation | 144
low haemoglobin | 144
mild neutrophilia | 144
high creatinine level | 144
high urea concentration | 144
normal troponin levels | 144
nasogastric tube insertion | 144
coffee-ground matter | 144
no active bleeding | 144
bedside TTE | 144
no differences from previous study | 144
presumptive diagnosis of mediastinitis | 144
AOF | 144
2000 cc of intravenous fluids | 144
0.5 mcg/kg/min of norepinephrine | 144
broad-spectrum antibiotics | 144
amoxicillin clavulanate | 144
fluconazole | 144
non-gated CT angiography | 144
multiple mediastinal lymph nodes | 144
small amount of fluid in the mediastinum and pericardium | 144
no extravasation of contrast medium | 144
no pneumomediastinum or pneumopericardium | 144
brain CT | 144
no focal lesion | 144
multiorgan failure | 168
low haemoglobin level | 168
high creatinine level | 168
intubation | 168
mechanical ventilation | 168
third TTE | 168
same amount of pericardial effusion | 168
preserved biventricular function | 168
no air in the cardiac cavities | 168
agitated saline injection | 168
bubbles in the left atrium and ventricle | 168
definitive diagnosis of AOF | 168
surgical repair | 168
left atrium necrotic rupture | 168
pericardial patch | 168
gastroscopy | 192
12 mm tear in the low oesophagus | 192
endoclips | 192
high-grade fever | 192
haemodynamic instability | 192
meropenem | 192
micafungin | 192
positive polymicrobial pleural fluid cultures | 192
discharged for rehabilitation | 720