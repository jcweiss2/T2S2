44 years old | 0
male | 0
admitted to the hospital | 0
dry cough | -120
fever | -120
hypoxia | -48
intubated | -48
COVID-19-related pneumonia | -48
hypertension | 0
type II diabetes mellitus | 0
previous stroke | 0
metformin | 0
alogliptin | 0
serum glucose 222 mg/dL | 0
azithromycin | -48
ceftriaxone | -48
hydroxychloroquine | -48
worsening hypoxemia | -24
cefepime | 0
vancomycin | 0
mechanically ventilated | 0
temperature of 102.8°F | 0
blood pressure of 138/77 mm Hg | 0
pulse of 114 beats per minute | 0
respirations of 16 | 0
oxygen saturation of 95% | 0
weight of 91 kilograms | 0
WBC of 17.1 | 0
lactate dehydrogenase of 570 | 0
C-reactive protein of 328 | 0
ferritin of 2043 | 0
d-dimer of 0.74 | 0
interleukin-6 of 21 | 0
procalcitonin of 5.59 | 0
dexamethasone | 120
fever resolution | 144
WBC of 24.9 | 240
piperacillin/tazobactam | 240
vancomycin | 240
possible aspiration pneumonia | 240
self-extubation | 240
reintubation | 240
tracheal aspirate negative | 240
blood cultures negative | 240
extubated | 384
BiPAP | 384
nasal cannula | 384
transferred to general medicine floor | 384
leukocytosis | 528
temperature of 101.1°F | 528
WBC of 14.7 | 528
altered mental status | 528
piperacillin/tazobactam | 528
vancomycin | 576
blood cultures negative | 576
urine cultures negative | 576
fungal cultures negative | 576
serum galactomannan negative | 576
beta-d-glucan negative | 576
urinalysis negative | 576
CXR showed patchy infiltrates | 576
sputum Gram stain showed Klebsiella pneumoniae | 576
Klebsiella pneumoniae resistant to piperacillin/tazobactam | 576
cefepime | 576
fever persisted | 576
leukocytosis persisted | 576
CT scan of chest and abdomen | 696
diffuse opacities | 696
consolidation in right lower lobe | 696
right hilar lymphadenopathy | 696
calcified subcarinal lymph nodes | 696
meropenem | 696
caspofungin | 696
vancomycin | 696
metronidazole | 696
caspofungin discontinued | 720
voriconazole | 720
leukocytosis | 720
intermittent fever | 720
sputum cultures negative | 720
CT scan showed increased multifocal cavitation | 840
blood cultures negative | 840
urine Legionella antigen negative | 840
serum galactomannan negative | 840
beta-d-glucan negative | 840
urine Histoplasma antigen negative | 840
Coccidioides immunoglobulin G antibody negative | 840
COVID-19 RT-PCR negative | 840
sputum smears positive for acid-fast bacilli | 840
Mycobacterium tuberculosis complex identified | 840
no rifampin resistance | 840
isoniazid | 840
rifampin | 840
ethambutol | 840
pyrazinamide | 840
vitamin B6 | 840
fever resolution | 876
leukocytosis resolution | 876
discharged | 1008
long-acting insulin | 0
rapid-acting insulin | 0
serum glucose levels ranged from 50 to 450 mg/dL | 0
positive purified protein derivative test | -8760
treated with isoniazid for 3 months | -8760
born in Haiti | 0
travels to Haiti regularly | 0