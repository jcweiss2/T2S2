25 years old | 0
female | 0
autoimmune hepatitis | 0
cirrhosis | 0
acute-onset excruciating bilateral lower extremity pain | 0
edema | 0
ascites | 0
fever | 0
chills | 0
nausea | 0
dizziness | 0
heavy menorrhagia | 0
unprotected sexual intercourse two weeks prior to presentation | -336
no history of tobacco use | 0
no history of alcohol use | 0
no history of substance use | 0
acetaminophen | 0
ibuprofen | 0
azathioprine | 0
prednisone | 0
not currently taking immunosuppressive medication | 0
prescriptions not filled in several months | 0
no follow-up with gastroenterology for over eight months | 0
no recent travel history | 0
influenza vaccination | 0
COVID-19 vaccination | 0
hemodynamically unstable | 0
blood pressure 67/39 mmHg | 0
heart rate 129 beats per minute | 0
respirations 33 per minute | 0
temperature 35.1 degrees Celsius | 0
jaundice | 0
scleral icterus | 0
abdominal ascites with fluid wave | 0
anasarca | 0
labia majora edema | 0
labia minora edema | 0
bilateral lower extremities edema | 0
erythematous vaginal vault | 0
minimal discharge | 0
no vesicles | 0
no lesions | 0
no retained foreign objects | 0
fine reticular violaceous patches on right proximal thigh | 0
lactic acidosis | 0
lactic acid 13.1 mmol/L | 0
creatinine 1.49 mg/dL | 0
aspartate transaminase 56 units/L | 0
alanine transaminase 62 units/L | 0
total bilirubin 3.7 mg/dL | 0
direct bilirubin 3.19 mg/dL | 0
alkaline phosphatase 213 units/L | 0
total protein 5.3 g/dL | 0
albumin 1.4 g/dL | 0
hemoglobin 5.2 g/dL | 0
leukocytes 1.3 k/uL | 0
platelets 90 k/uL | 0
prothrombin time 37.9 s | 0
international normalized ratio 3.9 | 0
beta-human chorionic gonadotropin test negative | 0
peripheral smear with occasional schistocytes | 0
paracentesis | 0
peritoneal fluid leukocyte count 9821 | 0
neutrophilic predominance (82%) | 0
CT angiography revealing cirrhosis | 0
portal hypertension | 0
large volume abdominal ascites | 0
splenomegaly | 0
generalized edematous wall thickening of the colon and rectum | 0
admitted to medical intensive care unit | 0
intubation due to labored breathing | 0
tachypnea | 0
early resuscitation with intravenous fluids | 0
blood products | 0
vasopressors | 0
broad-spectrum antibiotic therapy initiated | 0
vancomycin | 0
piperacillin-tazobactam | 0
doxycycline | 0
clindamycin | 0
concern for possible toxic shock syndrome | 0
received intravenous immunoglobulin | 0
large violaceous non-blanching ecchymoses extending from bilateral proximal thighs to calves | 16
several flaccid bullae developed | 16
skin over entire right leg dusky and violaceous with sharply demarcated borders | 36
left proximal thigh to mid-shin dusky and violaceous with sharply demarcated borders | 36
various-sized bullae up to greater than 10 cm filled with red to black-colored fluid | 36
lactate dehydrogenase 298 units/L | 0
fibrinogen 187 mg/dL | 0
D-dimer >20 mcg/mL | 0
urinalysis without signs of infection | 0
salicylate level negative | 0
acetaminophen level negative | 0
Chlamydia trachomatis nucleic acid amplification test negative | 0
Neisseria gonorrhea nucleic acid amplification test negative | 0
urine toxicology screen negative | 0
peritoneal fluid culture negative | 0
blood culture grew pan-susceptible Streptococcus pneumoniae | 0
progressive hypoxia | 0
shock despite maximal ventilator and vasopressor support | 0
passed away within 48 h of admission | 48
autopsy showed cirrhotic liver | 0
diffuse alveolar damage | 0
over five liters of serous fluid in the abdominal compartment | 0
no history of asplenia | 0
functional hyposplenia | 0
pneumococcal vaccination not received | 0
no health insurance | 0
limited access to healthcare system | 0
