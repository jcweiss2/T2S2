25 years old | 0
female | 0
presented to the Emergency Department | 0
epigastric pain | -1464
intermittent low-grade fever | -1464
multiple hospitalizations | -1464
postprandial vomiting | -1464
breathing difficulty on exertion | -1464
orthopnea | -1464
loss of appetite | -1464
weight loss | -1464
no typical chest pain | 0
no night sweats | 0
no limb edema | 0
no jaundice | 0
no decreased urine output | 0
severe shock | 0
tachycardia | 0
tachypnea | 0
unrecordable blood pressure | 0
epigastric tenderness | 0
left infrascapular crepts | 0
decreased breath sounds | 0
fluid resuscitation | 0
inotropes | 0
IV antibiotics | 0
azithromycin | 0
piperacillin/tazobactam | 0
blood culture | 0
portable chest radiograph | 0
pneumopericardium | 0
two-dimensional echocardiography | 0
cardiac tamponade | 0
echogenic materials | 0
pericardiocentesis | 0
pyo-pneumopericardium | 0
pus culture | 0
Candida species | 0
IV fluconazole | 0
clinical instability | 0
high inotropic support | 0
metabolic acidosis | 7
intubation | 7
mechanical ventilation | 7
clinical deterioration | 24
death | 24
