36 years old | 0
male | 0
admitted to the outpatient clinic | 0
swallowing difficulties | -72
plain chest radiography with a water soluble contrast swallow | -72
no pathological lesions | -72
PPI therapy | -72
Pantoprazol | -72
six food elimination diet | -72
noncompliant for follow-up | -72
swallowing complaints persisted | -72
presented to the emergency department | 8760
swallowing complaints | 8760
esophageal food bolus impaction | 8760
plain chest radiography with a water soluble contrast swallow | 8760
9 cm long stricture | 8760
food bolus impaction in the middle third of the esophagus | 8760
gastroscopy | 8760
food bolus impaction at 25 cm from dental arch | 8760
eosinophilic esophagitis | 8760
subcutaneous emphysema | 8760
thoracic computer tomography | 8760
pneumomediastinum | 8760
new upper GI endoscopy | 8760
esophageal perforation | 8760
general condition declined | 8760
transferred to surgical department | 8760
febrile | 8760
38.2°C | 8760
continuous chest pain | 8760
chest pain increases with motion | 8760
no emphysema | 8760
bilateral soft rough breathing sounds | 8760
hemodynamically stable | 8760
blood pressure 140/90mmHg | 8760
arterial pulse 85bpm | 8760
oxygen saturation 98% | 8760
increased inflammatory markers | 8760
mild eosinophilia | 8760
esophageal stricture | 8760
preoperative ICU evaluation | 8760
transhiatal esophagectomy | 8760
cervical esophagostomy | 8760
pyloromyotomy | 8760
feeding jejunostomy | 8760
eosinophilic esophagitis confirmed by histologic examination | 8760
eosinophilic gastritis | 8760
nutritional support | 8760
control contrast study | 8760
jejunostomy tube position confirmed | 8760
dextrose solution administered | 8760
Nutrison Advanced Peptisorb administered | 8760
rate increased to 80ml/h | 8760
no abdominal discomfort | 8760
discharged | 8880
hypoalbuminemia | 8880
poor enteral nutrition | 8880
cervical esophagogastrostomy | 17520
re-establish continuity of gastrointestinal tract | 17520
contrast imaging study | 17520
anastomotic integrity confirmed | 17520
clear fluids administered | 17520
enteral tube feeding decreased | 17520
diet changed to full fluid consistency | 17520
discontinued before discharge | 17520
discharged | 17544
correct oral nutrition | 17544
no swallowing disorders | 17544
no dysphagia | 17544
no esophageal food bolus impaction | 17544
no malabsorption syndrome | 17544
