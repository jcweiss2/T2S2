4 years old | 0
    male | 0
    admitted to the intensive care unit | 0
    malaise | -48
    lethargy | -48
    tachypnea | -48
    sore throat | -48
    abdominal pain | -48
    vomiting | -48
    dehydration | -48
    polyuria | -504
    polydipsia | -504
    4-kg weight loss in 3 weeks preceding admission | -504
    afebrile | 0
    tachypneic (46 breaths per minute) | 0
    Kussmaul respirations | 0
    heart rate 156 beats per minute | 0
    blood pressure 90/55 mm Hg | 0
    light drowsiness | 0
    no jugular distension | 0
    diffuse rhonchi in all lung areas | 0
    diabetic ketoacidosis confirmed | 0
    plasma glucose level 29.8 mmol/L | 0
    pH 6.788 | 0
    pO2 5.20 kPa | 0
    pCO2 4.43 kPa | 0
    bicarbonate 4.7 mmol/L | 0
    sodium 135 mmol/L | 0
    potassium 5.1 mmol/L | 0
    urine analysis revealed glucosuria | 0
    urine analysis revealed ketonuria |E0
    insulin infusion | 0
    intravenous saline | 0
    potassium replacement | 0
    symptomatic respiratory treatment | 0
    hypotension | 0
    volume expansion | 0
    vasopressors | 0
    inotropes | 0
    severe dyspnea | 24
    increased tachypnea | 24
    restlessness | 24
    cyanosis | 24
    diffuse crackles in all lung areas | 24
    diffuse rhonchi in all lung areas | 24
    hypoxemia confirmed | 24
    chest radiograph showed bilateral severe diffuse infiltrates | 24
    no cardiomegaly | 24
    acute respiratory failure secondary to ARDS diagnosed | 24
    transferred to the intensive care unit | 24
    oxygen by facemask | 24
    endotracheal intubation | 48
    mechanical ventilation required | 48
    throat culture positive for group A beta-hemolytic streptococci | 48
    cultures of urine negative | 48
    cultures of blood specimens negative | 48
    intravenous co-amoxiclav administered every 8 hours | 48
    clinical deterioration | 48
    transferred to our hospital | 48
    intubated on admission | 48
    mechanically ventilated by transport ventilator | 48
    FiO2 56% | 48
    arterial oxygen saturation 95% | 48
    respiratory rate 25 breaths per minute | 48
    heart rate 136 beats per minute | 48
    blood pressure 113/75 mm Hg | 48
    afebrile | 48
    sedated | 48
    diffusely edematous | 48
    leukocyte count 18.3 | 48
    neutrophils 67% | 48
    lymphocytes 25% | 48
    monocytes 7% | 48
    eosinophil 1% | 48
    prothrombin time normal | 48
    platelet count normal | 48
    troponin T level normal | 48
    liver function tests normal | 48
    serum amylase levels normal | 48
    urine amylase levels normal | 48
    urine analysis glucosuria noted | 48
    cultures of tracheal tube negative | 48
    cultures of urine negative | 48
    cultures of blood specimens negative | 48
    electrocardiography pattern normal | 48
    chest high-resolution computed tomography bilateral areas of patchy abnormalities | 48
    chest high-resolution computed tomography mixed ground-glass appearance | 48
    chest high-resolution computed tomography consolidation | 48
    predominantly in the right middle and left upper lobes | 48
    no cardiomegaly | 48
    no mediastinal lymphadenopathy | 48
    treatment with antibiotics continued for 10 days | 48
    subcutaneous injections of regular insulin replaced i.v. insulin | 72
    euglycemia maintained | 72
    weaned from ventilator | 96
    euglycemic | 96
    no ketonuria | 96
    subcutaneous regular insulin continued | 96
    good recovery | 168
    blood gas levels improved steadily | 168
    on room air after 7 days of hospital stay | 168
    all respiratory symptoms cleared | 168
    chest x-ray markedly improved | 168
    definitive diagnosis ARDS in association with DKA | 0
    type 1 diabetes mellitus diagnosed | 0
    survived without significant sequels | 168
    