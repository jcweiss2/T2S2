29 years old | 0
    female | 0
    native mitral valve endocarditis | 0
    native aortic valve endocarditis | 0
    active IVDU | 0
    presented to the Emergency Department | 0
    mother of two young children | 0
    poor social support network | 0
    underplayed severity of cardiac condition | 0
    no willingness to quit IVDU | 0
    no engagement in rehabilitation programs | 0
    initial decision for conservative treatment | 0
    antibiotic therapy | 0
    severe cardiogenic shock | -72
    severe aortic valve regurgitation | -72
    severe mitral valve regurgitation | -72
    referred for emergency inpatient cardiac surgery | -72
    obtained mother's consent | -72
    complex cardiac surgical procedure | -72
    aortic valve replacement | -72
    complex mitral valve repair | -72
    unable to wean off cardiopulmonary bypass | -72
    severe biventricular dysfunction | -72
    postcardiotomy venoarterial ECMO | -72
    clinical progress | 120
    failed attempt to wean off ECMO | 120
    mechanical circulatory support discontinued | 120
    remained in ICU | 120
    continuation of recovery | 120
    discharged to local convalescence center | 1800
    continuation of rehabilitation | 1800
    peak of COVID-19 pandemic | 0
    shortage of ICU beds | 0
    shortage of nurses | 0
    shortage of cardiac surgical operating rooms | 0
    ECMO machine unavailability | 0
    perfusionist unavailability | 0
    high-risk cardiac surgical procedure | 0
    unwilling to quit IVDU | 0
    high possibility of prosthetic valve endocarditis | 0
    lack of evidence for postcardiotomy ECMO | 0
    absence of bail-out strategies | 0
    contraindication for long-term mechanical support | 0
    contraindication for heart transplantation | 0
    rationing of resources | 0
    scarcity of resources | 0
    severe limitation on available resources | 0
    native valve endocarditis managed medically | 0
    valvular abscesses | 0
    large vegetation size | 0
    bradyarrhythmias | 0
    severe valve dysfunction | 0
    surgical intervention required | 0
    repeat surgical intervention | 0
    perioperative mortality | 0
    risk of prosthetic valve reinfection | 0
    prosthetic valve endocarditis | 0
    sepsis | 0
    renal failure | 0
    heart failure | 0
    patient-centered decision | 0
    tailored decisions to clinical goals | 0
    tailored decisions to social situation | 0
    emphasis on patient's wellbeing | 0
    respecting patient autonomy | 0
    beneficence | 0
    nonmaleficence | 0
    justice | 0
    curative treatment option | 0
    postoperative complications | 0
    massive consumption of resources | 0
    stewardship | 0
    deterioration | -72
    discussions regarding best mode of action | 0
    decision to perform surgery | 0
    contingency plan of rehabilitation | 0
    close community follow-up | 0
    organization support from Street Health | 0
    postoperative support | 0
    aid for substance use issues | 0
    plans to protect children | 0
    ECMO support required | -72
    no previous reports of postcardiotomy ECMO | 0
    limited experience with percutaneous ECMO | 0
    longer hospital stays | 0
    higher complication rates | 0
    ethical decision to use ECMO | 0
    allocation of perfusionist | 0
    reduction in cardiac operations | 0
    rationed ECMO use | 0
    stringent selection criteria | 0
    moral distress | 0
    consumption of resources | 0
    questioned patient's ability to appreciate harm | 0
    decision to pursue ECMO | 0
    survival | 0
    future rehabilitation | 0
    postcardiotomy ECMO as short-term support | 0
    high morbidity | 0
    high mortality | 0
    bridge to recovery | 0
    bridge to definitive therapy | 0
    long-term ventricular assist device | 0
    cardiac transplantation | 0
    limited evidence for patient selection | 0
    contraindication for long-term support | 0
    active substance abuse | 0
    need for social support | 0
    heart transplantation as high-risk procedure | 0
    immunosuppression required | 0
    satisfactory social support network required | 0
    no reports of heart transplants in active IVDU | 0
    infection spread risk | 0
    limited social support | 0
    options dependent on IVDU abstinence | 0
    potential LVAD | 0
    potential cardiac transplantation | 0
    allocation of scarce resources | 0
    COVID-19 pandemic strain | 0
    stringent eligibility criteria | 0
    active IVDU as contraindication | 0
    vast resource limitations | 0
    decision to pursue ECMO despite limitations | 0
    long recovery | 1800
    multidisciplinary team approach | 0
    postoperative abstinence from IVDU | 1800
    education on IVDU dangers | 1800
    intensive counseling | 1800
    changed patient's mind | 1800
    adamant promise to abstain | 1800
    one-month follow-up | 2160
    close follow-up | 2160
    conflict of interest declared | 0
    no financial support | 0