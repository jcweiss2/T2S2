69 years old | 0
female | 0
admitted to the ENT Department | 0
osteonecrosis involving upper and lower jaw | -1440
breast cancer surgery | -7920
zoledronic acid therapy | -6480
diabetes | 0
atrial fibrillation |
