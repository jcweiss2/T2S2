21 years old | 0
female | 0
admitted to the hospital | 0
premature rupture of membranes | 0
abdominal pain | 0
unplanned pregnancy | -2800
5 prenatal check-ups | -2800
alert | 0
normal vital signs | 0
fetal movement | 0
fetal heart rate 145 beats per minute | 0
cervix without cervical changes | 0
normal hemogram | 0
negative COVID-19 antigen test | 0
normal biophysical profile | 0
reactive fetal monitoring | 0
irregular uterine dynamics | 0
PROM in the prepartum phase | 0
vaginosis | 0
hospitalized for labor induction | 0
oxytocics | 0
failed labor induction | 23
bradycardia | 23
hypotension | 23
desaturation | 23
cardiorespiratory arrest | 23
advanced resuscitation maneuvers | 23
mechanical ventilation | 23
sulbactam ampicillin | 23
tranexamic acid | 23
dexamethasone | 23
newborn Apgar score 7 points at 1 minute | 23
newborn Apgar score 8 points at 5 minutes | 28
newborn Apgar score 9 points at 10 minutes | 33
fibrinogen 346 mg/dL | 24
arterial blood gasses without oxygenation disorders | 24
normal coagulation times | 24
lactate dehydrogenase 1.203 IU/L | 24
D-dimer >10,000 ng/mL | 24
pulmonary embolism | 24
pulmonary edema | 24
left pneumothorax | 24
respiratory infection | 24
polymerase chain reaction positive for SARS-CoV-2 | 24
elevated risk of pneumonia | 24
mild respiratory distress syndrome | 24
sepsis of pulmonary origin | 24
cardiogenic shock | 24
intensive care unit | 24
favorable clinical evolution | 120
mechanical ventilation withdrawn | 120
leukocytes 6250 × 103/mm3 | 120
neutrophils 60% | 120
procalcitonin <0.05 ng/mL | 120
blood cultures negative | 120
urine cultures negative | 120
orotracheal tube culture negative | 120
satisfactory recovery | 144
discharged from the hospital | 144