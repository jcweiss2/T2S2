72 years old | 0
male | 0
presented to the emergency department | 0
progressive shortness of breath | -72
intermittent chest pain | -72
altered level of consciousness | 0
significant respiratory distress | 0
heart rate of 122 beats/min | 0
blood pressure of 86/46 mmHg | 0
respiratory rate of 43 breaths/min | 0
oxygen saturations of 78% on room air | 0
temperature of 37.8°C | 0
sinus tachycardia | 0
thready central and peripheral pulses | 0
elevated jugular venous pressure | 0
S1 and S2 present | 0
absence of murmurs | 0
absence of extra heart sounds | 0
extremities mottled and cool | 0
bilateral peripheral edema | 0
breath sounds diminished at the lung bases | 0
diffuse crepitations bilaterally | 0
abdominal examination unremarkable | 0
mechanical ventilation | 0
hypertension | -inf
dyslipidemia | -inf
type 2 diabetes mellitus | -inf
oral anti-hyperglycemic medications | -inf
40 pack-year smoking history | -inf
atypical chest discomfort | -inf
myocardial perfusion imaging demonstrating mild ischemia in LAD territory | -inf
medical therapy | -inf
coronary angiogram scheduled | -inf
chest X-ray consistent with severe interstitial pulmonary edema | 0
inferolateral ST-segment elevation | 0
white blood cell count 8.4 × 10^9/L | 0
hemoglobin 104 g/L | 0
whole blood lactate 4.0 mmol/L | 0
creatinine kinase 1,178 μ/L | 0
high sensitivity troponin T 3,482 ng/L |,0
Killip IV inferolateral ST-segment elevation myocardial infarction | 0
intubated for hypoxemic respiratory failure | 0
emergency coronary angiogram | 0
culprit lesion in proximal to mid LAD | 0
revascularized with 2 drug-eluting stents | 0
chronic total occlusion of mid right coronary artery | 0
collaterals from LAD and left circumflex | 0
intra-aortic balloon pump | 0
transthoracic echocardiogram showing severe left ventricular dysfunction | 24
ejection fraction estimated at 20% | 24
akinesis of mid to distal anterior, apex, inferior, and lateral walls | 24
absence of left ventricular thrombus | 24
absence of hemodynamically significant valvular disease | 24
absence of pericardial effusion | 24
absence of myocardium abnormalities | 24
shock state persisted | 24
intra-aortic balloon pump requirement | 24
vasoactive medications | 24
inotropic medications | 24
norepinephrine | 24
vasopressin | 24
phenylephrine | 24
dobutamine | 24
oliguric renal failure | 24
continuous renal replacement therapy | 24
borderline fevers | 24
suspected mixed septic and cardiogenic shock | 24
broad spectrum antimicrobial therapy | 24
piperacillin/tazobactam | 24
vancomycin | 24
blood cultures positive for gram-negative bacilli | 36
Enterobacter cloacae | 36
antimicrobial therapy escalated to meropenem | 36
differential diagnoses considered | 24
mixed distributive/septic and cardiogenic shock | 24
recurrent ischemia secondary to stent complication | 24
evolving mechanical complication of ACS | 24
ventricular free wall rupture | 24
ventricular septal rupture | 24
papillary muscle rupture | 24
acute mitral regurgitation | 24
abrupt pulseless electrical activity cardiac arrest | 48
large circumferential pericardial effusion | 48
emergency pericardiocentesis | 48
arterial blood drained from pericardium | 48
pericardial effusion reaccumulated | 48
refractory cardiac tamponade | 48
mechanical circulatory support considered | 48
uncontrolled septicemia | 48
multiorgan dysfunction | 48
baseline frailty | 48
prohibitive surgical risk | 48
resuscitation unsuccessful | 48
left ventricular free wall rupture | 48
death | 48
autopsy showing large transmural myocardial infarction | 48
extensive necrosis | 48
multiple myocardial abscesses involving both ventricles | 48
gram-negative rods in myocardium | 48
left ventricular free wall rupture of mid inferior wall | 48
hemopericardium | 48
severe acute pyelonephritis of left kidney | 48
septic shock with E. cloacae bacteremia | 48
acute pyelonephritis | 48
acute myocardial ischemia | -inf
myocardial abscess formation | 48
tissue friability | 48
mechanical complications after AMI | 48
ventricular free wall rupture | 48
ischemic myocardial necrosis | 48
septic myocardial abscess | 48
myocardial abscess formation at site of ischemic myocardial necrosis | 48
metastatic spread into necrotic tissue | 48
respiratory infection source | 48
urinary tract infection source | 48
skin and soft tissue infection source | 48
Staphylococcus species | 48
Streptococcal species | 48
anaerobic myocardial abscess | 48
hypoxic postinfarction environment | 48
bacteremia | 24
persistent fever despite antimicrobials | 24
progressive hemodynamic deterioration | 24
focused application of echocardiography | 24
wall thickening | 24
honeycomb appearance to myocardium | 24
fistulous tracts draining into pericardium | 24
fatal clinical course | 48
contained rupture of abscess after AMI | 48
early identification of myocardial abscesses | 48
early identification of ventricular free wall rupture | 48
extracorporeal membrane oxygenation | 48
surgical repair | 48
mortality rate >50% | 48
left ventricular free wall rupture at site of septic myocardial abscess | 48
fatal outcome | 48
elevated jugular venous pressure |,0
high sensitivity troponin T 3,482 ng/L | 0
