57 years old | 0
male | 0
admitted to the emergency department | 0
right flank pain | 0
high fever | 0
poor health | 0
urosepsis | 0
referred to the urology department | 0
right nephrolithotomy | - (approximated as prior to admission, but exact timing not specified)
kidney stones | - (approximated as prior to admission, but exact timing not specified)
stenting | - (approximated as prior to admission, but exact timing not specified)
coronary heart disease | - (approximated as prior to admission, but exact timing not specified)
multiple kidney stones | 0
pyonephrosis | 0
renal cyst approximately 13 cm in size | 0
non-functional right kidney | 0
nephrostomy catheter insertion | 0
intravenous antibiotic therapy | 0
preoxygenation with 100% oxygen | 0
anesthesia induced with thiopental 400 mg | 0
anesthesia induced with rocuronium 50 mg | 0
anesthesia maintained with sevoflurane 1.5% | 0
N2O : O2 (50% : 50%) | 0
endotracheal intubation with 8.0 mm ID tube | 0
laparoscopy started | 0
converted to open surgery | 0
very adherent tissues | 0
kidney tissue removed | 0
cyst removed | 0
cyst ruptured at 50th minute of operation | 50
cyst content diffused to retroperitoneal area | 50
aspiration of retroperitoneal area | 50
irrigation of retroperitoneal area | 50
operation continued for 40 minutes after rupture | 50
duration of anaesthesia 100 minutes | 0
hemodynamic parameters stable | 0
extubated at end of surgery | 100
difficulty in breathing | 115
agitated | 115
blood gas analysis taken 18 minutes after extubation | 118
hypoxaemia | 118
pH: 7.49 | 118
pO2: 54 mmHg | 118
pCO2: 30 mmHg | 118
HCO3: 23 | 118
SpO2: 88 | 118
taken to intensive care unit | 115
conscious in ICU | 115
right lung sounds decreased | 115
serious respiratory distress | 115
chest X-ray revealed pleural effusion | 115
respiratory distress decreased after thoracentesis | 115
chest tube insertion | 115
cultures of pleural effusion | 115
cultures of cyst fluid | 50
Klebsiella pneumoniae | 115
imipenem 500 mg qid | 115
linezolid 600 mg bid | 115
metronidazole 500 mg tid | 115
intact diaphragm during surgery | 0
no defect on CT | 115
retroperitoneal fluid transition through diaphragmatic pores | 50
general condition improved | 115
antibiotic therapy | 115
drainage of pleural fluid | 115
pathology report indicated chronic pyelonephritis | 115
referred to urology department 4 days after surgery | 96
improvement in blood gas values | 96
pH: 7.35 | 96
pO2: 88 mmHg | 96
pCO2: 36 mmHg | 96
HCO3: 24 | 96
SpO2: 96 | 96
improvement in respiratory parameters | 96
improvement in chest radiography | 96
chest tube removed twelve days later | 288
discharged as healthy | 288
