71 years old | 0
female | 0
thyroid excision | -6720
spinal fusion | -6720
follicular thyroid cancer | -6720
metastasis to lungs | -6720
metastasis to cranial bones | -6720
metastasis to vertebrae | -6720
recurrence of spinal metastasis | -168
acetaminophen | -168
loxoprofen | -168
morphine | -168
dyspnea | 0
admitted to emergency department | 0
pulse 118 beats per minute | 0
blood pressure 121/86 mmHg | 0
respiratory rate 28 breaths per minute | 0
oxygen saturation level 96% | 0
no significant heart murmurs | 0
ST-segment elevation in leads I, aVL, and V2-5 | 0
cardiothoracic ratio 71% | 0
pulmonary congestion | 0
infiltrative shadow | 0
apical akinesis | 0
basal hyperkinesis | 0
leukocyte count 10,900 /μL | 0
C-reactive protein 27.7 mg/dL | 0
troponin T 0.16 mg/dL | 0
creatinine kinase 76 U/L | 0
N-terminal pro-brain natriuretic peptide 14,856 pg/mL | 0
left ventricular wall motion abnormalities | 0
Takotsubo syndrome | 0
treatment for heart failure | 0
treatment for pneumonia | 0
non-invasive positive pressure ventilation | 0
intravenous nitroglycerin | 0
furosemide | 0
heparin | 0
piperacillin tazobactam | 0
persistent ST-segment elevation in leads V2-5 | 48
worsening dyspnea | 216
harsh, loud, holosystolic murmur | 216
ventricular septal defect | 216
cardiac catheterization | 240
coronary angiography | 240
left ventriculography | 240
intra-aortic balloon pumping | 240
deeply inverted T-waves in leads V1-6 | 360
QT interval prolongation | 360
elective surgery | 384
extracorporeal circulation | 384
cardiac arrest | 384
VSP closed with Gore-Tex patch | 384
pathological examination | 384
loss of myocardial cells | 384
myocardial fibrosis | 384
lymphocyte and macrophage infiltration | 384
postoperative course uneventful | 384
cardiac magnetic resonance imaging | 1200
late gadolinium enhancement | 1200
discharged from hospital | 1512
follow-up electrocardiography | 8760
T-wave inversion in leads V1-5 | 8760
follow-up echocardiography | 8760
residual mild hypokinesis of apex | 8760