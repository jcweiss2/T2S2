5 weeks old | 0
infant | 0
congenital adrenal hyperplasia (CAH) | -792
admitted to the hospital | 0
fever | -24
fussiness | -24
cough | -96
runny nose | -96
hypoglycemia | -1152
respiratory distress | -1152
tachypnea | -1152
newborn screening test positive for CAH | -1152
cortisol level 1.2 mcg/dL | -1152
17-hydroxyprogesterone 813 ng/dL | -1152
ACTH stimulation test | -1152
post-stimulation 17 hydroxyprogesterone 17836 ng/dL | -1152
cortisol level 3.9 mcg/dL | -1152
hydrocortisone 30 mg/m²/day | -1152
fludrocortisone 0.1 mg daily | -1152
sodium chloride 2 grams | -1152
ER presentation | 0
no respiratory distress | 0
no diarrhea | 0
no vomiting | 0
no rash | 0
no decreased feeding | 0
afebrile | 0
oxygen saturation 100% | 0
irritable | 0
skin mottling | 0
no chest retractions | 0
no tachypnea | 0
no nasal flaring | 0
WBC 7.2 bil/L | 0
neutrophils 2.1 bil/L | 0
lymphocytes 2.5 bil/L | 0
monocytes 2 bil/L | 0
Na 136 mmol/L | 0
potassium 5.9 mmol/L | 0
HCO3 22 mmol/L | 0
glucose 110 mg/dL | 0
BUN 8 mg/dL | 0
creatinine 0.33 mg/dL | 0
CRP 1.9 mg/L | 0
SARS-CoV-2 detected | 0
blood culture negative | 0
urinalysis negative | 0
urine culture negative | 0
chest x-ray mild streaky bilateral perihilar streaks | 0
no focal consolidation | 0
no pleural effusions | 0
costophrenic angles clear | 0
unremarkable lung apices | 0
normal saline bolus | 0
maintenance IV fluids | 0
transferred to PICU | 0
hemodynamically stable | 0
fed appropriately | 0
no respiratory support | 0
discharged | 48
hydrocortisone weaned to home regimen | 48
doing well | 720
