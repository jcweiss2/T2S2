65 years old | 0
woman | 0
diagnosed with uveitis | -8760
bilateral cataracts | -8760
diabetes mellitus | -8760
palpitations | -25920
dizziness | -25920
sinoatrial block (SSS) | -25920
right bundle branch block | -25920
sinus arrest | -25920
dual-chamber pacemaker implantation | -25920
progressive dyspnoea | -26160
abnormal liver function | -26160
elevated brain natriuretic peptide (BNP) | -26160
decreased LVEF (62% to 51%) | -26160
heart failure with preserved ejection fraction | -26160
diuretics | -26160
angiotensin receptor antagonists | -26160
leg oedema | -26880
complete atrioventricular block | -26880
atrial-paced rhythm | -26880
ventricular-paced rhythm | -26880
hospitalized for worsening heart failure | -26880
junctional escape rhythm | -26880
atrial pacing failure | -26880
ventricular pacing failure | -26880
biventricular systolic dysfunction | -26880
giant right ventricular thrombus formation | -26880
anti-coagulant therapy with heparin | -26880
warfarin | -26880
pacemaker re-programming | -26880
cardiac arrest | -26880
temporary pacing electrode insertion into coronary sinus | -26880
transferred to hospital | -26880
ventricular pacing rhythm | 0
normal angiotensin converting enzyme | 0
normal calcium | 0
elevated soluble interleukin-2 receptor | 0
elevated BNP | 0
no significant stenosis on coronary angiography | 0
severe biventricular dysfunction | 0
reduced LVEF (30%) | 0
anteroseptal hypokinesis | 0
inferoseptal hypokinesis | 0
inferior wall dyskinesis | 0
severely dilated RV | 0
reduced TAPSE | 0
dilated tricuspid annulus | 0
severe tricuspid regurgitation | 0
right ventricular thrombus | 0
right atrial thrombus | 0
urgent thrombectomy | 24
removal of jugular vein pacemaker leads | 24
epicardial pacemaker implantation | 24
tricuspid annuloplasty | 24
endomyocardial biopsy confirming cardiac sarcoidosis | 24
cardiogenic shock | 48
intravenous dobutamine | 48
intravenous noradrenaline | 48
steroid pulse therapy | 48
maintenance steroid therapy | 48
LVEF improvement to 35% | 264
discharge | 1896
bisoprolol | 1896
enalapril | 1896
spironolactone | 1896
empagliflozin | 1896
warfarin | 1896
prednisolone | 1896
PET-CT showing no myocardial inflammation | 4368
sustained ventricular tachycardia | 10392
implantable cardioverter defibrillator | 10392
refractory ventricular electrical storm | 12720
mechanical ventilation | 12720
deep sedation | 12720
intravenous amiodarone | 12720
intravenous lidocaine | 12720
fever | 12720
arterial hypotension | 12720
leukocytosis | 12720
methicillin-resistant Staphylococcus epidermidis bacteraemia | 12720
Candida albicans bacteraemia | 12720
sepsis | 12720
death | 15528
