53 years old | 0
male | 0
admitted to the emergency department | 0
fever | -192
dry cough | -192
myalgia | -192
shortness of breath | -72
vomiting | -24
nonspecific epigastric discomfort | -24
denies chest pain | 0
Type-2 diabetes mellitus | 0
hypertension | 0
inferior MI in 2015 | -4824
coronary angiography refused | -4824
severe distress | 0
tachypneic | 0
tachycardiac | 0
normotensive | 0
O2 saturation of 93% | 0
body temperature normal | 0
severely breathless | 0
hypoxic | 0
crackles in both lung fields | 0
cardiac examination normal | 0
no significant repolarization abnormality | 0
1 mm ST elevation at lead V3 | 0
severe left ventricular systolic dysfunction | 0
estimated left ventricular ejection fraction of 35% | 0
segmental wall motion abnormalities | 0
bilateral patchy consolidative changes | 0
air space opacities | 0
intubated | 0
mechanical ventilation | 0
adult respiratory distress syndrome | 0
acute heart failure | 0
intravenous nitrates | 0
diuretics | 0
antibiotics | 0
oral aspirin | 0
clopidogrel | 0
enoxaparin | 0
noradrenaline | 0
polymerase chain reaction positive for CoV-2 | 0
biological inflammatory syndrome | 0
leukocytes 12.8 × 10^3/uL | 0
lymphocytes 0.5 | 0
C-reactive protein 150 mg/L | 0
ferritin 1979 ug/L | 0
troponin-T high sensitive 527 ng/L | 0
N-terminal-proB-type natriuretic peptide 722 pg/mL | 0
lactic acid 7.2 mmol/L | 0
admitted to intensive care unit | 0
serial ECG showed biphasic T wave | 0
inverted T waves | 0
peak cTn 1806 | 24
good response to medical therapy | 48
less oxygen requirement | 48
severely agitated | 72
hypotension | 72
severe bradycardia | 72
asystole | 72
return of spontaneous circulation | 72
worsening lactic acidosis | 72
pH 6.8 | 72
lactate concentration 19 mmol/L | 72
oxygen saturation 60% | 72
diffuse ST depression | 72
ST elevation in lead aVR | 72
taken to cath lab | 78
emergent coronary angiography | 78
tight stenosis of LAD | 78
normal flow | 78
tight ostial stenosis of obtuse marginal branch | 78
totally occluded mid-right coronary artery | 78
everolimus-eluting stent deployed | 78
ECG changes improved | 78
mechanical ventilation | 0
noradrenaline | 0
multiple antibiotics | 0
antivirals | 0
plasma protein fraction | 0
hydroxychloroquine | 0
acute kidney injury | 0
acute liver injury | 0
complete recovery of renal function | 408
complete recovery of liver function | 408
inflammatory markers normalized | 408
discharged home | 504