56 years old | 0
male | 0
type 2 diabetes mellitus | -8760
chronic obstructive pulmonary disease | -8760
obstructive sleep apnea | -8760
coronary artery disease | -8760
heart failure with preserved ejection fraction | -8760
tobacco abuse disorder | -8760
alcohol use disorder | -8760
admitted to the hospital | 0
septic shock | 0
left lower extremity osteomyelitis | 0
intubated | 0
drinking 5 beers daily on weekdays | -2160
drinking 5 to 10 beers on weekends | -2160
eating frozen meals | -2160
positive blood cultures for methicillin-sensitive Staphylococcus aureus | 0
treated with antibiotics | 0
vascular surgery consulted | 0
no surgical intervention | 0
infectious diseases consulted | 0
pressor support | 0
antibiotic treatment | 0
rash on presentation | 0
petechiae | 0
palpable hemorrhagic lesions | 0
vasculitis | 0
normal white blood cell count | 0
slightly low hemoglobin | 0
normal mean corpuscular volume | 0
normal platelet count | 0
elevated creatinine | 0
elevated erythrocyte sedimentation rate | 0
elevated C-reactive protein | 0
immunologic work up | 0
negative antinuclear antibody | 0
negative antineutrophil cycloplasmic antibody | 0
elevated Complement C3 | 0
normal Complement C4 | 0
negative HIV and hepatitis panel | 0
nutritional deficiency considered | 0
plasma vitamin C levels drawn | 0
started on 500 mg IV vitamin C daily | 0
low plasma vitamin C levels | 0
diagnosis of ascorbic acid deficiency | 0
skin findings improved | 24
mentation improved | 24
resolution of inflammatory markers | 24
resolution of elevated creatinine | 24
discharged | 168