5 years old | 0
male | 0
Crohn's disease | -720
brother with Crohn's disease | -720
history of bronchiolitis | -720
infliximab treatment | -96
protein-losing enteropathy | -96
recurrent intestinal pseudo-obstruction | -96
admitted to hospital | 0
abdominal pain | 0
bloody stool | 0
colectomy | 0
pneumonia | 24
acute respiratory distress syndrome (ARDS) | 24
ventilated | 24
fever | 24
hypotension | 24
tachycardia | 24
tachypnea | 24
bilateral crackles | 24
arterial blood pH: 7.10 | 24
pCO2: 55 | 24
pO2: 95 | 24
HCO3: 17 | 24
BE: −7 | 24
O2 saturation: 98% | 24
lactate: 6.8 | 24
hemoglobin: 9.9 g/dL | 24
white blood cell count: 19,300/mm3 | 24
platelets: 61,000/mm3 | 24
peripheral blood smear: Increased neutrophil band count | 24
C-reactive protein (CRP): 10 mg/dL | 24
procalsitonin: 100 ng/mL | 24
diffuse infiltration and consolidation on chest radiography | 24
antibiotics initiated | 24
vasopressors initiated | 24
Pseudomonas aeruginosa detected | 48
oliguric renal failure | 48
continuous venovenous hemodialysis | 48
fever subsided | 168
laboratory findings back to normal except CRP | 168
cultures sterile | 168
weaning attempt failed | 336
re-intubated | 336
ventilator settings showed restrictive pattern | 336
high-resolution computerized tomography (HRCT) | 336
interlobular septal thickening | 336
air bronchograms | 336
consolidated areas with bronchiectasia | 336
ground glass opacities | 336
cytological evaluation of deep tracheal aspirates | 336
neutrophilic infiltration | 336
tracheostomy | 552
prednisolone initiated | 552
clinical condition and pulmonary functions improved | 648
CRP returned to normal | 648
discharged from PICU | 768