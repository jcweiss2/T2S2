22 years old | 0 | 0 
male | 0 | 0 
admitted to the hospital | 0 | 0 
mild COVID-19 illness | -720 | -720 
sore throat | -720 | -720 
loss of sense of smell | -720 | -720 
positive COVID-19 PCR | -720 | -720 
recovery from COVID-19 | -720 | -336 
received first dose of inactivated SARS-CoV-2 vaccine | -336 | -336 
asymptomatic | -336 | -24 
received second dose of inactivated SARS-CoV-2 vaccine | -24 | -24 
headache | -24 | 0 
fatigue | -24 | 0 
fever | 0 | 168 
sore throat | 0 | 168 
abdominal pain | 0 | 168 
high-grade fever | 96 | 168 
myalgia | 96 | 168 
nausea | 96 | 168 
vomiting | 96 | 168 
diarrhea | 96 | 168 
faint erythematous non-itchy rash | 96 | 168 
dry irritant cough | 96 | 168 
no shortness of breath | 96 | 168 
no chest discomfort | 96 | 168 
no urinary symptoms | 96 | 168 
no pain or swelling of joints | 96 | 168 
temperature of 39°C | 0 | 0 
systolic blood pressure of 110 mm Hg | 0 | 0 
tachycardia | 0 | 168 
dry mucous membranes | 0 | 0 
congested throat | 0 | 0 
bilateral conjunctival injection | 0 | 0 
left conjunctival hemorrhage | 0 | 0 
generalised erythematous maculopapular rash | 0 | 168 
peripheral lymph nodes not enlarged | 0 | 0 
no audible cardiac murmurs | 0 | 0 
chest clear to auscultation | 0 | 0 
abdomen examination unremarkable | 0 | 0 
SARS-CoV-2 PCR negative | 0 | 0 
SARS-CoV-2 IgG positive | 0 | 0 
throat swab negative for group A streptococcus | 0 | 0 
sputum culture showed mixed flora | 0 | 0 
bacterial blood cultures negative | 0 | 0 
urinalysis showed significant proteinuria | 0 | 168 
ANA negative | 0 | 0 
dsDNA negative | 0 | 0 
c-ANCA negative | 0 | 0 
p-ANCA negative | 0 | 0 
C3 reduced | 0 | 0 
C4 reduced | 0 | 0 
WBC 15 | 0 | 0 
platelet 122 | 0 | 0 
creatinine 115 | 0 | 0 
AST 53 | 0 | 0 
ALT 81 | 0 | 0 
direct bilirubin 35 | 0 | 0 
albumin 16 | 0 | 0 
C reactive protein 249 | 0 | 168 
ferritin 4357 | 0 | 168 
D-dimer 14 | 0 | 168 
procalcitonin 9 | 0 | 168 
interleukin-6 90 | 0 | 168 
admitted to ICU | 0 | 0 
treated with ceftriaxone | 0 | 48 
treated with levofloxacin | 0 | 48 
treated with intravenous hydrocortisone | 0 | 48 
blood pressure stabilised | 48 | 48 
fever persisted | 48 | 168 
facial puffiness | 48 | 168 
generalised body oedema | 48 | 168 
tachycardia persisted | 48 | 168 
diarrhea persisted | 48 | 168 
myalgia | 48 | 168 
renal impairment | 48 | 168 
significant proteinuria | 48 | 168 
ECG showed sinus tachycardia | 48 | 48 
non-specific T-wave abnormalities | 48 | 48 
troponin-I raised | 48 | 48 
pro-BNP over 8000 | 48 | 48 
transthoracic echocardiogram showed severe tricuspid regurgitation | 48 | 48 
pulmonary hypertension | 48 | 48 
right atrium and ventricle moderately dilated | 48 | 48 
left ventricle cavity size normal | 48 | 48 
mildly reduced ejection fraction | 48 | 48 
thin rim of pericardial effusion | 48 | 48 
computed topography scan of chest showed bilateral moderate pleural effusion | 48 | 48 
basal atelectasis | 48 | 48 
discharged from ICU | 168 | 168 
treated with dexamethasone | 168 | 216 
generalised oedema subsided | 168 | 216 
skin rash resolved | 168 | 216 
conjunctivitis resolved | 168 | 216 
white blood cell count normalised | 168 | 216 
renal function improved | 168 | 216 
inflammatory markers came down to normal levels | 168 | 216 
repeat transthoracic echocardiography showed trace tricuspid regurgitation | 216 | 216 
right ventricular systolic function improved | 216 | 216 
pulmonary artery systolic pressure normalised | 216 | 216 
discharged from hospital | 216 | 216 
treated with oral prednisolone | 216 | 240 
follow-up in outpatient clinic | 240 | 240 
symptoms resolved | 240 | 240 
general weakness and fatigue | 240 | 240 
repeat echocardiogram completely normal | 240 | 240