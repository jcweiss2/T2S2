74 years old | 0
male | 0
height: 157.6 cm | 0
weight: 50.7kg | 0
squamous cell carcinoma | -720
neoadjuvant chemotherapy | -720
marginal mandibulectomy | 0
left supraomohyoid neck dissection | 0
reconstruction with reconstruction plate | 0
right radial forearm free flap | 0
general anesthesia | 0
no medical morbidities | 0
no hypertension | 0
no diabetes | 0
normal preoperative laboratory findings | 0
normal chest radiograph | 0
sinus arrhythmia | 0
low voltage in frontal leads | 0
ST elevation | 0
normal transthoracic echocardiogram | 0
hemodynamically stable | 0
transported to ICU | 0
nasotracheal tube | 0
ventilation with Ambu bagging | 0
oxygen 7 L/min | 0
100% peripheral oxygen saturation | 0
elevated blood pressure | 1
elevated heart rate | 1
pain | 1
analgesics administered | 1
opioids administered | 1
high blood pressure | 1
persistent pain | 1
agitating | 1
dexmedetomidine administered | 1
sedation | 1
respiratory rate dropped | 1
SpO2 dropped | 1
BP dropped | 1
ST elevation in ECG | 1
serial ECGs checked | 1
ST elevation in anterior and lateral leads | 1
elevated cardiac markers | 1
myoglobin measurements surged | 1
Troponin I measurements rose | 1
serum creatine kinase MB peaked | 1
referred to cardiology department | 2
TTE performed | 2
dilated left ventricular | 2
normal LV wall thickness | 2
akinesia of apical lateral | 2
inferior wall and mid-cavity | 2
severe systolic dysfunction | 2
LV ventriculogram | 2
estimated ejection fraction 25% | 2
ischemic insult of multivessel territory | 2
stress-induced cardiomyopathy suspected | 2
transferred to medical ICU | 2
inotropics administered | 2
chronotropics administered | 2
diuretics administered | 2
hemodynamic monitoring | 2
dopamine administered | 2
dobutamine administered | 2
norepinephrine administered | 2
rapid clinical improvement | 48
ST-segment elevations normalized | 48
extubated | 120
transferred to general ward | 120
Troponin I levels normalized | 720
laboratory test values normalized | 720
no clinical signs of heart failure | 720
consolidation radiotherapy | 720
oral cavity lesions healing | 720
complete dentures prepared | 720
good condition | 720