44 years old | 0
    woman | 0
    HER-2/Neu + score of +3 infiltrating ductal carcinoma | 0
    transferred from Kuwait | 0
    hyporesponsive | 0
    tachycardic | 0
    hypotensive | 0
    temperature of 101.8°F | 0
    mechanically ventilated | 0
    received multiple rounds of chemotherapy | -672
    received radiation | -672
    craniotomy for resection of a tumor | -672
    increased intracranial pressure | -48
    aspiration pneumonia | -48
    intubation | -48
    presumed pneumonia | 0
    possibly meningitis | 0
    continued meropenem 2 g every 8 hours | 0
    provided medical support for septic shock | 0
    magnetic resonance imaging of the brain revealed mild hydrocephalus | 0
    large enhancing cavitary lesion in the right hemisphere | 0
    craniotomy performed to place a ventricular drain | 96
    assist in monitoring intracranial pressures | 96
    epidural swabs performed intraoperatively | 96
    intracavitary swabs performed intraoperatively | 96
    CSF cultures revealed heavy growth of Enterococcus faecalis | 96
    initiated on therapeutic doses of vancomycin | 96
    initiated on meropenem | 96
    nonresponsive despite no use of analgesics or sedatives | 96
    changed from meropenem and vancomycin to ampicillin plus gentamicin | 168
    subsequent CSF cultures from August 13 through 27 remained positive | 168
    tried to open her eyes for the first time | 240
    began to regain her strength on the right side | 240
    extubated | 288
    began to verbally communicate | 288
    improvement in mental status | 288
    cultures remained positive | 288
    vancomycin administered intraventricularly via the ventriculostomy drain | 456
    CSF vancomycin concentrations could not be monitored | 456
    monitored closely for neurological changes | 456
    intraventricular vancomycin administered on August 27 | 456
    intraventricular vancomycin administered on August 30 | 480
    intraventricular vancomycin administered on September 3 | 504
    clinical status continued to improve | 504
    first CSF culture returned negative | 648
    subsequent cultures negative | 672
    deemed safe enough to restart chemotherapy | 672
    deemed safe enough for further treatments for her cancer | 672
    infection free at six months | 4320
    continues to undergo physical therapy | 4320
    positive improvements | 4320

    44 years old | 0  
    woman | 0  
    HER-2/Neu + score of +3 infiltrating ductal carcinoma | 0  
    transferred from Kuwait | 0  
    hyporesponsive | 0  
    tachycardic | 0  
    hypotensive |9 0  
    temperature of 101.8°F | 0  
    mechanically ventilated | 0  
    received multiple rounds of chemotherapy | -672  
    received radiation | -672  
    craniotomy for resection of a tumor | -672  
    increased intracranial pressure | -48  
    aspiration pneumonia | -48  
    intubation | -48  
    presumed pneumonia | 0  
    possibly meningitis | 0  
    continued meropenem 2 g every 8 hours | 0  
    provided medical support for septic shock | 0  
    magnetic resonance imaging of the brain revealed mild hydrocephalus | 0  
    large enhancing cavitary lesion in the right hemisphere | 0  
    craniotomy performed to place a ventricular drain | 96  
    assist in monitoring intracranial pressures | 96  
    epidural swabs performed intraoperatively | 96  
    intracavitary swabs performed intraoperatively | 96  
    CSF cultures revealed heavy growth of Enterococcus faecalis | 96  
    initiated on therapeutic doses of vancomycin | 96  
    initiated on meropenem | 96  
    nonresponsive despite no use of analgesics or sedatives | 96  
    changed from meropenem and vancomycin to ampicillin plus gentamicin | 168  
    subsequent CSF cultures from August 13 through 27 remained positive | 168  
    tried to open her eyes for the first time | 240  
    began to regain her strength on the right side | 240  
    extubated | 288  
    began to verbally communicate | 288  
    improvement in mental status | 288  
    cultures remained positive | 288  
    vancomycin administered intraventricularly via the ventriculostomy drain | 456  
    CSF vancomycin concentrations could not be monitored | 456  
    monitored closely for neurological changes | 456  
    intraventricular vancomycin administered on August 27 | 456  
    intraventricular vancomycin administered on August 30 | 480  
    intraventricular vancomycin administered on September 3 | 504  
    clinical status continued to improve | 504  
    first CSF culture returned negative | 648  
    subsequent cultures negative | 672  
    deemed safe enough to restart chemotherapy | 672  
    deemed safe enough for further treatments for her cancer | 672  
    infection free at six months | 4320  
    continues to undergo physical therapy | 4320  
    positive improvements | 4320