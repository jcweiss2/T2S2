36 years old|0
female|0
presented to the emergency department|0
fever|-168
hemoptysis|-168
left-sided chest pain|-168
breathlessness|-168
active hemoptysis|0
chest pain|0
transferred to Medical Intensive Care Unit|0
resuscitation|0
evaluated for coronary artery diseases|0
electrocardiography|0
two-dimensional echo|0
cardiac markers|0
tests for HIV|0
tests for hepatitis B virus surface antigen|0
tests for HCV|0
tests for autoimmune profile|0
chest X-ray revealed mass lesion|0
sputum examination|0
Gram staining|0
culture reports|0
CT scan thorax with contrast study|0
planned CT-guided FNAC|0
cytological examination|0
Gram staining (FNAC sample)|0
Ziehl–Neelsen staining|0
aerobic culture|0
negative for malignant cells|0
presence of Gram-positive branching filaments|0
coccoid elements|0
conventional Ziehl–Neelsen staining negative for acid-fast bacilli|0
modified Ziehl–Neelsen staining showed partially acid-fast branching filaments|0
blood agar plate after incubation|0
colonies on blood agar|0
empirically put on third-generation cephalosporin|0
empirically put on azithromycin|0
confirm diagnosis of pulmonary nocardiosis|0
cotrimoxazole started|0
rashes all over the body|0
antibiotic treatment changed to imipenem|0
imipenem for 10-day duration|0
oral linezolid|0
chest X-ray revealed gradual resolution of pneumonia|0
cavitation|0
complete resolution of left upper lobe lesion|4320
no significant history of diabetes|0
no significant history of malignancy|0
no significant history of drug intake|0
temperature 102°F|0
respiratory rate 32/min|0
blood pressure 100/76 mm Hg|0
heart rate 108/min|0
SpO2 92% in room air|0
breath sound decreased on left side|0
crepitation present on left infraclavicular|0
crepitation present on left axillary|0
crepitation present on left interscapular area|0
rest systems within normal limits|0
negative HIV test|0
negative hepatitis B virus surface antigen test|0
negative HCV test|0
negative autoimmune profile|0
no pathogenic organism in sputum Gram staining|0
no pathogenic organism in sputum culture|0
no respiratory distress|0
FNAC sample sent for cytological examination|0
FNAC sample sent for Gram staining|0
FNAC sample sent for Ziehl–Neelsen staining|0
FNAC sample sent for aerobic culture|0
dry whitish-to-tan colonies on blood agar|0
raised, chalky white appearance of colonies|0
characteristic earthy odor of Nocardia species|0
filamentous bacteria in culture|0
negative for malignancy|0
negative toxemia|0
