81 years old | 0
male | 0
admitted to the hospital | 0
distal wound abscess | -720
femoropopliteal composite bypass | -720
critical limb ischemia | -720
MRSA infection | -720
alcoholic liver disease | 0
atrial fibrillation | 0
left carotid stenting | 0
endovascular exclusion of left iliac aneurysm | 0
no fever | 0
hemoglobin 12 g/dL | 0
INR 1.38 | 0
blood cultures negative | 0
very thin and emaciated | 0
BMI 15 | 0
abdomen treatable | 0
no masses palpable | 0
physical and laboratory examinations of heart and chest normal | 0
femoral pulses palpable bilaterally | 0
popliteal and tibial pulses absent bilaterally | 0
right femoropopliteal bypass patent | 0
valid flow at Duplex-scan examination | 0
no exposure of graft through infected wound | 0
anticoagulation using low-molecular-weight heparin | 0
intravenous antibiotic therapy using Teicoplanin 400 mg daily | 0
acute limb ischemia | 96
bypass thrombosis | 96
increase of white blood cells count | 96
fever | 96
surgical exploration of popliteal artery | 96
no run-off from tibial vessels | 96
graft removal | 96
right thigh amputation | 96
postoperative course uneventful | 120
white blood cells count normalized | 120
fever disappeared | 120
no additional signs of infection | 120
wound of stump clean | 120
antibiotic therapy with Teicoplanin continued | 120
discharged on ninth postoperative day | 216
referred to clinic for rehabilitation | 216
pulsatile mass in right side of neck | 648
pulsatile mass in left groin | 648
dysphagia | 648
hemoptysis | 648
duplex ultrasound of neck and left groin | 648
angio-computed tomography scan | 648
right hypodense bulk at common carotid artery | 648
bifurcation 40 x 37 mm in diameter | 648
extended for 58 mm in length | 648
involved ICA | 648
dislocated right internal jugular vein | 648
invaded nearby parapharyngeal space | 648
small hematoma enveloping left iliac-femoral passage | 648
re-referred to IRCCS Policlinico's Operative Unit of Vascular Surgery | 648
no fever | 648
Teicoplanin 200 mg twice daily | 648
INR 5.5 | 648
leukocytosis | 648
anemia | 648
huge palpable tender pulsatile mass in right neck | 648
smaller mass in left groin | 648
trans-thoracic color-Doppler echocardiography | 648
normal preoperative heart ejection fraction | 648
referred to operating room | 648
selective right internal carotid angiography | 648
voluminous pseudoaneurysm arising from carotid bifurcation | 648
extending toward nearby parapharyngeal space | 648
0.035-in hydrophilic stiff wire placed into ICA | 648
short 5F sheath exchanged with long guiding 10F sheath | 648
Fluency PTFE-covered nitinol self-expanding stent placed | 648
angiographic control showed patency of ICA | 648
complete exclusion of lesion | 648
absence of signs of endoleaks | 648
mass no more pulsatile | 648
surgical right laterocervical incision | 648
hematoma evacuated | 648
PTFE graft wrapped around carotid wall | 648
incision closed in layers | 648
left femoral pseudoaneurysm excised | 648
vessel wall reconstructed using small pericardial patch | 648
admitted to intensive care unit for 24 h | 648
returned to ward | 672
culture samples of laterocervical mass and left femoral pseudoaneurysm | 672
MRSA presence | 672
postoperative blood samples negative | 672
urine culture revealed ESBL Escherichia coli | 672
antibiotic therapy with Ceftriaxone 2 g twice daily | 672
dual therapy continued for 4 weeks | 672
postoperative course uneventful | 720
laterocervical wound and both groin wounds healed completely | 720
no signs of infection recurrence | 720
discharged on POD 15th | 936
acetyl salicylic acid 100 mg daily | 936
low-molecular-weight heparin | 936
referred to clinic for further rehabilitation | 936
angio-CT scan of neck showed regular patency of covered stent | 936
no signs of endoleaks | 936
duplex ultrasound showed no flow impairment | 936
7 months follow-up | 3528
poor general condition | 3528
laterocervical and inguinal wounds healed well | 3528
stent still patent | 3528