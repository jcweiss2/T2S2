58 years old | 0
male | 0
hypertension | 0
diabetes mellitus | 0
admitted to Intensive care unit (ICU) | 0
septic shock | -312
coronary artery bypass grafting | -312
mitral valve replacement | -312
invasive mechanical ventilation | 0
norepinephrine infusion | 0
deteriorated renal function | 0
preserved urine output | 0
febrile | 0
central venous catheter (CVC) in internal jugular site | -144
culture of CVC tip | 0
blood samples from catheter and peripheral vein | 0
urine culture | 0
bronchoalveolar lavage | 0
absence of sternal instability | 0
computed tomography (CT) scan | 0
transthoracic echocardiography | 0
transesophageal echocardiography | 0
absence of valvular abnormality | 0
vancomycin | 0
imipenem | 0
colistin | 0
worsened clinical condition | 0
Klebsiella pneumoniae isolated from catheter culture | 0
Klebsiella pneumoniae isolated from blood samples | 0
intermediate to amikacin | 0
resistant to imipenem | 0
resistant to colistin | 0
resistant to tigecycline | 0
presence of blaOXA-48 gene | 0
presence of blaVIM-2 gene | 0
presence of blaCMY-2 gene | 0
presence of blaSHV-1 gene | 0
vancomycin stopped | 0
colistin stopped | 0
amikacin | 0
imipenem increased dose | 0
continuous venovenous hemodiafiltration (CVVHDF) | 1
amikacin administration with CVVHDF | 0
amikacin dose increased | 0
hemodynamic improvement | 0
norepinephrine stopped | 120
decreased CRP | 0
decreased procalcitonin | 0
decreased leukocytes | 0
treatment tolerated for 14 days | 336
discharged from ICU | 432
serum creatinine similar to pre-admission | 432
audiometric test excluded ototoxicity | 432
Klebsiella pneumoniae producing carbapenemase | 0
septic shock due to CR-Kp bloodstream infection | -312
successful treatment with amikacin and imipenem combined with CVVHDF | 0
high therapeutic failure | 0
high mortality | 0
limited number of agents available | 0
colistin as first-line regimen | 0
colistin resistance emergence | 0
combination therapy associated with improved mortality | 0
aminoglycoside monotherapy | 0
aminoglycoside combination therapy | 0
amikacin plus colistin | 0
aminoglycoside plus carbapenem | 0
amikacin renal toxicity | 0
renal uptake of amikacin | 0
CVVHDF for extrarenal clearance | 0
high peak concentrations | 0
increased antimicrobial efficacy | 0
rapid decrease in drug levels | 0
survival benefit of high dose combination | 0
CVVHDF prevention of nephrotoxicity | 0
CVVHDF increased antimicrobial activity | 0
