58 years old | 0
Hispanic female | 0
admitted to the hospital | 0
trigeminal neuralgia | -672
hyperlipidemia | -672
upper respiratory tract infection | -168
cough | -168
shortness of breath | -168
low-grade fevers | -168
decadron 40 mg i.m | -168
prescription for antibiotics | -168
did not fill the prescription for the antibiotics | -168
shortness of breath and cough were getting worse | -24
seen in the emergency | -24
diagnosed with an acute airway obstruction | -24
acute epiglottitis | -24
emergently intubated | -24
transferred to the intensive care unit | -24
hypotensive | -24
hypoxemic | -24
ventilator support | -24
vasopressors | -24
chest x-ray showed extensive bilateral peri-hilar consolidation and infiltrates | 0
computed tomography (CT) scan of the chest | 0
diffuse bilateral interstitial and alveolar infiltrates | 0
bilateral lower lobe air space consolidation | 0
CT scan of the neck | 0
diffuse swelling of the soft tissues | 0
loss of the fat planes throughout the pharyngeal region | 0
marked thickening of the retropharyngeal soft tissue | 0
minimal cervical adenopathy | 0
leukocytosis | 0
borderline hematocrit level | 0
normal platelet count | 0
normal sodium | 0
normal renal function | 0
normal liver function tests | 0
arterial blood gas showed significant acidosis | 0
pH of 7.03 | 0
PaCO2 level of 46 mmHg | 0
PaO2 of 46 mmHg | 0
blood cultures were negative | 0
remained intubated in the ICU | 24
endoscopic evaluation | 24
unremarkable for any unusual pathology | 24
started on intravenous solumedrol | 48
chest x-rays performed on multiple occasions | 48
continued to show bilateral infiltrates | 48
multiple workups for a source of infection | 48
all negative | 48
serology for influenza | 48
serology for parainfluenza | 48
serology for Brucella | 48
serology for tuberculosis | 48
serology for Bordetella pertussis | 48
serology for atypical pathogens | 48
all negative | 48
broad-spectrum antibiotics | 48
antifungal (fluconazole 400 mg daily) | 48
eventually extubated | 240
transferred to the medical floor | 240
developed recurrent respiratory distress | 264
reintubation | 264
ICU readmission | 264
bronchoscopy | 264
did not reveal any abnormalities | 264
bronchoalveolar lavage | 264
lung biopsy | 264
normal | 264
developed evidence of a lower GI hemorrhage | 288
upper endoscopy | 288
non-contributory | 288
biopsy was not done | 288
planned colonoscopy | 288
could not be performed | 288
developed hypotension | 288
KUB showed massive pneumoperitoneum | 288
emergent laparotomy | 288
evaluated by Pathology | 288
serosal surface of the bowel showed a variable green discoloration | 288
areas of adherent fibrinopurulent exudate | 288
multiple small bowel perforations | 288
4 cm long cecal perforation | 288
mucosa showed several shallow ulcers | 288
areas of edema | 288
marked thinning | 288
microscopic sections showed innumerable invasive fungal elements | 288
vascular invasion | 288
vascular thrombosis | 288
hemorrhage | 288
acute inflammation | 288
necrosis | 288
fungal morphology was most consistent with Mucormycosis | 288
started on liposomal amphotericin B | 288
micafungin | 288
discontinued fluconazole | 288
additional intestinal resections | 288
final laparotomy | 294
near complete intestinal infarction | 294
progressive multiorgan failure | 294
ongoing shock | 294
diffuse intestinal ischemia and infarction | 294
condition was deemed terminal | 294
discussions with her family | 294
DNR status | 294
withdrawal of care | 294
patient succumbed to the illness | 294