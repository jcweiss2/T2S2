37 years old | 0
male | 0
healthcare worker | 0
admitted to the hospital | 0
fever | -672
lethargy | -672
diarrhoea | -672
symptoms subsided | -667
recurrence of symptoms | -336
fever | -336
diarrhoea | -336
dizziness | -336
presented to the emergency department | 0
dizziness | 0
pre-syncope | 0
clinically shocked | 0
febrile | 0
tachypnoeic | 0
oxygen saturation level of 97% | 0
raised jugular venous pressure | 0
coarse crepitations on auscultation | 0
global moderate-to-severe left ventricular systolic dysfunction | 0
ejection fraction (EF) 35-40% | 0
transferred to critical care | 0
commenced on milrinone | 0
commenced on noradrenaline | 0
worsening of myocardial function | 24
intravenous immunoglobulin | 24
hydrocortisone | 24
anticoagulated with a heparin infusion | 24
high-dose Vitamin B & C | 24
leucocytosis | 24
lymphopenia | 24
elevated troponin | 24
brain natriuretic peptide | 24
ferritin | 24
D-dimer | 24
acute kidney injury | 24
coagulopathic | 24
transaminitis | 24
procalcitonin | 24
nasopharyngeal swab | 24
nasopharyngeal swab | 72
nasopharyngeal swab | 120
commenced on linezolid | 120
commenced on clarithromycin | 120
commenced on piperacillin-tazobactam | 120
serial echocardiograms | 120
worsening biventricular function | 120
reduction in global LV ejection fraction | 120
worsening of right ventricular function | 120
LV wall thickening | 120
bi-atrial dilatation | 120
increased pulmonary artery systolic pressures | 120
initial improvement in myocardial function | 120
commenced on prednisolone | 168
rapid recovery in myocardial function | 168
biochemical improvement in cardiac function | 240
radiological improvement in cardiac function | 240
cardiac magnetic resonance | 240
evidence of myocarditis | 240
LV wall thickening | 240
inhomogeneity of T1/T2 mapping values | 240
patchy non-infarct pattern late gadolinium enhancement | 240
recovery of overall LV systolic function | 240
normalization of RV volumes and function | 240
SARS-CoV-2 IgG positive | 312
commenced on an angiotensin-converting enzyme inhibitor | 312
commenced on a beta-blocker | 312
commenced on a mineralocorticoid receptor antagonist | 312
discharged from hospital | 336
repeat CMR | 696
resolution of ventricular function | 696
small areas of patchy LGE persisted | 696
on a slowly weaning regimen of prednisolone | 4992
on a beta-blocker | 4992
on an angiotensin-converting enzyme inhibitor | 4992
on a mineralocorticoid receptor antagonist | 4992