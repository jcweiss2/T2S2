28 years old | 0
male | 0
admitted to the hospital | 0
AML | -780
gingival swelling | -780
bone marrow aspiration | -780
diagnosed with AML | -780
peripheral blood stem cell transplantation | -624
busulfan | -624
cyclophosphamide | -624
cyclosporine A | -624
methotrexate | -624
grade I acute GVHD | -624
methylprednisolone | -624
CsA discontinued | -468
molecular relapse of AML | -364
azacitidine | -364
gemtuzumab ozogamicin | -364
donor lymphocyte infusion | -364
molecular complete remission | -260
second bone marrow transplantation | -260
tacrolimus | -260
short-term methotrexate | -260
skin and gut GVHD | -260
cytomegalovirus enterocolitis | -260
discharged | -156
bronchiolitis obliterans | -104
high-dose pulse mPSL therapy | -104
mycophenolate mofetil | -104
hematological relapse of AML | 0
recurrent pneumonia | 0
watery diarrhea | 0
maculopapular skin rash | 0
infiltrative shadow in the inferior lobe of the left lung | 0
meropenem | 0
vancomycin | 0
salvage chemotherapy | 4
mitoxantrone | 4
etoposide | 4
intermediate-dose cytarabine | 4
diarrhea worsened | 10
maculopapular skin rash expanded | 10
intestinal edema observed on CT | 10
mPSL increased | 10
beclomethasone dipropionate prescribed | 10
steroid pulse therapy | 13
colonoscopy not possible | 13
hemorrhagic diarrhea developed | 16
blood cultures positive for Gram-negative bacilli | 16
minocycline prescribed | 16
ciprofloxacin prescribed | 16
Gram-negative bacilli identified as S. maltophilia | 17
minocycline changed to trimethoprim-sulfamethoxazole | 17
patient died | 18
autopsy revealed erosion and petechial hemorrhaging | 18
Gram-negative bacilli found in all layers of the ileum | 18
hemorrhagic pneumonia caused by S. maltophilia | 18