33 years old | 0
male | 0
sub-Saharan African origin | 0
admitted to the intensive care unit | 0
severe hypotension | 0
persistent fever | 0
dyspnea | 0
chest pain | 0
diarrhea | 0
blood pressure 47/29 mm Hg | 0
tachycardia | 0
oxygen therapy | 0
hepatojugular reflux | 0
cardiogenic shock | 0
bilateral conjunctivitis | 0
cheilitis | 0
hypertension | -1008
fever episode | -1008
myalgia | -1008
dysgeusia | -1008
anosmia | -1008
coronavirus disease-2019 (COVID-19) | -1008
septic shock | 0
broad-spectrum antibiotics | 0
leukocytosis | 0
normocytic anemia | 0
elevated liver enzyme levels | 0
elevated creatine kinase levels | 0
acute kidney injury | 0
C-reactive protein (CRP) | 0
brain natriuretic peptide | 0
D-dimer | 0
troponin levels | 0
electrocardiogram | 0
sinus tachycardia | 0
transthoracic echocardiogram (TTE) | 0
global hypokinesis | 0
dilated inferior vena cava | 0
reduced ejection fraction | 0
acute myocarditis | 0
infectious work-up | 0
SARS-CoV-2 immunoglobulin G | 0
polymerase chain reaction (PCR) | 0
comprehensive etiological work-up | 0
coronary computed tomography (CT) scan | 336
multiple coronary aneurysms | 336
hemodynamic support | 0
norepinephrine infusion | 0
dobutamine infusion | 0
intravenous immunoglobulins (IVIG) | 120
prednisone | 120
aspirin | 120
resolution of all symptoms | 240
control TTE | 240
cardiac magnetic resonance imaging | 168
discharged | 288
partial regression of coronary aneurysms | 1440
complete disappearance of all aneurysms | 2160