38 years old | 0
woman | 0
abdominal discomfort | -24
nausea | -24
vomiting | -24
presented to the emergency room | 0
no fever | 0
no vaginal discharge | 0
initially evaluated in the Obstetric Emergency Department | 0
discharged home | 0
normal obstetric ultrasound | 0
returns to the ER | 144
persistent abdominal pain | 144
nausea (persistent) | 144
vomiting (persistent) | 144
tachycardic | 144
diffuse abdominal pain | 144
guarding on the right quadrants | 144
neutrophilia | 144
low prothrombinemia | 144
acute renal failure | 144
high procalcitonin | 144
high c-reactive protein | 144
abdominal ultrasound showed moderate fluid in all quadrants | 144
good foetal vitality | 144
worsening general condition | 144
surgical consultation obtained | 144
hypotension | 144
general abdominal guarding | 144
hyperlacticaemia | 144
hypokalaemia | 144
hyperglycaemia | 144
septic shock | 144
acknowledged | 144
emergency exploratory laparotomy | 144
generalised purulent peritonitis | 144
perforated acute appendicitis | 144
pus aspirated | 144
multiple interloop abscesses drained | 144
retrosplenic abscesses drained | 144
subfrenic abscesses drained | 144
pelvic abscesses drained | 144
retrouterine abscesses drained | 144
appendicectomy | 144
thorough abdominal washing | 144
generalised intraabdominal infection | 144
exuberant bowel distention | 144
possibility of abdominal compartment syndrome | 144
laparostomy performed | 144
admitted to the Intensive Care Unit | 144
septic shock (ICU admission) | 144
vasopressor therapy | 144
dialysis | 144
intravenous piperacillin-tazobactam antibiotherapy | 144
laparostomy revision | 192
marked bowel oedema | 192
distention (marked) | 192
mild intraabdominal soiling | 192
further peritoneal lavage | 192
new laparostomy with progressive closure technique | 192
recovered progressively | 192
taken to the Operating Room for surgical revision | 288
abdominal cavity primary closed | 288
no need of prosthesis | 288
antibiotherapy adjusted | 360
microbiological culture isolated Escherichia coli | 360
microbiological culture isolated Streptococcus orallis | 360
piperacillin-tazobactam suspended | 360
started amoxicillin with clavulanic acid | 360
remaining ICU stay uneventfully | 288
transferred to the obstetrics ward | 288
daily evaluated by obstetrics physicians | 288
good foetal viability observed | 288
discharged home | 336
kept obstetric follow-up | 336
remaining uncomplicated pregnancy | 336
admitted for an elective caesarean section | 984
gave birth to a healthy child | 984
ventral hernia needing correction | 984
thriving without neurological or other impairments | 984
