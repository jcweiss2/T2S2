3-day-old | 0
ex-full term male | 0
admitted to the emergency department | 0
multiple episodes of apnea | 0
born appropriate for gestational age | -72
birth weight 3065 g | -72
normal spontaneous vaginal delivery | -72
maternal polycystic ovarian syndrome | -672
metformin during the first trimester of pregnancy | -672
concerns for borderline gestational diabetes | -672
elevated glucose tolerance tests | -672
normal 3-h glucose test | -672
Group B Streptococcal infection | -672
adequate antibiotics provided before delivery | -672
difficulty with breastfeeding | -48
poor milk production | -48
supplemented with formula | -48
continued poor feeding | -24
apneic episodes | -24
ruddy in color | -24
going limp | -24
eyes rolling back | -24
vital signs were stable | 0
point-of-care glucose obtained | 0
undetectable glucose | 0
Dextrose 10% bolus | 0
D 10% infusion | 0
repeat glucose 18 mg/dL | 0
another D 10% bolus | 0
glucose infusion rate 13.85 mg/kg/min | 0
sepsis evaluation initiated | 0
urinalysis | 0
urine culture | 0
blood culture | 0
empiric treatment with ampicillin and gentamicin | 0
antibiotics discontinued | 48
chest X-ray normal | 0
COVID-19 negative | 0
screening complete blood count unremarkable | 0
comprehensive metabolic panel remarkable for hyperkalemia | 0
hypocalcemia | 0
transferred to the NICU | 0
glucose 44 mg/dL | 0
D 12.5% fluids continued | 0
weight at the 30th percentile | 0
length at the 25th percentile | 0
head circumference at the 55th percentile | 0
duplicated earlobes | 0
physical examination otherwise unremarkable | 0
glucose infusion rate weaned | 12
glucose stabilized | 12
Pediatric endocrinology consulted | 12
comprehensive evaluation for persistent hypoglycemia initiated | 12
serum glucose level 40 mg/dL | 12
normal ammonia level | 12
suppressed beta-hydroxybutyrate | 12
equivocal cortisol | 12
serum insulin level 6.0 µIU/mL | 12
Diazoxide initiated | 12
Chlorothiazide initiated | 12
Diazoxide increased | 48
Chlorothiazide dose increased | 96
pulmonary edema resolved | 96
repeat echocardiograms normal | 96
CH gene panel negative | 168
chromosome microarray revealed 1.46 Mb paternally inherited pathogenic duplication of chromosome 17q12 | 168
Diazoxide titrated down | 240
Chlorothiazide dose decreased | 240
discharged home | 240
serial cardiac examinations normal | 720
echocardiograms normal | 720
weaned off Diazoxide and Chlorothiazide | 720