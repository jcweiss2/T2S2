headache | -2160
blurred vision | -2160
kidney transplant | -5840
immunosuppression | -2160
methylprednisolone therapy | -2160
mycofenolate sodium | -2160
chronic kidney transplant disease | -2160
vascular rejection | -5840
chronic calcineurin-inhibitor toxicity | -5840
contrast-enhancing intracerebral lesions | -2160
perifocal edema | -2160
methylprednisolone stopped | -2159
dexamethasone administered | -2159
brain biopsy | -2158
cerebral PTLD diagnosed | -2158
diffuse large B-cell lymphoma | -2158
Epstein-Barr virus positive | -2158
chemotherapy | -2157
high-dose cytarabin | -2157
Rituximab | -2157
complete remission of PTLD | -2152
transplant function aggravated | -2152
eGFR 25.4 mL/min/1.73 m2 | -2152
cytomegalovirus reactivated | -2144
pneumocystis jirovecii pneumonia | -2144
chemotherapy changed | -2144
Rituximab dose increased | -2144
antiviral therapy | -2144
antibiotic therapy | -2144
mycofenolate sodium dose tapered | -2144
generalized seizure | -2128
cerebral MRI scan | -2128
recurrence of PTLD | -2128
HDMTX administered | 0
Leukovorine administered | 0
Rituximab administered | 0
vigorous hydration | 0
alkalinization of urine | 0
dialysis procedures started | 24
MTX-level measured | 24
dialysis session 1 | 24
dialysis session 2 | 36
dialysis session 3 | 48
dialysis session 4 | 72
nadir of leucocytes | 240
CMV- and E.coli pneumonia | 312
sepsis | 312
acute kidney transplant failure | 312
invasive ventilation | 312
sepsis managed | 312
cerebral MRI scan | 376
radiotherapy | 400
no response to radiotherapy | 400