68 years old | 0
male | 0
admitted to the hospital | 0
vomited | -96
consumed alcohol | -96
epigastralgia | -96
brought to the hospital by ambulance | -96
blood pressure 160/100 mm Hg | 0
pulse rate 105 beats/min | 0
respiratory rate 32 breaths/min | 0
body temperature 38.3°C | 0
SpO2 95% | 0
white blood cell count 5,900/μl | 0
red blood cell count 411 × 104/μl | 0
hemoglobin 12.3 g/dl | 0
neutrophils 81.7% | 0
platelets 9.7 × 104/μl | 0
total protein 6.1 g/dl | 0
albumin 2.4 g/dl | 0
blood urea nitrogen 34 mg/dl | 0
creatinine 1.2 mg/dl | 0
creatine phosphokinase 111 IU/l | 0
aspartate aminotransferase 28 IU/l | 0
alanine aminotransferase <10 IU/l | 0
total bilirubin 0.6 mg/dl | 0
Na 142 mEq/l | 0
Cl 108 mEq/l | 0
K 4.2 mEq/l | 0
C-reactive protein 40.2 mg/dl | 0
procalcitonin 12.5 ng/ml | 0
left pleural effusion | 0
cardiomegaly | 0
heart failure suspected | 0
chest X-ray | 0
diagnosed with spontaneous esophageal perforation | 48
chest tube drainage | 48
sepsis | 96
transferred to hospital | 96
emergent surgery | 96
perforated lesion covered with necrotic tissue | 96
food residue in left thoracic cavity | 96
pyothorax | 96
mediastinitis | 96
thoracic drainage | 96
nasoesophageal tube inserted | 96
transcervical mediastinal tube inserted | 96
feeding jejunostomy | 96
postoperative enteral nutrition | 96
blood laboratory data improved | 120
orally administered contrast medium seen as fistula | 1200
fistula diminished | 1392
lesion of esophageal perforation covered with regenerated epithelium | 1728
peroral intake started | 1824
discharged from hospital | 2064