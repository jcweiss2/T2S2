6 years old | 0
male | 0
admitted to the hospital | 0
fatigue | -120
looks pale | -120
fever | -120
abdominal pain | -120
shock | 0
altered consciousness | 0
Glasgow Coma Score 12 | 0
heart rate 135 beats per minute | 0
blood pressure 70/40 mmHg | 0
respiratory rate 40 breaths per minute | 0
temperature 36.5°C | 0
prolonged capillary refill time >2 s | 0
oxygen saturation 83% | 0
receiving oxygen 5 L/minutes via a simple mask | 0
no enlargement of the spleen and liver | 0
fluid resuscitation | 0
transfusion | 0
hemodynamic monitoring | 0
inotropic agent administration | 0
orotracheal intubation | 0
complete blood counts | 0
hemoglobin 2.9 g/dL | 0
hematocrit 9.3% | 0
leucocyte 18 × 10^3/μL | 0
basophil 0% | 0
eosinophil 0% | 0
neutrophil band 1% | 0
neutrophil segment 55% | 0
lymphocyte 33% | 0
monocyte 4% | 0
erythrocyte 1.13 × 10^12/L | 0
platelets counts 213 × 10^3/μL | 0
albumin 1.96 g/dL | 0
urea 46.2 g/dL | 0
serum creatinine 1.15 mg/dL | 0
aspartate transaminase 510 U/L | 0
alanine transaminase 173 U/L | 0
potassium 6 mmol/L | 0
sodium 123 mEq/L | 0
C-reactive protein 0.09 mg/dL | 0
procalcitonin 0.78 ng/mL | 0
blood gas analysis | 0
pH 6.8 | 0
pO2 24.2 mmHg | 0
pCO2 27.2 mmHg | 0
HCO3 4.8 mmol/L | 0
TCO2 5.6 mmol/L | 0
BE -2.78 mmol/L | 0
SO2 17.3% | 0
lactate dehydrogenase 10.6 mmol/L | 0
peripheral blood smear | 0
normochromic erythrocytes | 0
anisopoikilocytosis | 0
microcytic | 0
leukocytic hypersegmentation | 0
serum iron 157 mcg/dL | 0
Total Iron Binding Capacity 207 mcg/dL | 0
ferritin 3985 ng/mL | 0
SARS Cov-2 IgM reactive | 0
SARS Cov-2 IgG non-reactive | 0
Polymerase Chain Reaction SARS Cov-2 negative | 0
IgM anti-dengue reactive | 0
IgG anti-dengue non-reactive | 0
chest x-ray | 0
no abnormalities | 0
refractory septic shock | 0
aggressive fluid resuscitation | 0
broad-spectrum antibiotic | 0
inotropic agents | 0
multiple organ failure | 14
death | 14
coinfection with dengue | -120
no history of traveling | -120
no history of contact with COVID-19 patients | -120
no cough | -120
no breathing difficulties | -120
no bleeding | -120
no rashes | -120
active child | -48
symptoms abruptly worsened | -48
admitted to the pediatric emergency department | 0
discharged | - 
(Note: Since the patient died, there is no discharge event)