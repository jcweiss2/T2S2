23 years old | 0 | 0 
male | 0 | 0 
admitted to the hospital | 0 | 0 
history of methicillin-resistant Staphylococcus aureus (MRSA) impetigo | -8760 | -8760 
right tibia fracture | -8760 | -8760 
intramedullary fixation (IMN) | -8760 | -8760 
interlocking screws removed | -720 | -720 
skin irritation | -720 | -720 
pain | -720 | -720 
redness and swelling at the surgical site | -672 | -672 
stitch abscess | -672 | -672 
cultures from the surgical site were positive for MRSA | -672 | -672 
oral antibiotic treatment | -672 | -672 
discharged home | -672 | -672 
fever | -504 | -504 
right groin pain | -504 | -504 
discharged home with the diagnosis of viral infection | -504 | -504 
systemic fever | -336 | -336 
myalgia | -336 | -336 
difficult and painful ambulation | -336 | -336 
right forearm cellulitis | -336 | -336 
right sudden onset uveitis | -336 | -336 
systemic rash | -336 | -336 
right hip lymphadenopathy | -336 | -336 
increased CRP level | -336 | -336 
elevated WBC count | -336 | -336 
hepatic enzymes elevated | -336 | -336 
lactic dehydrogenase (LDH) elevated | -336 | -336 
creatine phosphokinase (CPK) elevated | -336 | -336 
radiograph of both hips in anterior-posterior view was unremarkable | -336 | -336 
treatment with intravenous (IV) antibiotics | -336 | -336 
medical condition continued to deteriorate | -336 | -168 
positron emission tomography-computed tomography (PET-CT) scan | -168 | -168 
OIM abscess with systemic manifestations | -168 | -168 
blood cultures were positive for MRSA bacteria | -168 | -168 
hemodynamic deterioration | -168 | -168 
fulminant MRSA sepsis | -168 | -168 
admitted to the intensive care unit (ICU) | -168 | -168 
ultrasound-guided drainage | -168 | -144 
full-body CT scan | -144 | -144 
abscesses diameter further enlarged | -144 | -144 
persistent fever | -144 | -144 
CRP level of 36 mg/dL | -144 | -144 
WBC count of 20,000 | -144 | -144 
surgical intervention | -144 | -144 
combined approach of Smith-Peterson and modified Stoppa | -144 | 0 
surgery | 0 | 0 
general anaesthesia with muscle relaxant | 0 | 0 
Stoppa approach | 0 | 0 
Smith-Peterson approach | 0 | 0 
drainage of the abscess | 0 | 0 
debridement of the OIM and adductor brevis muscle | 0 | 0 
lavage for the pelvic brim | 0 | 0 
improving general condition | 0 | 168 
less frequent fever spikes | 0 | 168 
decrease in CRP and WBC levels | 0 | 168 
additional antibiotic treatment support for 6 weeks | 0 | 504 
almost complete recovery | 504 | 504 
able to ambulate normally without any pain or functional limitations | 504 | 504 
returned to daily activities | 504 | 504