29 years old | 0
female | 0
admitted to the hospital | 0
sports-related injury | -2628
shoulder surgery | -2628
surgical revisions | -2628
Pseudomonas aeruginosa | -2628
Sphingomonas paucimobilis | -2628
Candida colliculosa | -2628
Staphylococcus aureus | -2628
shoulder infections | -2628
CRPS | -304
left shoulder tendon release | -304
revision | -304
asthma | 0
selective IgG3 deficiency | -730
electromyography | 0
brachial plexus injury | 0
oral medical management | 0
opioids | 0
antidepressants | 0
antispasmodics | 0
left stellate ganglion blockade | 0
continuous cervical epidural infusions | 0
placement of a left C6–C7 interlaminar epidural catheter | 0
fluoroscopic guidance | 0
preprocedure labs | 0
complete blood count | 0
complete metabolic panel | 0
creatinine phosphokinase | 0
antibiotic prophylaxis | 0
intravenous vancomycin | 0
epidural infusion | 0
0.25% bupivacaine | 0
hydromorphone | 0
clonidine | 0
oral home medications | 0
methadone | 0
hydromorphone | 0
diazepam | 0
baclofen | 0
amitriptyline | 0
decrease in pain | 24
improved sleep | 24
decrease in LUE spasms | 24
decrease in edema | 24
febrile | 120
increase in temperature | 120
wean the infusion | 120
remove the epidural catheter | 120
progressive headache | 126
neck pain | 126
increase in temperature | 126
neurological examination | 126
nontender to palpation | 126
blood and urine cultures | 126
chest x-ray | 126
increase in white count | 126
cephalosporin | 126
cefepime | 126
abatement of fever | 126
decrease in white count | 126
MRI | 130
cervical spine | 130
sagittal T1- and T2-weighted imaging | 130
sagittal inversion recovery | 130
axial fast spin echo | 130
gradient recall techniques | 130
epidural collection | 130
compression of the left C5 and C6 nerve roots | 130
effacement of the thecal sac | 130
interstitial edema | 130
left paraspinal muscles | 130
transfer to the neurosciences intensive care unit | 130
hourly neurological examination | 130
intractable nausea | 154
vomiting | 154
left arm weakness | 154
emergent decompression | 154
evacuation | 154
C3 to C7 cervical laminectomies | 154
C4–C5 and C5–C6 left foraminotomies | 154
intraoperative cultures | 154
P aeruginosa | 154
susceptible to cefepime | 154
resolution of arm weakness | 154
uneventful postoperative course | 154
discharged home | 216
intravenous cefepime | 216