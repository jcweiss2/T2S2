79 years old | 0
female | 0
hypertension | 0
severe aortic stenosis |==0
chronic heart failure | 0
elective transcatheter aortic valve replacement (TAVR) | 0
TAVR with 26 mm CoreValve™ | 0
general anesthesia | 0
temporary transvenous pacing (TVP) wires placed in the right ventricle (RV) | 0
fluoroscopic guidance | 0
left common femoral vein | 0
transferred to the Intensive Care Unit (ICU) | 0
extubated | 0
stable condition | 0
temporary pacemaker set as VVI | 0
rate of 50 beats/min | 0
threshold of 10 mA | 0
two-dimensional transthoracic echocardiography (TTE) | 24
POD 1 | 24
remove pacer wires | 24
became diaphoretic | 24.5
hypotensive (BP 40/25 mmHg) | 24.5
resuscitated with intravenous fluid boluses | 24.5
norepinephrine drip | 24.5
BP increased to 100/60 mmHg | 24.5
stat TTE | 24.5
moderate pericardial effusion around RV/right atrium | 24.5
excessive respiratory variation of the mitral inflow velocities | 24.5
mild RV collapse during diastole | 24.5
cardiac tamponade physiology | 24.5
emergency pericardiocentesis | 24.5
180 ml sanguineous fluid drained | 24.5
pericardial drain left in place | 24.5
RV rupture by temporary pacing wires | 24.5
POD 3 | 72
stable | 72
draining minimal fluid (15 ml in 24 h) | 72
repeat TTE | 72
no new pericardial effusion | 72
remove pericardial drain | 72
developed diaphoresis | 72.33
hemodynamically unstable | 72.33
emergent TTE | 72.33
reaccumulation of pericardial fluid | 72.33
pericardiocentesis | 72.33
200 ml frank blood drained | 72.33
coronary angiogram | 72.33
no obstruction | 72.33
aortic root aortogram | 72.33
no leakage or tear | 72.33
transesophageal echocardiography | 72.33
good valve function | 72.33
transferred back to ICU | 72.33
conservative management | 72.33
drain left in place for 72 h | 72.33
stable | 72.33
follow-up TTE | 72.33
computed tomography of the chest | 72.33
negative for fluid reaccumulation | 72.33
4th day after redrainage (POD 7) | 168
pericardial catheter clamped | 168
TTE 2 h postclamping | 168.08
no accumulation of pericardial fluid | 168.08
drain removed | 168.08
vital signs monitored continuously for 4 h | 168.08
after 24 h | 192
transferred from ICU to step-down | 192
