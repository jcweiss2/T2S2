29 years old | 0
male | 0
chest pain | 0
cough | 0
breathlessness | 0
breathlessness for 4 months | -2928
cough with white sputum for 2 months | -1440
loss of weight | -3624
loss of appetite | -3624
shooting pain in the right side of chest for 2 weeks | -336
blood pressure of 110/70 | 0
respiratory rate of 28/min | 0
oxygen saturation (SpO2) of 90% on room air | 0
chest X-ray revealed cardiomegaly | 0
pleural effusion with fissural extension | 0
underlying collapse on the right side | 0
fibrotic bands in right perihilar region | 0
total leucocyte count (TLC) count was 10,730 cells | 0
neutrophilic predominance | 0
pleural tap of 300 ml fluid | 0
exudative effusion | 0
intercostal drain (ICD) insertion | 0
diagnosis of lower respiratory tract infection | 0
treated with intravenous antibiotics (ceftriaxone/sulbactam and levofloxacin) | 0
nebulizations | 0
supportive measures | 0
pleural fluid analysis revealed sugars 75 mg/dl | 0
proteins <2 g/dl | 0
adenosine deaminase (ADA) 4.8 u/l | 0
pleural fluid cytology showed white blood cells of 950 cells | 0
predominantly lymphocytic (95%) | 0
reactive mesothelial cells | 0
two-dimensional Echo showed left atrial wall thickening | 0
infiltration or thrombus | 0
pulmonary vein obstruction | 0
good left ventricle function | 0
contrast-enhanced computed tomography (CT) chest showed homogeneous poorly enhancing soft tissue in subcarinal region indenting left atrium | 0
partial narrowing of right inferior pulmonary vein ostium extending along the interatrial groove | 0
encasing mass causing partial narrowing of the right main pulmonary artery | 0
encasing mass causing partial narrowing of azygous arch | 0
cervical mediastinoscopy | 0
biopsy of 4R lymph node station | 0
frozen section remained inconclusive | 0
patient's condition improved | 120
discharged at request on day 5 of admission | 120
advised to come back for VATS procedure | 120
underwent VATS and incisional biopsy after 10 days | 240
thoracotomy findings showed hard mass encasing heart and hilar structures infiltrating left atrium | 240
biopsy for histopathological examination | 240
biopsy for immunohistochemistry | 240
patient was extubated | 240
received noninvasive ventilation | 240
received oxygen (O2) support postoperatively | 240
patient developed tachypnea on postoperative day 4 | 240
shifted back to surgical intensive care unit | 240
procalcitonin levels raised (1.69 ng/ml) | 240
D-dimer levels within normal limits | 240
arterial blood gas showed partial pressure 54.5 | 240
SpO2 of 90% on bilevel positive airway pressure with O2 support of 10 L | 240
respiratory distress | 240
O2 desaturation | 240
intubated and connected to ventilator support on postoperative day 5 | 240
ET culture and sensitivity | 240
Gram stain | 240
fungal stain | 240
acid-fast bacilli stain | 240
Gram-negative coverage continued | 240
X-ray postintubation showed left lower lobe pneumonia | 240
basal crept bilaterally | 240
blood culture was negative | 240
endotracheal secretion culture grown pseudo hyphae | 240
hyaline septate with acute branching hyphae | 240
started on voriconazole 200mg BID therapy | 240
HPE report revealed epithelioid granulomas | 240
multinucleated giant cells | 240
areas of necrotising inflammation | 240
scattered acute branching fungal hyphae | 240
fungal hyphae amidst the inflammation | 240
fungal hyphae within the giant cells | 240
Periodic-acid-Schiff (PAS) staining | 240
Grocotts-methenamine-silver (GMS) staining | 240
septate, elongated, slender forms of fungal organisms morphologically resembling aspergillus | 240
diagnosis of acute respiratory distress syndrome | 240
diagnosis of invasive aspergillosis | 240
treated with low tidal volume strategy | 240
patient's condition worsened | 264
developed septic shock | 264
refractory hypoxemia | 264
serum creatinine increased to 3.1 mg/dl | 264
acute kidney injury | 264
started on renal replacement therapy | 264
hyperkalemia | 264
acidosis | 264
family refused further treatment | 264
left against medical advice | 264
expired on day 8 after suffering a cardiac arrest | 312
