37 years old | 0
    Afro-Caribbean | 0
    woman | 0
    admitted | 0
    three-week history of lethargy | -504
    three-week history of myalgia | -504
    three-week history of intermittent chest pain | -504
    uncomplicated pregnancy | -672
    acute kidney injury | 0
    severe hypercalcaemia | 0
    proteinuria | 0
    intravenous fluids | 0
    empirical antimicrobials | 0
    presumed sepsis | 0
    deteriorate | 24
    transferred to ICU | 24
    respiratory support | 24
    renal replacement therapy | 24
    differential diagnosis including vasculitis | 0
    differential diagnosis including autoimmune disease | 0
    differential diagnosis including sepsis | 0
    differential diagnosis including malignancy | 0
    relevant tests requested | 0
    leukocytosis | 0
    left shift | 0
    no abnormal cells | 0
    autoimmune screen negative | 0
    respiratory virus panel negative | 0
    human immunodeficiency virus negative | 0
    hepatitis B antibodies negative | 0
    hepatitis C antibodies negative | 0
    PTH level suppressed | 0
    recurrent episodes of narrow-complex tachycardia | 96
    recurrent episodes of broad-complex tachycardia | 96
    echocardiogram revealed poor global systolic function | 96
    no pericardial effusion | 96
    no obvious valvular abnormality | 96
    corrected serum calcium 3.3 mmol/L | 96
    DC cardioversion | 96
    antiarrhythmics | 96
    marked sensitivity to amiodarone | 96
    marked sensitivity to lignocaine | 96
    marked sensitivity to adrenaline | 96
    bradycardia | 96
    ventricular tachycardia | 96
    fatal brady-tachy arrhythmia | 96
    prolonged cardiac arrest | 96
    resuscitation unsuccessful | 96
    intracellular calcium deposition in cardiac myocytes | 96
    widespread calcification in medium-sized arteries | 96
    widespread calcification in small-sized arteries | 96
    intra-renal arteries micro-infarcts | 96
    infiltration of lymph nodes | 96
    infiltration of bone marrow | 96
    infiltration of lung | 96
    infiltration of liver | 96
    large lymphoid blasts | 96
    histiocytic haemophagocytosis | 96
    lymphoid blasts CD3 positive | 96
    lymphoid blasts CD25 positive | 96
    parathyroid glands normal | 96
    HTLV-1 antibodies positive | 96
    adult T-cell leukaemia-lymphoma | 96
    no malignant cells in peripheral blood film | 0
    
    
<|eot_id|>
