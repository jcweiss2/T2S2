48 years old | 0
    female | 0
    end-stage renal disease | -52560
    hypertensive | -61392
    maintenance hemodialysis twice a week | -4392
    hypertension well controlled with one antihypertensive agent | 0
    fasting blood sugar within normal limits | -72
    postprandial blood sugar within normal limits | -72
    glycated hemoglobin levels within normal limits | -72
    preoperative hemodialysis within 24 hours of scheduled surgery | -24
    standard monitoring applied | 0
    balanced general anesthesia administered | 0
    heart rate 94/min | 0
    mean arterial pressure 103 mmHg | 0
    SpO2 100% | 0
    central venous pressure 12 cm H2O | 0
    core temperature 98.6°F | 0
    arterial blood gas analysis after induction of anesthesia (10 AM) | 0
    lactate 1.9 mM/L | 0
    volume controlled ventilation adjusted | 0
    EtCO2 maintained between 35 mm and 40 mm Hg | 0
    hemodynamic parameters deteriorated three hours after induction | 3
    heart rate 122/min | 3
    mean arterial pressure 72 mmHg | 3
    central venous pressure 16 cm H2O | 3
    arterial blood gas analysis showed metabolic acidosis | 3
    elevated lactate levels | 3
    hyperglycemia | 3
    elevated anion gap | 3
    fall in hemoglobin | 3
    blood sample for ketone bodies tested negative | 3
    occult blood loss considered | 3
    IV fluids administered | 3
    two units of packed red blood cells transfused | 3
    noradrenaline infusion started | 3
    MAP maintained at 90 mmHg | 3
    sodium bicarbonate infusion started | 3
    insulin infusion started | 3
    allograft reperfused | 3
    urine output established 25 minutes after reperfusion | 3
    shifted to ICU 7 hours after induction | 7
    noradrenaline infusion (0.12 μg/kg/min) | 7
    elective ventilation | 7
    possible need for continuous renal replacement therapy | 7
    ABG analysis in ICU revealed progressively increasing lactic acidosis | 7
    hyperglycemia refractory to bicarbonate and insulin infusion | 7
    average urine output of 300 mL/h | 7
    possibility of sepsis considered | 7
    procalcitonin levels 14.6 ng/mL | 7
    empirical thiamine 300 mg administered intravenously 3 hours after surgery | 10
    ABG analysis 2 hours after thiamine administration | 12
    rapidly decreasing lactate levels | 12
    rapidly decreasing sugar levels | 12
    improvement in MAP | 12
    bicarbonate infusion stopped | 12
    insulin infusion stopped | 12
    noradrenaline infusion stopped | 12
    extubated 7 hours after completion of surgery |. 19
    thiamine injection 300 mg IV repeated | 19
    ABG analysis 8 hours after first dose of thiamine injection within normal limits | 20
    shifted to posttransplant isolation ward 12 hours after surgery | 12
    afebrile | 7
    normal total leukocyte counts | 7
    no significant hypotension when lactic acidosis was discovered | 7
    postoperative pro-calcitonin level high | 7
    T-cell antibody anti-thymocyte globulin received intraoperatively | 0
    surgical stress | 0
    accelerated glycolysis | 0
    enhanced pyruvate production | 0
    increased thiamine requirement | 0
    occult thiamine deficiency | 0
    defective thiamine activity | 0
    severe lactic acidosis with hyperglycemia | 0
    no proven adverse effects from excess thiamine dose | 19
    