65 years old|0
female|0
end-stage osteoarthritis of the right knee|0
progressively worsening joint pain|0
refractory to all non-operative measures|0
well-controlled hypertension|0
gastroesophageal reflux disease|0
remote history of DVT|0
right total knee arthroplasty|0
perioperative course uncomplicated|0
post-operative course uncomplicated|0
discharged home|48
enoxaparin|24
DVT prophylaxis|24
admitted|192
vague epigastric pain|192
lethargy|192
febrile episodes|192
decreased appetite|192
somnolence|192
anxiety|192
nausea|192
no vomiting|192
temperature 101.7 F|192
heart rate 111|192
respiration 20|192
blood pressure 123/87|192
oxygen saturation 92%|192
hyponatremia (126)|192
hypokalemia (2.6)|192
glucose (60)|192
hematocrit (25.3)|192
creatinine (0.8)|192
WBC count (14,900)|192
platelet count (161,000)|192
chest CT scan negative for pulmonary embolism|192
MRI of the brain negative for acute pathology|192
presumed sepsis|192
intravenous antibiotics|192
ceftriaxone|192
vancomycin|192
acyclovir|192
cultures obtained|192
deteriorated rapidly|192
transferred to intensive care unit|192
aggressive intravenous volume support|192
pressors|192
adrenal insufficiency|192
basal cortisol levels obtained|192
cosyntropin stimulation|192
cortisol levels 0.3 nmol/L|192
abdominal CT revealed bilateral adrenal hemorrhages|192
enoxaparin discontinued|192
high dose hydrocortisone|192
improved dramatically|216
left intensive care unit|216
glucocorticoid tapered|216
discharged without further complications|216
excellent range of motion|10560
X-rays demonstrate well-placed components|10560
no evidence of loosening|10560
returned to previous activity level|10560
bowling|10560
BAH|192
enoxaparin-induced BAH|192
adrenal hemorrhage|192
bilateral adrenal hemorrhage|192
acute adrenal insufficiency|192
hypotension|192
shock|192
no pulmonary embolism|192
no acute brain pathology|192
negative HIT antibody test|192
glucocorticoid administration|192
corticosteroid therapy|216
no long-term steroid therapy|10560
heparin-induced thrombocytopenia|192
chemoprophylaxis-related complications|192
bleeding risks|192
wound complications|192
adrenal insufficiency confirmed|192
cosyntropin stimulation test|192
glucocorticoid replacement therapy|216
improved clinically|216
returned to activity|10560
mechanical DVT prophylaxis|0
pharmacological DVT prophylaxis|0
anticoagulation prophylaxis|0
chemoprophylaxis|0
enoxaparin regimen|24
DVT prophylaxis regimen|24
post-operative enoxaparin|24
POD two discharge|48
enoxaparin started on POD one|24
discharged home with enoxaparin|48
POD eight admission|192
symptoms started on POD eight|192
metabolic encephalopathy|192
sepsis differential|192
adrenal insufficiency differential|192
CSF cultures|192
urine cultures|192
blood cultures|192
volume support|192
pressors administration|192
cosyntropin test|192
cortisol levels post stimulation|192
bilateral adrenal hemorrhages confirmed|192
enoxaparin cessation|192
hydrocortisone initiation|192
rapid improvement|216
ICU transfer|192
ICU discharge|216
glucocorticoid taper|216
post-discharge follow-up|10560
one-year visit|10560
activity resumption|10560
no complications|216
clinical suspicion for BAH|192
CT imaging|192
adrenal gland enlargement|192
hemorrhage confirmation|192
steroid treatment|216
diagnostic challenges|192
non-specific symptoms|192
early intervention|192
high clinical suspicion|192
steroid administration|216
no recurrence|10560
no loosening|10560
successful outcome|10560
