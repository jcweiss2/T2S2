71 years old | 0
female | 0
admitted to the hospital | 0
type 1 diabetes | -672
end-stage renal disease | -672
complete atrioventricular block | -672
previous myocardial infarction | -672
permanent pacemaker | -672
hemodialysis | -672
self-inflicted bite wound | -24
swelling of the left hand | -24
heat of the left hand | -24
redness of the left hand | -24
cellulitis | -24
intravenous cefazolin | -24
bacterial culture | -24
MRSA | -24
Kanavel’s cardinal signs of flexor tenosynovitis | -24
vancomycin infusion | -24
wound debridement | -24
partial amputation | -24
decompression of the median nerve | -24
purulent abscess | -24
abdominal pain | 120
gastrointestinal bleed | 120
systemic shock | 120
vasopressors | 120
elevated WBC count | 120
increased CRP | 120
increased creatinine | 120
reduced sodium | 120
reduced blood glucose | 120
reduced hemoglobin | 120
non-occlusive mesenteric ischemia | 120
small bowel resection | 120
norepinephrine | 120
COVID-19 exposure | 168
SARS-CoV-2 infection | 168
nasal swab test | 168
acute pneumonia | 192
chest radiograph | 192
CT scan | 192
consolidation of the lungs | 192
bilateral pleural effusions | 192
favipiravir | 192
intensive care unit | 192
hemodiafiltration | 192
necrotizing fasciitis | 216
septic shock | 216
mechanical respiration | 216
remdesivir | 216
hydrocortisone | 216
osteomyelitis | 240
vancomycin | 240
ARDS | 264
DIC | 264
ART-123 | 264
amputation of the distal forearm | 336
debridement | 336
lavage | 336
removal of infected tissue | 336
replacement of hemodialysis shunt | 336
septic shock | 744
cardiopulmonary arrest | 744