60 years old | 0
male | 0
Caucasian | 0
merchant ship captain | 0
presented to the emergency department | 0
headache | -24
dizziness | -24
disorientation | -24
ingestion of isopropanol | -24
ingestion of ethanol | -24
consumed ethanol | -24
consumed isopropanol | -24
brought empty bottle of rubbing alcohol | -24
label 70% volume per volume isopropyl alcohol | -24
capacity 473 mL | -24
patient consumed most of the liquid | -24
colleague consumed small amount | -24
no recent or past history of substance abuse | -24
disoriented | 0
clinical examination unremarkable | 0
unenhanced CT scan of the brain | 0
unenhanced CT scan unremarkable | 0
admitted for further investigations and management | 0
symptomatic treatment started | 0
collapsed in the hospital | 0.5
deeply comatose | 0.5
Glasgow Coma Scale score 3/15 | 0.5
developed hypotension | 0.5
blood pressure 80/40 mmHg | 0.5
pulse rate 65 per minute | 0.5
respiratory rate 8 per minute | 0.5
generalized hypotonia | 0.5
absent tendon reflexes | 0.5
no evidence of head trauma | 0.5
no evidence of cervical spine trauma | 0.5
administration of intravenous fluids | 0.5
endotracheal intubation | 0.5
admitted to intensive care department | 0.5
leukocytosis 26,000 white blood cells per μL | 0.5
hemoglobin 15.7 g/dL | 0.5
mean corpuscular volume 93 fl | 0.5
arterial blood gas pH 6.731 | 0.5
arterial blood gas pCO2 28.2 mmHg | 0.5
arterial blood gas pO2 141 mmHg | 0.5
arterial blood gas bicarbonate 3.5 mmol/L | 0.5
arterial blood gas oxygen saturation 95% | 0.5
blood urea nitrogen 9.5 mmol/L | 0.5
serum creatinine 157 μmol/L | 0.5
Na+ 141 mmol/L | 0.5
K+ 6 mmol/L | 0.5
Cl− 107 mmol/L | 0.5
HCO3 5 mmol/L | 0.5
capillary blood glucose 7.2 mmol/L | 0.5
severe metabolic acidosis | 0.5
acute renal failure | 0.5
blood lactic acid level 8.7 mmol/mL | 0.5
blood ketones negative | 0.5
blood ethanol negative | 0.5
blood isopropanol levels not obtained | 0.5
blood methanol levels not obtained | 0.5
blood ethylene glycol levels not obtained | 0.5
blood propylene glycol levels not obtained | 0.5
blood diethylene glycol levels not obtained | 0.5
liver enzymes normal | 0.5
serum amylase normal | 0.5
lipase levels normal | 0.5
increasing renal impairment | 2
hyperglycemia | 2
electrolyte imbalance | 2
low bicarbonate levels | 2
hyperkalemia | 2
follow-up arterial blood gas severe acidosis | 2
no growth on urine culture | 2
no growth on blood culture | 2
no crystals in urine | 2
serum pseudocholinesterase level 7,438 U/L | 2
calculated serum osmolarity 310 mOsmol/L | 2
received hemodialysis | 2
gradual improvement in blood pH | 2
gradual improvement in lactic acid levels | 2
treated with norepinephrine | 2
treated with intravenous fluids | 2
no improvement in blood pressure | 2
received 500 mL fractionated plasma protein stat | 2
received 2,000 mL normal saline | 2
kept on 200 mL/hour normal saline | 2
no response to intravenous fluids | 2
started on norepinephrine 10 μg per minute | 2
norepinephrine increased to 90 μg per minute | 2
blood pressure stabilized | 6
weaned off norepinephrine | 96
unenhanced MRI scans of the brain | 144
unenhanced MRI scans of the spine | 144
bilateral symmetrical hyperintensities on T2-weighted | 144
bilateral symmetrical hyperintensities on T1-weighted | 144
bilateral symmetrical hyperintensities on T2*-weighted | 144
bilateral symmetrical hyperintensities on FLAIR | 144
bilateral symmetrical hyperintensities on diffusion-weighted images | 144
cerebral cortex hyperintensities | 144
cerebellar cortex hyperintensities | 144
white matter hyperintensities | 144
basal ganglia hyperintensities | 144
thalami hyperintensities | 144
brainstem hyperintensities | 144
swollen and edematous cervical spinal cord | 144
T2-weighted hyperintensities in cervical spinal cord | 144
FLAIR hyperintensities in cervical spinal cord | 144
cerebellar tonsillar herniation 17 mm | 144
compression of proximal cervical cord | 144
petechial hemorrhages in brainstem | 144
petechial hemorrhages in gangliocapsular regions | 144
toxic brain damage | 144
toxic cervical spinal cord damage | 144
expired | 240
