61 years old | 0
male | 0
admitted to the hospital | 0
massive hemoptysis | 0
respiratory distress | 0
persistent cough | -2160
expectoration | -2160
COVID-19 pneumonia | -2160
tested positive for COVID-19 | -2160
streaky hemoptysis | -168
resolved spontaneously | -168
intravenous methylprednisolone | -2160
remdesivir | -2160
tocilizumab | -2160
prophylactic subcutaneous enoxaparin | -2160
high flow nasal oxygen | -2160
CRP mildly elevated | 0
D-dimer mildly elevated | 0
diabetic | 0
medication for diabetes | 0
HRCT of chest | -336
bilateral fibrotic sequelae of COVID pneumonia | -336
cavitary areas of breakdown in right lung | -336
tested negative for COVID-19 | 0
shifted to Respiratory intensive treatment unit | 0
low oxygen saturation | 0
Tranexamic acid | 0
Bilevel Positive Airway Pressure | 0
transfused with packed red blood cells | 0
CT Pulmonary Angiogram | 0
PAP in right lower lobe | 0
cavitating area in right lower lobe consolidation | 0
multiple ground glass alveolar infiltrates | 0
alveolar haemorrhage | 0
background fibro-reticular changes | 0
architectural distortion | 0
fibrotic sequelae of COVID-19 pneumonia | 0
endovascular embolization procedure | 0
pulmonary pseudoaneurysm | 0
Interventional Radiology Cath-lab suite | 0
right common femoral vein access | 0
ultrasound guidance | 0
6 French sheath | 0
right main pulmonary artery cannulated | 0
contrast pulmonary angiogram | 0
selective contrast angiograms | 0
bi-lobulated large PAP | 0
pseudoaneurysm embolised | 0
multiple coils deployed | 0
total embolization of aneurysm | 0
complete stasis of culprit branch | 0
optimal post-procedure angiographic result | 0
no further episodes of hemoptysis | 336
oxygen saturation improved | 336
superimposed fungal infection ruled out | 336
co-infection with mycobacterium tuberculosis ruled out | 336
interval contrast enhanced follow-up CT | 336
successful embolization of pseudoaneurysm | 336
discharged | 336