48 years old | 0
man | 0
medical history of smoking | 0
significant bowel resection 2 years previously | 0
presented to the emergency department | 0
intense headache | -48
abdominal pain | -48
dyspnoea | -168
generalized oedema | -168
asthenia | -168
decrease in urinary output | -168
no fever | 0
no neurological symptoms | 0
no respiratory symptoms | 0
no digestive symptoms | 0
no genitourinary symptoms | 0
worked as a hairdresser | 0
denied allergies | 0
denied exposure to new substances | 0
denied drugs | 0
denied ticks | 0
denied animals | 0
denied recent travels | 0
extensive small and large bowel partial resection 2 years previously | -17520
post-surgical short bowel syndrome | -17520
colostomy | -17520
non-specific abdominal pain | -17520
hypotension | -17520
elevated plasma lactate levels | -17520
elevated haematocrit | -17520
haemoconcentration | -17520
metabolic acidosis | -17520
normal plasma creatine phosphokinase levels | -17520
abdominal CT arteriography | -17520
exclusion of arterial occlusion | -17520
exclusion of venous thrombosis | -17520
intensive haemodynamic support | -17520
monitoring | -17520
emergent abdominal exploration | -17520
bowel resection | -17520
exclusion of cardiovascular disease | -17520
exclusion of sepsis | -17520
exclusion of drugs | -17520
non-occlusive mesenteric ischaemia | -17520
two more surgeries for partial bowel resection | -17520
post-surgery care | -17520
catheter-related superior vena cava thrombosis | -17520
implantation of a vascular access system | -17520
parenteral nutrition | -17520
3 months of hypocoagulation | -17520
three previous hospitalizations for oliguric acute renal injury | -26280
first episode 3 years previously | -26280
hypovolaemic shock | -26280
metabolic acidaemia | -26280
ICU admission | -26280
ionotropic support | -26280
renal replacement treatment | -26280
broad spectrum empiric antibiotics | -26280
unknown primary cause | -26280
2-day prodrome of intense headache | -26280
diffuse abdominal discomfort | -26280
physical exercise | -26280
heat exposure | -26280
haemodynamically unstable | 0
hypotension (85/45 mmHg) | 0
heart rate of 120 bpm | 0
no respiratory failure | 0
generalized oedema | 0
no skin flushing | 0
no urticaria | 0
no focal angioedema | 0
no stridor | 0
no lymphadenopathy | 0
normal abdominal evaluation | 0
normal neurological evaluation | 0
normal cardiac evaluation | 0
normal pulmonary evaluation | 0
severe metabolic acidaemia | 0
pH 7.27 | 0
HCO3 10.6 | 0
haemoconcentration | 0
Hgb 22.4 g/dl | 0
haematocrit 61% | 0
20.08 K/μl leucocytes | 0
uraemia (90 mg/dl) | 0
elevated creatinine (2.20 mg/dl) | 0
hypoalbuminaemia (2.0 g/dl) | 0
normal creatine phosphokinase | 0
normal coagulation | 0
normal liver function | 0
elevated BNP (222.5 pg/ml) | 0
normal troponin level | 0
normal electrocardiogram | 0
normal thoracic x-ray | 0
normal urinary study | 0
normal contrast-enhanced thoracoabdominal CT scan | 0
normal abdominal ultrasound | 0
normal renal ultrasound | 0
intensive fluid replacement therapy | 0
admitted to Internal Medicine Department | 0
haemodynamic stabilization | 0
renal function recovery | 0
normal inflammatory studies | 0
normal ESR | 0
normal CRP | 0
negative infectious study | 0
negative serologies | 0
negative blood cultures | 0
negative urinary cultures | 0
diagnosis of ISCLS | 0
prodromes of intense headache | 0
prodromes of abdominal pain | 0
association with heat exposure | 0
differential diagnosis sepsis | 0
differential diagnosis anaphylaxis | 0
differential diagnosis drug reactions | 0
exclusion of distributive shock | 0
exclusion of cardiogenic shock | 0
exclusion of hypovolaemic shock | 0
exclusion of obstructive shock | 0
normal thyroid function | 0
normal gonadal function | 0
normal adrenal steroid function | 0
normal immune function tests | 0
normal metabolic function tests | 0
normal complement studies | 0
normal C3 | 0
normal C4 | 0
normal CH50 | 0
normal C1 esterase inhibitor levels | 0
normal C1 esterase inhibitor function | 0
exclusion of hereditary angioedema | 0
normal cardiac study | 0
normal transthoracic echocardiography | 0
normal cardiovascular MRI | 0
normal whole endoscopic study | 0
exclusion of neuroendocrine tumours | 0
monoclonal gamma/lambda gammopathy | 0
IgG1 | 0
lambda light chains | 0
normal bone marrow biopsy | 0
IVIG administration (1 g/kg) | 0
clinical improvement | 0
nutritional supplementation | 0
discharged | 720
episodes of oedema | 720
fatigue | 720
partial leaks | 720
prophylactic treatment with terbutaline | 720
prophylactic treatment with theophylline | 720
periodic plasma level evaluations | 720
avoided physical exercise | 720
avoided heat exposure | 720
two more hospital admissions | 720
acute exacerbation | 720
subtherapeutic theophylline levels | 720
prophylactic IVIG (1 g/kg/month) | 720
maintained for 1 year | 720
good results | 720
