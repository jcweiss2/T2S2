21 years old | 0
male | 0
admitted to the hospital | 0
high-velocity motorcycle accident | -168
comminuted pelvic fractures | -168
multiple extremity fractures | -168
catastrophic degloving injury | -168
vascular injuries | -168
angioembolization of bilateral iliac arteries | -168
necrotizing soft tissue infection | -168
Acinetobacter spp. | -168
Pseudomonas spp. | -168
Stenotrophomonas maltophila | -168
Trichosporon asahii | -168
Saksenaea spp. | -168
Fusarium spp. | -168
aggressive surgical debridement | -168
antimicrobial therapy | -168
ceftazidime | -168
metronidazole | -168
trimethoprim-sulfamethoxazole | -168
micafungin | -168
amphotericin B | -168
posaconazole | -168
VERAFLO vac instillation | -168
multisystem organ failure | -168
shock | -168
lymphopenia | -168
neutrophilia | -168
IL-7 therapy | 59
informed consent | 59
test dose of IL-7 | 59
increased dosage of IL-7 | 60
improvement in clinical status | 63
decreased infectious spread | 63
decreased fungal proliferation | 63
improved wound healing | 63
healthier-appearing tissue margins | 63
improvement in fever curve | 63
improvement in tachycardia | 63
improvement in tachypnea | 63
increased absolute lymphocyte count | 63
decreased white blood cell count | 63
negative tissue cultures | 70
negative histology | 70
development of healthy granulation tissue | 70
skin grafting | 70
negative blood cultures | 70
negative wound cultures | 70
negative bone cultures | 70
exposed pelvic bone | 100
persistent perineal wound | 100
urethra disruption | 100
urine drainage | 100
isavuconazonium treatment | 100
biopsy of exposed pelvic bone | 100
biopsy of open wound margin | 100
Trichosporon asahii | 100
ELISpot assay | 59
increased T-cell function | 59
increased IFN-γ production | 59
increased lymphocyte adhesion molecules | 59
increased lymphocyte trafficking | 59
immunohistochemical staining | 59
increased CD3+ T cells | 59
mass cytometry | 59
increased pSTAT5 | 59
increased T-cell differentiation | 59
discharge from hospital | 120