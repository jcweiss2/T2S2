15 years old | 0
male | 0
admitted to the hospital | 0
vomiting | -48
lethargy | -48
left thigh swelling | -336
left femur shaft fracture | -336
orthopedic surgery | -324
discharged from the hospital | -312
poor oral intake | -48
elevated body temperature | -48
bilious vomiting | -24
lethargic | -24
decreased urine output | -24
dark urine | -24
dehydration | -24
gastrointestinal symptoms | 0
cerebral palsy | -6720
HSAN-IV | -6720
pain insensitivity | -6720
anhidrosis | -6720
recurrent orthopedic diseases | -6720
femur fractures | -6720
septic arthritis | -6720
osteomyelitis | -6720
mutilated fingertips | -6720
recurrent cellulitis | -6720
septic arthritis of fingers | -6720
impulse control disorder | -6720
unstable body temperature | -6720
autonomic dysregulation | -6720
unstable blood pressures | -6720
severe dry skin | -6720
hyperkeratosis | -6720
fissuring | -6720
xerotic eczema | -6720
wheelchair-bound | -6720
mentally retarded | -6720
hypokalemia | -6720
hypomagnesemia | -6720
Gitelman syndrome | -6720
anti-psychotics | -6720
psychostimulants | -6720
spironolactone | -6720
cachectic | 0
hip spica cast | 0
short stature | 0
low body weight | 0
blood pressure 130/88 mmHg | 0
pulse rate 97 beats/minute | 0
respiratory rate 21 times/minute | 0
body temperature 37.3°C | 0
anemic conjunctiva | 0
icteric sclera | 0
dehydrated lips and mucous membranes | 0
intact tympanic membranes | 0
non-palpable cervical lymph nodes | 0
symmetric chest wall expansion | 0
clear breath sounds | 0
regular heartbeat | 0
soft and flat abdomen | 0
no tenderness or rebound tenderness | 0
hyperactive bowel sounds | 0
no shifting dullness | 0
non-palpable liver or spleen | 0
no peripheral edema | 0
no digital clubbing | 0
no cyanosis | 0
mutilated fingertips | 0
dry skin | 0
no rash | 0
no petechia | 0
sodium 138 mmol/L | 0
potassium 3.2 mmol/L | 0
AST 23 IU/L | 0
ALT 12 IU/L | 0
total bilirubin 1.0 mg/dL | 0
BUN 29 mg/dL | 0
creatinine 0.41 mg/dL | 0
CRP <0.03 mg/dL | 0
serum magnesium 1.6 mg/dL | 0
supportive treatment | 0
high fever | 72
temperature 41.8°C | 72
no response to antipyretic drugs | 72
low blood pressure 50/17 mmHg | 72
seizure-like movements | 72
upward eyeball deviation | 72
loss of consciousness | 72
generalized clonic movement | 72
fixed pupils | 72
WBC count 19.4×10^3/µL | 72
hemoglobin level 9.6 g/dL | 72
platelet count 90×10^3/µL | 72
sodium level 137 mmol/L | 72
potassium level 2.6 mmol/L | 72
AST level 454 IU/L | 72
ALT level 258 IU/L | 72
total bilirubin level 4.3 mg/dL | 72
direct bilirubin level 2.6 mg/dL | 72
amylase level 228 IU/L | 72
lipase level 888 IU/L | 72
creatinine phosphate kinase level 1,258 IU/L | 72
lactate dehydrogenase level 985 IU/L | 72
BUN level 49 mg/dL | 72
creatinine level 1.62 mg/dL | 72
CRP level 0.6 mg/dL | 72
acute liver failure | 72
acute pancreatitis | 72
disseminated intravascular coagulation | 72
rhabdomyolysis | 72
acute kidney injury | 72
anemia | 72
plasma hemoglobin level 27.5 mg/dL | 72
serum ferritin level 250 ng/mL | 72
weakly positive antinuclear antibody | 72
repeated blood testing | 72
AST 492 IU/L | 72
ALT 545 IU/L | 72
total bilirubin 10.8 mg/dL | 72
direct bilirubin 5.1 mg/dL | 72
amylase 520 IU/L | 72
lipase 5,071 IU/L | 72
PT INR 3.1 | 72
aPTT 52.7 seconds | 72
fibrinogen 160 mg/dL | 72
D-dimer 17.62 µg/mL | 72
alkaline phosphatase 126 IU/L | 72
γ-glutamyltranspeptidase 98 IU/L | 72
aggressive management | 72
fluid resuscitation | 72
intravenous inotropes | 72
antibiotics | 72
gabexatemesilate | 72
transfer to PICU | 72
ventilator care | 72
seizure-like movements | 96
lorazepam | 96
mannitol | 96
abdominal computed tomography | 96
multiple filling defects in both kidneys | 96
brain magnetic resonance imaging | 96
hypoxic ischemic encephalopathy | 96
low serum ceruloplasmin level | 120
excessive urine copper level | 120
liver biopsy | 120
centrilobular confluent necrosis | 120
marked copper deposition | 120
hepatic copper dry weight 74 µg/g | 120
ophthalmologic examination | 120
Kayser–Fleischer rings | 120
gene studies | 120
NTRK1 gene sequencing | 120
c.2002G>T, p.Asp668Tyr heterozygote | 120
c.360-1G>A, (IVS3) heterozygote | 120
compound heterozygote mutation | 120
SLC12A3 gene sequencing | 120
heterozygote c.1216A>C | 120
ATP7B gene sequencing | 120
negative results | 120
trientine treatment | 168
low copper diet | 168
clinical improvement | 168
WBC count 8.66×10^3/µL | 360
hemoglobin level 12.9 g/dL | 360
platelet count 364×10^3/µL | 360
sodium level 137 mmol/L | 360
potassium level 4.0 mmol/L | 360
AST level 128 IU/L | 360
ALT level 127 IU/L | 360
total bilirubin level 1.3 mg/dL | 360
BUN level 25 mg/dL | 360
creatinine level 0.1 mg/dL | 360
PT INR 1.15 | 360
aPTT 52.3 seconds | 360
tracheostomy | 432
percutaneous endoscopic gastrostomy | 432
home ventilator care | 432
gastrostomy feeding | 432
trientine treatment | 432
copper restriction diet | 432