74 years old | 0
male | 0
hospitalized for wide excision of squamous cell carcinoma on the left mandible | 0
received neoadjuvant chemotherapy twice | -720
underwent marginal mandibulectomy | 0
underwent left supraomohyoid neck dissection | 0
underwent reconstruction with reconstruction plate | 0
underwent reconstruction with right radial forearm free flap | 0
general anesthesia | 0
no medical morbidities including hypertension or diabetes | 0
preoperative laboratory findings normal | 0
preoperative chest radiograph normal | 0
ECG finding of sinus arrhythmia | 0
ECG finding of low voltage in frontal leads | 0
ECG finding of ST elevation | 0
TTE normal | 0
hemodynamically stable throughout the perioperative time | 0
transported to ICU | 0
NTT remained in airway | 0
ventilation assisted with Ambu bagging | 0
oxygen 7 L/min | 0
SpO2 100% | 0
vital signs taken | 0
elevated BP | 0
elevated HR | 0
complained of pain | 0
analgesics administered | 0
opioids administered | 0
BP remained high (259/115 mmHg) | 0
HR surged (168 beats/min) | 0
complained of persistent pain | 0
complained of agitating | 0
dexmedetomidine administered | 0
respiratory rate dropped to 7 breaths/min | 0
SpO2 dropped to 89% | 0
BP dropped due to sedatives | 0
ST elevation in ECG monitor | 0
serial ECGs checked | 0
ST elevation in anterior and lateral leads | 0
elevated cardiac markers | 0
myoglobin surged to 1275.8 ng/ml | 0
Troponin I rose to 6.32 ng/ml | 0
serum creatine kinase MB peaked at 55.6 ng/ml | 0
referred to cardiology department | 0
TTE performed | 0
dilated left ventricular | 0
normal LV wall thickness | 0
akinesia of apical lateral | 0
akinesia of inferior wall | 0
akinesia of mid-cavity | 0
severe systolic dysfunction | 0
LV ventriculogram showed EF of 25% | 0
ischemic insult of multivessel territory | 0
stress-induced cardiomyopathy suspected | 0
transferred to medical ICU | 0
managed conservatively with inotropics | 0
managed conservatively with chronotropics | 0
managed conservatively with diuretics | 0
hemodynamic monitoring | 0
dopamine 5 µg/kg/min administered | 0
dobutamine 5 µg/kg/min administered | 0
norepinephrine 0.1 µg/kg/min administered | 0
rapid clinical improvement | 0
ST-segment elevations normalized by third postoperative day | 72
extubated on fifth postoperative day | 120
transferred to general ward in dental hospital | 120
Troponin I levels normalized | 72
all laboratory test values within normal ranges | 72
TTE showed no evidence of cardiac ischemia | 720
TTE showed left ventricular EF of 63% | 720
no clinical signs of heart failure | 720
received consolidation radiotherapy (total dose: 5040 cGy) | 720
oral cavity lesions healing well | 720
complete dentures being prepared | 720
patient in good condition | 720
Takotsubo cardiomyopathy diagnosis | 0
transient hypokinesis | 0
akinesis | 0
dyskinesis of left ventricular mid-segments | 0
hyperkinetic base | 0
akinetic apex | 0
absence of obstructive coronary artery disease | 0
absence of acute plaque rupture | 0
new electrocardiographic abnormalities | 0
absence of pheochromocytoma | 0
absence of myocarditis | 0
clinical symptoms of TTC | 0
angina | 0
dyspnea | 0
ischemic changes on ECG | 0
patent coronary arteries | 0
no abnormal findings in periodic follow-up | 720
surgery-induced stress | 0
medication-induced stress | 0
BP and HR elevation in ICU | 0
surgical site pain | 0
discomfort from NTT | 0
hypertension | 0
tachycardia | 0
transfer between hospitals | 0
cold temperature exposure | 0
lengthy surgery (14 hours) | 0
general anesthesia stress | 0
patient's advanced age (74 years) | 0
male gender | 0
physical stress trigger | 0
ST elevation | 0
T wave inversion | 0
modest elevation in cardiac troponin | 0
reversible heart failure | 0
transient form of heart failure | 0
emotional stress association | 0
physiologic stress association | 0
extended operation time | 0
early recognition of TTC | 0
proper postoperative care | 0
complete recovery | 720
