16 years old| 0
    male | 0
    admitted to the hospital | 0
    fatigue | 0
    epistaxis | 0
    dyspnea | 0
    white cell count of 1900 per cubic millimeter | -720
    absolute neutrophil count 90 per cubic millimeter | -720
    hemoglobin 5.3 g per deciliter | -720
    platelets 36 000 per cubic millimeter | -720
    hospitalized | -672
    bone marrow biopsy | -360
    aplastic anemia | -360
    discharged | -720
    packed red blood cells | -720
    pooled platelet transfusions | -720
    intravenous antibiotics | -720
    admitted to the US National Institute of Health Clinical Center | 0
    fever | -168
    dysphagia | -168
    odynophagia | -168
    cough | -168
    scant hemoptysis | -168
    body temperature 38.2oC | 0
    blood pressure 126/91 mm Hg | 0
    heart rate 88 beats per minute | 0
    respiratory rate 18 breaths per minute | 0
    oxygen saturation 98% | 0
    thin | 0
    lethargic | 0
    spitting blood@-@tinged saliva | 0
    denied dyspnea | 0
    phonating normally | 0
    tender diffusely around the neck | 0
    white cell count of 1430 per cubic millimeter | 0
    absolute neutrophil count 0 per cubic millimeter | 0
    hemoglobin 10.7 g per deciliter | 0
    platelets 33 000 per cubic millimeter | 0
    radiographic imaging showed classic "thumbprint" sign | 0
    direct laryngoscopy showed erythematous, enlarged, posteriorly ptotic epiglottis | 0
    intravenous piperacillin/tazobactam | 0
    vancomycin | 0
    micafungin | 0
    intravenous dexamethasone | 0
    nebulized racemic epinephrine | 0
    clinically improved | 0
    no need for definitive airway management by intubation | 0
    blood cultures showed no growth | 0
    endoscopically directed cultures isolated Enterobacter cloacae | 0
    resistant to cefazolin | 0
    cefoxitin | 0
    ceftazidime | 0
    ceftriaxone | 0
    co@-@amoxiclav | 0
    ampicillin | 0
    aztreonam | 0
    piperacillin/tazobactam | 0
    prescribed meropenem | 0
    clinically improved | 0
    follow@-@up laryngoscopy 17 days later showed significant improvement | 408
    