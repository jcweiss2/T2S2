86 years old | 0
    female | 0
    presented to the Emergency Department (ED) in acute respiratory distress | 0
    discharged from the inpatient unit | -24
    hospitalized for a complicated urinary tract infection | -672
    hypothyroid disorder | -105120
    mild dementia from traumatic brain injury | -105120
    complained of substernal chest pain | 0
    complained of shortness of breath | 0
    blood pressure of 105/74 mm Hg | 0
    heart rate 132 | 0
    respiratory rate 26 | 0
    oral temperature of 36.7 °C | 0
    oxygen saturation of 88% on room air | 0
    rapid heart rate | 0
    bilateral crackles on auscultation of the lungs | 0
    12-lead electrocardiogram (EKG) showed sinus tachycardia | 0
    ST-segment depressions in the precordial leads V2 to V5 | 0
    arterial blood gas significant for hypoxemia | 0
    arterial blood gas significant for mild metabolic acidosis | 0
    chest radiography demonstrated moderate pulmonary edema | 0
    chest radiography demonstrated small pleural effusions bilaterally | 0
    white blood cell count of 26.89 × 10∗3/μL | 0
    initial troponin I of 0.38 ng/mL | 0
    subsequent rise to 64.50 ng/mL | 0
    treatment instituted for flash pulmonary edema | 0
    treatment instituted for non-ST segment elevation myocardial infarction | 0
    placed on non-invasive ventilation | 0
    initiated on aspirin | 0
    initiated on clopidogrel | 0
    initiated on atorvastatin | 0
    initiated on antibiotics | 0
    initiated on furosemide | 0
    initiated on nitroglycerin | 0
    initiated on heparin | 0
    admitted to the intensive care unit | 0
    underwent transthoracic echocardiography | 24
    transthoracic echocardiography showed moderate mitral valve regurgitation | 24
    transthoracic echocardiography showed stenosis | 24
    subsequent left heart catheterization | 48
    left heart catheterization revealed a large saddle embolism involving two vessels of non-dominant circumflex coronary artery | 48
    left heart catheterization revealed no associated stenosis | 48
    intensive medical management recommended per cardiology consultation | 48
    respiratory status continued to deteriorate | 72
    not a candidate for invasive mechanical ventilation | 72
    previously expressed do-not-resuscitate instructions | -105120
    previously expressed do-not-intubate instructions | -105120
    sustained cardiopulmonary arrest | 96
    death | 96
    
    <|eot_id|>
  