75 years old | 0
    woman | 0
    visited emergency room | 0
    dyspnea | -168
    idiopathic thrombocytopenic purpura | -672
    corticosteroids | -672
    prednisolone | -672
    tapered 10 mg/day | -672
    blood pressure 156/122 mmHg | 0
    heart rate 180 beats/min | 0
    respiratory rate 44 breaths/min | 0
    oxygen saturation 56% | 0
    body temperature 37.7°C | 0
    increased high-sensitivity C-reactive protein | 0
    white blood cell count 15.340/μL | 0
    neutrophils 89.0% | 0
    negative influenza antigen | 0
    negative respiratory virus test | 0
    negative bacterial PCR | 0
    P. jirovecii PCR test | 0
    aspergillosis antigen test | 0
    chest radiography | 0
    diffuse ground-glass opacities | 0
    infiltration in both lungs | 0
    chest computed tomography | 0
    diffuse geographic consolidations | 0
    ground-glass opacities in both lungs | 0
    two cavitary lesions in both lower lungs | 0
    admitted to intensive care unit | 0
    empirical treatment for community-acquired pneumonia | 0
    intravenous piperacillin/tazobactam | 0
    azithromycin | 0
    possible PCP infection | 0
    sulfamethoxazole/trimethoprim | 0
    methylprednisolone | 0
    endotracheal intubation | 72
    mechanical ventilator support | 72
    antibiotics switched to meropenem | 72
    levofloxacin | 72
    hospital day 7 | 168
    fraction of inspiration O2 reduced to 45% | 168
    clinical improvement | 168
    initial serology positive | 168
    PCP PCR positive | 168
    aspergillus antigen test positive | 168
    itraconazole initiated | 168
    follow-up chest CT | 168
    newly formed ground-glass opacities | 168
    cavitary changes in right middle lobe | 168
    hospital day 9 | 216
    bronchoscopy | 216
    bronchoalveolar lavage | 216
    aspergillus antigen tests performed | 216
    hospital day 11 | 264
    aspergillosis reported in BAL fluid cytology | 264
    IA diagnosed | 264
    antifungal agent changed to voriconazole | 264
    hospital day 13 | 312
    percutaneous dilatational tracheostomy | 312
    bronchoscopy with BAL | 312
    BAL fluid cytology (second) | 312
    aspergillosis again | 312
    condition deteriorated | 312
    family declined aggressive management | 312
    hospital day 15 | 360
    PCP PCR positive in BAL fluid | 360
    fungus culture no growth | 360
    hospital day 16 | 384
    died | 384
    multi-organ failure | 384
    septic shock | 384
    