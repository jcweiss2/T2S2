84 years old | 0
    male | 0
    presented to the hospital | 0
    progressively worsening lethargy | -96
    worsening fatigue | -96
    weakness | -96
    bloody urine | -24
    denied nausea | 0
    denied vomiting | 0
    denied abdominal pain | 0
    intermittent fevers | 0
    ischemic cardiomyopathy | 0
    heart failure | 0
    atrial fibrillation | 0
    Coumadin | 0
    hepatosplenomegaly | 0
    petechial rash | 0
    elevated total bilirubin (2.8 mg/dL) | 0
    elevated alkaline phosphatase (159) | 0
    elevated AST (42) | 0
    elevated ALT (51) | 0
    INR 4.7 | 0
    albumin 3.2 | 0
    white blood count 5.1 | 0
    hemoglobin 11.3 g/dL | 0
    platelet count 109,000 | 0
    ascites | 0
    CBD diameter 0.5 cm | 0
    fresh frozen plasma | 0
    vitamin K | 0
    INR remained >3 | 0
    intermittent fevers (up to 103.2°F) | 0
    negative blood cultures | 0
    bilirubin increased to 15.1 g/dL | 120
    direct bilirubin 11.5 g/dL | 120
    paracentesis | 120
    ascites albumin 1.2 g/dL | 120
    serum albumin 2.4 g/dL | 120
    ascites neutrophil count 91 | 120
    low haptoglobin | 120
    worsening encephalopathy | 120
    continued fevers | 120
    piperacillin-tazobactam | 120
    hypotension | 120
    transferred to ICU | 120
    peripheral smear obtained | 120
    intravenous clindamycin | 120
    quinine | 120
    bilirubin increased to 24 g/dL | 120
    negative Lyme serology | 120
    negative Ehrlichia serology | 120
    negative Anaplasmosis serology | 120
    passed away | 120
    acute liver failure | 120
    fulminant liver failure | 120
    Babesiosis diagnosis | 120
    <|eot_id|>
    