47 years old | 0
female | 0
Caucasian | 0
cigarette smoking | -3120
alcohol consumption | -8760
untreated chronic psoriasis vulgaris | -8760
unconscious | -2
found on the floor | -2
interhospital transfer | -2
admitted to OMFS department | 0
normal temperature | 0
tachypnea | 0
tachycardia | 0
hypotension | 0
tumefaction in the right area of her face and neck | 0
bilateral palpebral microabscesses | 0
large occipital psoriatic plaque | 0
massive crepitations in the occipital and posterior cervical regions | 0
emergency surgery | 1
wide posterior cervical incision | 1
right submandibular incision | 1
extensive necrosis | 1
necrectomy | 1
sterile dressing | 1
oxygenated water and povidone-iodine solution | 1
postoperative contrast-enhanced computed tomography scan | 2
empirical antibiotic therapy | 2
vancomycin | 2
imipenem | 2
metronidazole | 2
limited right lateral cervical and supraclavicular necrectomy | 72
excision of the platysma muscle | 72
partial excision of the lateral cervical skin flap | 72
total necrectomy of the splenius capitis muscles | 72
partial necrectomy of the semispinalis capitis muscles | 72
leukocytosis | 72
fever | 72
bacteriological wound drainage | 96
drug sensitivity testing | 96
Staphylococcus epidermidis | 96
Klebsiella sp. | 96
Acinetobacter sp. | 96
colistin | 96
necrectomy of the entire epicranial galea | 168
necrectomy of the right temporal fascia | 168
edema of the entire face | 168
clean wounds with granulation tissue | 1080
plastic reconstruction | 1080
multiple reconstructions with flaps | 1080
free skin grafts | 1080
discharged | 1824