48 years old | 0
female | 0
admitted to the hospital | 0
cardiopulmonary resuscitation | -48
loss of consciousness | -48
pale face | -48
salivation at the corners of the mouth | -48
urinary incontinence | -48
no nausea | -48
no vomiting | -48
no limb twitching | -48
high blood pressure | -48
low heart rate | -48
third-degree atrioventricular block | -48
low serum potassium | -48
diarrhea | -72
temporary pacemaker implanted | -48
chest CT scan | -48
exudative lesions in the lungs | -48
head CT scan | -48
no abnormality in head CT scan | -48
transferred to ICU | -24
stable vital signs | -24
fever | 0
high blood pressure | 0
heart rate | 0
respiratory rate | 0
trachea intubation | 0
mechanical ventilation | 0
appendectomy incision | 0
temporary cardiac pacing catheter | 0
left femoral vein catheterization | 0
high white blood count | 0
high procalcitonin | 0
high pro-B type natriuretic peptide | 0
high hypersensitive troponin T | 0
high ALT | 0
high AST | 0
cardiac respiratory arrest | 0
post-CPR syndrome | 0
third-degree atrioventricular block | 0
broad empirical therapy with imipenem and vancomycin | 0
temperature rose | 72
inflammation indexes elevated | 72
left femoral vein catheter removed | 72
catheter blood and venous blood cultures sent | 72
gram-negative rods detected | 86
colistin applied | 86
strains isolated from blood, chocolate, and MacConkey Agar | 96
initial identification of Myroides spp. | 96
definitive identification of Myroides odoratimimus | 96
catheter-related bloodstream infection diagnosed | 96
septic shock | 96
antimicrobial susceptibility tests | 96
resistant to most agents | 96
susceptible to cefoperazone/sulbactam | 96
treatment changed to cefoperazone/sulbactam and levofloxacin | 96
infection under control | 120
no causative organism detected in blood culture | 120
cardiac respiratory arrest again | 120
temporary pacemaker reinstalled | 120
coronary angiography | 120
coronary myocardial bridge | 120
permanent cardiac pacemaker considered | 120
transferred to local hospital for rehabilitation | 120