68 years old | 0
female | 0
admitted to the hospital | 0
dyspnea | -72
wheezing | -72
productive cough | -72
albuterol | -72
corticosteroid regimen | -672
gained 30 pounds | -672
COPD exacerbations | -720
treated with antibiotics | -720
treated with inhaled bronchodilators | -720
treated with systemic corticosteroids | -720
last hospitalization | -5760
no previous history of intubation | 0
no previous history of stridor | 0
no previous history of reflux symptoms | 0
mMRC symptom score 3 | 0
150 pack-year smoking history | -26280
quit smoking | -720
sleeps in a seated position | 0
dyspnea occurs when lies flat | 0
chairbound | 0
hypertension | 0
depression | 0
obstructive sleep apnea | 0
end-stage renal disease | 0
hemodialysis | 0
fluticasone/salmeterol | 0
tiotropium | 0
albuterol | 0
prednisone | 0
3 L oxygen by nasal cannula | 0
CPAP at night | 0
simvastatin | 0
diltiazem SR | 0
sertraline | 0
pulmonary rehabilitation program | -17520
temperature 98.6 F | 0
blood pressure 150/72 | 0
pulse rate 90/min | 0
respiratory rate 26/min | 0
body mass index 36 kg/m2 | 0
oxygen saturation 96% | 0
Cushingoid facies | 0
centripetal obesity | 0
rapid regular rhythm | 0
no murmur | 0
bilateral expiratory wheezing | 0
no pedal edema | 0
chest radiograph showed no infiltrates or congestion | 0
ECG showed sinus tachycardia | 0
non-specific ST changes | 0
hemoglobin 11 g/dL | 0
glucose 147 mg/dL | 0
potassium 4.7 mEq/L | 0
creatinine 9.1 mg/dL | 0
exacerbation of COPD | 0
intravenous glucocorticoids | 0
albuterol nebulizer treatments | 0
bi-level positive airway pressure | 0
broad-spectrum antibiotics | 0
hemodialysis | 0
oxygenation improved | 24
symptoms improved | 24
PFT showed FEV1/ FVC ratio of 62% | 24
FEV1 of 41% predicted | 24
GOLD 3 | 24
transthoracic echocardiogram | 24
left ventricular ejection fraction of 70% | 24
normal right ventricular function | 24
Grade 1 diastolic dysfunction | 24
normal valves | 24
workup for thrombophilia | 24
negative | 24
CT soft tissue neck | 24
unremarkable | 24
non-contrast dynamic expiratory chest CT | 24
diffuse pulmonary emphysema | 24
11 mm right upper lobe pulmonary nodule | 24
greater than 50% collapse in the distal trachea/multiple central bronchi | 24
complete collapse of the bronchus intermedius | 24
tracheobronchomalacia | 24
declined lung biopsy | 24
silicone stent placement | 24
bronchoscopy | 24
dynamic Y Boston scientific tracheobronchial stent | 24
went home | 48
stable condition | 48
arterial blood gases | 48
pH 7.35 | 48
pCO2 47 | 48
PO2 85 | 48
inhaler technique good | 48
found hypotensive | 72
found unresponsive | 72
acute hypoxic respiratory failure | 72
admitted to ICU | 72
endotracheal intubation | 72
intravenous vasopressors | 72
systemic corticosteroids | 72
broad-spectrum antibiotics | 72
nebulized bronchodilator treatment | 72
mucolytic agents | 72
chest radiograph showed no infiltrates or edema or pneumothorax | 72
normal position of the tracheobronchial stent | 72
sepsis ruled out | 72
myocardial ischemia ruled out | 72
COPD exacerbation improved | 96
wanted to be placed on home hospice | 96
discharged | 96