58 years old | 0
    woman | 0
    admitted to the intensive care unit | 0
    fever | -240
    fatigue | -240
    generalized body aches | -240
    diarrhea | -72
    chest tightness | -72
    shortness of breath | -72
    visited two local hospitals | -240 to -72
    leukopenia | -240 to -72
    thrombocytopenia | -240 to -72
    antibiotics (cephalosporin) | -240 to -72
    antipyretics | -240 to -72
    symptoms not relieved | -240 to -72
    farmer | -240
    engaged in agriculture | -240
    no history of tick bite | -672
    temperature 36.5 ℃ | 0
    heart rate 117/min | 0
    respiratory rate 45/min | 0
    blood pressure 170/100 mmHg | 0
    conscious state | 0
    crackles in both lungs | 0
    scattered skin petechiae | 0
    swollen lymph node | 0
    leukopenia (WBC 3.1 ×109/L) | 0
    thrombocytopenia (platelets 24 ×109/L) | 0
    elevated liver enzymes | 0
    elevated muscle enzymes | 0
    elevated aspartate aminotransferase | 0
    elevated alanine aminotransferase | 0
    elevated creatine kinase | 0
    elevated lactic dehydrogenase | 0
    slightly elevated procalcitonin | 0
    slightly elevated C-reactive protein | 0
    positive urine occult blood | 0
    positive urine protein | 0
    chest CT multiple patchy infiltrations | 0
    chest CT ground-glass opacities | 0
    bronchoscopy edema of airway mucosa | 0
    bronchoscopy white mold | 0
    arterial blood gas PH 7.233 | 0
    arterial blood gas PaO2 91.8 mmHg | 0
    arterial blood gas PaCO2 55.6 mmHg | 0
    arterial blood gas SaO2 95.8% | 0
    preliminary diagnosis pulmonary infection | 0
    preliminary diagnosis sepsis | 0
    empiric antibiotic treatment | 0
    biapenem | 0
    voriconazole | 0
    blood culture | 0
    BALF culture | 0
    mNGS | 0
    mental confusion | 24
    PaCO2 increased 79.4 mmHg | 24
    endotracheal intubation | 24
    mechanical ventilation | 24
    serological tests negative | 24
    serum galactomannan positive | 24
    serum 1,3-β-d-glucan positive | 24
    mNGS Aspergillus fumigatus | 24
    mNGS Aspergillus flavus | 24
    mNGS Aspergillus terreus | 24
    mNGS SFTSV | 24
    confirmed SFTS | 24
    confirmed invasive pulmonary aspergillosis | 24
    no pathogens isolated from culture | 24
    oral ribavirin | 24
    plasma transfusion | 24
    persistent thrombocytopenia | 24
    platelet transfusion | 24
    acute renal failure | 48
    heart failure | 48
    CRRT | 48
    metaraminol therapy | 48
    fever 37.8 ℃ | 168
    increased WBC count 10.44 ×109/L | 168
    increased procalcitonin 2.66 ng/ml | 168
    chest X-ray multiple patchy infiltrations | 168
    Acinetobacter baumannii isolated | 168
    tigecycline | 168
    pulmonary function improved | 168 to 312
    radiological findings improved | 312
    thrombocytopenia (platelets 40 ×109/L) | 408
    anemia (RBC 2.41 ×1012/L) | 408
    elevated creatine kinase 1534 IU/L | 408
    prolonged APTT 63.2 s | 408
    bronchoscopy uncontrolled white mold | 408
    mNGS Aspergillus fumigatus (DNA) | 432
    SFTSV not detected | 432
    discharged | 432
    died | 456
    
    
    <|eot_id|>