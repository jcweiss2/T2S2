57 years old | 0
male | 0
admitted to the hospital | 0
unconscious | 0
alcohol abuse | -672
alcohol dementia | -672
arterial hypertension | -672
fully conscious | -24
increasingly confused | -12
unresponsive | -6
Glasgow coma scale 3/15 | 0
cyanotic | 0
hypothermic | 0
temperature 34.7°C | 0
Kussmaul breathing | 0
breathing frequency 28 breaths per min | 0
blood pressure 150/90 mmHg | 0
heart rate 75-150 beats per min | 0
atrial fibrillation | 0
ECG frequency 92 beats per min | 0
rigid limbs | 0
pupils with absent light reflex | 0
computed tomography of the cerebrum | 0
chest X-ray | 0
hyperkalemia | 0
high anion gap | 0
elevated lactic acid | 0
high anion gap metabolic acidosis | 0
pH 7.07 | 0
HCO3− 6.4 mmol/L | 0
bladder catheterization | 0
clear urine | 0
urine drug screening positive for benzodiazepines | 0
intubated | 0
transmitted to the Intensive Care Unit (ICU) | 0
treatment with bicarbonate | 0
electrolyte correction | 0
intravenous ethyl alcohol infusion | 0
treatment with intravenous antibiotics | 0
increasing creatinine values | 6
decreasing urine production | 6
hyperkalemia | 6
worsening of acidosis | 6
pH 6.90 | 6
increased anion gap | 6
hemodialysis | 6
hypotension | 6
increased heart rate | 6
treated according to local guidelines | 6
new urine sample sent for examination | 6
multiple COM crystals | 6
supporting the diagnosis of ethylene glycol poisoning | 6
extubated | 48
hemodialysis discontinued | 48
ethyl alcohol infusion discontinued | 48
regained acceptable urine production | 48
furosemide stimulation | 48
normalized creatinine | 48
normalized calcium | 48
acidosis corrected | 48
lactate decreasing | 48
transferred from the ICU to the medical ward | 48
discharged to home | 72
ethylene glycol poisoning | -24
previous hospitalization with similar picture | -672
previous intake of antifreeze coolant | -672
previous diagnosis of ethylene glycol poisoning | -672
previous confirmation of ethylene glycol poisoning | -672