44 years old | 0
female | 0
postpartum | -840
vaginal delivery | -840
endometritis | -720
treated with cephalexin | -720
treated with metronidazole | -720
hypertension | 0
asthma | 0
admitted to the hospital | 0
severe chest pain | 0
chest pain radiating to back | 0
tachycardic | 0
hemodynamically stable | 0
blood pressure 142/57 mm Hg | 0
heart rate 99 beats per minute | 0
respiration rate 16 breaths per minute | 0
oxygen saturation 100% | 0
first and second heart sounds appreciated | 0
no aortic regurgitation murmur | 0
complete blood count normal | 0
kidney function normal | 0
electrolytes normal | 0
D-dimer negative | 0
high-sensitivity troponin levels elevated | 0
electrocardiogram showed sinus tachycardia | 0
no ST-segment changes | 0
chest radiograph unremarkable | 0
computed tomography of the chest | 0
splenic aneurysm | 0
splenic infarct | 0
pulmonary edema | 0
dilated pulmonary arteries | 0
no acute aortic dissection | 0
transthoracic echocardiogram | 0
masses on the tricuspid aortic valve | 0
severe aortic regurgitation | 0
mildly dilated left ventricle | 0
moderate eccentric hypertrophy | 0
dilated atria | 0
elevated atrial pressure | 0
moderate mitral regurgitation | 0
mild pulmonary hypertension | 0
coronary angiography | 0
luminal filling defect in the distal left main lesion | 0
no other angiographic coronary artery disease | 0
surgical thrombectomy | 12
aortic valve replacement | 12
vegetation removed | 12
aortic valve replaced with mechanical prosthesis | 12
transferred to intensive care unit | 12
sent to the ward | 120
repeat angiography | 120
culture results negative | 120
antibiotics continued | 120
discharged home | 360
intravenous vancomycin | 360
ceftriaxone | 360
follow-up with cardiac surgery | 720
follow-up with infectious diseases | 720
echocardiogram | 1008