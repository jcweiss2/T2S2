38 years old | 0
male | 0
non-smoker | 0
teetotaler | 0
diagnosed with PSC | -1096
without inflammatory bowel disease | -1096
colonoscopy-directed mucosal biopsy | -1096
ursodeoxycholic acid | -1096
developed three episodes of BC | -432
last episode requiring intensive care unit admission | -432
septic shock | -432
mucosal irregularities in the right and left hepatic duct | -432
areas of beading in segments 3, 6 and 8 of the liver | -432
no dominant strictures | -432
normal immunoglobulin type G4 serum level | -432
normal carbohydrate antigen 19-9 level | -432
no cholangiocarcinoma | -432
listed for LT | -216
persistent pruritus | -72
jaundice | -72
fourth episode of BC | -72
Escherichia coli bacteremia | -144
sensitive to cephalosporins | -144
Enterococcus fecalis | -72
sensitive to linezolid | -72
FMT | 0
informed consent | 0
nephew as donor | 0
standard screening protocol | 0
stool sample collection | 0
homogenization | 0
endoscopic FMT | 0
weekly for 4 weeks | 0
withheld antibiotics | 0
continued UDCA | 0
blood biochemistries | 0
stool microbial community analyses | 0
afebrile | 24
anicteric | 48
pruritus worsened | 24
pruritus decreased | 72
improvements in liver functions | 168
circulating total and toxic bile acids | 168
modification of bacterial communities | 168
relative abundance of Proteobacteria decreased | 168
relative abundance of Bacteroidetes increased | 168
relative abundance of Firmicutes increased | 168
Bifidobacterium increased | 168
Coprococcus increased | 168
Megamonas increased | 168
Bacteroides increased | 168
Enterobacter decreased | 168
Catenibacterium decreased | 168
Dialister decreased | 168
Fecalibacterium decreased | 168
Oscillopsira decreased | 168
Lachnospira decreased | 168
cholangitis recurred | 876
broad spectrum antibiotics | 876
pathogenic changes in gut microbial communities | 876
emergence of pathogenic species | 876
second cycle of FMT declined | 876
referred to LT center | 876