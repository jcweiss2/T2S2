8 years old | 0
    male | 0
    admitted to the hospital | 0
    severe abdominal pain | -24
    ALL (L3) diagnosis | -35040
    bone marrow transplant | -26280
    second relapse | -26280
    last chemotherapy | -504
    high dose methotrexate | -504
    no vaccination against chickenpox | 0
    normal body temperature | 0
    hepatosplenomegaly | 0
    periumbilical tenderness | 0
    hemoglobin 12.1 g/dL | 0
    WBC 3,490/mm3 | 0
    segmented neutrophils 80.0% | 0
    platelet 135,000/mm3 | 0
    increased AST 78 U/L | 0
    increased ALT 135 U/L | 0
    normal chest x-ray | 0
    normal abdomen x-ray | 0
    normal abdomen and pelvis CT | 0
    fever up to 39.0℃ | 24
    empirical IV antibiotics started | 24
    persistent abdominal pain | 24
    multiple erythematous vesicles on trunk | 72
    acyclovir 1,500 mg/m2/day started | 72
    vesicles spread across whole body | 120
    dyspnea | 120
    chest x-ray showing numerous small nodules | 120
    varicella pneumonia diagnosis | 120
    WBC 5,090/mm3 | 120
    platelet 32,000/mm3 | 120
    AST 931 U/L | 120
    ALT 788 U/L | 120
    LDH 3,196 U/L | 120
    DIC profile positive | 120
    IV acyclovir continued | 120
    IV antibiotics changed | 120
    IVIG 500 mg/kg/day added | 120
    single donor platelets | 120
    fresh frozen plasma | 120
    antithrombin III | 120
    transfer to ICU | 120
    drowsy mental state | 144
    aggravated dyspnea | 144
    chest x-ray total haziness | 144
    ARDS diagnosis | 144
    intubation | 144
    mechanical respiratory support | 144
    IVIG increased to 1 g/kg/day | 144
    chest x-ray marked improvement | 168
    cardiomegaly | 168
    platelet 69,000/mm3 | 168
    AST 224 U/L | 168
    ALT 280 U/L | 168
    recovery from DIC | 168
    IVIG total four days | 168
    persistent fever | 168
    unchanged vesicular skin lesions | 168
    normal cardiac function on echocardiography | 168
    increased BP up to 150/125 mm/Hg | 216
    IV labetarol started | 216
    no effect from labetarol | 216
    VZV detected in serum | 216
    IVIG extended two more days | 216
    generalized tonic-clonic seizure | 264
    hypertensive crisis suspected | 264
    VZV CNS involvement suspected | 264
    IV nitroprusside added | 264
    CSF tapping | 264
    normal CSF results | 264
    VZV antibody negative in CSF | 264
    VZV PCR negative in CSF | 264
    antihypertensives increased | 264
    IV phenytoin added | 264
    no further seizures | 264
    pulmonary condition stable | 312
    ventilator removed | 312
    no fever | 312
    skin lesions scarring stage | 312
    transfer to general ward | 408
    vital signs stable | 408
    improved laboratory data | 408
    lymphocyte subset CD3 87.0% | 408
    CD4 14.8% | 408
    CD8 70.6% | 408
    CD19 9.6% | 408
    CD56 3.0% | 408
    cellular immunity not recovered | 408
    brain MRI performed | 408
    EEG performed | 408
    brain MRI showing VZV-induced encephalitis | 408
    normal EEG | 408
    phenytoin stopped | 408
    IV antibiotics ceased | 456
    acyclovir ceased | 456
    no symptoms | 456
    discharged | 456
    chemotherapy resumed | 720
    follow-up brain MRI three months later | 2160
    VZV-induced encephalitis lesions disappeared | 2160
