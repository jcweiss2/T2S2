74 years old | 0
male | 0
hypertension | 0
diabetes mellitus | 0
presented to emergency department | 0
intermittent subjective fever | -96
rigors | -96
generalized headache | -96
altered mentation | -96
body malaise | -96
nausea | -96
vomiting | -96
no history of loss of consciousness | 0
no abdominal pain | 0
no change in stool habits | 0
no change in urine color | 0
denied recent trauma | 0
denied falls | 0
resides in malaria-endemic region | 0
previous uncomplicated malarial infections | 0
oral anti-malarials | 0
febrile (38.7 °C) | 0
tachypneic | 0
disoriented | 0
good nutritional status | 0
not jaundiced | 0
not cyanosed | 0
pulse rate of 103 beats/min | 0
sinus rhythm | 0
respiratory rate of 23 breaths/min | 0
blood pressure 96/60 mmHg | 0
oxygen saturation 98% | 0
normal vesicular breath sounds | 0
normal abdominal examination | 0
intravenous resuscitation | 0
analgesia | 0
WBC 8.2 × 10³/μL | 0
hemoglobin 11.5 g/dL | 0
thrombocytopenia 46,000/mm³ | 0
creatinine 117 μmol/L | 0
BUN 10.5 mmol/L | 0
sodium 131 mmol/L | 0
normal serum electrolytes | 0
normal liver profile | 0
normal coagulation profile | 0
normal chest X-ray | 0
P. falciparum with high parasitemia | 0
admitted to ICU | 0
intravenous artesunate-based regimen | 0
supportive measures | 0
shifted to general ward | 72
acute abdomen | 120
progressive dull constant generalized abdominal pain | 120
left upper quadrant pain | 120
nausea | 120
non-bilious vomiting | 120
lying still in bed | 120
anxious | 120
afebrile | 120
diaphoretic | 120
tachycardic | 120
tachypneic | 120
hypotensive | 120
saturating well on room air | 120
distended abdomen | 120
tender on superficial palpation | 120
inaudible bowel sounds | 120
Hb 7.1 g/dL | 120
ultrasound hypoechoic nodular cystic area | 120
splenomegaly | 120
CT scan hyperdense intrasplenic hematoma | 120
hypodense subcapsular hematoma | 120
splenic laceration | 120
intraperitoneal free fluid | 120
grade 3 splenic injury | 120
spontaneous splenic rupture | 120
resuscitation | 120
explorative laparotomy | 120
splenectomy | 120
evacuated 2.5 L frank blood | 120
enlarged spleen | 120
firm spleen | 120
splenic laceration on upper pole | 120
uneventful postoperative period | 168
discharged home | 168
