63 years old | 0
female | 0
admitted to the Emergency Department | 0
fever | -240
diarrhea | -240
confused | 0
febrile | 0
wet | 0
heart rate 121 bpm | 0
blood pressure 85/50 mmHg | 0
SpO2 95% | 0
fluid challenge with normal saline | 0
leukopenia | 0
low neutrophil count | 0
low lymphocyte count | 0
thrombocytopenia | 0
high levels of C-reactive protein | 0
high levels of D-dimers | 0
high levels of lactic dehydrogenase | 0
mild renal insufficiency | 0
rapid serology testing positive for SARS-CoV-2 | 0
nasopharyngeal swab test negative | 0
pulmonary CT scan showed diffuse pulmonary basal lobe opacifications | 0
empiric antibiotic therapy with meropenem and gentamycin | 0
admitted to the COVID-19 intensive care unit | 0
decrease in leukocytes and platelets | 24
coagulation tests indicating a diffuse intravascular coagulation | 24
blood and fresh frozen plasma transfusions | 24
sedated | 48
intubated | 48
mechanical ventilation | 48
extubated | 72
mental confusion | 72
unresponsiveness to external stimuli | 72
non-convulsive status epilepticus | 72
EEG recording | 72
benzodiazepine I.V. bolus | 72
ineffective benzodiazepine I.V. bolus | 72
I.V. levetiracetam | 72
SE resolution | 96
cerebral spinal fluid examination | 96
brain MRI | 96
discharged from ICU | 240
discharged home | 480
worsening mental slowing | 528
aphasia | 528
afebrile | 528
motor seizure | 528
right upper limb jerks | 528
bilateral tonic-clonic seizure | 528
confused | 528
partially oriented | 528
hypertonic and hyposthenic left lower limb | 528
focal convulsive SE | 528
STESS rating of 5 | 528
admitted to Neurology Unit | 528
brain MRI showed signal alterations | 528
diffuse intravascular coagulation | 528
second CSF examination | 528
polymerase chain reaction testing for SARS-CoV-2 and neurotropic viruses | 528
autoimmune panel for encephalitis | 528
serology test for SARS-CoV-2 antibodies | 528
nasopharyngeal swab | 528
cytokine levels | 528
whole-body positron emission tomography-computed tomography scan | 528
I.V. lacosamide | 544
motor signs ceased | 544
confusion persisted | 544
psychiatric symptoms | 544
behavioral disturbances | 544
persecutory ideation | 544
aggressiveness | 544
levetiracetam withdrawn | 550
treatment with valproic acid and dexamethasone | 550
clinically improved | 556
EEG monitoring showed SE resolution | 556
control brain MRI | 572
discharged home | 608
alert | 608
oriented to herself | 608
able to follow commands | 608
compliant | 608
no focal neurological deficits | 608
repetitive and fatuous | 608
lacosamide | 608
valproic acid | 608
slightly improved | 653
no further seizures | 653
new EEG | 653
mild diffuse slowing | 653
no epileptiform activity | 653