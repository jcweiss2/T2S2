53 years old | 0
male | 0
admitted to the emergency room | 0
fever | -72
myalgia | -72
confusion | -24
severe frontal headache | -24
no history of sick contacts | 0
no recent travels | 0
no recreational use of drug | 0
no history of chronic alcoholism | 0
no diabetes | 0
no chronic kidney disease | 0
no cardiac disease | 0
no recent throat infection | 0
no skin infection | 0
confused and lethargic | 0
Glasgow Coma Scale score of 10 | 0
could not follow commands | 0
neck rigidity on flexion | 0
rigidity in the left upper extremity | 0
increased tone on the left side | 0
white blood cell count of 10×10^9/L | 0
hemoglobin level of 13.4 g/dl | 0
thrombocytopenia with a platelet count of 54×10^9/L | 0
sodium level of 134 mEq/l | 0
calcium level of 8.4 mg/dl | 0
magnesium level of 1.7 mg/dl | 0
phosphorus level of 3.2 mg/dl | 0
bicarbonate level of 24 mEq/l | 0
blood glucose level of 142 mg/dl | 0
troponin level increased from 0.16 ng/ml–0.38 ng/ml | 0
electrocardiogram showed normal sinus rhythm | 0
ammonia level of 47 mcmol/l | 0
thyroid-stimulating hormone level within normal limits | 0
liver function tests within normal limits | 0
tested negative for flu | 0
tested negative for respiratory syncytial virus | 0
tested negative for coronavirus disease 2019 | 0
urine analysis negative | 0
urine toxicology screen negative | 0
salicylate and alcohol levels negative | 0
lumbar puncture performed | 0
elevated white blood cell count of 682×10^9/l | 0
neutrophil 81% | 0
red blood cell count of 10×10^9/l | 0
protein level of 117 mg/dl | 0
glucose level of 58 mg/dl | 0
possible bacterial meningitis | 0
admitted to the MICU | 0
received empirical therapy for meningitis | 0
vancomycin | 0
cefepime 2 g every 8 h | 0
ampicillin 2 g every 4 h | 0
new-onset left-sided weakness | 24
stroke team called | 24
computed tomography scan showed no evidence of intracranial hemorrhage | 24
incidental finding of a 778 mm mass concerning an aneurysm | 24
neurosurgery recommended a neuro interventional radiology consultation | 24
blood grew Methicillin-sensitive staphylococcal aureus | 24
antibiotics deescalated to Oxacillin 2 g | 24
steroid stopped | 24
transesophageal echo showed vegetation in the aortic valve | 24
intubated for respiratory distress | 48
persistently bacteremic and febrile | 48
ceftaroline added | 48
MRI showed a large posterior cerebral artery infarct | 48
cardiothoracic surgery team consulted for aortic valve replacement | 72
surgery not deemed appropriate | 72
repeat computed tomography head scan showed an intraparenchymal bleed | 96
lactic acid level started rising | 96
worsening kidney function | 96
bicarbonate administered | 96
oxygen saturation levels decreased to 40% | 120
cardiac arrest | 120
cardiopulmonary resuscitation initiated | 120
advanced life support measures employed | 120
patient could not be revived | 120
pronounced dead | 120