58 years old | 0
female | 0
alcoholism | -672
chronic obstructive pulmonary disease (COPD) | -672
tobacco abuse | -672
shortness of breath | 0
cough | 0
respiratory rate of 32 breaths/min | 0
temperature of 38.0°C | 0
heart rate of 115 bpm | 0
blood pressure of 73/40 mmHg | 0
oxygen saturation of 72% on room air | 0
lethargic but arousable to voice | 0
tachycardic but with regular rhythm and no murmurs | 0
mild respiratory distress with coarse rhonchi on auscultation of the lungs | 0
warm extremities with strong pulses | 0
white blood cell count (WBC) of 12.4×103 cells/uL | 0
arterial blood gas demonstrated a pH of 7.07 | 0
pCO2 of 106 mmHg | 0
pO2 of 80 mmHg | 0
bicarbonate of 30 mmol/L | 0
Chest X-ray (CXR) on admission did not demonstrate any acute pathology | 0
computed tomography (CT) imaging of the chest revealed evidence of multifocal pneumonia | 0
diagnosed with septic shock secondary to community-acquired pneumonia (CAP) | 0
started on ceftriaxone and azithromycin | 0
fluid resuscitated with 3 liters of lactated ringers | 0
started on norepinephrine | 0
intubated | 0
improved after a 5-day course of ceftriaxone and azithromycin | 120
liberated from norepinephrine on hospital day 2 | 48
fraction of inspired oxygen (FiO2) and positive end expiratory pressure (PEEP) were 40% and 5 cm H2O on hospital day 5 | 120
fraction of inspired oxygen (FiO2) and positive end expiratory pressure (PEEP) were 30% and 5 cm H2O on hospital day 6 | 144
successfully extubated in the morning on hospital day 6 | 144
developed respiratory distress with a respiratory rate of 28 breaths/min | 144
temperature of 38.2°C | 144
heart rate of 112 bpm | 144
blood pressure of 80/55 mmHg | 144
oxygen saturation of 85% on 60 L of heated high-flow oxygen therapy | 144
re-intubated and restarted on norepinephrine | 144
FiO2 and PEEP needs at this time were 100% and 5 cm H2O | 144
new left lower lobe infiltrate on CXR | 144
started on vancomycin and cefepime for treatment of VAP | 144
MRSA nasal swab taken from the bilateral nares after re-intubation was negative | 144
vancomycin was discontinued on hospital day 7 | 168
continued on cefepime monotherapy | 168
fevers up to 38.2°C | 168
up-trending leukocytosis | 168
ongoing vasopressor need | 168
culture from an endotracheal tube aspirate, collected from the day of re-intubation, tested positive for 3+ MRSA bacteria | 216
vancomycin was re-prescribed | 216
improved and was liberated from both norepinephrine and the ventilator | 240
transferred out of the ICU | 240
completed a total of 7 days of intravenous vancomycin | 288