54 years old | 0
female | 0
admitted to the hospital | 0
shortness of breath | 0
drowsiness | 0
type 2 diabetes mellitus | -8760
stopped metformin | -8760
stopped subcutaneous insulin | -8760
started lifestyle modifications | -8760
started traditional Chinese medications | -8760
polydipsia | -4320
back and thigh aches | -4320
weight loss | -4320
muscle atrophy | -4320
leg muscle atrophy | -4320
slow gait | -4320
difficulty climbing stairs | -4320
dehydration | 0
sinus tachycardia | 0
tachypnoea | 0
heart rate 125 | 0
respiratory rate 28 | 0
blood pressure 157/113 | 0
Glasgow Coma Scale 6 | 0
afebrile | 0
saturating well on room air | 0
cachexic | 0
malnourished | 0
equal and reactive pupils | 0
no pink skin | 0
no bright red lips | 0
no signs of pancreatitis | 0
lipaemic blood | 0
strawberry pink blood | 0
high anion gap metabolic acidosis | 0
lactic acidosis | 0
ketosis | 0
hyperkalaemia | 0
hypokalaemia | 0.5
severe hypertriglyceridaemia | 0
hypercholesterolaemia | 0
diabetic ketoacidosis | 0
sepsis | 0
intubated | 0
fluid resuscitation | 0
intravenous insulin | 0
discharged | 432
total serum cholesterol 47.07 mmol/L | 0
serum triglycerides 267.66 mmol/L | 0
high-density lipoprotein 0.28 mmol/L | 0
low-density lipoprotein 3.85 mmol/L | 0
glycated haemoglobin 8.2% | 0
urine full examination positive for glucose 4+ | 0
urine full examination positive for ketones 4+ | 0
urine full examination positive for proteins 4+ | 0
ECG sinus tachycardia | 0
CXR grossly normal | 0
abdominal X-ray grossly normal | 0
CT brain imaging grossly normal | 0
blood cultures positive for E. coli | 72
urine cultures negative | 72
started on statins | 96
started on fibrates | 96
started on omega-3 fish oil | 96
lactic acidosis resolved | 48
ketoacidosis resolved | 72
weaned off intravenous insulin | 96
extubated | 96
transferred out of ICU | 96
total serum cholesterol 11.69 mmol/L | 432
serum triglycerides 0.78 mmol/L | 432
random urine protein <0.04 mg/dL | 744
UFEME negative for glucose and ketones | 744