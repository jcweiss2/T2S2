48 years old | 0
woman | 0
sleeve gastrectomy for obesity | -480
referred to the ophthalmology clinic | 0
blurred vision in right eye | -72
reoperated 6 days after gastrectomy | -528
wound evisceration | -528
intensive care unit for 13 days | -528
systemic hypertension | 0
type 2 diabetes mellitus | 0
chronic obstructive pulmonary disease | 0
sleep apnea syndrome | 0
intravenous cefazolin for prophylaxis initiated | -528
recurrent fever | 0
blood cultures negative | 0
urine cultures negative | 0
rectal swab cultures negative | 0
Klebsiella pneumonia in catheter tip cultures | 0
Acinetobacter baumannii in catheter tip cultures | 0
colistin 150 mg IV 3 times a day | 0
clinical improvement not observed | 0
cultures repeated | 0
meropenem 2 g IV 3 times a day added | 0
referred for blurred vision in right eye persisting for 3 days | -72
visual acuity of light perception in right eye | 0
0.00 logMAR in left eye | 0
anterior segment examination normal | 0
light reaction results normal | 0
vitreous clear | 0
central hemorrhagic hypopigmented lesion in right fovea | 0
bulging from retina | 0
3 or 4 small hypopigmented lesions in both peripheral retinas | 0
SD-OCT showed hyperreflective vitreous dots | 0
elevated subfoveal lesion | 0
hyperreflective foveal lesion originated in choroidea | 0
hyperreflective dots in nearby vitreous | 0
fluorescein angiography revealed early hypofluorescence | 0
late phase leakage in foveal lesion | 0
suspected fungal chorioretinitis | 0
IV voriconazole maintenance dose 200 mg 2 times a day | 0
loading dose 6 mg/kg 2 times a day for 48 hours | 0
no deterioration in daily follow-up | 0
improvement in ocular findings on third day | 72
visual acuity counting fingers from 1 meter in right eye | 72
significant decrease in retinal lesions after 1 week | 168
no growth in final cultures | 168
IV voriconazole for 10 days | 0
oral voriconazole for 4 weeks | 240
first-month control visit | 720
right eye vision 0.20 logMAR | 720
left eye vision 0.00 logMAR | 720
anterior segment of both eyes natural | 720
pigment changes in right eye fovea | 720
SD-OCT revealed disruption of retinal pigment epithelium layer | 720
inner segment/outer segment junction disruption | 720
window defect in FA images | 720
