36 years old | 0
male | 0
admitted to the hospital | 0
splenectomy | -9360
abdominal pain | -24
vomiting | -24
septic shock | -24
norepinephrine | -24
peripheral ischemia of four extremities | -24
right knee disarticulation | -56
left trans-femoral amputation | -56
right elbow disarticulation | -56
skin flap operation of the right knee | -44
skin flap operation of the left hand | -41
joint range of motion exercise | -41
isometric exercise | -41
admitted to the Severance Rehabilitation Hospital | 0
prostheses measurement | 0
rehabilitation | 0
psychiatric consultation | -24
depression | -24
antidepressant medication | -24
anorexia | -24
sociophobia | -24
negative body image | -24
accepted situation | 0
got over with negative body image | 0
wanted active rehabilitation | 0
motivation increased | 0
short-term goals | 0
long-term goals | 0
multidisciplinary team approach | 0
right elbow disarticulation prosthesis | 168
elbow disarticulation socket | 168
elbow flexion device control unit | 168
elbow lock control cable | 168
outside locking hinge | 168
constant friction wrist unit | 168
figure of 8 harness | 168
artificial hand | 168
bimanual activity training | 168
left hand function test | 168
pinch power | 168
Box and Block Test | 168
limitation of using left hand as dominant hand | 168
motion of left wrist limited | 168
skin condition thin and fragile | 168
contracture of left hand | 168
decided right hand as dominant hand | 168
trained each hand proportionally | 168
wheelchair measurement | 168
ADL training on wheelchair level | 168
improve independency | 168
use walking aid more efficiently | 168
sitting balance good | 0
ADL training | 0
Functional Independence Measure score | 0
self-care subunit | 0
intensive ADL training | 168
don upper prosthesis by himself | 168
dressing | 168
eating | 168
grooming | 168
minimal assistance | 168
occupational therapy | 168
spoon use | 168
drinking with a cup | 168
buttoning and unbuttoning | 168
follow-up FIM score | 744
upper dressing by himself | 744
left hand muscle power improved | 744
hip joint muscle power improved | 744
strengthening exercise | 744
Cybex isokinetic training | 744
deconditioning | 0
impaired pulmonary function | 0
vital capacity | 0
peak cough flow | 0
Ambu bag | 168
air stacking exercise | 168
vital capacity improved | 744
peak cough flow improved | 744
right knee disarticulation prosthesis | 504
end bearing socket | 504
polycentric knee | 504
endoskeletal shank | 504
dynamic solid ankle cushion heel foot | 504
left trans-femoral amputation prosthesis | 672
quadrilateral socket | 672
polycentric knee | 672
endoskeletal shank | 672
dynamic SACH foot | 672
parallel bar weight shift training | 756
gait training with anterior walker | 840
gait pattern analyzed | 840
left leg dragged on swing phase | 840
shortened left leg | 840
improved gait pattern | 840
multidisciplinary team approach | 0
prostheses fitting | 0
hand function recovery | 0
gait pattern | 0
cane gait difficult | 840
walker indoors | 840
electronic wheelchair outdoors | 840
family education | 840
stump site management | 840
occupational rehabilitation program | 840
ADL training | 840
computer training | 840
car training | 840
rented a car for disabled people | 840
trained to move to driver's seat | 840
drive short distance | 840
universal cuff | 840
typing speed improved | 840
discharge | 1008
ADL independency improved | 1008
Functional Independence Measure score | 1008
Modified Barthel Index score | 1008
functional level status improved | 1008
absolute bed rest | 0
come to sit by himself | 1008
gait with anterior walker | 1008
follow-up | 1008
went back to work | 1008
used electronic wheelchair | 1008
performed ADL by himself | 1008
without help | 1008
on wheelchair level | 1008