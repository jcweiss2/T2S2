80 years old | 0
female | 0
non-smoker | 0
hypertension | 0
admitted to the hospital | 0
acute dyspnea | 0
fecal incontinence | -12
left hemiplegia | -12
dextroversion | -12
dysarthria | -12
vomiting | -12
impaired consciousness | 0
Japan coma scale score of Ⅱ-10 | 0
right thalamus and putamen bleeding | 0
conservative treatment | 0
Glasgow coma scale score 12 | 0
systolic blood pressure 91 mmHg | 0
respiratory rate 24/min | 0
oxygen saturation of arterial blood (SpO2) 86% | 0
poor oral hygiene | 0
diminished breath sounds on the left side | 0
coarse crackles in the right lung | 0
decrease in breath sounds in the front of the chest | 0
respiratory condition deteriorated | 0
endotracheal intubation | 0
mechanical ventilation | 0
bilateral infiltration | 0
admitted to the intensive care unit (ICU) | 0
decreased leukocyte count | 0
mildly elevated C-reactive protein (CRP) level | 0
respiratory failure | 0
partial pressure of oxygen in arterial blood (PaO2) 64 mmHg | 0
hepatorenal function normal | 0
extensive infiltration shadows on chest radiography | 0
hematoma extending from the right basal ganglia and putamen to the thalamus | 0
cerebral edema | 0
consolidations admixture with ground-glass opacities on chest CT | 0
A-DROP score corresponded to patient age | 0
increased blood urea nitrogen | 0
decreased SpO2 | 0
impaired consciousness | 0
antigen test for coronavirus disease 2019 negative | 0
Mendelson's syndrome | 0
aspiration of gastric contents | 0
chemical pneumonitis | 0
bacterial aspiration pneumonia | 0
sputum culture showed Streptococcus agalactiae and Klebsiella oxytoca | 0
leukocytopenia | 0
low serum CRP level | 0
respiratory viral pneumonia | 0
management in the ventilator mode started | 0
meropenem | 0
levofloxacin | 0
partial pressure of oxygen in arterial blood/fraction of inspired oxygen (PaO2/FiO2) 128.75 | 0
prednisolone started at 1 mg/kg/day | 0
infiltration shadows improved by Day 12 | 288
extubated on Day 12 | 288
transferred to the Department of Neurosurgery on Day 22 | 528
transferred to a rehabilitation hospital for sequelae of stroke | 528