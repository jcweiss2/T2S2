73 years old | 0
female | 0
hypertension | 0
diabetes mellitus type 2 | 0
diabetic nephropathy | 0
chronic renal impairment | 0
dual pacemaker | 0
sick sinus syndrome | 0
ST elevation myocardial infarction | -8760
three drug-eluting stents | -8760
PEG | -4320
refusal to eat | -4320
possibility of true bulbar palsy | -4320
early signs of Alzheimer's disease | -4320
furosemide 80 mg twice daily | 0
carvedilol 6.25 mg twice daily | 0
spironolactone 50 mg once daily | 0
clopidogrel 75 mg once daily | 0
admitted with hypotension | 0
pulmonary edema | 0
ventilator support | 0
tracheal intubation | 0
inotropes | 0
renal replacement therapy | 0
improvement | 0
extubated | 72
acute on chronic renal failure | 72
restart of renal replacement therapy | 72
severe global hypokinesia of the left ventricle | 0
low ejection fraction (< 20%) | 0
bilateral lung ultrasonic B lines | 0
bilateral mild pleural effusions | 0
low cardiac output | 0
generalized edema | 0
improved initially | 0
noradrenaline infusion discontinued | 0
dobutamine infusion discontinued | 0
hemodialysis | 168
hypotension episode (85/42 mm Hg) | 168
noradrenaline infusion during procedure | 168
tachypnea (33 breaths/min) | 168
vague abdominal pain | 168
blood pressure 105/45 mm Hg | 168
heart rate 93 beats/min | 168
abdomen slightly distended | 168
nontender abdomen | 168
hypoactive bowel sounds | 168
elevated alanine aminotransferase (360.1 U/L) | 168
elevated aspartate aminotransferase (577.3 U/L) | 168
elevated lactate dehydrogenase (381 U/L) | 168
elevated white blood cell count (16.00 × 10^3/L) | 168
elevated C-reactive protein (83.4 mg/L) | 168
anion gap metabolic acidosis | 168
lactate rising from 1.8 to 8.6 mmol/L | 168
pH 7.00 | 168
lactic acidosis | 168
restart of noradrenaline infusion | 168
restart of dobutamine infusion | 168
reintubated | 168
POCUS showed sluggish intestinal movement | 168
echocardiography showed impaired systolic function | 168
hyperechoic dot artifacts in liver | 168
portal venous gas | 168
pneumatosis intestinalis | 168
CT showed portal venous gas | 168
gas in superior mesenteric vein | 168
gas in stomach walls | 168
gas in right colon | 168
gas in small bowel loops | 168
atherosclerotic changes in aorta | 168
attenuated hepatic artery | 168
attenuated superior mesenteric artery | 168
attenuated celiac trunk | 168
nonvisualized inferior mesenteric artery | 168
minimal pelvic fluid | 168
no occlusive thrombosis | 168
no significant luminal narrowing | 168
diagnosed with nonocclusive diffuse intestinal ischemia | 168
family counseled | 168
no further interventions recommended | 168
passed away | 216
ST elevation myocardial infarction | -7200
three drug-eluting stents | -7200
hemodialysis | 240
hypotension episode (85/42 mm Hg) | 240
