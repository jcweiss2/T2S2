72 years old| 0
female| 0
known diabetic for last 16 years| 0
admitted to the intensive care unit| 0
sudden onset unconsciousness| -12
oral hypoglycemic drugs| 0
poor glycemic control| 0
hypertensive| 0
controlled on medication| 0
no history of convulsions| 0
no history of fever| 0
no history of vomiting| 0
no history of headache| 0
no history of trauma| 0
no history of neurodeficit| 0
neurological score 5/15| 0
pulse 88/min| 0
blood pressure 140/80 mm Hg| 0
respiratory rate 16/min| 0
irregular bilateral vesicular breath sounds| 0
capillary blood glucose 28 mg/dL| 0
total leukocyte count 16,200/mm3| 0
neutrophil predominance| 0
serum alanine aminotransferase 31 IU/mL| 0
serum aspartate aminotransferase 71 IU/mL| 0
alkaline phosphatase 22 IU/L| 0
total protein 4.8 g/dL| 0
albumin 2.4 g/dL| 0
urea 54 mg/dL| 0
creatinine 1.2 mg/dL| 0
total bilirubin 0.6 mg/dL| 0
conjugated bilirubin 0.3 mg/dL| 0
computerized tomographic scan showed focal ischemia| 0
hypoglycemic encephalopathy| 0
hypoxic brain damage| 0
intubated| 0
ventilator support| 0
glycemic status restored| 0
piperacillin + tazobactam| 0
day 3 of treatment| 72
response to painful stimulus| 72
blood sugar uncontrolled| 72
day 4 of treatment| 96
low grade fever| 96
endotracheal secretions culture| 96
Acinetobacter baumanii isolated| 96
significant colony count (>106 CFU)| 96
sensitive to netilmicin| 96
sensitive to polymixin B| 96
blood cultures sent| 72
no growth| 72
chest X-ray mild right sided basal opacity| 72
netilmicin| 96
cefepime| 96
day 7 of treatment| 168
high grade fever| 168
total leukocyte count 8400/mm3| 168
neutrophilic predominance| 168
serum creatinine 2 mg/dL| 168
catheterized urine sample culture| 168
blood culture sent| 168
urine culture Escherichia coli| 168
sensitive to meropenem| 168
sensitive to polymyxin B| 168
sensitive to cotrimoxazole| 168
sensitive to nitrofurantoin| 168
meropenem added| 168
general condition deteriorated| 168
total leukocyte count 4000/mm3| 168
blood cultures sent on day 7| 168
blood cultures sent on day 8| 168
Enterococcus faecium growth| 168
standard laboratory procedures| 168
antibiotic susceptibility by Kirby Bauer disc diffusion| 168
sensitive to vancomycin| 168
resistant to linezolid| 168
disk diffusion testing| 168
E-test linezolid strips| 168
no zone of inhibition| 168
MIC >256 μg/mL| 168
agar dilution method| 168
MIC 1024 μg/mL| 168
automated susceptibility testing by Vitek 2| 168
vancomycin started| 168
condition deteriorated| 168
declared dead| 360
other ICU patients cultures| 168
no similar organisms| 168
no previous history of linezolid medication| 0
linezolid resistant enterococci| 168
vancomycin susceptible| 168
ampicillin susceptible| 168
tetracycline susceptible| 168
aminoglycosides susceptible| 168
teicoplanin susceptible| 168
nosocomial spread| 168
fatal case| 360
