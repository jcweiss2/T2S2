39 years old | 0
female | 0
partial pancreaticoduodenectomy due to periampullary neuroendocrine tumor | -25920
periampullary neuroendocrine tumor with locoregional extension | -25920
9/12 metastatic lymph nodes | -25920
neuroendocrine tumor | -25920
immunohistochemically positive for gastrin | -25920
Ki 67 5% | -25920
Grade 2 | -25920
liver metastases | -21600
monthly dose of 120 mg lanreotide | -21600
progression of liver metastases | -19440
sunitinib | -19440
discontinued sunitinib | -19440
extreme fatigue | -19440
muscle weakness | -19440
delirium | -19440
moon face | 0
hirsutism | 0
severe proximal weakness | 0
anemia | 0
hyperglycemia | 0
severe hypokalemia | 0
24-h urinary free cortisol: 2152 nmol/day | 0
morning serum cortisol 4883.4 nmol/L | 0
plasmatic ACTH 127.3 pmol/L | 0
SCS due to EAS | 0
ketoconazole | 0
acute upper gastrointestinal bleeding | 0
hemodynamic instability | 0
subendocardial ischemia | 0
atrial fibrillation | 0
Forrest Ib gastric ulcer | 0
intravenous fluconazole 400 mg/day | 0
mental state improved | 48
morning cortisol decreased 25% | 48
fluconazole titrated to 600 mg/day | 72
cortisolemia decreased 55% | 168
liver transaminases increased 3 times over normal limit | 168
fluconazole decreased to 400 mg/day | 168
bilirubin and albumin levels remained normal | 168
prothrombin time remained normal | 168
baseline cortisol decreased by 65% | 168
hypokalemia | 0
metabolic alkalosis | 0
acetazolamide 250 mg/day | 0
spironolactone | 0
amiloride | 0
severe thrombocytopenia | 0
multiple platelet transfusions | 0
intravenous Gamma globulin | 0
bone marrow biopsy | 0
marked hypocellularity | 0
viral serology tests negative | 0
Eltrombopag | 0
bilateral adrenalectomy | 360
hydrocortisone | 360
fludrocortisone | 360
lanreotide 120 LAR | 360
prolonged hospitalization in ICU | 360
sepsis | 360
emphysematous cystitis | 360
disseminated Herpes Zoster infection | 360
antibiotics | 360
intravenous acyclovir | 360
chemoembolization of liver metastases | 432
liver metastases decreased in size | 432
rehabilitation therapy program | 17520
depression | 0
physical and psychological impairment | 0
