67 years old | 0
female | 0
admitted to the hospital | 0
right loin pain | -12
vomiting | -12
denies urinary symptoms | -12
denies haematuria | -12
autoimmune liver cirrhosis | 0
atrophic gastritis | 0
Type 2 diabetes mellitus | 0
hysterectomy | -1560
coronary artery bypass surgery | -1560
metformin | 0
non-anaphylactic reactions to penicillin | 0
non-anaphylactic reactions to IV contrast | 0
pale | 0
temperature of 36.8 °C | 0
BP 141/72 | 0
pulse of 81 beats per minute | 0
generalised right sided tenderness | 0
right upper quadrant tenderness | 0
loin tenderness | 0
no crepitus | 0
anaemia | 0
Hb 9.8 g/dL | 0
impaired renal function | 0
urea 13.2 mmol/L | 0
creatinine 183 μmol/L | 0
HbA1c of 5.3% | 0
normal liver function tests | 0
prothrombin time 17.5 s | 0
activated partial thromboplastin time 37.4 s | 0
absence of neutrophil leucocytosis | 0
WCC 9 × 10^9/L | 0
urinalysis displaying trace of blood | 0
Urology referral | 0
CTKUB | 0
gas outlining the pelvicalyceal system of the right kidney | 0
perifascial gas tracking along the right ureter | 0
no discrete fluid collections | 0
no calculi | 0
intravenous antibiotics | 0
intravenous fluids | 0
blood cultures | 0
urine cultures | 0
Escherichia coli | 0
sensitive to Meropenem | 0
Metronidazole | 0
anaerobic cover | 0
pyrexia | 12
tachycardia | 12
hypotension | 12
oliguria | 12
high dependency unit | 12
C-reactive protein 8 mg/L | 0
C-reactive protein 109 mg/L | 24
leucocyte count 6 g/dL | 12
platelet count 198 × 10^9/L | 0
platelet count 100 × 10^9/L | 12
kidney function deterioration | 12
creatinine 258 μmmol/L | 12
severe sepsis | 12
end-organ failure | 12
emergency right nephroureterectomy | 24
open approach | 24
right loin incision | 24
peritoneum opened | 24
free peritoneal fluid | 24
cirrhosis of the liver | 24
abdominal viscera normal | 24
necrosis of the right renal pelvis | 24
necrosis of the right ureter | 24
oedema in the retroperitoneum | 24
peri-ureteric gas | 24
no perinephric abscess | 24
no collection | 24
right nephrectomy | 24
ligation of the renal vessels | 24
kidney specimen | 24
ureter specimen | 24
retroperitoneal space | 24
inferiorly towards the pelvis | 24
main wound closed | 24
second incision | 24
diseased distal ureter excised | 24
en bloc with the kidney specimen | 24
retroperitoneal drain | 24
urethral catheter | 24
intensive care unit | 24
histopathology analysis | 48
microscopic parenchymal abscesses | 48
perinephric fat | 48
haemorrhagic infarction of the ureteric mucosa | 48
serositis | 48
pyrexia | 96
CT of the abdomen and pelvis | 96
small bilateral pleural effusions | 96
normal post-operative changes | 96
no significant retroperitoneal collections | 96
IV antibiotics | 0
7 days of IV antibiotics | 168
smooth recovery | 168
discharged | 312
follow-up | 336
no early complications | 336
admission with worsening renal function | 744
conservatively managed | 744
long term nephrology follow-up | 744