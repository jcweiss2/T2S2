74 years old | 0
male | 0
non-traumatic acute subdural hematoma | -24
emergency cranial trepanation | -24
mechanical ventilation | -24
ventilator-associated pneumonia | -24
CT scan | 0
soft-tissue infection of the craniotomy wound | 0
purulent secretion | 0
erythema | 0
swelling | 0
cerebral herniation | 0
elevated intracranial pressure | 0
midline shift | 0
external ventricular drain | 0
surgical revision | 0
intraoperative exploration | 0
old hematoma | 0
deep purulent secretion | 0
intracranial abscess formation | 0
empirical antibiotic therapy | 0
meropenem | 0
rifampicin | 0
vancomycin | 0
intraoperative swabs | 0
blood culture series | 0
bronchoalveolar lavage | 0
diagnosis of intracranial abscess | 24
leucocyte count | 0
C-reactive protein level | 0
fever | 0
septic shock | 24
norepinephrine therapy | 24
Gram-negative pathogens | 48
MDR Acinetobacter baumannii | 48
MDR Klebsiella pneumoniae | 48
intravenous fosfomycin | 48
intravenous meropenem | 48
intravenous colistin | 48
intraventricular colistin | 48
chest radiography | 192
tracheal aspirates | 192
normothermia | 192
de-escalation strategy | 192
TDM | 240
colistin levels | 240
renal function | 240
acute renal insufficiency | 312
continuous venovenous hemodialysis | 312
intermittent dialysis | 336
oliguria | 336
urine output increased | 432
dialysis weaned | 432
sufficient renal function | 432
quantitative resistance testing | 240
sensitivity to colistin | 240
repetitive drainage of CSF | 240
lumbar Tuohy catheter | 240
intrathecal colistin stopped | 624
intravenous colistin monotherapy | 624
colistin serum levels | 624
CSF levels | 624
sterile microbiological analyses | 624
ICU treatment | 1920
neurological rehabilitation facility | 1920
follow-up | 4320
neurological side effect | 4320
intraventricular colistin therapy | 4320