35 years old | 0
female | 0
admitted to the emergency room | 0
generalized tonic-clonic seizures | -3
urinary incontinence | -3
altered sensorium | -3
headache | -3
unsafe abortion | -240
severe fatigue | -240
shortness of breath | -240
pedal edema | -240
severe anemia | -240
ongoing blood loss | -240
blood transfusion | -240
drowsy | 0
not obeying commands | 0
withdraws limbs to painful stimuli | 0
deep tendon reflexes sluggish | 0
withdrawal response in plantar reflex | 0
normal hemoglobin | 0
neutrophilic leukocytosis | 0
urinary tract infection | 0
elevated C-reactive protein | 0
normal ESR | 0
normal liver function tests | 0
normal renal function tests | 0
dimorphic anemia | 0
normal coagulation profile | 0
normal autoantibodies | 0
normal neoplastic markers | 0
increased cerebrospinal fluid protein | 0
normal chest radiography | 0
normal arterial blood gas analysis | 0
MRI brain findings | 0
electroencephalography epileptiform discharges | 0
incomplete right bundle branch block | 0
admitted to intensive care unit | 0
intravenous fluids | 0
antibiotics | 0
antiepileptics | 0
blood pressure monitoring | 0
normal sensorium | 168
normal leukocyte counts | 168
normal vital signs | 168
discharged | 168
uneventful follow-up | 240
35 years old|0
female|0
admitted to the emergency room|0
generalized tonic-clonic seizures|-3
urinary incontinence|-3
altered sensorium|-3
headache|-3
unsafe abortion|-240
severe fatigue|-240
shortness of breath|-240
pedal edema|-240
severe anemia|-240
ongoing blood loss|-240
blood transfusion|-240
drowsy|0
not obeying commands|0
withdraws limbs to painful stimuli|0
deep tendon reflexes sluggish|0
withdrawal response in plantar reflex|0
normal hemoglobin|0
neutrophilic leukocytosis|0
urinary tract infection|0
elevated C-reactive protein|0
normal ESR|0
normal liver function tests|0
normal renal function tests|0
dimorphic anemia|0
normal coagulation profile|0
normal autoantibodies|0
normal neoplastic markers|0
increased cerebrospinal fluid protein|0
normal chest radiography|0
normal arterial blood gas analysis|0
MRI brain findings|0
electroencephalography epileptiform discharges|0
incomplete right bundle branch block|0
admitted to intensive care unit|0
intravenous fluids|0
antibiotics|0
antiepileptics|0
blood pressure monitoring|0
normal sensorium|168
normal leukocyte counts|168
normal vital signs|168
discharged|168
uneventful follow-up|240
