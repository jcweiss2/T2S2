65 years old | 0
male | 0
family history of diabetes mellitus | 0
prostatic hyperplasia | 0
simple umbilical hernia repaired | 0
admitted to the hospital | 0
diffuse abdominal pain | -120
nausea | -120
vomiting | -120
abdominal distension | -120
inability to pass flatus | -24
inability to evacuate | -24
tachycardia | 0
hypotension | 0
diffuse abdominal tenderness | 0
peritoneal irritation | 0
severe distension | 0
leukocytosis | 0
hemoglobin 18.1 g/dL | 0
platelet count 207 × 10^3 | 0
acute renal failure | 0
serum creatinine 3 mg/dL | 0
blood urea nitrogen 60 mg/dL | 0
urea 210 mg/dL | 0
dilated loops | 0
no free air | 0
thick and irregular fibrous capsule at the base of the appendix | 0
central low-attenuation necrotic component | 0
surrounding inflammatory changes | 0
periappendiceal reactive nodal enlargement | 0
pneumoperitoneum | 0
dilated large bowel | 0
appendix enlarged | 0
perforation at the tip of the appendix | 0
bowel perforation | 0
peritonitis | 0
emergency laparotomy | 0
massive bowel dilatation | 0
purulent intraperitoneal fluid | 0
appendectomy | 0
postoperative care | 0
moderate pain | 24
oral intake reintroduced | 72
discharged | 168
follow-up examination | 720
follow-up examination | 4320
inflammatory myofibroblastic tumor | 0
fibroblastic proliferation | 0
dense inflammatory infiltrate | 0
myxoid changes | 0
spindle cells | 0
polyclonal plasma cells | 0
lymphocytes | 0
vimentin positive | 0
smooth muscle actin positive | 0
anaplastic lymphoma kinase negative | 0
septic shock | 0
visceral perforation | 0
tumor-like lesion | 0
histological examination | 0
immunohistochemistry | 0