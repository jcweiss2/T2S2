50 years old | 0
    woman | 0
    admitted for altered mental status | 0
    acute alcohol intoxication | 0
    binge drinking an unknown quantity of wine | -12
    blood pressure of 88/58 mm Hg | 0
    drowsy | 0
    arousable | 0
    partially oriented | 0
    blood alcohol level of 353 mg/dl | 0
    anion gap of 17 | 0
    lactate of 4.5 mmol/L | 0
    beta hydroxybutyrate of 0.7 mmol/L | 0
    positive urine ketones | 0
    serum glucose of 80 mg/dl | 0
    serum osmolality of 383 mOsm/kg | 0
    normal serum osmolal gap | 0
    elevated ethanol | 0
    undetectable levels of methanol | 0
    undetectable levels of isopropanol | 0
    undetectable levels of acetone | 0
    received 7 L of normal saline | 0
    hypotension | 0
    serum alcohol normalized | 12
    anion gap normalized | 12
    lactate normalized | 12
    serum ketones normalized | 12
    hypotension normalized | 12
    mental status normalized | 12
    workup for sepsis | 12
    unresponsive | 24
    blood pressure of 93/60 mm Hg | 24
    Glasgow Coma Score of 3 | 24
    required fluid resuscitation | 24
    intubation for airway protection | 24
    CT of the head unremarkable | 24
    lactate increased to 4.5 mmol/L | 24
    anion gap increased to 17 | 24
    extubated | 48
    serum lactate normalized to 1.4 mmol/L | 48
    anion gap normalized to 7 | 48
    mental status returned to alert | 48
    mental status returned to fully oriented | 48
    unresponsive | 72
    next to an open and empty bottle of ethanol based hospital hand sanitizer | 72
    vital signs normal | 72
    Glasgow Coma Score of 3 | 72
    repeat head CT unremarkable | 72
    lactate of 3.9 mmol/L | 72
    anion gap of 15 | 72
    serum ethanol of 362 mg/dl | 72
    methanol of 0 mg/dl | 72
    acetone of 11 mg/dl | 72
    isopropanol of 14 mg/dl | 72
    arterial blood gas pH of 7.32 | 72
    PaCO2 43 mm Hg | 72
    PaO2 73 mm Hg | 72
    bicarbonate 22 mmol/L | 72
    admitted to the intensive care unit | 72
    required nasopharyngeal airway | 72
    required supportive care | 72
    mental status gradually returned to normal | 78
    elevated lactate levels gradually returned to normal | 78
    metabolic acidosis gradually returned to normal | 78
    admitted to drinking ethanol based hospital hand sanitizer | 78
    denied suicidality | 78
    hand sanitizers removed from her room | 78
    placed on one-to-one monitoring | 78
    discharged | 78
    in-patient alcohol treatment program | 78