45 years old | 0
male | 0
admitted to the hospital | 0
upper abdominal pain | -72
nausea | -72
vomiting | -72
tender abdomen | 0
no muscle guarding | 0
high-grade infection | 0
no pneumoperitoneum | 0
widespread thickening of the gastric wall | 0
diffuse erythema | 0
edema of the gastric wall | 0
gastric ischemia | 0
malignancy | 0
H2-blocker therapy | 0
antibiotic therapy with cefuroxime and metronidazole | 0
septic shock | 24
multiple organ failure | 24
high serum lactate | 24
diagnostic laparoscopy | 24
laparotomy | 24
total gastrectomy | 24
intensive care unit admission | 24
hemodynamic support | 24
continuous veno-venous hemofiltration | 24
Roux-Y esophagojejunostomy | 48
streptococcal toxic shock syndrome | 48
group A Streptococcus | 48
phlegmonous gastritis | 48
discharged | 336
leukocytes 21.5 10E9/L | 0
C-reactive protein (CRP) 281 mg/L | 0
creatinine 83 μmol/L | 0
urea 6.1 mmol/L | 0
lactate - | 24
leukocytes 25.8 10E9/L | 24
C-reactive protein (CRP) 366 mg/L | 24
creatinine 424 μmol/L | 24
urea 17.4 mmol/L | 24
lactate 9.2 mmol/L | 24