60 years old | 0
male | 0
Saudi | 0
admitted to King Khalid University Hospital | 0
erythroderma | -1300
pruritic | -1300
erythematous lesions | -2600
trunk | -2600
retroauricular area | -2600
misdiagnosed as severe eczema | -2600
treated with oral prednisolone | -2600
treated with oral cyclosporine | -2600
no improvement | -2600
confluent lichenified erythromelanotic plaques | 0
greasy scales | 0
face | 0
neck | 0
trunk | 0
genitalia | 0
upper extremities | 0
lower extremities | 0
palms | 0
soles | 0
sparing of the nails | 0
sparing of the scalp | 0
bilateral lower lid ectropion | 0
skin punch biopsies | 0
lower back | 0
left buttock | 0
right upper extremity | 0
epidermotropism | 0
atypical lymphocytes | 0
lymphocytic band infiltrate | 0
dermal fibrosis | 0
immunofluorescence study | 0
negative for fibrinogen | 0
negative for C3 | 0
negative for IgA | 0
negative for IgM | 0
negative for IgG | 0
tumor cells positive for CD3 | 0
tumor cells positive for CD45RO | 0
tumor cells negative for CD4 | 0
tumor cells negative for CD8 | 0
tumor cells negative for CD7 | 0
CD30 positive | 0
peripheral blood count normal | 0
peripheral blood smear normal | 0
no Sézary cells | 0
flow cytometry of peripheral blood | 0
no evidence of monoclonality | 0
CT scan of abdomen and pelvis | 0
enlarged bilateral external iliac lymph nodes | 0
enlarged inguinal lymph nodes | 0
no solid organ involvement | 0
CT scan of chest | 0
no lymphadenopathy | 0
ultrasound-guided incisional lymph node biopsy | 0
atypical cells | 0
negative for clonal T-cell receptor gene rearrangement | 0
diagnosis of double-negative CD4/CD8 MF | 0
advanced stage | 0
referred to hematology and oncology unit | 0
plan of further staging | 0
excisional lymph node biopsy | 0
septic shock | 720
admitted to intensive care unit | 720
passed away | 1440
1.5 months after diagnosis | 1440 
5 years after the start of symptoms | -1300