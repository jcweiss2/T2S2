59 years old | 0
male | 0
non-obstructive hypertrophic cardiomyopathy | 0
hospitalized | 0
cardiac insufficiency | 0
inotropic therapy | 0
worsening of clinical picture | 0
use of intra-aortic balloon | 0
prioritized for cardiac transplantation | 0
pre-transplant period | 0
infectious complications | 0
blood cultures | -48
blood cultures | -24
bicaval-bipulmonary heart transplantation | 0
surgery | 24
hemostasis | 24
mechanical ventilation | 0
vasoactive drugs | 0
intra-aortic balloon | 0
good clinical condition | 0
mycophenolate mofetil | 0
cyclosporine | 0
prednisone |A 59-year-old male patient with non-obstructive hypertrophic cardiomyopathy was hospitalized to manage cardiac insufficiency with inotropic therapy. The worsening of his clinical picture required the use of an intra-aortic balloon, and he was prioritized for cardiac transplantation. During the pre-transplant period, the patient did not develop any infectious complications. Blood cultures collected 24 and 48 h before transplantation were negative.
