69 years old | 0
female | 0
admitted to the emergency department | 0
oral ingestion of Roundup | -2
vomiting | -2
lethargy | -2
conscious and disoriented | 0
Glasgow coma scale of 12 | 0
blood pressure 91/56 mmHg | 0
SpO2 of 91% | 0
tenderness throughout the abdomen | 0
gastric lavage | 0
transferred to the emergency ICU | 0
hydrated with normal saline | 0
correction of acidosis with sodium bicarbonate | 0
arterial blood gas analysis | 0
elevated serum lactate level | 0
hemoperfusion | 0
decreased consciousness level | 6
required ventilatory support | 6
vasoactive support | 6
high total leukocyte count | 6
elevated creatinine | 6
elevated glutamic oxalacetic transaminase | 6
elevated alanine aminotransferase | 6
elevated alkaline phosphatase | 6
elevated creatine kinase | 6
uncontrolled seizures | 8
elevated lactate levels | 8
worsening metabolic acidosis | 8
administering multiple high-dose vasoactive agents | 8
structured fat emulsion injection | 8
large amount of fluid | 8
low blood pressure | 8
CRRT initiated | 8
infusion of large amounts of plasma | 8
albumin infusion | 8
glucocorticoids | 8
ulinastatin | 8
increased urine output | 8
stabilized blood pressure | 8
pulmonary effusion | 8
massive fluid accumulation in the intestinal wall and lumen | 8
edema in the interstitial spaces | 8
capillary leak syndrome | 8
CRRT discontinued | 72
extubated | 168
transferred out of the intensive care unit | 240
discharged | 480
no abnormal signs and symptoms at 3 months | 744