67 years old | 0
    male | 0
    hypertension | 0
    schizophrenia | 0
    shortness of breath | -24
    generalized weakness | -24
    nausea | -24
    diarrhea | -24
    abrupt onset | -24
    denies splenectomy | 0
    nonsmoker | 0
    denies illicit drug use | 0
    denies heavy alcohol consumption | 0
    resides in group home | 0
    denies sick contacts | 0
    refused pneumococcal vaccination | 0
    refused influenza vaccination | 0
    hypotension | 0
    blood pressure 80/30 mm Hg | 0
    fever 101.1°F | 0
    clear lungs | 0
    regular heart sounds | 0
    no hepatosplenomegaly | 0
    no peritoneal signs | 0
    normal neurologic examination | 0
    denies headache | 0
    denies cough | 0
    denies chest pain | 0
    watery non-bloody diarrhea | 0
    WBC 42.3/nL | 0
    neutrophils predominance | 0
    hemoglobin 10 g/dL | 0
    platelet count 78/nL | 0
    BUN 47 mg/dL | 0
    creatinine 5.5 mg/dL | 0
    bicarbonate 19.2 mEq/L | 0
    anion gap 23 | 0
    lactic acid 4.3 mmol/L | 0
    alkaline phosphatase 162 U/L | 0
    AST 210 U/L | 0
    total bilirubin 2 mg/dL | 0
    direct bilirubin 0.4 mg/dL | 0
    CK 5750 U/L | 0
    fibrinogen 170 mg/dL | 0
    LDH 5490 U/L | 0
    D-dimer >69,000 ng/mL | 0
    microangiopathic hemolytic anemia | 0
    schistocytes | 0
    CT chest negative | 0
    CT abdomen negative | 0
    CT pelvis negative | 0
    no pulmonary infiltrates | 0
    no colitis | 0
    no intraabdominal infection | 0
    diagnosed severe sepsis | 0
    admitted to ICU | 0
    fluid resuscitation 30 mL/kg | 0
    vancomycin | 0
    piperacillin-tazobactam | 0
    developed retiform violaceous patches | 0
    central dusky necrosis | 0
    upper extremities involvement | 0
    thighs involvement | 0
    back involvement | 0
    lower legs involvement | 0
    dorsal feet involvement | 0
    abdomen involvement | 0
    retiform purpura | 0
    ischemic changes | 0
    gangrene | 0
    required norepinephrine | 24
    blood cultures Gram positive cocci | 24
    discontinued piperacillin-tazobactam | 24
    initiated ceftriaxone | 24
    initiated clindamycin | 24
    identified S. pneumoniae | 24
    antibiotics narrowed to ceftriaxone | 24
    Legionella negative | 24
    Clostridioides difficile negative | 24
    oliguric renal failure | 24
    hemodialysis initiated | 24
    echocardiogram no vegetations | 24
    preserved ejection fraction | 24
    repeat blood cultures negative | 24
    weaned off norepinephrine | 72
    β-D-Glucan Assay negative | 72
    Strongyloides serology negative | 72
    antiphospholipid antibodies negative | 72
    anti-cardiolipin antibodies negative | 72
    C-ANCA negative | 72
    PANCA negative | 72
    complement C3 normal | 72
    complement C4 normal | 72
    cryoglobulin negative | 72
    HIV negative | 72
    HBV negative | 72
    HCV negative | 72
    renal function improved | 168
    liver function improved | 168
    weaned off hemodialysis | 168
    rash nearly resolved | 168
    septic shock | 0
    multiorgan failure | 0
    disseminated intravascular coagulation | 0
    PF | 0
    <|eot_id|>
    