48 years old | 0
postmenopausal female | 0
lateral neck pain | -240
diabetic | -6720
oral hypoglycemic medication | -96
skipped medication | -96
hypothyroidism | 0
hypertension | 0
thyroxine | 0
liraglutide | 0
repaglinide | 0
aspirin | 0
atorvastatin | 0
alcohol | 0
admitted to hospital | 0
neck examination | 0
localized ill-defined area | 0
tender | 0
local rise in temperature | 0
crepitations | 0
distal neurovascular status intact | 0
lymph nodes palpable | 0
total leukocyte count | 0
neutrophils | 0
hemoglobin level | 0
platelets count | 0
random blood sugar level | 0
serum urea | 0
serum creatinine | 0
serum sodium | 0
serum potassium | 0
urine examination | 0
serum protein | 0
serum albumin | 0
arterial blood gas analysis | 0
diagnosis of diabetic ketoacidosis | 0
neck abscess | 0
insulin | 0
intravenous fluids | 0
piperacillin | 0
tazobactam | 0
ultrasonography neck | 12
large ill-defined mass | 12
neck exploration | 24
wound swab | 24
pseudomonas aeruginosa | 24
ciprofloxacin | 24
amikacin | 24
histopathology report | 24
necrotizing fasciitis | 24
daily dressing | 24
oral feeding | 48
lab reports | 168
hematological parameters | 168
renal function | 168
blood sugar | 168
wound healing | 168
discharged home | 168
regular dressing | 168
blood sugar monitoring | 168