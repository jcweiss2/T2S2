3 years 2 months old | 0
    female | 0
    admitted to the hospital | 0
    personality changes | -336
    behavioral regression | -288
    unsteady gait | -288
    headache | -288
    irritable crying | -288
    catatonia-like response | -288
    generalized choreoathetoid movements | -288
    orofacial dyskinesia | -288
    collapsed lung | -288
    transferred to pediatric intensive care unit | -288
    cerebrospinal fluid pleocytosis | 0
    lymphocytes predominance | 0
    leptomeningeal enhancement | 0
    nodular enhancement along tentorium | 0
    tiny white-matter lesions | 0
    global cortical dysfunction | 0
    no epileptiform discharge | 0
    empiric treatment with acyclovir | 0
    empiric treatment with azithromycin | 0
    positive NMDA receptor antibody | 0
    intravenous immunoglobulin | 0
    pulse methylprednisolone therapy | 0
    maintenance oral prednisolone | 0
    aripiprazole | 0
    midazolam sedation | 0
    choreoathetosis | 0
    orofacial dyskinesia | 0
    episodic sepsis | 0
    autonomic instability | 0
    gastrointestinal bleeding | 0
    plasmapheresis | 1680
    anaphylactic reactions | 1680
    bilateral pneumonia | 1680
    collapsed lung | 1680
    rituximab | 1680
    cyclophosphamide pulse therapy | 1680
    azathioprine | 1680
    passive range-of-motion exercise | 0
    generalized choreoathetosis | 0
    facilitation training | 0
    postural training | 0
    percutaneous endoscopic gastrostomy | 0
    discharged | 5040
    maximal assistance in mobility | 5040
    maximal assistance in self-care | 5040
    maximal assistance in cognition | 5040
    physical therapy | 5040
    occupational therapy | 5040
    speech therapy | 5040
    developmental age 6–8 months gross-motor | 8760
    developmental age 6–8 months fine-motor | 8760
    developmental age 9–12 months cognition | 8760
    simple verbal orders | 8760
    mutism | 8760
    cognitive deficits | 8760
    gross-motor skills 24–27 months | 17520
    fine-motor skills 20–23 months | 17520
    cognition 24–29 months | 17520
    simple self-care tasks | 17520
    occasional incontinence | 17520
    speak more than five words | 17520
    tricycle riding | 17520
    balance-beam exercise | 17520
    cognitive-behavioral therapy | 26280
    attention improvement | 26280
    memory improvement | 26280
    emotion regulation | 26280
    full IQ 62 | 26280
    performance IQ 58 | 26280
    verbal IQ 71 | 26280
    full gross-motor development | 50400
    continence sphincter control | 50400
    complete sentences | 50400
    improved reasoning | 50400
    performance IQ 64 | 61200
    mild mental retardation | 61200
    impulsive personality | 61200
    easily distracted | 61200
    