66 years old | 0
female | 0
admitted to the hospital | 0
chills | -48
fever | -48
pharynx pain | -48
chest tightness | -48
headache | -48
no cough | -48
no sputum | -48
no wheezing | -48
no dysphagia | -48
no hoarseness | -48
no weight loss | -48
no edema of lower extremities | -48
diagnosed with acute upper respiratory tract infection | 0
type 2 diabetes mellitus | -0
no history of respiratory disease | -0
no history of trauma | -0
no history of foreign-body ingestion | -0
temperature 39.1 °C | 0
pulse rate 125 beats per min | 0
respiratory rate 24 breaths/min | 0
blood pressure 110/68 mmHg | 0
no clubbing | 0
no icterus | 0
no generalized lymphadenopathy | 0
leukocyte count 9900/μL | 0
segmented neutrophils 88% | 0
elevated erythrocyte sedimentation rate 79 mm/h | 0
increased C-reactive protein 42.9 mg/dL | 0
CT of the lung normal | 0
MRI of the brain normal | 0
ultrasonic study of the heart and liver normal | 0
treatment with intravenous amoxicillin | 24
treatment with levofloxacin | 24
treatment with ribavirin | 24
body temperature 39.0 °C | 48
preliminary result of blood culture gram-positive cocci | 48
antibiotics changed to teicoplanin | 48
antibiotics changed to moxifloxacin | 48
dyspnea worsened | 120
respiratory and cardiac arrest | 120
lost consciousness | 120
systemic cyanosis | 120
arterial blood gas analysis | 120
cardiopulmonary resuscitation | 120
intravenous epinephrine | 120
emergency tracheal intubation | 120
simple breathing bag | 120
transferred to the Respiratory Intensive Care Unit | 120
penicillin-sensitive Kocuria kristinae isolated from blood samples | 120
diagnosis of sepsis | 120
intravenous antibiotic therapy changed to vancomycin | 120
intravenous antibiotic therapy changed to piperacillin-tazobactam | 120
mechanical ventilation withdrawn | 144
extubated | 144
bedside chest radiograph normal | 144
evaluation of arterial blood gas analysis met the weaning criteria | 144
dyspnea again | 192
heart and respiratory rates slowed | 192
lost consciousness again | 192
arterial blood gas analysis | 192
emergency tracheal intubation | 192
mechanical ventilation | 192
acute airway obstruction | 192
lumbar puncture | 192
analysis of cerebrospinal fluid | 192
high leukocyte count | 192
lymphocytes 75% | 192
no Cryptococcus | 192
increased protein level | 192
cerebrospinal fluid culture negative | 192
CT scan of the neck | 216
soft tissue swelling of the nasopharyngeal and oropharyngeal wall | 216
occlusion of the nasopharyngeal and oropharyngeal cavity | 216
bedside flexible bronchoscopy | 216
edema of the nasopharynx and oropharynx mucosa | 216
MRI | 312
obvious soft tissue swelling and thickening in the anterior region of the neck | 312
stenosis of the nasopharynx, oropharynx, and upper airway | 312
diagnosis of RPA | 312
incision and drainage of the RPA | 336
histopathology of surgical specimens | 336
inflammatory necrosis with granulation tissue | 336
culture of pus negative | 336
MRI demonstrated stenosis of the upper airway alleviated after surgery | 336
discharged from hospital | 504
asymptomatic | 504
no recurrence of RPA | 504