32 years old | 0
male | 0
white | 0
mediastinal lymphoma | 0
EPOCH-R | 0
etoposide | 0
vincristine | 0
adriamycin | 0
cyclophosphamide | 0
rituximab | 0
oral prednisone | 0
Neulasta | 0
dyspnea | -168
worsening dyspnea | -168
CLS suspected | -168
third cycle without Neulasta | -96
sudden-onset dyspnea | 0
tachypnea | 0
tachycardia | 0
hypotension | 0
diffuse interstitial infiltrate | 0
fluid bolus | 0
broad-spectrum antibiotics | 0
meropenem | 0
vancomycin | 0
intubated | 24
pressor support | 24
recovered | 48
extubated | 48
weaned off pressor support | 48
moved out of ICU | 48
bilateral pleural effusion | 72
consolidation | 72
broad-spectrum antibiotic therapy | 72
ventilator-associated pneumonia | 72
Staphylococcus epidermidis growth | 72
positron emission tomography/CT scan | 168
excellent remission of lymphoma | 168
resolution of abnormalities | 168
CHOP | 168
cyclophosphamide | 168
vincristine | 168
adriamycin | 168
prednisone | 168
leukocytosis | 0
thrombocytosis | 0
elevated hematocrit | 0
normal BUN | 0
normal creatinine | 0
normal electrolytes | 0
normal liver enzymes | 0
low serum albumin | 0
elevated lactic acid | 0
elevated procalcitonin | 0
exudative pleural effusion | 0
elevated leukocyte count | 0
albumin 4.2 g/dL | -168
hematocrit 36.2% | -168
albumin 4.1 g/dL | -168
hematocrit 37.6% | -168
albumin 3.8 g/dL | -168
hematocrit 35.9% | -168
albumin 3.7 g/dL | -168
hematocrit 37.7% | -168
albumin 3.9 g/dL | -24
hematocrit 34.6% | -24
albumin 3.3 g/dL | 0
hematocrit 49.9% | 0
albumin 3.3 g/dL | 24
hematocrit 51.4% | 24
albumin 2.3 g/dL | 48
hematocrit 44.0% | 48
albumin 2.6 g/dL | 72
hematocrit 44.9% | 72
albumin 3.1 g/dL | 96
hematocrit 31.9% | 96
hematocrit 25.5% | 120
hematocrit 28.1% | 144
albumin 4.0 g/dL | 168
hematocrit 33.9% | 168
albumin 4.5 g/dL | 216
hematocrit 36.7% | 216
albumin 4.0 g/dL | 264
hematocrit 38.8% | 264
albumin 4.0 g/dL | 312
hematocrit 41.2% | 312