85 years old | 0
male | 0
farmer | 0
active lifestyle | 0
admitted to the geriatric medicine unit | 0
transferred to the rehabilitation unit | 0
atrial fibrillation | -672
benign prostatic hypertrophy | -672
trismus | -336
hypertonia | -336
injured his leg | -336
admitted to a local hospital | -336
treated with immunoglobulins | -336
tetanus vaccination | -336
metronidazole | -336
transferred to the intensive care unit | -336
tracheostomy | -336
mechanical ventilation | -336
vasoactive support | -336
respiratory failure | -336
seizures | -336
baclofen | -336
midazolam | -336
diazepam | -336
electroencephalography | -336
slow cerebral activity | -336
opacity on chest radiography | -336
peripheral leukocytosis | -336
ventilator-associated pneumonia | -336
blood cultures | -336
tracheal secretion samples | -336
Klebsiella pneumoniae | -336
methicillin-sensitive Staphylococcus aureus | -336
piperacillin-tazobactam | -336
transferred to a geriatric unit | -336
coma | -336
breathed spontaneously | -336
supplemental oxygen | -336
tracheal cannula | -336
antibiotic therapy | -336
linezolid | -336
meropenem | -336
septic shock | -336
cholestasis | -336
acute edematous pancreatitis | -336
endoscopic treatment | -336
urinary tract infection | -336
multidrug-resistant organisms | -336
K. pneumoniae | -336
Acinetobacter baumannii | -336
Enterococcus faecalis | -336
colistin | -336
amoxicillin-clavulanate | -336
MDRO isolation | -336
tracheal supplemental oxygen | -336
bladder catheter | -336
pressure ulcers | -336
sarcopenic | -336
low handgrip strength | -336
appendicular skeletal mass | -336
rehabilitative evaluations | -336
Clostridioides difficile infection | -336
oral vancomycin | -336
atrial fibrillation | -336
third-degree atrioventricular block | -336
heart rate | -336
single-chamber pacemaker implantation | -336
hyperkinetic delirium | -336
Pseudomonas aeruginosa bloodstream infection | -336
ceftazidime-avibactam | -336
amikacin | -336
SARS-CoV-2 | -336
remdesivir | -336
droplet isolation | -336
second recurrence of C. difficile | -336
fidaxomicin | -336
bloodstream infection | -336
Candida parapsilosis | -336
MSSA | -336
Candida tropicalis | -336
intravenous catheter | -336
caspofungin | -336
cefazolin | -336
bloodstream infection | -336
P. aeruginosa | -336
piperacillin-tazobactam | -336
aztreonam | -336
ceftazidime-avibactam | -336
cefepime | -336
tracheostomy closure | -336
ENT specialist | -336
pulmonologist | -336
nutritional supplementation | -336
malnutrition | -336
sarcopenia | -336
motor rehabilitation | -336
respiratory reconditioning | -336
postural transition | -336
aided transfers | -336
axial stability | -336
balance improvement | -336
standing position | -336
breath-movement coordination | -336
thoracic expansion | -336
girdle opening | -336
inhalation-exhalation | -336
wheelchairs | -336
walkers | -336
mobility deficit | -336
safe postural transitions | -336
rehabilitation | -336
ENT | -336
geriatric follow-up | -336
discharged | 720