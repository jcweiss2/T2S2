63 years old | 0
female | 0
168 cm height | 0
53 kg weight | 0
papillary thyroid carcinoma | -9720
resection | -9720
radiotherapy | -9720
stenosis of the esophagus | -8760
repeated aspiration | -8760
respiratory insufficiency | -8760
pneumonia | -8760
purulent pleurisy | -8760
pleurectomy | -8760
restrictive ventilation pattern | -8760
recurrent nerve palsy | -8760
percutaneous endoscopic gastrostomy | -8760
tracheostoma | -8760
home ventilation | -8760
secondary depression | -8760
mobility decreased | -8760
stopped talking | -8760
mandible nearly fixed | -8760
could not open mouth | -8760
left axis vertebralis stented | -4380
stenosis of the internal axis carotis | -4380
arterial hypertension | -4380
secondary lactase deficiency | -4380
esophageal stenosis dilated | -120
fistula between esophagus and tracheal membrane | -120
referred to University of Erlangen | -120
decreasing general condition | -120
examined by chiefs and consultants | -120
deemed too unstable for open surgery | -120
inability to open mouth | -120
recurrent nerve palsy | -120
minimal invasive orthograde approach impossible | -120
referred to hospital | 0
suffering from pneumonia | 0
4-multiresistente gramnegative Pseudomonas aeruginosa | 0
veno-venous extracorporeal membrane oxygenation | 0
partial thromboplastin time 60 seconds | 0
preseptic status | 0
ventilated through tracheostoma | 0
low ventilation forces | 0
thoracic computed tomography | 24
big fistula of tracheal membrane | 24
tracheal cannula ended shortly beneath lower limit of mediastinal fistula | 24
decision to try endobronchial stenting | 48
plan to close fistula with pedicled omentum majus replacement | 48
abutment and secured continuous airway replacement | 48
procedure performed | 72
vv-ECMO partly ineffective | 72
rising septical issues | 72
high volume input of physiological saline | 72
oral approach only allowed small flexible bronchoscope | 72
approach for upper part of trachea had to be performed through percutaneous tracheostoma | 72
retrograde stenting | 72
Dumon and one-hybrid self expandable metalic y-stent | 72
Freitag stent | 72
mandatory additional ventilation | 72
nasal jet catheter | 72
double-lumen endotracheal tube exchange catheter | 72
ventilation line introduced orally or through tracheostoma | 72
placed distally below main carina | 72
successful retrograde stenting performed in four steps | 72
Step I | 72
regular bronchoscopes | 72
jagwires | 72
jet-catheters | 72
DLETs | 72
manually compressed y of FS pushed downward | 72
main carina | 72
Step II | 96
frontal surface of stent cut | 96
new stoma for regular tracheal cannula created | 96
lower new edge of stoma fixed subcutaneously | 96
Step III | 120
jagwire introduced through mouth into trachea | 120
running out of new FS stoma | 120
leaving dorsal membrane of cut FS behind | 120
soft-tip stiff DLET introduced | 120
dragged out of new stoma of cut FS | 120
distal jagwire introduced into oral orifice of FS | 120
bended up curve | 120
FS flipped with upper part over soft-tip stiff DLET | 120
into upper third of trachea | 120
whole fistula bridged by FS | 120
up to level of vocal cords | 120
upper edge of new FS stoma fixed subcutaneously | 120
Step IV | 144
regular tracheal cannula introduced | 144
for ventilation | 144
lungs not aerated | 144
vv-ECMO running | 144
high volume input of physiological saline | 144
spontaneous breathing work increased | 168
vv-ECMO support reduced | 168
lungs became re-aerated | 168
patient woke up | 168
could communicate with family | 168
by writing | 168
by eyes | 168
infections continued | 168
severe | 168
spontaneous work of breathing never exceeded tidal ventilation of 170 mL per breath | 168
reduction of intravenous saline injection limited | 168
mandatory but reduced vv-ECMO support | 168
patient and family decided to reduce vv-ECMO support | 240
with risk of death | 240
patient died | 360
pulmonary infection | 360