23 years old | 0
male | 0
admitted in the ICU | 0
sudden onset of pain abdomen | -72
respiratory distress | -72
intestinal perforation | 0
blood pressure 110/60 mm Hg | 0
pulse 86 beats/min | 0
respiratory rate 22 breaths/min | 0
SpO2 99% on room air | 0
afebrile | 0
urgent laparotomy | 0
asymptomatic for next 2 days after surgery | 72
blood pressure fall up to 84 mmHg (systolic) | 72
CVC in right subclavian vein | 72
administration of drugs | 72
administration of intravenous fluid | 72
right subclavian vein cannulated | 72
7.5F triple lumen CVP catheter (Edward) | 72
standard Seldinger technique | 72
USG guidance | 72
aseptic precautions | 72
lateral approach | 72
needle inserted longitudinally | 72
guide wire confirmed well in position | 72
guide wire movement free at insertion | 72
guide wire movement free during removal | 72
all channels of CVC aspirated for blood | 72
CVC fixed at 15 cm | 72
CVP waveform appeared dampened | 72
CVP waveform not improved | 72
chest radiograph performed | 72
catheter migrated to left subclavian vein | 72
right subclavian CVC removed | 72
CVC reintroduced under color Doppler guidance | 72
modified Seldinger technique | 72
guide wire traced much beyond subclavian vein | 72
repeat chest radiograph confirmed correct placement | 72
normal CVP tracing | 72
