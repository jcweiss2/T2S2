22 years old | 0
male | 0
white | 0
admitted to the hospital | 0
gastroesophageal reflux disease | -8760
past cholecystectomy | -8760
intermittent esophageal dysphagia | -8760
omeprazole | -8760
EGD evaluation | 0
esophageal dysphagia | 0
procedural sedation | 0
propofol | 0
intravenous propofol | 0
total of 150 mg of intravenous propofol | 0
mild esophageal stricture | 0
esophagogastric junction | 0
balloon dilator | 0
dilated to 20 mm | 0
esophageal mucosal changes | 0
ringed esophagus | 0
feline appearance | 0
longitudinal furrows | 0
middle and lower third of the esophagus | 0
eosinophilic esophagitis | 0
biopsies | 0
upper GI tract | 0
unremarkable | 0
tolerated the procedure | 0
anesthesia well | 0
sudden onset of severe epigastric pain | 1.5
emesis | 1.5
after a meal | 1.5
emergency department | 2
elevation of lipase | 2
14,000 U/L | 2
total leukocyte count | 2
30,000 cells per liter | 2
no eosinophilia | 2
high neutrophils | 2
normal lymphocyte counts | 2
triglycerides level | 2
79 mg/dL | 2
abdominal and pelvic computed tomography | 2
peripancreatic fluid | 2
no evidence of cyst | 2
abscess | 2
necrosis | 2
general medical floor | 2
intravenous fluid hydration | 2
pain control | 4
intensive care unit | 4
deterioration | 4
hypoxia | 4
hemodynamic instability | 4
acute hypoxic respiratory failure | 6
acute respiratory distress syndrome | 6
intubation | 6
mechanical ventilation | 6
septic shock | 8
vasopressor support | 8
broad-spectrum antibacterial | 8
antifungal agents | 8
pleural effusion | 10
thoracentesis | 10
chest tube placement | 10
acute kidney injury | 12
repeat abdominal and pelvic computed tomography | 12
pancreatic necrosis | 12
extensive peripancreatic fluid | 12
post-pararenal space | 12
retroperitoneal fluid collection | 12
percutaneous drain placement | 14
pancreatic necrosectomy | 16
ischemic colitis | 18
shock | 18
subtotal colectomy | 20
prolonged course of hospitalization | 24
ICU setting | 24
multiple medical and surgical specialties | 24
rehab facility | 168
doing well | 168
cholecystectomy | -720
gallstone pancreatitis | -720
pancreatic divisum | -720
alcohol use | -720
infectious pathogens | -720
nasopharyngeal respiratory viral polymerase chain reaction | -720
human rhinovirus | -720
serum testing | -720
viral cause | -720
autoimmune etiology | -720
immunoglobulin levels | -720
normal serum triglyceride level | -720
elevated lipase level | -720
total white count | -720
omeprazole | -720
previous trauma | -720
exposure to drugs | -720
toxins | -720
cystic fibrosis | -720
myotonic dystrophy | -720
vascular disease | -720
vasculitis | -720
drug allergies | -720
environmental allergies | -720
propofol administration | 0
acute pancreatitis | 2
multiorgan failure | 12
idiosyncratic reaction | 12
pancreatitis awareness | 168
life-threatening adverse event | 168
propofol sedation | 168
abdominal pain | 168
periprocedural air insufflation | 168
cost | 168
risks | 168
benefits | 168
propofol-induced deep sedation | 168
benzodiazepines | 168
opioid-induced conscious sedation | 168
GI endoscopic procedures | 168
alternative sedatives | 168