16 years old|0
male|0
presented with fever|0
fatigue|0
scleral icterus|0
jaundice|0
dark urine|0
right abdominal pain|0
right shoulder pain|0
diagnosed with ulcerative colitis (UC) 2 years prior|-17520
no significant medical history|-17520
corticosteroid-dependent course|-17520
experienced several acute exacerbations|-17520
escalation of therapy from aminosalicylates to immunomodulators|-17520
completed a three-dose induction course of infliximab|-720
latest UC flare| -504
colonoscopy showing pancolitis| -504
treated with IV corticosteroids| -504
another dose of infliximab| -504
improved| -504
alkaline phosphatase (ALP) at that time was 88 U/L| -504
leukocytosis (16,000/µL)|0
anemia (6.9 g/dL)|0
thrombocytopenia (53,000/µL)|0
transaminitis (AST 570 U/L, ALT 296 U/L)|0
highly elevated ALP (426 U/L)|0
hyperbilirubinemia (3.1 mg/dL)|0
CRP 20.4 mg/dL|0
CT showed multiple multi-loculated abscesses in the right hepatic lobe|0
largest abscess in segment 7 measured approximately 10 cm|0
presence of gas|0
extensive intrahepatic thrombosis of the right portal vein|0
splenomegaly|0
bilateral pleural effusions|0
diffuse colonic wall thickening|0
no megacolon|0
no free intraperitoneal air|0
no other signs of perforation|0
appendix was normal|0
abscess drained by interventional radiology|0
cultures positive for Peptostreptococci|0
cultures positive for skin flora (Gram-positive cocci in clusters and pairs)|0
cultures positive for Escherichia coli|0
acid-fast bacilli stain negative|0
bacteremic with Streptococcus viridans|0
bacteremic with E. coli|0
surgical drainage required due to abscess size|0
repeat wound cultures showed same organisms|0
developed septic shock post-operatively|24
required ICU management|24
antimicrobial therapy changed from vancomycin and meropenem to ceftriaxone and metronidazole|24
repeat CT 10 days after initial study|240
continued improvement in abscess size|240
repeat CT 20 days after initial study|480
therapy de-escalated to oral amoxicillin-clavulanate|480
completed 2-week course of amoxicillin-clavulanate|480
symptomatically improved|480
CRP down-trending|480
discharged|480
amino acid-based formula via nasogastric tube|480
advancing oral diet|480
liver loculations improved|2016
liver loculations resolved on ultrasonography|2016
normalization of liver enzymes|2016
normalization of inflammatory markers|2016
no UC therapy other than exclusive enteral nutrition|480
not consistently compliant with enteral nutrition|480
remained without signs or symptoms of UC|480
developed severe pancolitis 11 months from admission| -720
underwent total colectomy| -720
surgical gross pathology showed moderately to severely active chronic pancolitis| -720
mural abscesses| -720
mucosa diffusely tan-red and hyperemic| -720
scattered diffuse areas of ulceration| -720
nodularity| -720
pseudopolyps| -720
ileum without significant abnormalities| -720
appendix without significant abnormalities| -720
no evidence of ischemia| -720
no evidence of dysplasia| -720
no granulomas| -720
findings compatible with UC| -720
