13 years old | 0
male | 0
admitted to the hospital | 0
uncontrolled bleeding at the operation site of the right thenar muscle | 0
swelling of the right thenar muscle | -4032
fall | -4032
hematoma | -4032
no treatment | -4032
no improvement | -4032
excision of the lesion | -2016
no bleeding tendency | -2016
normal coagulation screening tests | -2016
two additional operations | -1440
bleeding continued | -1440
pathologic finding suggested malignancy | -1440
transferred to our hospital | 0
poor general state | 0
pallor | 0
weakness | 0
bruising at the intravenous site | 0
purpura on the operation site | 0
continuous bleeding | 0
lymph node in the right axillary area | 0
hepatosplenomegaly | 0
decreased platelet levels | 0
decreased hemoglobin levels | 0
features suggestive of DIC | 0
white blood cell count 9900 /µL | 0
hemoglobin 4.8 g/dL | 0
platelets 28000 /µL | 0
prothrombin time 1.47 INR | 0
activated partial thromboplastin time 45.4 sec | 0
fibrinogen 87 mg/dL | 0
fibrin/fibrinogen degeneration product 656.4 µg/mL | 0
D-dimer 16.17 mg/L | 0
normal coagulation factors II, VII, IX, fibrinogen, von Willebrand factor | 0
factor V 30% | 0
factor VIII 40% | 0
hypermetabolic lesions in the right thenar muscle | 0
hypermetabolic lesions in the right axillary space | 0
post-operative inflammation in the right thenar muscle | 0
metastatic lymphadenopathy in the right axillary space | 0
massive bleeding worsened | 72
gross hematuria | 72
alveolar rhabdomyosarcoma diagnosis | 96
transferred to intensive care unit | 96
VAC chemotherapy administered | 96
repeated transfusions | 96
synthetic protease inhibitor | 96
antithrombin-III substitution | 96
massive epistaxis | 240
hematemesis | 240
transfusions of RBCs, PCs, FFP, cryoprecipitate | 240
cauterization | 240
improvement in DIC laboratory findings | 336
BM section biopsy | 336
axillary LN biopsy | 336
rhabdomyosarcoma involvement in BM | 336
rhabdomyosarcoma involvement in axillary LN | 336
blood transfusions total 311 units | 480
discharged | 672
combination chemotherapy every 3 weeks | 672
decrease in right axillary LN size | 1512
BM disappearance of rhabdomyosarcoma | 3528
nodule in the right forearm | 4536
biopsy revealing alveolar rhabdomyosarcoma | 4536
salvage chemotherapy | 4536
palliative radiation therapy | 4536
disease progression to liver and brain | 4536
death | 4536
