49 years old | 0
female | 0
low back pain | -72
right leg pain | -72
intractable cough | -504
productive green sputum | -504
no chest pain | -504
no shortness of breath | -504
no fevers | -504
no paraesthesia | -504
no weakness of lower limbs | -504
no urinary symptoms | -504
no bowel symptoms | -504
oral cephalexin | -504
hypertension | -504
chronic low-back pain | -504
smokes 20 cigarettes per day | -504
15 pack year smoking history | -504
no respiratory distress | 0
normal vital signs | 0
bronchial breath sounds in right lung mid to lower zones | 0
coarse crepitations | 0
soft abdomen | 0
non-tender abdomen | 0
antalgic gait | 0
normal sensation in lower limbs | 0
normal power in lower limbs | 0
normal reflexes in lower limbs | 0
white cells 19.2 × 10^9/L | 0
neutrophilia | 0
chest radiograph obscured right heart border | 0
infective consolidation of right middle lobe | 0
community acquired pneumonia | 0
low back pain precipitated by cough | 0
benzyl penicillin | 0
doxycycline | 0
analgesics | 0
admitted under medical team | 0
medical emergency team review | 48
hypotension | 48
presyncope | 48
new onset epigastric pain | 48
new onset chest pain | 48
back pain | 48
pale appearance | 48
heart rate 78 bpm | 48
blood pressure 66/38 mmHg | 48
unchanged chest examination | 48
soft abdomen | 48
haemoglobin drop from 115 g/L to 77 g/L | 48
shock | 48
haemorrhagic shock | 48
suspected aortic dissection | 48
suspected aortic aneurysm rupture | 48
suspected haemorrhage from peptic ulcer | 48
differential diagnosis sepsis | 48
differential diagnosis pulmonary embolism | 48
bilateral large bore intravenous access | 48
fluid resuscitation | 48
red blood cell transfusion | 48
intravenous ceftriaxone | 48
moved to high dependency unit | 48
surgical review | 48
haemodynamically responsive to resuscitation | 48
urgent CT scan with contrast | 48
ruptured spleen | 48
large perisplenic haematoma | 48
large haemoperitoneum | 48
active bleeding in portal venous sequences | 48
bilateral pulmonary consolidation | 48
no pulmonary embolism | 48
splenic rupture secondary to repeated coughing | 48
emergency laparotomy | 48
vertical midline upper abdominal laparotomy | 48
large haematoma removed | 48
ongoing bleeding | 48
spleen nearly avulsed | 48
incomplete splenophrenic ligament | 48
partial rupture of spleen under ligament | 48
absent splenonephric ligament | 48
mobile spleen with medial lie | 48
Ligasure division of short gastric arteries | 48
Ligasure division of splenic arteries | 48
Ligasure division of splenic veins | 48
spleen removed | 48
satisfactory haemostasis | 48
splenic artery oversewn | 48
Blake’s drain placed in left subdiaphragmatic space | 48
abdomen closed | 48
transfusion of six units red blood cells | 48
transfusion of two units fresh frozen plasma | 48
transfer to intensive care unit | 48
extubated | 144
discharged home | 192
pneumonia resolved | 192
surgical wounds healing well | 192
resumed nearly all activities | 192
persisting back pain | 192
immunized against Pneumococcus | 192
immunized against Meningococcus | 192
immunized against Haemophilus influenza type b | 192
declined trivalent influenza vaccine | 192
prophylactic amoxicillin | 192
added to splenectomy register | 192
uncomplicated recovery | 336
investigations negative for influenza A | 192
investigations negative for influenza B | 192
investigations negative for RSV | 192
negative respiratory virus PCR | 192
negative sputum microscopy | 192
negative sputum culture | 192
negative legionella urinary antigen | 192
negative pneumococcus urinary antigen | 192
negative chlamydia serology | 192
negative EBV serology | 192
negative legionella serology | 192
spleen histopathology | 192
preserved pulp architecture | 192
no evidence of malignancy | 192
atraumatic splenic rupture | 48
community acquired pneumonia | -504
