35 years old | 0
woman | 0
gravida 3 | 0
para 0 | 0
adenomyosis | 0
infertility | 0
IVF-ET | 0
amnion cavity acrinol-induced labor | 0
menstrual period | 0
slow-release gonadotropin-releasing hormone agonist | 0
HP-HMG 225 IU/day | 0
oocyte retrieval | 0
vaginal progesterone 0.6 g/day | 0
triplet (monozygotic twin and singleton) | 35
ultrasound-guided selective pregnancy reduction | 35
fetal nuchal translucency 4.6 mm | 13*7*24
abnormal forearms and wrist joints | 13*7*24
single umbilical artery | 13*7*24
hospitalization for genetic testing | 18*7*24
umbilical cord blood sampling attempted | 18*7*24
rivanol injection into amniotic cavity attempted | 18*7*24
failure due to fetal position and oligohydramnios | 18*7*24
fever (highest 40°C) | (18*7*24) + 36
right upper quadrant tenderness | (18*7*24) + 36
antibiotic administration | (18*7*24) + 36
carboprost administration | (18*7*24) + 36
postpartum hemorrhage | (18*7*24) + 36 + delivery time
febrile | (18*7*24) + 36 + delivery time
hypotension | (18*7*24) + 36 + delivery time
HBG 84 g/L | (18*7*24) + 36 + delivery time
white blood cell 14.61 × 10^9/L | (18*7*24) + 36 + delivery time
platelet 81 × 10^9/L | (18*7*24) + 36 + delivery time
D-D 135,337 ng/ml | (18*7*24) + 36 + delivery time
blood pressure 79/41 mmHg | (18*7*24) + 36 + delivery time
septic shock | (18*7*24) + 36 + delivery time
DIC | (18*7*24) + 36 + delivery time
hemorrhagic shock | (18*7*24) + 36 + delivery time
transfer to ICU | (18*7*24) + 36 + delivery time
total abdominal hysterectomy | (18*7*24) + 36 + delivery time
endometritis | (18*7*24) + 36 + delivery time
uterus cellulitis | (18*7*24) + 36 + delivery time
antibiotics continuation | (18*7*24) + 36 + delivery time
abdominal debridement | (18*7*24) + 36 + delivery time + recovery time
suturing | (18*7*24) + 36 + delivery time + recovery time
discharge | (18*7*24) + 36 + delivery time + recovery time + 16*24
no postoperative problems | (18*7*24) + 36 + delivery time + recovery time + 16*24
Escherichia coli in vaginal discharge | (18*7*24) + 36 + delivery time
Escherichia coli in uterine discharge | (18*7*24) + 36 + delivery time
missed abortion history | 0
curettage history | 0
spontaneous abortion history (two-time) | 0
PID risk | 0
tubo8-ovarian abscess risk | 0
adenomyosis-related risks | 0
repeated pelvic operations | 0
transvaginal oocyte retrieval | 0
transvaginal selective pregnancy reduction | 0
transabdominal umbilical cord blood sampling | 0
amniotic cavity rivanol injection | 0
failed amniocentesis | 0
adenomyosis-related risks |>
