10 years old | 0
male | 0
admitted to the hospital | 0
papulovesicular skin lesions | -240
fever | -96
altered sensorium | -24
malena | -24
respiratory rate 32/min | 0
heart rate 173/min | 0
capillary refill time 4 seconds | 0
blood pressure 90/50 mmHg | 0
SpO2 93% | 0
poor peripheral pulses | 0
severe pallor | 0
crusted pus discharging lesions | 0
Glasgow Coma Scale score of E4M4V4 | 0
generalized hypotonia | 0
elicitable deep tendon reflexes | 0
flexor plantar reflex | 0
no cranial nerve palsies | 0
absent meningeal signs | 0
resuscitated with normal saline boluses | 0
intravenous infusion of adrenaline | 0
intravenous infusion of noradrenaline | 0
intravenous infusion of vasopressin | 0
intravenous infusion of dobutamine | 0
PRBCs transfusion | 0
intravenous antibiotics | 0
mechanical ventilation | 0
shifted to pediatric intensive care unit | 6
developed acute kidney injury | 48
started on peritoneal dialysis | 48
deranged liver function tests | 48
inotropes tapered and stopped | 96
extubated | 144
severe anemia | 168
hypotensive shock | 168
multiple episodes of massive malena | 168
resuscitated with fluid boluses | 168
PRBCs transfusions | 168
vasoactive drugs | 168
UGI endoscopy | 168
bleeding lesion in the first part of duodenum | 168
computed tomography angiography | 168
GDA pseudoaneurysm | 168
digital subtraction angiography | 168
coil embolization | 168
transiently controlled bleeding | 168
massive episodes of malena | 180
second endovascular cyanoacrylate glue embolization | 192
life-threatening UGI bleeding | 192
received massive PRBC transfusion | 192
received fresh frozen plasma | 192
received platelet concentrates | 192
amylase levels normal | 192
ANA normal | 192
ANCA normal | 192
HBsAg normal | 192
HCV normal | 192
HIV normal | 192
laparotomy | 216
duodenostomy | 216
ligation of GDA aneurysm | 216
UGI bleeding stopped | 216
inotropes tapered | 216
respiratory support tapered | 216
extubated | 264
developed critical illness neuromyopathy | 264
discharged | 600
follow-up | 4320
ambulatory | 4320
no recurrence of symptoms | 4320