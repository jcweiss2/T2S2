19 years old | 0
male | 0
army officer | 0
fever | -120
arthralgia | -120
myalgia | -120
headache | -120
productive cough | -120
yellowish sputum | -120
chest heaviness | -120
dyspnea | -120
diarrhea | -120
reduced oral intake | -120
dehydrated | 0
cold peripheries | 0
febrile | 0
hypotensive | 0
tachycardic | 0
tachypnoeic | 0
oxygen saturation 75–80% | 0
coarse crepitation | 0
tenderness at epigastric region | 0
palpable liver | 0
haemoglobin 11.3 g/dL | 0
low white blood cell | 0
neutrophil predominance | 0
platelet count 80 × 10^6/L | 0
C-reactive protein 28.28 mg/dL | 0
acute kidney injury | 0
serum sodium 137 mmol/L | 0
potassium 3.7 mmol/L | 0
urea 14 mmol/L | 0
creatinine 206 μmol/L | 0
liver function tests normal | 0
serum albumin 22 g/dL | 0
creatinine kinase 351 IU/L | 0
arterial blood gases | 0
pH 7.378 | 0
pCO2 37 mmHg | 0
pO2 52.7 mmHg | 0
O2 saturation 89% | 0
HCO3 21.7 mmol/L | 0
Dengue NS-1 Antigen negative | 0
IgG and IgM antibody negative | 0
chest radiograph | 0
consolidation of right upper lobe | 0
left lower lobes | 0
diagnosis of severe community acquired pneumonia | 0
acute kidney injury | 0
resuscitated with normal saline | 0
non-invasive ventilation | 0
inotropic support | 0
intravenous ceftriaxone | 0
azithromycin | 0
intubation | 12
mechanical ventilation | 12
persistent type 2 respiratory failure | 12
bronchoscopy | 48
copious amount of haemoserous | 48
greenish secretion | 48
repeated chest radiograph | 48
worsening consolidation | 48
early changes of abscess formation | 48
intravenous meropenem | 48
cloxacillin | 48
antiviral oseltamivir | 48
continuous venous-venous haemofiltration | 48
severe metabolic acidosis | 48
oliguric acute kidney injury | 48
persistent spiking of temperature | 48
worsening of septic parameters | 48
refractory hypotension | 48
multiple inotropic agents | 48
deteriorated further | 48
blood cultures negative | 72
atypical bacterial and Leptospiral serologies negative | 72
Hepatitis B/C and HIV serologies undetected | 72
Respiratory viruses screening negative | 72
tracheal aspiration positive for MDR Acinetobacter baumannii | 72
bronchoalveolar lavage positive for MDR Acinetobacter baumannii | 72
MDR Acinetobacter baumannii susceptible only to polymyxin B | 72
minimum inhibitory concentration 0.5 μg/ml | 72
MDR Acinetobacter baumannii resistant to penicillin group | 72
ampicillin/sulbactam | 72
third generation cephalosporins | 72
fluoroquinolone | 72
carbapenem group | 72
PCR for carbapenemases genes NDM, OXA-23, OXA 24 or OXA-58 not performed | 72
died | 72