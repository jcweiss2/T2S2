48 years old| 0
male| 0
sudden fever| 0
tachycardia| 0
hypotension| 0
right neck swelling| 0
right neck redness| 0
right neck tenderness| 0
right neck warmth| 0
headache| 0
coma| -4
emergency decompressive craniotomy| 0
CVC insertion through right subclavian vein| 0
absence of ultrasound assistance for CVC insertion| 0
absence of chest X-ray for CVC tip assessment| 0
transfer to ICU| 48
septic shock| 0
leukocytosis| 0
elevated C-reactive protein| 0
elevated procalcitonin| 0
elevated alanine aminotransferase| 0
elevated aspartate aminotransferase| 0
pH 7.30| 0
PaCO2 33 mmHg| 0
PaO2 108 mmHg| 0
lactate 3.8 mmol/L| 0
HCO3- 16.8 mmol/L| 0
thrombosis in right internal jugular vein| 0
CVC misplaced into right internal jugular vein| 0
gas bubbles surrounding CVC| 0
hyperechoic lines with dirty shadowing| 0
comet-tail artifacts| 0
septic emphysematous thrombophlebitis diagnosis| 0
CVC removal| 0
peripheral venous blood culture| 0
CVC blood culture| 0
fluid resuscitation| 0
intravenous noradrenaline| 0
vancomycin administration| 0
imipenem-cilastatin administration| 0
low-molecular-weight heparin administration| 0
methicillin-resistant Staphylococcus cohnii isolation| 96
redness subsiding| 168
swelling subsiding| 168
left limb weakness due to stroke| 168
transfer to general ward| 168
discharge| 240
right internal jugular vein thrombus organization| 720
stable blood flow| 720
