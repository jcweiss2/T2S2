57 years old | 0
female | 0
severe rheumatic mitral stenosis | -672
severe aortic stenosis | -672
severe tricuspid regurgitation | -672
chronic atrial fibrillation | -672
hypertension | -672
pacemaker placement for sick sinus syndrome | -672
warfarin | -672
no history of bleeding | -672
implantation of a 25 mm mitral and a 19 mm aortic On-X valve | 0
de Vega tricuspid annuloplasty | 0
Maze procedure | 0
cardiopulmonary bypass | 0
aortic cross-clamp | 0
intubated | 0
high infusion rates of inotropic and vasopressor agents | 0
epinephrine | 0
norepinephrine | 0
vasopressin | 0
milrinone | 0
severely hypocoagulable | 0
thrombocytopenia | 0
hypofibrinogenemia | 0
elevated international normalized ratio (INR) | 0
subcutaneous heparin 5000 IU every 12 h | 192
prophylaxis against deep vein thrombosis | 192
removal of the epicardial pacing wires | 216
pericardial tamponade | 216
emergent opening of the sternum | 216
progressive worsening of pulmonary hypertension | 216
severe right heart failure | 216
biventricular failure | 216
intra-aortic balloon pump | 216
inhalational epoprostenol therapy | 216
renal failure | 216
continuous renal replacement therapy | 216
consumptive thrombocytopenia | 216
thrombocytopathia | 216
disseminated intravascular coagulopathy (DIC) | 504
multiple blood component transfusions | 504
desmopressin | 504
cryoprecipitate | 504
factor VII | 504
waxing and waning coagulopathy | 504
thrombocytopenia | 504
profuse, life-threatening bleeding | 1008
respiratory and upper gastrointestinal tracts | 1008
natural orifices | 1008
attempts to initiate anticoagulation | 1008
prophylactic doses of heparin | 1008
diagnostic bronchoscopy | 1008
upper and lower gastrointestinal endoscopies | 1008
extensive arteriovenous malformations (AVMs) | 1008
respiratory and gastrointestinal tracts | 1008
no anticoagulation | 1008
frequent transthoracic and transesophageal echocardiographic examinations | 1008
no valve thrombi | 1008
discharged to a long-term acute care facility | 4008
aspirin | 4008
warfarin | 4008
subtherapeutic INR of 1.6 | 4008
no history of thromboembolism | 4008
no further bleeding episodes | 4008
died | 4320
pulmonary aspiration | 4320
sepsis | 4320