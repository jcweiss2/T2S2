78 years old | 0
    female | 0
    myasthenia gravis (MG) | -3360
    worsening right shoulder pain | -72
    intermittent right shoulder pain | -2160
    persistent right shoulder pain | -168
    worsening severity | -168
    hypertension | -3360
    chronic kidney disease | -3360
    obesity | -3360
    proctosigmoidectomy for rectal cancer | -1464
    L3-L4 laminectomy and foraminotomy for spinal stenosis | -1752
    percutaneous spinal cord stimulator implantation | -1464
    myasthenic crisis | -1440
    dysphagia | -1440
    ptosis | -1440
    dysarthria | -1440
    intubated | -1440
    plasma exchange | -1440
    prednisone 60 mg daily | -1440
    pyridostigmine | -1440
    discharged home on pyridostigmine and prednisone | -1440
    mycophenolate | -336
    prednisone 40 mg daily | -336
    left hand and wrist purulent cellulitis | -720
    contrasted CT of left upper extremity | -720
    soft tissue ulceration | -720
    cellulitis | -720
    ill-defined intramuscular abscess | -720
    hand surgery evaluation | -720
    no surgical intervention | -720
    ceftaroline for three days | -720
    discharged home on doxycycline | -720
    trimethoprim-sulfamethoxazole (TMP-SMX) | -720
    Pneumocystis jirovecii prophylaxis | -720
    chronic steroid use | -720
    culture of purulence grew Nocardia farcinica | -720
    right shoulder pain | -72
    denied recent trauma | 0
    denied fevers | 0
    denied chills | 0
    denied sweats | 0
    resolved left-hand cellulitis | 0
    temperature of 35.8°C | 0
    heart rate of 88 bpm | 0
    respiratory rate of 18 bpm | 0
    blood pressure of 135/85 mmHg | 0
    oxygen saturation of 97% | 0
    right shoulder pain with passive range of motion | 0
    limited active range of motion | 0
    no erythema | 0
    no warmth | 0
    no swelling | 0
    white blood cell count of 14,300/µL | 0
    absolute neutrophil count of 11,930/µL | 0
    CRP of 7.63 mg/dL | 0
    ESR of 45 mm/h | 0
    unremarkable comprehensive metabolic panel | 0
    contrasted CT of right shoulder | 0
    multiloculated collections | 0
    abscesses | 0
    moderate subacromial bursa fluid | 0
    bursitis | 0
    moderate glenohumeral joint effusion | 0
    septic arthritis | 0
    bedside arthrocentesis of right shoulder synovium | 24
    synovial fluid WBC count of 107,865/µL | 24
    95% neutrophilic | 24
    1% lymphocytic | 24
    5% monocytic | 24
    no crystals | 24
    Gram stain revealed gram positive beaded bacilli | 24
    culture grew N. farcinica | 24
    CRP of 26.32 mg/dL | 24
    ESR of 71 mm/h | 24
    operative debridement of right shoulder | 48
    intra-operative purulent material | 48
    foul smell | 48
    organized loculations | 48
    chronic infection | 48
    evacuated 15 cc intra-articular purulence | 48
    evacuated 40 cc extra@-articular purulence | 48
    periscapular fluid culture grew N. farcinica | 48
    meropenem 2g twice daily | 72
    TMP-SMX 320–1600 mg three times daily | 72
    improved leukocytosis (8400/µL) | 240
    CRP 0.5 mg/dL | 240
    ESR 23 mm/h | 240
    repeat CT showed decreased fluid collections | 240
    evaluate pulmonary and intracranial disease | 240
    chest CT: bibasilar effusions | 240
    chest CT: bibasilar infiltrates | 240
    chest CT: scattered nodularity | 240
    no brain MRI due to spinal cord stimulator | 240
    head CT no intracranial abscesses | 240
    dual antimicrobial therapy with meropenem and TMP-SMX | 240
    meropenem discontinued due to resistance | 240
    continued on TMP-SMX for two months | 240
    severe thrombocytopenia | 1464
    transitioned to amoxicillin-clavulanate | 1464
    admitted for altered mentation | 1464
    failure to thrive | 1464
    transitioned to hospice care | 1464
    <|eot_id|>
    