78 years old | 0
man | 0
acute strangulated small bowel obstruction | 0
pacemaker implantation 17 years ago | -149304
advanced atrioventricular block | -149304
transient loss of pacing capture 5 months before presentation | -3600
ICU stay for septic cholangitis | -3600
pacemaker interrogation 5 months before presentation | -3600
pulse generator upgraded 2 months before presentation | -1440
battery depletion | -1440
Medtronic Advisa pacemaker programmed to DDD mode | -1440
lower rate limit 70 beats/min | -1440
previous gastrectomy for gastroduodenal ulcer | 0
type 2 diabetes mellitus | 0
medications glargine | 0
medications vildagliptin | 0
moderate distress | 0
blood pressure 176/73 mm Hg | 0
abdominal tenderness right upper quadrant | 0
electrocardiogram dual-chamber pacing and capture 70 beats/min | 0
hematocrit 32.5% | 0
anesthesia induced with remifentanil | 0
anesthesia induced with propofol | 0
muscle relaxation with rocuronium | 0
anesthesia maintained with sevoflurane | 0
anesthesia maintained with remifentanil | 0
pacemaker interrogated after anesthesia induction | 0
DDD mode lower rate 70 beats/min | 0
DDD mode upper rate 120 beats/min | 0
complete atrioventricular block | 0
slow ventricular escape rhythm | 0
ventricular pacing threshold 1.5 V | 0
ventricular pacing duration 0.4 ms | 0
ventricular pacing output 2.5 V | 0
battery impedance acceptable | 0
lead impedance acceptable | 0
sensing amplitudes acceptable | 0
capture management not enabled | 0
pacing mode changed to DOO | 0
lower rate limit 70 beats/min | 0
adhesiolysis for small bowel obstruction | 0
cholecystectomy | 0
uneventful surgery | 0
no pacing issues | 0
ultrasound-guided rectus sheath block | 0
levobupivacaine 40 mL 0.25% | 0
pacemaker reinterrogated | 0
pacemaker reprogrammed to DDD mode | 0
ventricular pacing threshold 1.25 V | 0
emergence from anesthesia uneventful | 0
extubated 30 minutes after rectus sheath block | 30
asystole confirmed post-extubation | 30
cardiopulmonary resuscitation started | 30
ventricular pacing output increased to 3.5 V | 30
ventricular pacing duration 0.4 ms | 30
stable hemodynamics achieved | 30
ventricular pacing threshold rechecked 3.0 V | 30
arterial blood gas pH 7.29 | 30
arterial blood gas Pco2 46 mm Hg | 30
arterial blood gas Po2 112 mm Hg | 30
arterial blood gas HCO3 22.5 mmol/L | 30
sodium 142 mmol/L | 30
potassium 4.4 mmol/L | 30
transthoracic echocardiography good LV function | 30
no regional wall motion abnormalities | 30
transferred to ICU | 30
ventricular pacing threshold 1.75 V at 8 hours ICU | 8
full recovery | 240
discharged home postoperative day 12 | 288
ventricular pacing threshold 0.75 V | 288
ventricular pacing duration 0.6 ms | 288
ventricular pacing output 2.5 V | 288
ventricular pacing duration 0.9 ms | 288
no acid-base disturbance | 0
no electrolyte disorder | 0
no myocardial ischemia | 0
no antiarrhythmic drugs administered | 0
local anesthetic plasma concentration elevation | 0
sodium channel inhibition by levobupivacaine | 0
