26 years old| 0
male | 0
admitted to the emergency room | 0
gastrointestinal obstructive symptoms | -24
aspiration pneumonia | -24
septic shock | -24
chronic pancreatitis | *
alcoholism | *
Type 1 diabetes mellitus | *
schizophrenia | *
epilepsy | *
severely malnourished | 0
body mass index 15.7 kg/m² | 0
abdomen distended | 0
abdomen tympanic | 0
abdomen non-tender | 0
diminished breath sounds at lower base of right lung | 0
transferred to intensive care unit | 0
refractory shock | 0
started on vasopressors | 0
started on broad-spectrum antibiotics | 0
nasogastric tube placed | 0
bilious output 1.8 L | 0
computed tomography scan | 24
distended stomach | 24
distended first and second portion of duodenum | 24
extrinsic compression of third portion of duodenum | 24
narrow aortomesenteric angle 14.3° | 24
diagnosis of SMA syndrome | 24
extrinsic compression of left renal vein | 24
esophagogastroduodenoscopy performed | 48
Candida esophagitis | 48
antibiotic treatment initiated | 48
post-obstruction Dobhoff tube placed | 48
improved | 72
discharged | 72
enteric nutrition | 72
oral antibiotics | 72
denied hematuria | 0
denied decreased urine output | 0
denied flank pain | 0
denied low back pain | 0
BMI 18 kg/m² at follow-up | 1488
resolution of gastrointestinal obstructive symptoms | 1488
no recurrence of abdominal pain | 1488
denied hematuria at follow-up | 1488
denied oliguria | 1488
denied flank pain at follow-up | 1488
denied low back pain at follow-up | 1488
CT imaging avoided | 1488
26 years old|0
male|0
admitted to the emergency room|0
gastrointestinal obstructive symptoms|-24
aspiration pneumonia|-24
septic shock|-24
chronic pancreatitis|*
alcoholism|*
Type 1 diabetes mellitus|*
schizophrenia|*
epilepsy|*
severely malnourished|0
body mass index 15.7 kg/m²|0
abdomen distended|0
abdomen tympanic|0
abdomen non-tender|0
diminished breath sounds at lower base of right lung|0
transferred to intensive care unit|0
refractory shock|0
started on vasopressors|0
started on broad-spectrum antibiotics|0
nasogastric tube placed|0
bilious output 1.8 L|0
computed tomography scan|24
distended stomach|24
distended first and second portion of duodenum|24
extrinsic compression of third portion of duodenum|24
narrow aortomesenteric angle 14.3°|24
diagnosis of SMA syndrome|24
extrinsic compression of left renal vein|24
esophagogastroduodenoscopy performed|48
Candida esophagitis|48
antibiotic treatment initiated|48
post-obstruction Dobhoff tube placed|48
improved|72
discharged|72
enteric nutrition|72
oral antibiotics|72
denied hematuria|0
denied decreased urine output|0
denied flank pain|0
denied low back pain|0
BMI 18 kg/m² at follow-up|1488
resolution of gastrointestinal obstructive symptoms|1488
no recurrence of abdominal pain|1488
denied hematuria at follow-up|1488
denied oliguria|1488
denied flank pain at follow-up|1488
denied low back pain at follow-up|1488
CT imaging avoided|1488
