10 years old | 0
male | 0
born by caesarean section | 0
birth weight 2100 g | 0
birth length 48 cm | 0
Apgar score 8 | 0
prominent forehead | 0
relative macrocephaly | 0
limb asymmetry | 0
5th finger clinodactyly | 0
2/3 toe syndactyly | 0
SRS suspected | 0
genetic examination | 0
hypomethylation of 11p15 region | 0
SRS confirmed | 0
delayed motor development | 0
walked independently at 16 months | -120
hepatic dysfunction suspected | -14
increased AlAT | -14
increased AspAT | -14
increased creatine kinase | -14
DMD considered | -14
genetic test performed | -21
DMD confirmed | -21
exon deletion 49-50 detected | -21
DMD diagnosed in asymptomatic phase | -21
frequent falling | -21
tiptoed gait | -21
Achilles tendon contractures | -21
Gover's syndrome positive | -21
calf enlargement | -21
prednisone treatment | -48
deflazacort treatment | -24
slower height velocity observed | -48
G-CSF treatment started | -48
G-CSF administered 5 days monthly | -48
improvement in 6MWT | -48
sepsis hospitalization | -48
intensive care treatment | -48
severe hypoglycemia | -48
neurological symptoms | -48
glucose level 14 mg/dl | -48
hypospadias | 0
cardiological diagnostics | 0
sinus tachycardia | 0
heart murmur | 0
cardiomyopathy excluded | 0
propranolol treatment | 0
height deficiency | 0
weight deficiency | 0
growth hormone deficiency excluded | 0
rhGH qualification | 0
physical examination at admission | 0
hypotonia | 0
malocclusion | 0
Tanner stage 1 | 0
height 115.9 cm | 0
weight 19.9 kg | 0
BMI 14.8 kg/m² | 0
target height SDS 0.61 | 0
height velocity 4.3 cm/year | 0
OGTT normal | 0
IGF-1 231 ng/ml | 0
IGFBP-3 7.29 µg/ml | 0
MRI transparent septum cyst | 0
rhGH treatment started | -13
height velocity increased to 6.9 cm/year | 12
IGF-1 increased | 12
BMI increased to 21.9 kg/m² | 18
impaired glucose tolerance | 12
insulin resistance | 12
HOMA-IR 9.66 | 12
HbA1c elevated | 12
6MWT distance decreased | 12
gait abnormality | 12
rhGH dose reduced | 12
lifestyle modification recommended | 12
rhGH discontinued | 18
bone density Z-score -2.2 | 12
body composition assessed | 12
reduced muscle mass | 12
high fat content | 12
scoliosis not developed | 18
conflict of interest none | 0
