58 years old | 0
female | 0
admitted to the hospital | 0
lethargy | -48
fever | -48
watery, non-bloody diarrhea | -48
confusion | -48
hypertension | 0
rheumatoid arthritis | 0
chronic kidney disease | 0
chronic obstructive pulmonary disease | 0
current smoker | 0
20 pack-year smoking history | 0
no history of alcohol or illicit drug use | 0
temperature of 39.4 °C | 0
heart rate of 112 beats per minute | 0
respiratory rate of 20 per minute | 0
blood pressure of 127/75 mm Hg | 0
oxygen saturation of 85% on room air | 0
oxygen saturation of 100% on 3 L nasal cannula | 0
drowsy | 0
oriented to place and person but not to time | 0
no focal neurological deficits | 0
no neck rigidity | 0
no meningeal signs | 0
no rashes | 0
white blood cells 17,400 cells per μL | 0
neutrophils 87% | 0
hemoglobin 10.7 g/dL | 0
platelet count 235,000 per μL | 0
sodium 126 mEq/L | 0
potassium 3.0 mEq/L | 0
bicarbonate 19.3 mEq/L | 0
blood urea nitrogen 32 mg/dL | 0
creatinine 2 mg/dL | 0
aspartate aminotransferase 260 Units/L | 0
alanine aminotransferase 40 Units/L | 0
Creatine kinase 347,700 units/liter | 0
hepatitis A IgM antibody negative | 0
hepatitis B surface antigen negative | 0
hepatitis B core IgM antibody negative | 0
hepatitis C antibodies negative | 0
stool studies showed no WBC in stools | 0
normal osmolality | 0
normal calprotectin | 0
urine, blood and stool cultures negative | 0
urine legionella pneumophila serogroup 1 antigen positive | 0
urinalysis showed 51–100/hpf of WBC | 0
urinalysis showed 6–10/hpf of red blood cells | 0
urinalysis showed 3+ occult blood | 0
new bibasilar densities on chest X ray | 0
patchy right basilar opacities on CT chest | 0
small right pleural effusion on CT chest | 0
colonic diverticulosis | 0
no evidence of diverticulitis | 0
started on broad spectrum antibiotics | 0
switched to azithromycin | 24
improvement in mental status | 24
improvement in diarrhea | 24
worsening renal function | 24
worsening creatine kinase | 24
anuria | 48
volume overload | 48
started on hemodialysis | 48
transferred to intensive care unit | 48
received 14 day course of azithromycin | 168
weaned off pressors | 168
weaned off supplementary oxygen | 168
started on midodrine | 168
rhabdomyolysis started to resolve | 168
discharged | 408
follow up hemodialysis as an outpatient | 408
complete renal recovery | 1440