29 years old | 0
male | 0
previous history of right knee fracture | -672
admitted to the hospital | 0
persistent fever | -336
fever with chills | -336
swelling and pain of right knee joint | -240
shortness of breath | -240
fatigue after physical activity | -240
oliguria | -240
frothy and foul-smelling urine | -240
hypothermia | 0
heart rate 100 beats/min | 0
respiratory rate 20 breaths/min | 0
blood pressure 138/80 mmHg | 0
infection | 0
cavity effusion and synovial thickening in right knee joint | 0
pneumonia | 0
hepatic cyst in S7 segment | 0
empiric antibiotic therapy | 0
piperacillin/tazobactam | 0
blood cultures | 0
cavity effusion sample | 24
yellow color of cavity effusion | 24
white blood count (WBC) (+++/HP) | 24
red blood count (RBC) (1–3/HP) | 24
turbidity | 24
persistent fever | 48
peak temperature at 39.5 °C | 48
carbapenems (biapenem) | 72
empiric gram positive coverage | 72
IV vancomycin | 72
Klebsiella pneumoniae | 120
hypermucoviscosity phenotype | 120
antibiotic sensitivity testing | 120
levofloxacin | 120
cefotaxime | 120
piperacillin/tazobactam | 120
carbapenems | 120
voriconazole | 144
urine culture Candida albicans | 144
meropenem | 168
RFP | 168
vancomycin discontinued | 168
voriconazole discontinued | 168
clinically improved | 192
afebrile | 192
discharged | 336
meropenem combined with RFP | 168
treated for 10 days | 168
hyperglycemia | 0
high blood glucose concentration | 0
diabetes mellitus | -672
independent risk factor | -672
hyperglycemia | -672
inhibited chemotaxis and adhesion of leukocytes | -672
damaged intestinal barrier | -672
promoted formation of liver abscess | -672
changed structure and function of vascular intima | -672
Klebsiella pneumoniae transported to blood | -672
caused liver abscess | -672
capsular polysaccharide | -672
increased virulence | -672
protected strain against human defense activities | -672
rmpA gene | -672
magA gene | -672
most important virulence factor of hvKP | -672
related to migration, adhesion, and proliferation of hvKP | -672
produced more capsular polysaccharide | -672
explained why treatment was not effective | -672
RFP | -672
inhibited transcription of rmpA gene | -672
inhibited capsular polysaccharide biosynthesis | -672
reduced capsular thickness | -672
exerted strong mucoviscosity-suppressing activity | -672
enabled RFP to fight against hvKP effectively | -672
benefited patient | -672