56 years old | 0
male | 0
admitted to the hospital | 0
neck mass detected while shaving | 0
heterogeneous ovoid mass in the left submandibular region | 0
enlarged left paramedial submental lymph node | 0
biopsy of the neck mass | 0
EMC staining positive for CK7, CKAE1/AE3, CK903, S100, and smooth muscle actin | 0
negative for CK20, PAX8, GATA, CDX2, GFAP | 0
infiltrates into soft tissue | 0
fragments of salivary gland with fibrosis and atrophy | 0
resected in piecemeal fashion | 0
final pathology report confirming EMC | 0
Hodgkin lymphoma | -262080
mantle field RT | -262080
chemotherapy | -262080
splenectomy | -262080
no evidence of recurrence | -262080
diffuse large B cell lymphoma | -17520
PET scan displaying diffuse disease | -17520
treatment with denosumab | -17520
six cycles of rituximab, cyclophosphamide, doxorubicin, vincristine, and prednisone | -17520
dizziness | -17520
ataxia | -17520
memory loss | -17520
brain MRI showing two ring-enhancing lesions | -17520
whole brain radiation therapy | -17520
intrathecal cytarabine | -17520
coronary artery disease | -17520
hypertension | -17520
hypothyroidism | -17520
gastroesophageal reflux disease | -17520
mini-stroke | -17520
coronary artery bypass grafting x 4 vessels | -17520
right carotid endarterectomy | -17520
appendectomy | -17520
aortic valve replacement | -17520
maternal grandfather with lung cancer | -17520
maternal uncle with colon cancer | -17520
paternal grandfather with lung cancer | -17520
no first degree relatives with a history of cancer, heart disease, alcoholism, asthma, bleeding disorder, diabetes, or thyroid disease | -17520
32-pack year smoking history | -17520
asbestos exposure | -17520
no alcohol or illicit drug use | -17520
bilateral dense fibrosis | 0
revision surgery with additional neck dissection | 0
resection of the left submandibular gland | 0
dissection of level IA, IB, and suprahyoid neck nodes | 0
histologic examination revealed EMC in 1/2 left level IB lymph nodes | 0
0/3 left level IA lymph nodes | 0
pT2pN1M0 | 0
extensive lymphovascular invasion | 0
positive margins on the primary mass | 0
adjuvant chemoradiation | 0
intensity-modulated radiation therapy | 0
5040 cGy in 28 fractions | 0
3D-boost of 1620 cGy in 9 fractions | 0
cumulative dose totaled 6660 cGy in 37 fractions | 0
concurrent chemotherapy with weekly carboplatin and paclitaxel | 0
no evidence of EMC disease | 0
xerostomia | 0
fibrosis of the neck tissues | 0
restaging PET scan demonstrated mild to moderate FDG uptake in right upper lobe lung nodule | 240
interval growth of the nodule | 240
bronchoscopy with biopsy revealed neuroendocrine tumor | 240
tumor positive for CAM 5.2, TTF1, synaptophysin, and chromogranin | 240
Ki67 immunoperoxidase stain with low proliferation rate | 240
denied any cough | 240
denied shortness of breath | 240
denied diarrhea | 240
denied flushing | 240
denied weight loss | 240
elected for observation | 240
intensely FDG focus in left thyroid lobe | 240
thyroid ultrasound with Doppler | 240
fine needle aspiration revealed follicular lesion of undetermined significance | 240
predominantly Hurthle cells | 240
benign nodular hyperplasia | 240
elected to proceed with chemoradiation | 240
hemithyroidectomy | 240
follow-up CT scan displayed interval growth of right upper lobe NET | 2400
several new bilateral pulmonary nodules | 2400
PET scan noted new intensely FDG avid focus in left pterygoid muscle | 2400
intensely avid hilar lymphadenopathy | 2400
moderately avid mediastinal lymph nodes | 2400
biopsy of pulmonary nodules and mediastinal lymph nodes negative for malignancy | 2400
elected for SBRT to right lung | 2400
5250 cGy over 5 fractions | 2400
developed pneumonia | 2400
sepsis | 2400
vasopressor requirement | 2400
bilateral pleural effusions | 2400
flow cytometry of pleural fluid notable for CD10-positive lambda-skewed B cell population | 2400
negative peripheral blood flow cytometry | 2400
transfer to palliative care unit | 2400
inpatient hospice | 2400
expired | 2400
