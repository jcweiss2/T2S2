56 years old| 0
    male| 0
    admitted to the hospital| 0
    chronic left leg ulcer| 0
    liver cirrhosis| 0
    congestive heart failure| 0
    substance use disorder| 0
    bacteremia| 0
    leg infection| 0
    non-healing wound on left leg| 0
    pain in both legs| 0
    chills| 0
    subjective fevers| 0
    febrile| 0
    heart rate 98| 0
    respiratory rate 16| 0
    oxygen saturation 99| 0
    mean arterial pressure 100| 0
    alert and oriented| 0
    no cardiorespiratory distress| 0
    no murmur| 0
    no friction rub| 0
    clear breath sounds| 0
    soft abdomen| 0
    no guarding| 0
    no rigidity| 0
    tenderness on deep palpation at left lower quadrant| 0
    bilateral chronic venous stasis changes| 0
    hyperpigmentation| 0
    dryness| 0
    superficial scaling| 0
    edema| 0
    left leg ulcer| 0
    clean margins| 0
    clean base| 0
    no drainage| 0
    no crepitus| 0
    pedal pulses appreciated| 0
    grossly intact sensation| 0
    grossly intact motor function| 0
    able to move knees| 0
    able to move feet| 0
    able to move toes| 0
    right knee suprapatellar effusion| 0
    not tender| 0
    unremarkable rest of examination| 0
    cellulitis of the right leg| 0
    qSOFA score zero| 0
    hypertension| 0
    hyperlipidemia| 0
    stroke 12 years ago| -105120
    left sided residual weakness| -105120
    Childs Pugh A liver cirrhosis| 0
    untreated hepatitis C| 0
    heart failure with ejection fraction 40-45| 0
    polysubstance use| 0
    methadone maintenance program| 0
    aspirin 81 mg daily| 0
    atorvastatin 40 mg daily| 0
    ferrous sulfate 325 mg daily| 0
    folic acid 1 mg daily| 0
    gabapentin 300 mg twice daily| 0
    metoprolol succinate 50 mg daily| 0
    mirtazapine 15 mg nightly| 0
    sacubitril 24 mg twice daily| 0
    valsartan 26 mg twice daily| 0
    thiamine 100 mg daily| 0
    misses medications on occasion| 0
    multiple emergency room visits| 0
    multiple admissions for chronic left leg ulcer| 0
    previous wound cultures grew Streptococcus epidermidis| 0
    previous wound cultures grew Streptococcus pyogenes| 0
    admitted two weeks prior| -336
    blood culture no growth| -336
    completed 10 days intravenous vancomycin| -336
    discharged to shelter| -336
    wheelchair bound| 0
    lives in shelter| 0
    started drinking alcohol at 14| -153528
    drinking 10 tall cans beer daily| 0
    last drink one day prior| -24
    denied smoking cigarettes| 0
    opioid use disorder with heroin since age 24| -281856
    intranasal administration| -281856
    intravenous method| -281856
    last heroin use two days prior| -48
    normocytic anemia| 0
    normochromic anemia| 0
    chronic thrombocytopenia| 0
    white blood cells within normal limits| 0
    elevated C-reactive protein| 0
    normal lactic acid| 0
    sinus tachycardia| 0
    no acute ischemic changes| 0
    blood cultures obtained| 0
    loaded with intravenous vancomycin| 0
    started on ampicillin-sulbactam| 0
    persistence of abdominal tenderness| 0
    urinalysis significant hematuria| 0
    otherwise unremarkable urinalysis| 0
    no deep venous thrombosis| 0
    normal chest radiograph| 0
    right lower extremity radiography severe joint space narrowing| 0
    right lower extremity radiography small suprapatellar joint effusion| 0
    left lower extremity radiography moderate degenerative changes| 0
    left lower extremity radiography suprapatellar joint effusion| 0
    left lower extremity radiography subcutaneous emphysema| 0
    bibasilar atelectasis| 0
    coronary artery atherosclerosis| 0
    cardiomegaly| 0
    nodular liver contour| 0
    liver enlargement| 0
    mild splenomegaly| 0
    splenorenal varices| 0
    gastric varices| 0
    degenerative changes L5-S1| 0
    blood cultures positive Empedobacter falsenii/tilapiae| 96
    multidrug resistance| 96
    urine culture no growth| 96
    swab culture left leg ulcer grew vancomycin-resistant Enterococcus faecalis| 96
    received vancomycin| 0
    received ampicillin-sulbactam| 0
    started on piperacillin-tazobactam| 0
    urology consulted| 0
    urine cytology recommended| 0
    prostate specific antigen levels recommended| 0
    tamsulosin started| 0
    wound care recommended cleansing| 0
    XeroForm occlusive gauze| 0
    foam dressing| 0
    Kerlix wrap daily| 0
    orthopedics consulted| 0
    compressive knee support recommended| 0
    ice packs recommended| 0
    elevation of lower extremities recommended| 0
    careful weight bearing recommended| 0
    shifted to cefepime| 96
    fever defervesced on day 2| 48
    stayed afebrile| 48
    continued improvement| 96
    discharged home| 168
    oral trimethoprim-sulfamethoxazole| 168
    missed follow up| 720
    admitted one month later| 720
    left lower extremity cellulitis| 720
    urinary tract infection| 720
    urine culture grew Klebsiella pneumoniae| 720
    levofloxacin recommended| 720
    discharged after antibiotics| 720
    admitted two months later| 1464
    acute hypoxemic respiratory failure| 1464
    pneumonia| 1464
    septic shock| 1464
    encephalopathy| 1464
    blood culture grew Klebsiella pneumoniae| 1464
    bronchial aspirate culture grew multidrug resistant Staphylococcus aureus| 1464
    