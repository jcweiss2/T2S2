75 years old | 0
female | 0
habit of taking vinegar daily | -43800
hypertension | -8760
amlodipine 10 mg daily | -8760
vomiting | -1
loss of consciousness | -1
unconscious | 0
hypotensive | 0
respiratory failure | 0
sinus tachycardia | 0
oxygen saturation 90% | 0
no subcutaneous emphysema | 0
no signs of peritoneal irritation | 0
white blood count 3500 | 0
C-reactive protein level 8.7 mg/dL | 0
renal dysfunction | 0
electrolytes normal | 0
liver function normal | 0
urinalysis normal | 0
computed tomography of thoracic and abdomen | 0
poor contrast in middle intrathoracic esophagus | 0
mediastinal emphysema | 0
right pneumothorax | 0
pleural effusion | 0
septic shock due to esophageal rupture | 0
emergency surgery | 0
esophageal rupture | 0
esophagectomy | 0
intrathoracic lavage drainage | 0
esophageal fistula | 15
enteric fistula | 15
intensive care | 0
vitals stable | 15
esophageal and enteric fistulae | 15
esophageal mucosa blackened | 15
esophageal fistula mucosa normalized | 120
esophageal reconstruction | 1440
posterior sternal pathway cervical esophagogastric anastomosis | 1440
cholecystectomy | 1440
oral intake | 1552
discharged | 1620