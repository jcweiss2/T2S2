13 years old | 0
male | 0
admitted to the hospital | 0
electric burn | -720
electric burn over the right arm | -720
electric burn over the right axilla | -720
electric burn over the right-sided thoracic and abdominal region | -720
electric burn over the left foot | -720
debridement | -720
amputation of the right great toe | -720
amputation of the 4th and 5th toes of the left foot | -720
skin grafting | -720
post-burn contracture release | 0
difficulty in extension of arm | -2160
contracture release of right axillary region | -720
skin grafting | -720
multiple blood transfusions | -720
vegetarian diet | 0
weight loss | -216
reduced appetite | -216
feeling tired | -216
feeling weaker | -216
wounds taking a long time to heal | -216
poor concentration | -216
feeling cold | -216
restriction of exertional activity | 0
BMI 12.9 | 0
underweight | 0
able to go to school | 0
able to walk at normal speed | 0
weight 32 kg | 0
normal chest X-ray | 0
normal electrocardiogram | 0
informed consent | 0
monitors attached | 0
preoperative vitals noted | 0
heart rate 94/min | 0
BP 104/62 mmHg | 0
SpO2 98% | 0
premedicated with Inj. Glycopyrrolate | 0
premedicated with Inj. Ondansetron | 0
premedicated with Inj. Midazolam | 0
premedicated with Inj. Fentanyl | 0
preoxygenated with 100% oxygen | 0
anesthesia induced with Inj. Propofol | 0
relaxed with Inj. Atracurium | 0
intubated orally with cuffed ET tube | 0
anesthesia maintained with Sevoflurane | 0
intraoperative monitoring | 0
tachycardia | 1
hypotension | 1
HR 150/min | 1
BP 70/30 mmHg | 1
SpO2 84% | 1
pink frothy secretions | 1
bilateral crepitations | 1
FiO2 increased to 100% | 1
Inj. Furosemide given | 1
positive pressure ventilation | 1
deeper plane of anesthesia | 1
Inj. Atracurium given | 1
Inj. Noradrenaline started | 1
arterial blood gas analysis | 1
hypoxia | 1
decreased PaO2/FiO2 ratio | 1
lactate level 4.5 mmol/l | 1
surgery completed | 45
reversed with Inj. Neostigmine | 45
reversed with Inj. Glycopyrrolate | 45
extubated | 45
O2 support | 45
shifted to intensive care unit | 45
cardiac status evaluated | 45
LVEF 20% | 45
global LV hypokinesia | 45
dilated LV | 45
mild MR/TR | 45
thiamine deficiency suspected | 45
Inj. Thiamine started | 45
Tab. Carvedilol started | 45
Tab. Spironolactone + Furosemide started | 45
Tab. Enalapril started | 45
chest X-ray | 45
pulmonary edema | 45
IV fluid restricted | 45
urine output measured | 45
total input/output | 93
vasopressor requirement decreased | 69
vasopressor requirement stopped | 69
oxygen requirement decreased | 69
repeat ABGA | 69
improved PaO2/FiO2 ratio | 69
air entry equal and clear | 69
repeat 2D echo | 93
LVEF 50% | 93
fair LV function | 93
normal-sized cardiac chambers | 93
no MR/TR | 93
discharged | 168
follow up after six weeks | 168
thiamine rich diet | 168