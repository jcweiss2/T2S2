8 years old|0
    female spayed|0
    domestic shorthair cat|0
    acute onset of lethargy|0
    acute onset of pain|0
    indoor/outdoor cat|0
    not up to date with vaccinations|0
    no known history of trauma|0
    no recent medication administration|0
    elevated body temperature|0
    hypotensive|0
    blood pressure 80 mmHg|0
    tachypneic|0
    respiratory rate 60 breaths per min|0
    painful at thoracolumbar spine|0
    three small puncture wounds on back|0
    mild hyperglycemia|0
    complete blood count normal|0
    white blood cell count 17.27 × 109/l|0
    PCV 41%|0
    total protein 7.5 g/dl|0
    negative retroviral disease|0
    radiographs of thorax and abdomen|0
    mild diffuse bronchointerstitial pulmonary pattern|0
    normal abdomen|0
    normal skeletal structures|0
    soft tissue swelling and gas dorsal to lumbar spine|0
    cellulitis|0
    intravenous crystalloid fluid boluses|0
    lactated Ringer’s solution|0
    blood pressure increased to 98 mmHg|0
    IV lactated Ringer’s solution|0
    IV buprenorphine|0
    hospitalization declined|0
    discharged|0
    oral transmucosal buprenorphine|0
    oral amoxicillin/clavulanic acid|0
    culture of wound declined|0
    lethargic at home| -23
    anorexic at home| -23
    re-presented to hospital| -23
    obtunded| -23
    body temperature 37.7°C| -23
    respiratory rate 50 breaths per min| -23
    heart rate 180 beats per min| -23
    IV catheter placed in right cephalic vein| -23
    severely hypotensive| -23
    blood pressure 30 mmHg| -23
    hypoglycemic| -23
    blood glucose 1.9 mmol/dl| -23
    focused assessment with ultrasound for trauma negative| -23
    skin on dorsum warm| -23
    subcutaneous fluid pocket suspected| -23
    fine-needle aspirate| -23
    cytology consistent with septic suppurative inflammation| -23
    fluid sample for aerobic culture| -23
    abdominal ultrasound negative| -23
    PCV 43%| -23
    total protein 6.3 g/dl| -23
    venous blood gas normal| -23
    admitted to intensive care unit|0
    treated with ampicillin–sulbactam|0
    treated with enrofloxacin|0
    treated with metronidazole|0
    treated with vitamin C|0
    treated with maropitant citrate|0
    treated with famotidine|0
    fentanyl constant rate infusion|0
    dextrose bolus|0
    LRS with dextrose and potassium chloride|0
    sedated with fentanyl and midazolam|0
    wound opened surgically|0
    wound debrided|0
    wound lavaged with saline|0
    wet-to-dry tie over bandage placed|0
    double-lumen catheter placed in left jugular vein|0
    indwelling urinary catheter placed|0
    unsuccessful arterial catheter placement|0
    hypotension persisted|0
    norepinephrine constant rate infusion started|0
    dopamine constant rate infusion started|0
    vasopressin constant rate infusion started|0
    arterial cut-down performed|0
    arterial catheter placed in right dorsal pedal artery|0
    MAP 30 mmHg|0
    dopamine dose increased|24
    MAP 40 mmHg|24
    vasopressin dose unchanged|24
    hydrocortisone CRI started|24
    dextrose supplementation discontinued|24
    dopamine discontinued|24
    norepinephrine dose decreased|24
    vasopressin CRI discontinued|24
    third day of hospitalization|72
    able to maintain sternal recumbency|72
    ate small amount of food|72
    motor function present|72
    pain sensation present|72
    unable to stand or walk|72
    less painful|72
    fentanyl CRI decreased|72
    wet-to-dry bandage changed|72
    norepinephrine and vasopressin doses decreased|72
    MAP 70-80 mmHg|72
    day 5 hospitalization|120
    anesthetized|120
    Jackson-Pratt drain placed|120
    wound closed|120
    hypotension during surgery|120
    MAP 45 mmHg|120
    treated with dopamine|120
    hypotension resolved|120
    dopamine discontinued|120
    PCV 19%|120
    anemia suspected|120
    blood type A|120
    packed red blood cells transfusion|120
    eating readily|120
    transitioned to oral antibiotics|120
    wound culture scant growth|120
    enrofloxacin discontinued|120
    day 6|144
    right thoracic limb swollen|144
    right pelvic limb swollen|144
    limbs cold to touch|144
    IV catheters removed|144
    central venous catheter maintained|144
    day 7|168
    paws cold to touch|168
    paws painful|168
    paws discolored|168
    skin sloughing on paw pads|168
    line of demarcation noted|168
    strong pedal pulses|168
    clopidogrel started|168
    clopidogrel continued until healing|168
    normotensive|168
    MAP >70 mmHg|168
    continued wound care|168
    hydrotherapy|168
    discharged after 11 days|264
    soft padded bandages|264
    paws fully healed|264
    necrotic skin debrided|264
    bandage changes over 2 weeks|264
    ambulatory with mild pelvic limb weakness|264