36 years old| 0
female | 0
admitted to the hospital | 0
abdominal pain | -216
diarrhea | -216
mucus blood | -216
pus | -216
recurrent tenesmus attacks | -216
fecal microbiota transplantation | -216
anuria | -144
vomiting | -144
severe diarrhea | -144
UC (diagnosed ten years ago) | -87600
mesalazine | -87600
prednisone | -87600
dark colored urine (100 mL) | 0
bloody fluid discharged from urethral catheter | 0
dyspneic | 0
cold clammy limbs | 0
increased pulse rate | 0
abdominal cavity pressure 25 mmHg | 0
grade IV abdominal hypertension | 0
total colonic wall thickening | 0
erosions in luminal surface of colon | 0
hyperemia | 0
friability | 0
bleeding | 0
ulcerations | 0
white blood count 40.77 × 109/L | 0
red blood count 2.41 × 1012/L | 0
hemoglobin 60 G/L | 0
sequential organ failure assessment score 10 | 0
suspicious thin perforations at rectosigmoid colon | 0
massive ascites | 0
septic shock | 0
colonic perforation | 0
UC (active) | 0
acute renal failure | 0
disseminated intravascular coagulation | 0
severe anemia | 0
total proctocolectomy | 0
ileostomy | 0
massive ascites (observed during surgery) | 0
total colonic necrosis | 0
edema | 0
dilatation of small intestine | 0
no obvious perforation | 0
no arterial thrombosis | 0
ascites culture negative | 0
mucosal inflammation (histopathology) | 0
necrosis (histopathology) | 0
hemorrhage (histopathology) | 0
transferred to ICU | 24
symptoms alleviated | 24
urine excretion normal | 24
maintenance of renal perfusion | 24
ascites fluid drained (1880&ndash;3880 mL daily for 7 d) | 24
possibility of thrombosis considered | 24
anticoagulant therapy | 24
ascites volume reduced | 24
condition improved | 24
computed tomography angiography | 72
thrombosis in trunk of portal vein | 72
thrombosis in intrahepatic branches | 72
thrombosis in superior mesenteric vein | 72
thrombosis in splenic vein | 72
recovered | 72
discharged | 72
antibacterial treatment | 72
anticoagulant treatment | 72
nutritional support treatment | 72
