37 years old | 0
male | 0
unmarried | 0
lived with a cousin | 0
worked in a plastics factory | 0
admitted to the hospital | 0
fever | -96
vomiting | -24
loose stools | -24
abdominal cramps | -24
headache | -24
tachycardia | 0
mild tachypnea | 0
blood pressure 100/70 mmHg | 0
macular erythematous rash | 0
Glasgow coma scale score 15 | 0
no neck stiffness | 0
thrombocytopenia | 0
high serum concentrations of creatinine | 0
high serum concentrations of urea | 0
high serum concentrations of total bilirubin | 0
high serum concentrations of aspartate aminotransferase | 0
high serum concentrations of alanine aminotransferase | 0
high serum concentrations of C-reactive protein | 0
mild bilateral haziness on chest X-rays | 0
started on empirical treatment with ceftriaxone | 0
provisionally diagnosed with acute gastroenteritis | 0
provisionally diagnosed with acute kidney injury | 0
admitted to the hospital | 0
continued to receive fluids and antibiotics | 0
became more tachypneic | 48
became more tachycardic | 48
fever spike of 38.3°C | 48
episode of hypoglycemia | 48
transferred to the Intensive Care Unit | 72
started on treatment with piperacillin/tazobactam | 72
intubated and ventilated | 72
required vasopressors | 96
required higher positive end-expiratory pressure | 96
blood culture positive for S. moniliforms | 120
diagnosed with RBF | 120
started on intravenous penicillin G | 120
showed rapid improvement | 144
weaned off the ventilator | 144
vasopressor tapered | 144
renal functions improved | 144
acidosis improved | 144
extubated | 144
discharged from the hospital | 240
rats may have been present in his house | -96
rats may have been present in his workplace | -96
frequently leaves food uncovered at both sites | -96
no history of rat bite | 0
no shortness of breath | 0
no chest pain | 0
no heart failure | 240
no infective endocarditis | 240
normal findings on echo-cardiography | 240