21 years old | 0
woman | 0
consulted the emergency department | 0
38 weeks of gestation | 0
premature rupture of membranes | 0
occasional contraction-type abdominal pain | 0
pregnancy | 0
5 prenatal check-ups | 0
alert | 0
normal vital signs | 0
fetal movement | 0
fetal heart rate of 145 beats per minute | 0
cervix without cervical changes | 0
normal hemogram | 0
negative COVID-19 antigen test | 0
normal biophysical profile | 0
reactive fetal monitoring | 0
irregular uterine dynamics | 0
pregnancy at term | 0
vaginosis | 0
whitish vaginal discharge | 0
hospitalized for labor induction with oxytocics | 0
after 23 hours without cervical changes | 23
34 hours of PROM | 34
induction failure | 34
bradycardia | 34
hypotension | 34
desaturation | 34
cardiorespiratory arrest | 34
resuscitation maneuvers | 34
return of spontaneous circulation | 34
required mechanical ventilation | 34
sulbactam ampicillin | 34
3 doses of tranexamic acid | 34
dexamethasone | 34
newborn Apgar score 7 at 1 minute | 34
Apgar score 8 at 5 minutes | 34
Apgar score 9 at 10 minutes | 34
fibrinogen 346 mg/dL | 34
normal arterial blood gasses | 34
normal coagulation times | 34
PT 13 seconds | 34
TPT 28 seconds | 34
lactate dehydrogenase 1.203 IU/L | 34
D-dimer >10,000 ng/mL | 34
angiotomography showed pulmonary embolism | 34
pulmonary edema | 34
respiratory infection | 34
asymptomatic SARS-CoV-2 infection | 34
elevated risk of pneumonia | 34
mild ARDS | 34
sepsis | 34
cardiogenic shock | 34
intensive care unit stay for 6 days | 168
mechanical ventilation withdrawn | 168
leukocytes 6250 × 103/mm3 | 168
neutrophils 60% | 168
procalcitonin <0.05 ng/mL | 168
negative blood cultures | 168
negative urine cultures | 168
negative orotracheal tube culture | 168
satisfactory recovery | 168
discharged | 168
21 years old| 0
woman| 0
consulted the emergency department| 0
38 weeks of gestation| 0
premature rupture of membranes| 0
occasional contraction-type abdominal pain| 0
pregnancy| 0
5 prenatal check-ups| 0
alert| 0
normal vital signs| 0
fetal movement| 0
fetal heart rate of 145 beats per minute| 0
cervix without cervical changes| 0
normal hemogram| 0
negative COVID-19 antigen test| 0
normal biophysical profile| 0
reactive fetal monitoring| 0
irregular uterine dynamics| 0
pregnancy at term| 0
vaginosis| 0
whitish vaginal discharge| 0
hospitalized for labor induction with oxytocics| 0
after 23 hours without cervical changes| 23
34 hours of PROM| 34
induction failure| 34
bradycardia| 34
hypotension| 34
desaturation| 34
cardiorespiratory arrest| 34
resuscitation maneuvers| 34
return of spontaneous circulation| 34
required mechanical ventilation| 34
sulbactam ampicillin| 34
3 doses of tranexamic acid| 34
dexamethasone| 34
newborn Apgar score 7 at 1 minute| 34
Apgar score 8 at 5 minutes| 34
Apgar score 9 at 10 minutes| 34
fibrinogen 346 mg/dL| 34
normal arterial blood gasses| 34
normal coagulation times| 34
PT 13 seconds| 34
TPT 28 seconds| 34
lactate dehydrogenase 1.203 IU/L| 34
D-dimer >10,000 ng/mL| 34
angiotomography showed pulmonary embolism| 34
pulmonary edema| 34
respiratory infection| 34
asymptomatic SARS-CoV-2 infection| 34
elevated risk of pneumonia| 34
mild ARDS| 34
sepsis| 34
cardiogenic shock| 34
intensive care unit stay for 6 days| 168
mechanical ventilation withdrawn| 168
leukocytes 6250 × 103/mm3| 168
neutrophils 60%| 168
procalcitonin <0.05 ng/mL| 168
negative blood cultures| 168
negative urine cultures| 168
negative orotracheal tube culture| 168
satisfactory recovery| 168
discharged| 168
