43 years old | 0
male | 0
pedestrian accident | -1
admitted to the hospital | 0
comatose | 0
Glasgow coma score of 3 | -1
nonreactive pupils 5 mm in diameter | -1
ventilated | 0
hemodynamically stable condition | 0
bilateral otorrhea | 0
rhinorrhea | 0
bruising in face and jaw | 0
bruising on right side of the scalp | 0
diffuse brain injury | 0
severe cerebral swelling | 0
right-side acute subdural hemorrhage | 0
ring fracture around the foramen magnum | 0
clivus fracture | 0
petrous temporal bones fracture | 0
posterior part of the foramen magnum fracture | 0
no signs of atlanto-occipital dislocation | 0
cervical spine intact | 0
admitted to the neurosurgical intensive care unit | 0
no subsequent neurological changes | 0
brain death suspected | 0
healthy before the accident | -1
Glasgow coma scale score of 3 | 0
fixed, nonreactive pupils 6 mm in diameter | 0
no signs of brain stem activity | 0
stable vital signs | 0
magnetic resonance imaging | 648
swelling of the brain stem | 648
cerebellum swelling | 648
transtentorial herniation | 648
foraminal herniation | 648
pontomedullary laceration | 648
comatose for 34 days | 816
died of pneumonia | 816
sepsis | 816