36 years old | 0
female | 0
gravida 1 para 1001 | 0
admitted to the hospital | 0
labial pain | -72
swelling | -72
fevers | -72
hypertension | -672
body mass index (BMI) 56 kg/m2 | -672
polysubstance abuse | -672
intravenous drug use | -672
opioid abuse | -672
tobacco | -672
asthma | -672
bipolar disorder | -672
obsessive-compulsive disorder | -672
chronic pain syndrome | -672
homelessness | -672
prior cesarean section | -672
body temperature 38.4 °C | 0
blood pressure 135/69 | 0
heart rate 121 beats per minute (bpm) | 0
respiratory rate 18 | 0
large right labial and mons abscess | 0
small opened wound with drainage | 0
mild leukocytosis 16.5 | 0
lactic acid 0.6 mmol/L | 0
hemoglobin A1C 5.6 | 0
Streptococcus viridians | 0
Staphylococcus aureus | 0
Enterococcus faecalis | 0
Actinomyces species | 0
Corynebacterium species | 0
CT abdomen and pelvis showed moderate soft-tissue inflammatory stranding | 0
subcutaneous gas overlying the pubis and extending into the right labia majora | 0
started on standard sepsis protocol | 0
aggressive IV fluids | 0
empiric antibiotics (vancomycin, piperacillin-tazobactam, and clindamycin) | 0
desired to leave against medical advice | 0
four-point restraints were placed | 0
combative behavior | 0
security and local police department were involved | 0
Benign gynecology and general surgery teams were consulted | 0
two-attending consent | 0
emergent surgical debridement | 17
skin-sparing debridement | 17
vulvar and mons NSTI | 17
fascia was not involved | 17
care was taken to avoid major underlying vasculature and clitoris | 17
second-stage debridement | 24
wound dressings were changed daily | 24
Veraflow wound vacuum was placed | 240
Plastic surgery was consulted | 720
delayed-primary closure | 720
mons pubis panniculectomy | 720
#19 Blake drain was placed | 720
#19 Blake drain was removed | 744
infectious disease team transitioned her broad-spectrum antibiotics | 240
Augmentin twice daily | 240
severe agitation | 0
maladaptive personality | 0
emotional dysregulation | 0
additional four-point restraints were utilized | 24
IV access was commonly lost | 24
attempts to leave from the hospital were made | 24
wound disruptions | 24
vacuum changes | 24
pain exacerbations | 24
IV narcotics | 24
Psychiatry and palliative care team were essential | 24
haloperidol and lorazepam | 24
olanzapine and quetiapine | 24
trazadone and hydroxyzine | 24
scheduled acetaminophen and non-steroidal anti-inflammatory agents | 24
gabapentin | 24
oral narcotics | 24
suboxone regimen | 240
multidisciplinary meetings | 240
safe and appropriate discharge planning | 240
transferred to jail | 720
loss to follow-up with gynecology | 720