70 years old | 0
male | 0
obstructive sleep apnea | 0
type 2 diabetes | 0
hypertension | 0
admitted to the hospital | 0
BCG instillation | -4
traumatic catheter placement | -4
hemorrhagic catheter placement | -4
flu-like syndrome | 0
fever | 0
chills | 0
oliguric acute kidney injury (AKI) | 0
liver failure | 0
thrombocytopenia | 0
sepsis | 0
amoxicillin-clavulanic acid | 0
inflammatory syndrome | 0
hepatic cytolysis | 0
cholestasis | 0
sediment and urinary cultures negative | 0
blood cultures for mycobacteria | 0
empirical anti-tuberculous treatment | 0
isoniazid | 0
rifampicin | 0
vitamin B6 | 0
night fever peaks | 0
prostatic encapsulated abscess | 24
ceftazidime | 24
aerobic and anaerobic blood cultures negative | 24
positron emission tomography scanner (pet-scan) | 168
pelvic magnetic resonance imagery | 168
no improvement in patient’s condition | 168
liver deterioration | 168
stop antimicrobial treatment | 168
lung symptoms | 168
cough | 168
grade II dyspnea | 168
bilateral pneumonia | 168
pleural effusion | 168
bronchoscopy | 168
bronchoalveolar lavage (BAL) | 168
Ziel and auramine colorations | 168
trans-bronchial biopsies | 168
mycobacterial research negative | 172
cytology highlighted inflammatory trails | 172
granulocytes | 172
anti-tuberculous treatment restarted | 172
isoniazid | 172
moxifloxacin | 172
corticosteroids | 172
clinical and biological improvement | 180
no more fever | 180
no more chills | 180
normalization of inflammatory and hepatic markers | 180
regression of lung infiltrates | 180
positive blood cultures | 360
discharged from ICU | 360
rehabilitation ward | 360
returned home | 360