24 years old | 0
male | 0
admitted to the hospital | 0
diabetes mellitus type 1 | 0
hyperlipidemia | 0
nausea | -24
nonbilious vomiting | -24
hematemesis | -24
subjective fevers | -24
fatigue | -24
dry cough | -24
chills | -24
denied dyspnea | -24
denied chest pain | -24
denied diarrhea | -24
denied constipation | -24
denied recent ill contacts | -24
denied recent travel | -24
noncompliant with medications | -24
temperature 36.4°C | -24
pulse rate 122 beats/min | -24
blood pressure 141/84 mmHg | -24
respiratory rate 16 breaths/min | -24
oxygen saturation 95% | -24
hypothermic (32.9°C rectally) | -24
Foley probe temperature 36.8°C | -24
mild distress | -24
lethargic | -24
delayed responses | -24
alert and oriented | -24
dry mucous membranes | -24
unremarkable physical examination | -24
blood glucose 507 mg/dL | -24
hemoglobin A1c 15.8% | -24
bicarbonate 2 mEq/L | -24
ketonuria 160 mg/dL | -24
creatinine 1.4 mg/dL | -24
anion gap 30.6 mEq/L | -24
blood cultures | -24
urine culture | -24
SARS-CoV-2 RT-PCR test | -24
chest X-ray no cardiopulmonary disease | -24
sinus tachycardia | -24
assessed for DKA | -24
metabolic encephalopathy | -24
sepsis | -24
vancomycin | 0
cefepime | 0
sodium bicarbonate 150 mEq | 0
potassium repletion 100 mL | 0
insulin infusion 6 units/h | 0
lethargic | 24
fell asleep during examination | 24
diagnosed DKA | 24
anion gap metabolic acidosis | 24
acute kidney injury | 24
oxygen saturation 99% | 24
leukocyte count 12.4 | 24
negative cardiac troponins | 24
respiratory distress | 48
febrile 38.3°C | 48
tachypneic | 48
SARS-CoV-2 positive | 48
intubated | 48
mechanical ventilation | 48
respiratory rate 14 breaths/min | 48
tidal volume 500 mL | 48
FiO2 80% | 48
PEEP 15 cm H2O | 48
arterial blood gas improvement | 48
chest X-ray COVID-19 pneumonia | 48
febrile 40°C | 72
azithromycin added | 72
hydroxychloroquine added | 72
blood glucose stabilized | 96
febrile | 96
tachycardic 118 beats/min | 96
attempted FiO2 60% | 96
oxygen saturation 86% | 96
FiO2 increased to 80% | 96
blood pH 7.40 | 96
oxygen desaturation | 168
febrile | 168
leukocyte count increased | 168
sputum culture | 168
vancomycin discontinued | 168
cefepime discontinued | 168
meropenem added | 168
voriconazole added | 168
yeast isolates | 192
chest X worsening infiltrates | 192
febrile | 216
FiO2 titration failed | 216
desaturations | 216
hypercapnia pCO2 61 mmHg | 216
chest X-ray ARDS | 216
desaturation 50% | 216
hypotensive 40/20 mmHg | 216
bradycardic | 216
pulseless | 216
advanced cardiovascular life support | 216
death | 216
hypoxic respiratory failure | 216
SARS-CoV-2-induced COVID-19 | 216
ARDS | 216
