76 years old|0
woman|0
presented with shortness of breath|0
presented with dysphagia|0
presented with nausea|0
presented with neck discomfort|0
eating| -1
morbid obesity| -148,920
underwent laparoscopic adjustable gastric band| -148,920
LAGB complicated by esophageal dilation| -148,920
intermittent dysphagia| -148,920
band removed| -35,064
noncontrast computed tomography of the chest|0
dilated esophagus|0
right lateral diverticulum|0
impacted food bolus|0
diverticulum not apparent on abdominal CT| -35,064
LAGB still in place| -35,064
underwent endoscopy|0
intubated|0
partial removal of food bolus|0
massive food bolus found in diverticulum|0
GIF-190 scope not advanced into true esophageal lumen|0
GIF-XP scope not advanced into true esophageal lumen|0
compression of lumen by diverticulum|0
unable to tolerate entire procedure|0
transferred to medical intensive care unit|0
stayed in ICU for 1 month|0
inability to wean off mechanical ventilation|0
severe sepsis|0
acute respiratory distress syndrome|0
no surgical intervention|0
tracheostomy placed|0
surgical gastrostomy tubes placed|0
discharged to long-term acute care hospital|720
achalasia|0
outflow tract obstruction|0
mass lesion|0
paraesophageal hernia|0
bariatric procedure|0
pseudoachalasia|0
Zenker diverticulum|0
high esophageal lumen pressure|0
tight LAGB at gastroesophageal junction|0
subsequent esophageal musculature weakness|0
continued dysphagia|0
impactions|0
removal of LAGB| -35,064
no identification of mass lesion|0
no identification of hernia|0
manometry not completed|0
fluoroscopy not completed|0
definitive diagnosis difficult|0
no shortness of breath|0
denies chest pain|0
