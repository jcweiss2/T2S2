42 years old | 0
female | 0
diagnosed with relapsing-remitting MS | -7224
treated with methotrexate | -7224
discontinued methotrexate | -7224
treated with interferon beta 1-a | -7224
discontinued interferon beta 1-a | -4680
treated with fingolimod | -3360
major depression disorder | 0
hypothyroidism | 0
recurrent urinary tract infection | 0
histories of pulmonary embolism | 0
myasthenia gravis | -7224
thymectomy | -7224
expanded disability status scale score was 1.0 | -168
positive Babinski sign | -168
moderate disease burden in the brain | -168
2 right-sided cervical cord lesions | -168
lymphocyte count was 842.4/μL | -168
experienced symptoms | -4
sought medical attention | 0
decreased sensation | 0
reduced muscle strength | 0
brisk reflexes | 0
right positive Babinski sign | 0
EDSS of 4 | 0
admitted for a relapse workup and treatment | 0
afebrile | 0
vital signs within normal limits | 0
C-reactive protein of 76 mg/L | 0
erythrocyte sedimentation rate of 46 mm | 0
decrease in absolute lymphocyte count | 0
methylprednisolone IV 1,000 mg/d | 0
chest X-ray showed a ground glass opacity | 0
started on azithromycin 500 mg daily | 0
developed dry cough | 48
developed dyspnea | 48
developed fever | 48
tachycardia | 48
increased respiratory rate | 48
decrease in blood pressure | 48
decrease in oxygen saturation | 48
decrease in lymphocyte counts | 48
fingolimod was stopped | 48
ceftriaxone 1 g twice daily | 48
started on oxygen via a nasal cannula | 48
chest CT was performed | 72
ground glass opacities | 72
COVID-19 was suspected | 72
nasopharyngeal swab was obtained | 72
transferred to the special COVID ward | 72
received a combination of hydroxychloroquine, oseltamivir, and piperacillin/tazobactam | 72
ceftriaxone and azithromycin were discontinued | 72
felt well | 120
vital signs were stabilized | 120
became afebrile | 120
lymphocyte counts increased | 120
COVID-19 test was reported positive | 144
all other medications except hydroxychloroquine were discontinued | 144
symptoms of cough and dyspnea gradually improved | 168
neurologic symptoms gradually improved | 168
discharged | 312
started on glatiramer acetate | 312
lymphocyte count was 1,000.5/ul | 312
self-quarantined at home | 384
no respiratory or neurologic symptoms | 384