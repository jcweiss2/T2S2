69 years old | 0
male | 0
hyperlipidemia | 0
hypertension | 0
bioprosthetic mitral valve replacement | -8760
admitted to the hospital | 0
left parietal hemorrhage | 0
left middle cerebral artery stroke | -336
thrombectomy | -336
sedated | 0
intubated | 0
external ventricular drain | 0
mild fatigue | -24
headache | -24
warfarin | -336
aspirin | -336
rosuvastatin | -336
III/IV holosystolic murmur | 0
transesophageal echocardiogram | 0
mobile echodensities on the posterior mitral valve leaflet | 0
cefepime | 0
gentamicin | 0
vancomycin | 0
Aspergillus galactomannan antigen | 0
1,3-β-D-glucan | 0
Karius cell-free DNA plasma quantitative test | 0
liposomal amphotericin B | 0
voriconazole | 0
fungal blood cultures | 144
Aspergillus fumigatus | 144
right eye fungal endophthalmitis | 0
intravitreal voriconazole | 0
valve repair surgery | 0
combined antifungal therapy | 0
isavuconazole | 504
prolonged QTc | 504
renal insufficiency | 1200
micafungin | 1200
generalized weakness | 1680
failure to thrive | 1680
white blood cell count elevation | 1680
splenic infarcts | 1680
splenic abscess | 1680
wedge-shaped renal infarcts | 1680
septic emboli | 1680
hypotensive | 1692
vasopressor initiation | 1692
persistent mobile echodensity | 1692
acute embolic occlusions | 1692
worsening hypoxemia | 1692
intubation | 1692
mechanical ventilation | 1692
increased vasopressor requirements | 1692
transitioned to comfort measures | 1698
died | 1698