26 years old | 0
African American | 0
woman | 0
hospitalization for possible rheumatic fever | -672
pyrexia | -672
polyserositis | -672
cardiac tamponade requiring pericardial drainage | -672
pericarditis | -672
presented on July 19, 2013 | 0
progressive abdominal pain | -72
nausea | -72
vomiting | -72
diarrhea | -72
quit smoking | -672
family history of mild hypertension | -672
treated with colchicine 0.6 mg | 0
lisinopril 20 mg | 0
omeprazole 20 mg | 0
pantoprazole 40 mg | 0
ranitidine 150 mg | 0
tramadol 50 mg daily | 0
penicillin G 2.5 million units | 0
albuterol for shortness of breath | 0
tachycardia | 0
112 beats per minute | 0
2/6 systolic murmur | 0
severe leukocytosis | 0
hemoglobin 107 g/L | 0
serum albumin 28 g/L | 0
serum creatinine level 53 µmol/L | 0
urinalysis revealed 1+ protein | 0
severe abdominal pain | 0
pelvic pain | 0
computed tomography notable for colitis | 0
stable mild ascites | 0
sepsis | 0
Clostridium difficile colitis | 0
intravenous metronidazole | 0
fluids | 0
oral vancomycin | 0
admitted to the transitional intensive care unit | 0
nephrology consultation | 96
potential oliguric acute tubular necrosis | 96
possibly vasculitis | 96
serum creatinine level increased to 159 µmol/L | 96
leukocyte count increased to 60×109/L | 96
platelet count decreased to 71×109/L | 96
stable hemoglobin level | 96
prepped for percutaneous renal biopsy | 96
new-onset anemia | 96
hemolytic anemia | 96
schistocytes present on peripheral smear | 96
elevated lactate dehydrogenase | 96
diagnosis of thrombotic thrombocytopenic purpura | 96
initiated high-dose steroids | 96
daily plasma exchange | 96
ADAMTS13 level drawn | 168
transferred | 312
continued daily plasma exchange | 312
dialysis initiated | 312
mycophenolate mofetil initiated | 312
developed seizure disorder | 312
levetiracetam initiated | 312
vision loss | 312
bilateral retinal damage | 312
disc hemorrhages | 312
macular hemorrhages | 312
retinal hemorrhages in all four quadrants | 312
mid-periphery hemorrhages | 312
presumed irreversible damage | 312
considered vitrectomy | 312
considered injection of vascular endothelial growth factor inhibitors | 312
discharged | 312
receive dialysis | 312
plasma exchange three times weekly | 312
follow-up with retinal specialist | 312
bilateral central artery occlusion | 312
bilateral central vein occlusion | 312
vitreous hemorrhage | 312
blindness | 312
best-noted acuity of 1–2 feet | 312
received plasma exchange every other day | 936
dialysis three times weekly | 936
no improvement | 936
ADAMTS13 activity level 61% | 936
diagnosis of aHUS | 936
eculizumab initiated | 1224
renal indices began to improve | 1224
little interdialytic weight gain | 1224
increased urinary output | 1224
hemodialysis discontinued | 1704
plasma exchange discontinued | 1704
presented to emergency department with hypertensive emergency | 20208
altered mental status | 20208
potential TMA complication | 20208
eculizumab dosing schedule shortened to 12 days | 20208
retinal specialist noted eyes clearing | 13416
no additional therapies planned | 13416
improvement in sight | 13416
improvement in functional status | 13416
walked without assistance | 13416
continues to receive eculizumab 1200 mg every 12 days | 13416
platelet count 527×109/L | 13416
normal hemoglobin levels | 13416
normal LDH levels | 13416
serum creatinine level 139 µmol/L | 13416
