43 years old | 0
man | 0
admitted to the hospital | 0
ACTH-secreting pituitary carcinoma | 0
cerebellar metastases | 0
cervical drop metastases | 0
COVID-19 infection | 0
surgery | - multiple treatment modalities (assigned timestamp - weeks based on previous therapies, approximated to -672)
radiotherapy | -672
ketoconazole | -672
pasireotide | -672
cabergoline | -672
bilateral (subtotal) adrenalectomy | -672
temozolomide chemotherapy | -672
immune checkpoint inhibitors (ipilimumab and nivolumab) | -672
maintenance nivolumab | -672
ketoconazole 800 mg daily | -672
stabilized disease | 0
surgical resection of left adrenal remnant (planned but not done) | 0
consulted emergency department for severe respiratory complaints | 0
upper respiratory tract symptoms | -168 (1 week before admission)
progressive dyspnoea | -72 (3 days before admission)
tested positive for SARS-CoV-2 | -24 (day before admission)
O2 saturation 72% | 0
tachypnoea (40/min) | 0
bilateral pulmonary crepitations | 0
temperature 37.2°C | 0
blood pressure 124/86 mmHg | 0
pulse rate 112 bpm | 0
high-flow oxygen therapy | 0
O2 saturation 89% | 0
tachypnoea 35/min | 0
urgent intubation | 0
type 1 respiratory insufficiency | 0
PaO2 52.5 mmHg | 0
PaCO2 33.0 mmHg | 0
pH 7.47 | 0
P/F ratio 65.7 | 0
elevated C-reactive protein (275.7 mg/L) | 0
white blood cell count 7.1 × 10⁹/L | 0
72.3% neutrophils | 0
ACTH 213 ng/L | -672 (3 weeks prior)
cortisol 195 µg/L | -672
increased cortisol 547 µg/L | +504 (3 weeks after admission)
decreased ACTH 130 ng/L | +504
high-dose dexamethasone | 0
broad-spectrum antibiotics | 0
Serratia in sputum | 0
methicillin-susceptible Staphylococcus aureus | 0
Haemophilus influenzae | 0
thromboprophylaxis with tinzaparin | 0
block-replacement regimen | 0
ketoconazole restarted day 11 | +264
hydrocortisone supplementation | 0
metabolic acidosis | varies (multiple organ involvement)
acute renal failure | varies
continuous venovenous hemofiltration | varies
acute coronary syndrome type 2 | varies
septic thrombophlebitis | varies
critical illness polyneuropathy | varies
ventilator-associated pneumonia | + (readmission)
central line-associated bloodstream infection | + (readmission)
discharged | varies
