2-month-old | 0
male | 0
admitted to the hospital | 0
mild cough | -24
fever | -24
malaise | -24
close contact with brother | -24
born very preterm | -6720
low birth weight | -6720
hospitalized for neonatal pneumonia | -6720
coagulation dysfunction | -6720
intracranial hemorrhage | -6720
neonatal pathological jaundice | -6720
vaccinated with Bacillus Calmette-Guerin | -6720
symptomatic treatments | 0
mask oxygen inhalation | 0
piperacillin tazobactam | 0
ambroxol | 0
budesonide + ipratropium bromide atomization | 0
tachypnea | 24
low oxygen saturation | 24
transferred to PICU | 24
body temperature 37.3°C | 0
heart rate 172 beats per minute | 0
respiratory rate 56 breaths per minute | 0
blood pressure 96/50 mmHg | 0
puffy nose | 0
triple concave signs | 0
mild cyanosis of the lips | 0
Glasgow Coma Score 13 | 0
oxygen saturation 93% | 0
rough breath sounds | 0
wheezing in both lungs | 0
umbilical hernia | 0
anterior fontanelle bulge | 0
low response | 0
screaming after stimulation | 0
computed tomography scan of the chest | 0
multiple plaques, streaks, solid shadows, and indistinct reticular shadows in both lungs | 0
magnetic resonance imaging of the brain | 0
bilateral frontal, parietal, and temporal extracranial spaces slightly wider | 0
no obvious abnormality in the brain parenchyma | 0
echocardiography | 0
no abnormalities | 0
hemoglobin level 84 g/L | 0
red blood cell count 3.05 × 10^12/L | 0
white blood cell count 6.5 × 10^9/L | 0
neutrophil count 3.59 × 10^9/L | 0
lymphocyte count 2.16 × 10^9/L | 0
platelet count 280 × 10^9/L | 0
liver and kidney function tests normal | 0
diagnosed with respiratory failure | 0
diagnosed with severe pneumonia | 0
diagnosed with septic shock | 0
diagnosed with encephalopathy | 0
antibiotic therapy with meropenem, vancomycin, and levetiracetam | 0
worsening dyspnea | 3
groans | 3
gray face | 3
cold limbs | 3
speckles all over the body | 3
bilateral crackles | 3
capillary refill time 5 seconds | 3
oxygen saturation dropped to 54% | 3
lactate level 7.07 mmol/L | 3
procalcitonin 14.29 ng/mL | 3
invasive ventilator-assisted ventilation | 3
norepinephrine | 3
mannitol | 3
fructose glycerol | 3
immunoglobulin | 3
fresh frozen plasma | 3
viral nucleic acid extracted from BALF specimens | 0
multiplex quantitative real-time PCR assay for respiratory viruses | 0
negative results for respiratory viruses | 0
serological tests of Mycoplasma pneumonia, Chlamydia trachomatis, and cytomegalovirus | 0
negative results for Mycoplasma pneumonia, Chlamydia trachomatis, and cytomegalovirus | 0
sputum bacterial cultures | 0
negative results for sputum bacterial cultures | 0
tuberculin test | 0
negative results for tuberculin test | 0
detection of Bordetella from nasopharyngeal specimen | 0
Bordetella pertussis positivity | 0
confirmation of B pertussis by testing for ptxS1 | 0
CSF assay | 0
normal CSF assay results | 0
CSF cultures | 0
negative results for CSF cultures | 0
m-NGS of blood and CSF | 0
detection of B pertussis in blood and CSF by m-NGS | 0
intravenous levofloxacin | 48
chest x-ray | 48
inflammation in the lungs gradually absorbed | 312
weaned off mechanical ventilation | 312
discharged | 888
full recovery | 888