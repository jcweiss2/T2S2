73 years old | 0
male | 0
admitted to the emergency department | 0
previous history of bioprosthetic aortic valve replacement | -3600
bioprosthetic aortic valve replacement | -3600
active endocarditis | 0
cardiogenic shock | 0
prosthetic heart valve failure | 0
acute aortic regurgitation | 0
infective endocarditis | 0
B-cell lymphoma | 0
ongoing chemotherapy | 0
evaluation of the acute clinical situation | 0
pre-existing comorbidities | 0
heart team recommendation | 0
TAVR as the treatment option of choice | 0
time window of at least 72 hours after negative blood culture results | 0
negative blood culture results | -72
transfemoral valve-in-valve TAVR | 168
balloon-expandable Edwards Sapien 3 heart valve | 168
general anesthesia | 168
excellent immediate procedural result | 168
full recovery | 168
prolonged suppressive antibiotic therapy | 168
management of patients with infective endocarditis | 0
multidisciplinary approach | 0
infectious disease specialists | 0
cardiologists | 0
cardiac surgeons | 0
identification of patients at specific risk | 0
embolic stroke | 0
systemic embolization | 0
septic shock | 0
intensive care treatment | 0
pathoanatomical presentation of infective endocarditis | 0
microorganism involved | 0
valves affected by minor bacterial colonization | 0
mobile and floating vegetations | 0
abscess or fistula formation | 0
leaflet or cusp destruction | 0
prosthetic heart valve disease | 0
diagnosis and decision making | 0
specialized reference centers | 0
local and experienced endocarditis expert team | 0
distinct differentiation between destructive infective heart valve endocarditis and prosthetic heart valve failure | 0
concomitant septicemia of a different origin | 0
refined imaging technologies | 0
dedicated algorithm for the diagnosis of prosthetic heart valve endocarditis | 0
transthoracic echocardiography | 0
transesophageal echocardiography | 0
first-line imaging technologies | 0
sensitivity of these tools for a conclusive evaluation | 0
exclusion of infective endocarditis | 0
multidetector-row computed tomography (CT) | 0
functional imaging with fluorine-18–fluoro-2-deoxyglucose (FDG) positron emission tomography (PET)/CT | 0
diagnosis of infective endocarditis | 0
inflammatory cells | 0
morphologic changes | 0
Duke criteria | 0
possible infective endocarditis | 0
radiolabeled white blood cell single-photon emission CT | 0
perivalvular lesions | 0
interdisciplinary decision to perform TAVR | 0
clinical parameters | 0
2020 joint American College of Cardiology and American Heart Association guideline | 0
management of patients with valvular heart disease | 0
optimal therapy for cardiac device–related infective endocarditis | 0
complete device extraction | 0
prolonged course of parenteral antibiotic therapy | 0
incomplete removal and sterilization of affected valvular structures | 0
relapsing infections | 0
recurrent endocarditis | 0
deep tissue infection | 0
TAVR as bailout strategy | 0
rescue therapy | 0
short-term setting of confirmed infective endocarditis | 0
cardiogenic shock secondary to severe aortic regurgitation | 0
inoperable patients | 0
bridge to definitive surgical repair | 0
initiation of TAVR as early as possible | 0
multiorgan failure | 0
reversible | 0
maximal clinical and prognostic benefit | 0
right timing | 0
central challenge of the heart team | 0
sterile blood culture results | 0
procedural considerations | 0
use of cerebral filter devices | 0
procedural safety measure | 0
septic cerebral embolism | 0
frequent monitoring | 0
prolonged antibiotic treatment | 0
cardiac radionuclide imaging | 0
duration of suppressive antibiotic therapy | 0
monitor treatment success | 0
international guideline recommendations | 0
treatment of prosthetic heart valve failure secondary to active infective endocarditis | 0
transcatheter heart valve technologies | 0
well-selected patients | 0
success story of this case report | 0
fortune favors the bold or brave | 0
new chapter in the success story of TAVR | 0
literature needs to advise future guideline recommendations | 0
research grants to the institution | 0
Edwards Lifesciences | 0
Medtronic | 0
Abbott Vascular | 0
Guerbet AG | 0
Boston Scientific | 0
consultant to Boston Scientific | 0
BTG | 0
Teleflex | 0
human studies committees | 0
animal welfare regulations | 0
Food and Drug Administration guidelines | 0
patient consent | 0