19 years old | 0
male | 0
admitted to the hospital | 0
alcohol addiction | -8760
Tourette syndrome | -8760
sleepiness | 0
unclear speech | 0
drinking bout | -72
pneumonia | 0
intubation | 0
mechanical ventilation | 0
numerous vegetations on the heart valves | 0
transfer to intensive care unit | 0
midazolamum | 0
fentanyl | 0
grade 4 mitral insufficiency | 0
vegetation on the anterior cusp | 0
rupture of the tendinous cords | 0
vegetation on the posterior cusp | 0
marginal thickening of the aortic valve | 0
grade 1 insufficiency of the aortic valve | 0
tricuspid valve insufficiency | 0
central regurgitation jet | 0
suspected vegetation on the tricuspid valve | 0
empiric antibiotic therapy | 0
imipenem | 0
vancomycin | 0
clindamycinum | 0
sterile bacteriological analysis | 0
dental consultation | 0
inflammatory foci in the oral cavity | 0
extraction of 8 carious teeth | 0
mobile vegetations on the valves | 168
embolization risk | 168
surgical procedure | 168
extracorporeal circulation | 168
median sternotomy | 168
aortic cross-clamping | 168
cardioplegic solution | 168
tricuspid valve removal | 168
mitral valve removal | 168
aortic valve removal | 168
implantation of valve bioprostheses | 168
Medtronic Hancock II Porcine 29 | 168
Edwards Lifesciences C-E Perimount 21 | 168
Medtronic Hancock II Porcine 33 | 168
recovery room | 340
hemodynamically stable | 340
moderate doses of catecholamines | 340
mediastinal drains removal | 72
intensive care unit | 72
antibiotic therapy | 72
sterile cultures from blood and valves | 72
extubation | 336
sepsis | 552
high fever | 552
Pseudomonas aeruginosa | 552
central venous catheter | 552
urine | 552
bronchial secretions | 552
targeted antibiotic therapy | 552
imipenem | 552
Brulamycin | 552
no clinical improvement | 552
vegetation on the aortic valve bioprosthesis | 552
transesophageal echocardiography | 552
computed tomography | 552
X-ray | 552
reoperation | 1104
aortic valve bioprosthesis replacement | 1104
Edwards Lifesciences C-E Perimount 21 | 1104
recovery room | 1144
extubation | 1163
antibiotic therapy | 1163
Pseudomonas aeruginosa | 1163
sterile bacteriological tests | 1163
cardiac rehabilitation hospital | 1264
oral anticoagulation | 1264
antibiotic therapy | 1264
control echocardiographic examination | 1456
normal function of all bioprostheses | 1456