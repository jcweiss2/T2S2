35 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
gave birth to healthy twins | -24 | -24 | Factual
in vitro fertilization | -280 | -280 | Factual
facial nerve paresis | -672 | 0 | Factual
severe headache | 24 | 24 | Factual
generalized tonic–clonic seizures | 24 | 26 | Factual
loss of consciousness | 24 | 26 | Factual
arterial blood pressure 195/110 mmHg | 24 | 24 | Factual
heart rate 120 beats/min | 24 | 24 | Factual
eclampsia | 24 | 24 | Factual
antihypertensive therapy | 24 | 120 | Factual
magnesium sulphate | 24 | 24 | Factual
ebrantil | 24 | 24 | Factual
20% manitol | 24 | 24 | Factual
diazepam | 24 | 24 | Factual
bilateral vision loss | 48 | 48 | Factual
proteinuria 2+ | 48 | 48 | Factual
normal complete blood count | 48 | 48 | Factual
normal liver function tests | 48 | 48 | Factual
normal clotting parameters | 48 | 48 | Factual
normal electrocardiogram | 48 | 48 | Factual
cortical blindness | 48 | 120 | Factual
mild right-sided facial nerve paresis | 48 | 120 | Factual
hypodensity of the posterior white matter | 72 | 72 | Factual
vasogenic edema | 72 | 120 | Factual
T2- and fluid-attenuated inversion recovery-weighted images hyperintense signals | 72 | 72 | Factual
hyperintense signals in the white matter | 72 | 72 | Factual
parietal and occipital regions | 72 | 72 | Factual
junctions of vascular watershed zones of the brain | 72 | 72 | Factual
stabilization of the general condition | 72 | 120 | Factual
oral antihypertensive medication | 120 | 192 | Factual
enalapril maleate | 120 | 192 | Factual
methyldopa | 120 | 192 | Factual
human albumin | 120 | 120 | Factual
bilateral improvement of the visual function | 120 | 120 | Factual
best-corrected visual acuity 1.0 | 120 | 120 | Factual
peripheral relative scotoma | 120 | 120 | Factual
depressed sensitivity of the paracentral left visual field | 120 | 120 | Factual
regression of the edema | 192 | 192 | Factual
discrete residual changes over the posterior horns of the side ventricles | 192 | 192 | Factual
discharge from the clinic | 216 | 216 | Factual
oral antihypertensive therapy | 216 | 0 | Factual
physical therapy for the paresis of the facial nerve | 216 | 0 | Factual