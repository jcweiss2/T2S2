42 years old | 0
male | 0
admitted to the hospital | 0
generalized weakness | -2160
fever | -2160
cough | -2160
weight loss | -2160
HIV-antibody test positive | -2160
sputum AFB smear positive | -2160
lived in Guatemala | -8760
HIV-1 Western blot test positive | -40
CD4 cell count 10/µL | -40
HIV RNA titer 18,000 copies/mL | -40
anti-tuberculosis medications started | -40
fluconazole started | -40
trimethoprim/sulfamethoxazole started | -40
generalized weakness persisted | 0
fever persisted | 0
oral thrush | 0
hepatosplenomegaly | 0
ascites | 0
hemoglobin 10.6g/dL | 0
white blood cell 2,700/µL | 0
platelet 58,000/µL | 0
total bilirubin 2.4mg/dL | 0
AST/ALT 131/48IU/L | 0
ALP 114IU/L | 0
GGT 133 IU/L | 0
costophrenic angle blunting | 0
fluid shifting in the right hemithorax | 0
mild pneumonic infiltration in left lung | 0
disseminated tuberculosis suspected | 0
anti-retroviral agents started | 0
pancytopenia progressed | 24
hemoglobin 7.4g/dL | 24
white blood cell 1,070/µL | 24
platelet 13,000/µL | 24
rifampin discontinued | 24
zidovudine discontinued | 24
trimethoprim/sulfamethoxazole discontinued | 24
new pulmonary infiltrates | 120
septic shock | 120
empirical antibiotic therapy started | 120
piperacillin/tazobactam started | 120
mechanical ventilator support started | 144
bone marrow aspiration and biopsy performed | 216
Histoplasma capsulatum identified | 216
died | 240
refractory septic shock | 240
hypoxia | 240