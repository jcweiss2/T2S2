63 years old | 0
male | 0
presented to emergency department | 0
right sided hemiparesis | -78
altered mental status | -78
NIH stroke scale 18 | 0
stroke alert called | 0
driving | -102
became confused | -102
aphasic | -102
right upper and lower extremity hemiparesis | -102
non-contrast CT scan of the brain negative | 0
chronic opacification of left mastoid air cells | 0
fluid in mastoid air spaces bilaterally | 0
CT angiography head and neck | 0
no hemodynamically significant findings | 0
no flow limiting arterial stenosis | 0
contrast-enhanced perfusion CT brain negative | 0
tissue plasminogen activator not given | 0
worsening encephalopathy | 0
intubated for airway protection | 0
fever 103 degrees Fahrenheit | 2
heart rate increased to 120 bpm | 2
dilated non-reactive right pupil | 2
repeat NCCT scan of the brain | 2
rapidly developing white matter edema | 2
pons edema | 2
no specific etiology | 2
cranial nerve III involvement | 2
lumbar puncture attempted | 2
lumbar puncture not completed | 2
consult interventional radiology | 2
cerebrospinal fluid obtained | 2
intravenous vancomycin | 2
ceftriaxone | 2
ampicillin | 2
acyclovir | 2
white blood cell count 15,200/μL | 2
lactic acid 3.2 mmol/L | 2
severe sepsis | 2
admitted to ICU | 2
intubated and sedated | 2
cerebrospinal fluid analysis 3,278 WBC/μL | 2
neutrophils 98% | 2
glucose <1 mg/dL | 2
total protein 670 mg/dL | 2
gram-positive cocci in chains | 2
Streptococcus pneumoniae | 2
acute on chronic mastoiditis | 2
consult otolaryngology | 2
left myringotomy with tympanostomy tube | 2
cranial nerve palsy resolved | 2
sensitivities reported | 72
ceftriaxone 2g twice a day | 72
dexamethasone four days | 72
follow-up NCCT improved | 72
weaned off sedation | 96
neurologically stable for extubation | 96
encephalopathy resolved | 96
right sided motor weakness resolved | 96
transferred to general medical floor | 96
diabetes mellitus 2 | 0
bilateral mastoidectomies | -8760
progressive left ear pain | -72
acute left-sided mastoiditis | 0
sustained full neurologic recovery | 0
discharged | 96
