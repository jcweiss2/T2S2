54 years old | 0
female | 0
type 2 diabetes | 0
hypertension | 0
peripheral vascular disease | 0
right-foot transmetatarsal amputation | -26208
lisinopril | 0
metoprolol succinate | 0
pravastatin | 0
aspirin | 0
hydrochlorothiazide | 0
metformin | 0
insulin detemir | 0
insulin lispro discontinued | -24
hypoglycemia | 0
glucagon administered | 0
confusion | 0
hypotension | 0
blood pressure 70/39 mmHg | 0
disorientation | 0
dry oral mucosa | 0
decreased bowel sounds | 0
unresponsive | 0
cardiopulmonary arrest | 0
pulseless electrical activity | 0
cardiopulmonary resuscitation | 0
endotracheal intubation | 0
mechanical ventilation | 0
spontaneous circulation | 3
norepinephrine infusion | 0
blood pressure 98/37 mmHg | 0
arterial pH 6.57 | 0
HCO3- 2 mEq/L | 0
anion gap 30 mmol/L | 0
osmolar gap 21 | 0
lactate 16.3 mmol/L | 0
glycosylated hemoglobin 7.3 mg/dL | 0
creatinine 8.07 mg/dL | 0
computed tomography scan | 0
gallbladder wall thickening | 0
vasopressin infusion | 0
differential diagnosis | 0
suspected sepsis | 0
suspected acute coronary event | 0
metformin toxicity diagnosis | 0
impaired renal function | 0
mechanical ventilation continued | 0
norepinephrine continued | 0
vasopressin continued | 0
hemodialysis initiated | 0
acidemia resolved | 0
hemodynamics improved | 0
norepinephrine reduced | 0
vasopressin reduced | 0
blood culture negative | 0
stool culture negative | 0
elevated troponin 4.42 ng/mL | 0
serial electrocardiograms negative | 0
echocardiogram | 24
ejection fraction 50% | 24
norepinephrine discontinued | 96
vasopressin discontinued | 96
extubation | 144
metformin concentration 42 mcg/mL | 168
discharged from ICU | 216
discharged from hospital | 360
dialysis discontinued | -720
serum creatinine 0.86 mg/dL | -1440
grandson's gastroenteritis | -72
nuclear stress test abnormal | 360
coronary angiography | 360
three-vessel disease | 360
coronary artery bypass graft | 360
Pressors discontinued on day 4 (96 hours), extubated on day 6 (144), metformin level back on day 7 (168), ICU discharge on day 9 (216), hospital discharge on day 15 (360). Dialysis discontinued within a month post-discharge, so that's after hospital discharge, timestamp 360 + (up to 720), but the assistant uses -720. Wait, the assistant's entry has "dialysis discontinued | -720", which doesn't make sense because discontinuation happened after discharge. Maybe it's a mistake. Alternatively, the serum creatinine two months prior was 0.86, which is -1440 hours (2 months ≈ 8 weeks, 8*7*24=1344, but 2 months is approx 8.67 weeks, so 1440 hours). So that's timestamp -1440.
hypertension |2 0
HCO36 2 mEq/L | 0
