36 years old | 0
    male | 0
    hypertension | -26208
    systemic lupus erythematosus | -26208
    systemic vasculitis | -26208
    coronary artery disease | -26208
    3-vessel coronary artery bypass graft | -26208
    seizure disorder | -26208
    superior vena cava syndrome | -26208
    end-stage renal disease | -26208
    hemodialysis | -26208
    multiple dialysis catheter placements | -26208
    transhepatic central catheter | -26208
    infected multiple times | -26208
    multiple intensive care unit admissions | -26208
    sepsis | -26208
    disseminated intravascular coagulation | -26208
    bacteremia | -26208
    vancomycin-resistant Enterococcus | -26208
    extended-spectrum beta-lactamase-producing Klebsiella | -26208
    required multiple antibiotics | -26208
    cefepime | -26208
    linezolid | -26208
    syncopal episode | 0
    complete heart block | 0
    junctional escape rhythm | 0
    heart rate 35 beats per minute | 0
    transesophageal echocardiogram | 0
    mildly sclerosed mitral and aortic valves | 0
    mild-to-moderate mitral regurgitation | 0
    mild-to-moderate tricuspid regurgitation |9 0
    normal LV function | 0
    no regional wall motion abnormalities | 0
    attempted Micra leadless pacemaker implantation | 0
    right ventricle access attempt | 0
    common iliac veins completely occluded | 0
    right internal jugular vein access attempt | 0
    superior vena cava chronically occluded | 0
    computed tomography scan confirmation | 0
    transhepatic approach discussed | 0
    transhepatic catheter infection history | 0
    methicillin-resistant Staphylococcus aureus | -26208
    vancomycin-resistant enterococcus | -26208
    multiple transhepatic catheter infections | -26208
    surgical epicardial pacing decision | 0
    left anterolateral minithoracotomy | 0
    fifth intercostal space incision | 0
    sixth rib resection | 0
    epicardial leads placed | 0
    no capture | 0
    frailty of myocardium | 0
    suture-on bipolar lead placed | 0
    acceptable thresholds (~2 mV) | 0
    lead failure next day | 24
    complete heart block persisted | 24
    junctional escape rhythm persisted | 24
    temporary transvenous pacing wire placed | 24
    transhepatic RV pacing | 24
    FDA compassionate use plea | 24
    institutional review board approval | 24
    WiSE-CRT device provided | 24
    transmitter and battery implantation | 24
    general anesthesia | 24
    fourth intercostal space incision | 24
    midaxillary incision | 24
    subcutaneous tunnel created | 24
    WiSE-CRT transmitter placement | 24
    battery pocket creation | 24
    hemostasis achieved | 24
    electrode insertion phase | 24
    right femoral artery access | 24
    12F sheath insertion | 24
    retrograde LV access | 24
    transesophageal echocardiogram guidance | 24
    heparinization | 24
    activated coagulation time maintenance | 24
    deflectable sheath insertion | 24
    LV lateral wall placement | 24
    receiver electrode deployment | 24
    barb deployment confirmation | 24
    sheath withdrawal | 24
    device programming | 24
    pacing capture confirmed | 24
    heparin reversal | 24
    arterial access closure | 24
    LV pacing success | 24
    intra-abdominal infection | 336
    sepsis secondary | 336
    death | 336