50 years old | 0
female | 0
severe lower abdominal pain | -120
nausea | -120
vomiting | -120
fever | -120
constipation | -120
history of hypertension | 0
history of dyslipidemia | 0
history of heart failure | 0
history of rheumatologic disease | 0
taking furosemide | -6720
taking captopril | -6720
taking spironolactone | -6720
taking prednisone | -14400
taking sodium diclofenac | -24
admitted to the hospital | 0
ill-looking cushingoid and pale patient | 0
cyanotic extremities | 0
decreased tissue perfusion | 0
marked lower limbs edema | 0
slightly disoriented | 0
blood pressure = 50/30 mmHg | 0
pulse = 110 beats/minute | 0
respiratory rate = 24 respiratory movements/minute | 0
axillary temperature = 37 °C | 0
abdomen distended and diffusely tender | 0
bowel sounds decreased | 0
rebound tenderness test negative | 0
liver palpable up to 1 cm below the right costal margin | 0
extracellular volume repletion with saline | 0
ceftriaxone | 0
metronidazole | 0
hydrocortisone | 0
noradrenaline | 0
referred to the intensive care unit (ICU) | 0
initial laboratory workup | 0
Hemoglobin = 12.6 g/dL | 0
Creatinine = 2.9 mg/dL | 0
Hematocrit = 37.4% | 0
Potassium = 4.7 mEq/L | 0
Leucocytes = 19100/mm3 | 0
Sodium = 110 mEq/L | 0
Bands = 17% | 0
ALT = 28 U/L | 0
Segmented = 72% | 0
AST = 44 U/L | 0
Eosinophils = 1% | 0
LDH = 336 U/L | 0
Basophils = 0% | 0
CK = 933 U/L | 0
Lymphocytes = 8% | 0
Amylase = 11 U/L | 0
Monocytes = 2% | 0
Lipase = 15 U/L | 0
Platelets = 382.103/mm3 | 0
Total protein = 4.9 g/dL | 0
CRP = 142 mg/L | 0
Albumin = 2.3 g/dL | 0
BUN = 62 mg/dL | 0
PT (INR) = 1.21 | 0
abdominal ultrasound | 0
minimal amount of free fluid in the abdominal cavity | 0
diffuse and marked decrease of the small bowel peristaltic movements | 0
liquid distention | 0
anti-HIV serology negative | 0
hemodynamically unstable | 0
continuous administration of norepinephrine | 0
continuous administration of vasopressin | 0
petechiae and ecchymoses on the abdomen and upper limbs | 72
mental status worsened | 72
orotracheal intubation | 72
mechanical ventilation | 72
Multi sensitive E. coli isolated in the blood culture | 72
died on the fourth day of hospitalization | 96
autopsy | 96
petechial skin lesions on abdominal wall and limbs | 96
generalized edema of the limbs | 96
mild ascites | 96
larvae of S. stercoralis in the dermis of the skin lesions | 96
foci of hemorrhage | 96
diffuse alveolar damage | 96
septic shock | 96
multiple areas of recent and previous alveolar hemorrhage | 96
hemosiderin-laden macrophages | 96
S. stercoralis larvae in the interstitium of the lung | 96
giant cell granulomatous reaction | 96
flat lesions consistent with healing ulcers in small bowel mucosa | 96
petechial foci of hemorrhage in small bowel mucosa | 96
multiple small foci of hemorrhage on abdominal serous surfaces | 96
S. stercoralis larvae in duodenal mucosa | 96
S. stercoralis larvae in omentum | 96
acute hematogenous pyelonephritis | 96
multiple small subcapsular abscesses | 96
bacterial hematogenous spread in the spleen | 96
acute inflammation | 96
septic emboli | 96
areas of acute infarction | 96
systemic findings of sepsis and shock | 96
lipid depletion and hemorrhagic foci in adrenal glands | 96
necrosis on zone 3 in liver | 96
acute tubular necrosis in renal cortex | 96
foci of ischemic pancreatitis | 96
diffuse dilatation of chambers and softening of the myocardium | 96
focal hyaline thrombi | 96
disseminated intravascular coagulation | 96
S. stercoralis hyperinfection syndrome | 96
Gram-negative bacterial septicemia | 96
septic shock | 96