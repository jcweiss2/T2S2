63 years old | 0
female | 0
smoker | 0
chronic obstructive pulmonary disease | 0
admitted to the emergency department | 0
dyspnea | 0
dysphasia | 0
vaccinated with 3rd dose of BNT162b2mRNA | -360
SARS-CoV-2 PCR positive | 0
percutaneous transluminal angioplasty | -192
left anterior tibial posterior occlusion | -192
conscious but not cooperative | 0
lower extremity pulses could not be obtained | 0
arterial blood pressure 120/60 mm Hg | 0
heart rate 120/min | 0
respiratory rate 24/min | 0
body temperature 36.5℃ | 0
O2 saturation 90% | 0
sinus tachycardia | 0
diffuse atherosclerosis | 0
thrombotic events | 0
multiple embolic infarcts in the left temporal and bilateral frontal lobes | 0
stenosis of bilateral internal carotid arteries less than 50% | 0
embolism in the right lower lobe and segmental pulmonary artery branches | 0
minimal consolidation area in the left lung lower lobe | 0
pericardial effusion | 0
left ventricular ejection fraction 60% | 0
acute thrombosis of the ulnar vein in the proximal right upper extremity | 0
crural artery circulation could not be clearly defined | 0
subacute deep vein thrombosis in the bilateral main femoral vein | 0
non-invasive mechanical ventilation support | 0
pleural fluid drained through the catheter | 0
enoxaparin sodium 6,000 IU administered twice a day | 0
iloprost and asetilsalisilik asit treatment | 0
high D-Dimer | 0
normal platelets | 0
vasculitis markers negative | 0
cardiovascular surgeon stated acute arterial thrombosis and necrosis in both lower extremities | 0
both lower extremities amputated below the knee | 0
transferred to the service | 0
discharged home from the ward | 0
readmitted to another hospital 2 days later | 48
died on the 13th day of hospitalization | 312