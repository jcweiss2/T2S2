23 years old | 0
male | 0
asthma | 0
remote substance abuse | 0
seizures | -1
vaping | -1
tachycardic | 0
tachypneic | 0
hypoxic | 0
altered mental status | 0
inability to follow commands | 0
subcostal retractions | 0
diffuse rhonchi | 0
respiratory acidosis | 0
intubated | 0
leukocytosis | 0
creatinine 1.69 | 0
sinus tachycardia | 0
bilateral upper lobe collapse | 0
sepsis | 0
systemic inflammatory response syndrome (SIRS) | 0
extubated | 24
electroencephalogram unremarkable | 24
treated with levetiracetam | 24
renal function improved | 96
discharged | 120
vaping use | -1
EVALI | 0
bilateral upper lobe collapse/atelectasis | 0
respiratory failure | 0
ventilator support | 0 
midazolam administered | -1 
non-rebreather mask | 0 
afebrile | 0 
CT chest confirmed bilateral upper lobe collapse | 0 
CT brain unremarkable | 0 
blood cultures negative | 0 
cerebral spinal fluid cultures negative | 0 
viral tests negative | 0 
seizure activity free | 24 
intravenous fluids | 0 
no infectious etiology identified | 0 
high index of suspicion of vaping/e-cigarette use | 0 
young age | 0 
lack of prior lung injury | 0 
lack of comorbidities | 0 
extensive workup | 0 
diagnosis of exclusion | 0 
cessation and patient education | 120 
lung injuries | 0 
younger patients using vaping products | 0 
continued discussion between patient and physician | 120