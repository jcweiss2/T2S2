77 years old | 0
male | 0
schizophrenic | 0
admitted to the hospital | 0
abdominal distension | -168
diarrhea | -168
incontinence | -24
infrequent vomiting | -168
weight loss | -168
anorexia | -168
no abdominal pain | 0
mild metabolic alkalosis | 0
elevation of C-reactive protein | 0
normal complete blood count | 0
normal electrolytes panel | 0
normal liver function tests | 0
computed tomography (CT) of the abdomen | 0
contracted gallbladder | 0
gallstones | 0
gas bubbles in gallbladder | 0
suspected cholecystocolonic fistula | 0
admitted for observation | 0
serial abdominal examination | 0
persistent abdominal distension | 0
persistent diarrhea | 0
Hepatobiliary Imino-Diacetic Acid (HIDA) scan | 120
occlusion of the cystic duct | 120
Endoscopic Retrograde Cholangiography (ERC) | 120
sphincterotomy | 120
pancreatic stent placement | 120
fevers | 20
hypotension | 20
tachycardia | 20
transferred to Intensive Care Unit (ICU) | 20
CT scan of the abdomen | 20
free intraabdominal fluid | 20
normal Serum Amylase and Lipase levels | 20
open abdominal exploration | 24
fistulous tract between gallbladder and hepatic flexure | 24
division of fistulous tract | 24
retrieval of two stones from gallbladder | 24
biopsy of exposed colonic mucosa | 24
frozen section analysis | 24
absence of neoplastic changes | 24
partial cholecystectomy | 24
fulguration of remaining mucosa | 24
tangential resection of hepatic flexure | 24
external drainage tube placement | 24
hospitalization for two weeks | 168
episodic nocturnal desaturation | 168
central sleep apnea | 168
discharge from hospital | 168
right upper quadrant abscess | 504
treatment with antibiotics | 504
percutaneous drainage | 504
uneventful follow-up | 876