39 years old| 0
woman| 0
systemic lupus erythematosus (SLE)| -8760
immune thrombocytopenic purpura| -8760
fatigue| -8760
abdominal pain| -8760
severe thrombocytopenia (platelets 5 × 10^9/L)| -8760
multiple platelet transfusions| -8760
intravenous methylprednisolone| -8760
intravenous immunoglobulin (IVIg)| -8760
splenectomy| -8760
refractory thrombocytopenia| -8760
intra-abdominal hematoma| -8760
ischemic left foot| -8760
below-the-knee amputation| -8760
SLE exacerbation| -8760
enterocolitis| -8760
sepsis| -8760
transfer to intensive care unit| -8760
deterioration| -8760
sloughing| -8760
profound hypotension| -8760
transfer to our hospital at day 36| 0
temperature 31.5°C| 0
heart rate 87| 0
blood pressure 90-100/405-50 mm Hg| 0
blood oxygen saturation 99% (FiO2 40%)| 0
admitted to burn intensive care unit| 0
confluent dusky Nikolsky-positive plaques on face| 0
confluent dusky Nikolsky-positive plaques on neck| 0
confluent dusky Nikolsky-positive plaques on breasts| 0
confluent dusky Nikolsky-positive plaques on arms| 0
upper chest denudation| 0
abdomen denudation| 0
mons pubis denudation| 0
upper left leg denudation| 0
right leg dusky patches in reticulate pattern| 0
crusted erosions on lips| 0
crust on conjunctiva| 0
greater than 90% total body surface area denuded or Nikolsky positive| 0
severe lactic acidosis| 0
anemia (hemoglobin 5.3g/dL)| 0
thrombocytopenia (platelets 42 × 10^9/L)| 0
coagulopathy| 0
international normalized ratio 1.3| 0
prothrombin time 15.1| 0
partial thromboplastin time 60.5| 0
decreased protein S level (27%)| 0
right femoral vein deep venous thrombosis| 0
multifocal renal cortical infarctions| 0
started on IV methylprednisolone| 0
continuous renal replacement therapy| 0
mitral valve thickening| 0
noninfectious mitral valve thickening| 0
started on ciprofloxacin| 0
started on gentamycin| 0
started on vancomycin| 0
started on prophylactic heparin| 0
biopsy showing full-thickness epidermal necrosis| 0
biopsy showing microvascular thrombi| 0
additional samples showing resolving interface dermatitis| 0
thrombotic vasculopathy| 0
acute SLE flare| 0
concern for catastrophic anti-phospholipid antibody syndrome| 0
concern for acute lupus flare| 0
started on plasma exchange| 0
started on IVIg| 0
started on mycophenolate mofetil| 0
negative anticardiolipin antibodies| 0
negative anti-β2 glycoprotein I antibodies| 0
negative antiphosphatidylserine antibodies| 0
fever| 0
ventilator-associated pneumonia| 0
increasing ventilator requirements| 0
vancomycin-resistant Enterococcus bacteremia| 0
withdrawal of life-sustaining therapies| 0
autopsy determined cause of death as refractory hypotension| 0
third spacing from massive fluid losses| 0
toxic epidermal necrolysis involving >90% total body surface area| 0
acute hemorrhagic pancreatitis| 0
extensive necrosis| 0
fat necrosis along bowel mesentery and omentum| 0
widespread vesiculobullous dermatitis| 0
hypercoagulability| 0
anti-nuclear antibody-like syndrome| 0
received amphotericin B| -8760
received piperacillin/tazobactam| -8760
received cefazolin| -8760
Nikolsky-positive lesions| 0
denudation encompassing >90% total body surface area| 0
lower extremity livedo reticularis| 0
potential antiphospholipid antibody syndrome| 0
multiple thrombotic events| 0
renal infarctions| 0
ischemic leg requiring amputation| 0
deep venous thrombosis| 0
microvascular thrombi| 0
thrombotic storm| 0
lack of response to treatment| 0
ASAP (acute syndrome of apoptotic pan-epidermolysis)| 0
full-thickness epidermal necrosis| 0
rapid progression of ASAP| 0
concurrent severe hypercoagulability| 0
