24 years old | 0
female | 0
primiparous | 0
no significant medical history | 0
normal delivery | -504
depressive mood | -168
emotional incontinence | -168
auditory hallucination | -168
abnormal behavior | -168
hospitalized | -168
diagnosed with postpartum psychosis | -168
treated with antipsychotic drugs | -168
somnolence | -160
unstable breathing | -160
generalized seizure | -160
status epilepticus | -160
hyperthermia | -160
transferred to intensive care unit | -160
treated with methylprednisolone | -160
treated with intravenous immunoglobulin | -160
involuntary movements | -144
orofacial dyskinesia | -144
athetoid movement | -144
fever | -144
inflammatory reaction | -144
mild liver dysfunction | -144
lymphocytic pleocytosis | -144
elevated protein level | -144
normal glucose level | -144
anti-NMDAR antibody positive | -144
diffuse beta activity | -144
high-voltage rhythmic delta bursts | -144
abdominal computed tomography | -144
ovarian cystic tumor | -144
diagnosed with anti-NMDAR encephalitis | -144
laparoscopic removal of ovarian tumor | 1008
treated with IVIg | 1008
treated with mPSL pulse therapy | 1008
treated with plasma exchange | 1008
treated with double filtration plasmapheresis | 1008
involuntary movements improved | 1344
respiratory failure improved | 1344
transferred to rehabilitation hospital | 1344
severe cognitive dysfunction | 1344
memory disturbance | 2016
mental juvenility | 2016
independent gait | 2016
verbal communication | 2016
no brain atrophy | 2016
no abnormal signals | 2016