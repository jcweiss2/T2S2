83 years old | 0
male | 0
admitted to the hospital | 0
prostatic cancer | -8760
diabetes mellitus | -8760
hypertension | -8760
hyperuricemia | -8760
compression fracture of L2 vertebra | -840
taking painkillers | -840
lower back pain | -840
tenderness in left thigh | 0
stabbing pain in left thigh | 0
erythematous rash | 0
heart rate of 140 beats/min | 0
respiratory rate of 39 breaths/min | 0
percutaneous arterial oxygen saturation of 89 % | 0
oxygen therapy via nasal cannula at 2 L/min | 0
white blood cell count of 30,600 cells/mm3 | 0
neutrophils of 92.9 % | 0
hemoglobin of 10.9 g/dL | 0
creatinine of 2.48 mg/dL | 0
C-reactive protein of 42.72 mg/dL | 0
procalcitonin of 29.69 ng/mL | 0
glucose level of 156 mg/dL | 0
glycated hemoglobin level of 6.1 % | 0
massive pleural effusion in left thoracic cavity | 0
fluid retention in left iliopsoas muscle | 0
air extending to lower limb | 0
inflammation in retroperitoneal cavity | 0
Sequential Organ Failure Assessment (SOFA) score of 6 | 0
rapid infusion | 0
pressor agents | 0
intravenous meropenem | 0
thoracotomy tube insertion | 0
pleural effusion drainage | 0
abscess incision and drainage | 0
catheter insertion into retroperitoneal cavity | 0
continuous hemodiafiltration | 0
ventilator control | 0
meropenem | 0
clindamycin | 0
died of multiple organ failure | 72
necrotizing fasciitis | 72
myositis | 72
neutrophil infiltration | 72
gram-positive bacteria | 72
anaerobic culture of pleural effusion | 24
blood culture | 72
gene sequencing | 96
identification of P. micra | 96
P. micra infection | 0