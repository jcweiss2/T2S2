30 years old | 0
primigravida | 0
intrauterine fetal death | -672
induction of labor | 0
amniotic fluid embolism | 0
acute STEMI | 0
mifepristone administration | 0
misoprostol administration | 0
epidural catheter placement | 0
dizziness | 1
emesis | 1
convulsive seizure | 1
magnesium administration | 1
cardiorespiratory arrest | 1
cardiopulmonary resuscitation | 1
pulseless electrical activity | 1
return of spontaneous circulation | 2
ST-elevation in II, III, aVF, and V6 | 2
forceps extraction | 2
postpartum hemorrhage | 2
suspected diagnosis of AFE | 2
echo-cardiography | 2
transesophageal echocardiography | 3
globally hyperkinetic left ventricle | 3
hypokinesia to akinesia of the inferior wall | 3
normal right ventricle | 3
no signs of aortic dissection or valvular heart disease | 3
coagulation and fibrinolysis markers | 3
thromboelastometry | 3
coagulation essays | 3
completely abolished clotting | 3
fulfilled criteria for DIC | 3
platelets 97×10^9/L | 3
D-dimers 4154 ng/L | 3
prothrombin time not quantifiable | 3
fibrinogen level 0.35 g/L | 3
infusion of high doses of fibrinogen | 4
infusion of human coagulation factor XIII | 4
infusion of prothrombin concentrate complex | 4
antifibrinolytic therapy | 4
tranexamic acid | 4
transfusion of thrombocytes | 4
transfusion of packed red blood cells | 4
oxytocin administration | 4
Bakri balloon installation | 4
full-body computed tomography scan | 5
no occult bleeding complications | 5
no pulmonary embolism | 5
ST-segment elevations resolved | 6
cardiac bio-markers peaked | 11.5
low-dose aspirin administration | 12
angiotensin converting enzyme inhibitor administration | 12
prophylactic heparin therapy | 12
extubation | 12
normal oxygenation | 12
recovery from disorientation | 12
no residual neurological impairment | 12
vasoactive agents tapered off | 12
transthoracic echocardiography | 48
normal LV chamber dimension | 48
mildly reduced biplane ejection fraction | 48
akinesia of the inferior wall | 48
hypokinesia in the basal and midventricular inferolateral segments | 48
normal right ventricle | 48
no signs of pulmonary hypertension | 48
cardiac magnetic resonance imaging | 2160
preserved LVEF | 2160
inferior and inferolateral akinesia | 2160
late gadolinium enhancement | 2160
myocardial scarring | 2160
adenosine stress and rest perfusion imaging | 2160
no inducible ischemia | 2160
aspirin and lisinopril continued | 2160
cardiac rehabilitation | 4320
regular physical exercise | 4320
free from symptoms | 4320
echocardiography | 4320
improved systolic LV function | 4320
small mid inferolateral hypokinetic area | 4320
pregnancy | 6480
uneventful pregnancy and delivery | 6480