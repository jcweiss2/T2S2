53 years old | 0
male | 0
admitted to the hospital | 0
chief complaint of sudden loss of vision in his left eye | -120
feeling unwell | -120
shortness of breath | -120
generalized body pains | -120
fever | -120
chills | -120
denies headache | -120
denies extremity weakness or numbness | -120
denies chest pain | -120
denies cough | -120
denies abdominal pain | -120
denies nausea | -120
denies vomiting | -120
history of IV drug use | -6720
history of chronic obstructive lung disease | -6720
exploratory laparotomy | -8760
temperature 36.8ºC | 0
heart rate 92 bpm | 0
blood pressure 91/55 mmHg | 0
respiratory rate 18 breaths/min | 0
oxygen saturation 92% on 2 L of oxygen | 0
moderate respiratory distress | 0
diffuse bilateral rhonchi | 0
regular heart rate and rhythm | 0
ejection murmur in the tricuspid area | 0
soft and nontender abdomen | 0
left eye endophthalmitis | 0
intubated | 0
fluid resuscitation | 0
vasopressor therapy | 0
vitreous tap | 0
injection of vancomycin | 0
injection of ceftazidime | 0
empiric antibiotic therapy | 0
elevated white blood cell count | 0
hemoglobin 8.4 g/dL | 0
platelet count 210 000/mm3 | 0
creatinine 1.45 mg/dL | 0
urine drug screen positive for benzodiazepine | 0
urine drug screen positive for opiates | 0
blood cultures obtained | 0
HIV antigen/antibody testing nonreactive | 0
chest X-ray showed left upper lobe reticulonodular infiltrates | 0
chest X-ray showed prominent pulmonary arteries | 0
chest X-ray showed coarse left basilar and right upper lung zone markings | 0
CT scan showed multiple scattered cystic-like areas of opacity | 0
CT scan showed consolidation mainly in the upper lungs and periphery | 0
CT scan of the orbit showed minimal edema of the left preseptal soft tissues | 0
CT scan of the orbit showed subtle thickening of the sclera of the left globe | 0
CT scan of the orbit showed slight intraconal fat stranding | 0
transthoracic echocardiogram showed a large mobile echo density | 0
transthoracic echocardiogram showed a small echo density | 0
blood cultures revealed S. marcescens | 48
switched from cefepime to meropenem | 48
gentamicin added to the regimen | 48
vancomycin continued | 48
tricuspid valve replacement | 48
left upper lung/pleural abscess drainage | 48
tricuspid valve heavily encased in endocarditic vegetation | 48
severe regurgitation | 48
Epic porcine tissue valve placed | 48
tissue cultures from the tricuspid valve showed S. marcescens | 48
tissue cultures from the lung abscess showed S. marcescens | 48
dark red blood coming out of his nasogastric tube | 72
low hemoglobin level | 72
gastrointestinal bleeding suspected | 72
esophagogastroduodenoscopy showed esophagitis | 72
large amount of clotted blood in the fundus of the stomach | 72
four ischemic ulcers | 72
hemoclips placed | 72
culture of vitreous taken from the patient’s left eye grew S. marcescens | 96
ophthalmological examination showed stable eye | 96
no hypopyon | 96
switched to ciprofloxacin | 96
IV vancomycin discontinued | 96
follow-up blood cultures became negative | 192
Epsilometer test showed S. marcescens susceptible to ciprofloxacin | 192
gentamicin switched to IV ciprofloxacin | 192
follow-up ophthalmological examination showed persistent chemosis | 192
anterior chamber cloudy | 192
repeat CT scan of the orbit showed minimal asymmetric preseptal swelling | 192
repeat intravitreal injection of ceftazidime | 192
B-scan ultrasound showed increased vitreous debris | 336
pars plana vitrectomy | 360
subconjunctival pus noted | 360
conjunctival peritomy performed | 360
lens removed by phacofragmentation | 360
infection eroded through the sclera | 360
purulent intraocular drainage | 360
vitreous biopsy and anterior chamber paracentesis performed | 360
iris membrane removed | 360
vitreous injection of vancomycin and ceftazidime | 360
posterior perforation found | 360
left eye enucleation | 456
antibiotic therapy continued for 6 weeks | 840
discharged to a nursing home | 840
readmitted to the hospital with Staphylococcus aureus bacteremia | 2160