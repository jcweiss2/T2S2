44 years old | 0
    male | 0
    presented to the emergency department | 0
    persisting fever over 39°C | -216
    productive cough | -216
    chest pain | -216
    treatment with amoxicillin–clavulanate | -216
    treatment with paracetamol | -216
    no GI symptoms | 0
    clinical history was negative | 0
    no smoking history | 0
    no drugs use | 0
    isolated anal fissure | -175200
    sometimes slightly bleeding | -175200
    diagnosed 20 years ago | -175200
    COVID-19 diagnosed by RT-PCR | 0
    chest plain film showed right infrahilar opacity | 0
    chest plain film showed bilateral peripheral reticular pattern | 0
    CRP 16.64 mg/dL | 0
    PCT 0.29 ng/mL | 0
    ferritin 1966 ng/mL | 0
    D-dimer 1248 ng/mL | 0
    INR 1.53 | 0
    LDH 380 U/L | 0
    minimal neutrophilia | 0
    blood count normal | 0
    interleukin-6 levels <3.0 pg/mL | 0
    AST 38 UI/L | 0
    ALT 28 UI/L | 0
    bilirubin 1.20 mg/dL |-
    