58 years old | 0
male | 0
high grade fever | -336
chills | -336
bilateral loin pain | -336
left thigh pain | -336
diabetes mellitus | 0
recurrent urinary tract infection | 0
creatinine 917 mmoL/L | 0
hemoglobin 6.5 g/dL | 0
total leucocytic count 40.7 × 103 | 0
INR 1.8 | 0
creatinine kinase 447 | 0
random blood sugar 8.45 mmol/L | 0
E. coli in urine culture | 0
bilateral emphysematous pyelonephritis | 0
right kidney hydronephrosis | 0
right ileopsoas muscle infiltration | 0
left kidney small with stones | 0
septic shock | 0
ICU admission | 0
broad spectrum antibiotics | 0
bilateral nephrostomy tubes fixation | 0
retroperitoneal drains | 0
total leucocytic count 16.6 | 48
creatinine 663 mmol/L | 48
hemoglobin 8.2 g/dL | 48
follow-up CT showing improvement | 48
deterioration | 72
profuse rectal bleeding | 72
colonoscopy showing mucosal bleeding | 72
inotropes | 72
death | 168
