23 years old | 0
male | 0
admitted to the hospital | 0
right thigh swelling | -1560
draining sinus | -1560
skin changes | -1560
no history of fever | -1560
no systemic symptoms | -1560
past medical history unremarkable | 0
no regular medications | 0
life-long non-smoker | 0
denies alcohol or illicit substance use | 0
closed midshaft fracture of the right femur | -18240
motorbike accident | -18240
intramedullary fixation | -18240
surgical site infection | -8760
hardware removal | -8760
two-week course of antibiotics | -8760
asymptomatic for several years | -8760
migrated to Australia | -6240
experienced symptoms in right thigh | -1560
hemodynamically stable | 0
afebrile | 0
body mass index of 19 kg/m2 | 0
prolonged difficulty gaining weight | 0
able to weight bear with minimal pain | 0
right thigh swollen | 0
scaly skin discoloration | 0
draining sinus on the posterolateral aspect of the distal thigh | 0
neurovascular status of the limb intact | 0
preserved tone, power and range of motion | 0
minimally elevated white cell count | 0
C-reactive protein elevated | 0
erythrocyte sedimentation rate elevated | 0
electrolytes and liver function tests within normal range | 0
computed tomography scan | 0
united right femur fracture | 0
intramuscular collection within the vastus intermedius | 0
non-specific bony changes | 0
magnetic resonance imaging | 0
radiological findings suggestive of chronic osteomyelitis | 0
bone scintigraphy scan | 0
technetium-99m and gallium-67 study | 0
punch biopsy of the skin | 0
chronic spongiotic tissue reaction | 0
superimposed lichen simplex chronicus | 0
long-term dermatitis | 0
ultrasound-guided aspiration of the sinus | 0
culture yielded multi-resistant A. xylosoxidans | 0
initial sinus tract excision and drainage | 0
soft tissue and bone samples confirmed presence of A. xylosoxidans | 0
co-infection with S. aureus | 0
debridement of the medullary canal | 168
reamer-irrigator-aspirator technique | 168
systemic sepsis | 168
transferred to the Intensive Care Unit | 168
intravenous fluid resuscitation | 168
transfusion of 2 units of packed red blood cells | 168
vasopressor support with noradrenaline | 168
haemodynamic stability restored | 168
commenced on intravenous antibiotic therapy | 168
flucloxacillin | 168
meropenem | 168
blood cultures taken on post-operative day 1 | 192
positive for methicillin-sensitive S. aureus | 192
repeat sample 48 hours later returned a negative result | 240
discharged to the ward | 336
treated with intravenous antibiotics for one month | 720
transitioned to oral flucloxacillin | 720
co-trimoxazole | 720
asymptomatic after one month of oral antibiotics | 1680
weight bearing with no pain | 1680
full range of motion in right hip and knee | 1680
intact neurovascular status | 1680
surgical wound healed | 1680
no sign of infection | 1680
hyperpigmentation persisted around the wound site | 1680
successful ongoing weight gain | 1680
no adverse effects from antibiotic therapy | 1680
mild gastrointestinal discomfort | 1680
full recovery at six-month follow-up | 4320
CRP and leukocyte counts within normal limits | 4320
skin changes resolved | 4320
returned to full function | 4320
no reports of pain | 4320
full recovery at one-year follow-up | 8760
CRP and leukocyte counts within normal limits | 8760
no clinical evidence of infection | 8760
plain radiograph of the affected femur showed no residual disease | 8760
discharged from services | 8760