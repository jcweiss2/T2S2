60 years old | 0
male | 0
admitted to the emergency department | 0
acute anaemia | -48
fever | -48
diabetes mellitus | 0
laparoscopic radical cystectomy | -720
bilateral pelvic lymph node dissection | -720
urinary diversion | -720
discharged one month prior | -720
septic shock | 0
haemorrhagic shock | 0
enhanced abdominal CT | 0
diffuse extravasation of the contrast medium | 0
right external iliac artery disruption | 0
broad-spectrum antibiotics (imipenem) | 0
open exploratory operation | 0
extensive adhesion formation | 0
inflammation around the ileal bladder | 0
inflammation around the external iliac artery | 0
vessel split of the right external iliac artery | 0
vascular stent insertion | 0
transferred to the intensive care unit | 0
Klebsiella pneumoniae subsp. Pneumoniae (KPSP) isolated in blood culture | 72
drug susceptibility test | 72
sensitive to tigecycline | 72
sensitive to imipenem | 72
antibiotics (tigecycline plus imipenem) | 72
vital signs normalized | 504
blood tests normalized | 504
repeat enhanced CT | 720
no effusion of the contrast medium | 720
discharged | 792
follow-up every 3 months | 0
follow-up every 6 months | 0
no relapse | 0
