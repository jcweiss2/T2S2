66 years old | 0
male | 0
sick sinus syndrome | -3.6
paroxysmal atrial fibrillation | -3.6
severe lumbar back pain | 0
mental status changes | 0
hypotension | 0
acute renal failure | 0
hypoxemic respiratory failure | 0
intubated | 0
sepsis | 0
vasopressin | 0
norepinephrine | 0
methicillin-sensitive Staphylococcus aureus | 0
vancomycin | 0
nafcillin | 0
left ventricular ejection fraction 55% | 0
patent foramen ovale | 0
osteomyelitis of the lower spine | 0
multiple small, 2- to 3-mm, acute infarctions | 0
septic emboli to the distal extremities | 0
repeat blood cultures | 0
transesophageal echocardiogram | 0
vegetation in the right atrium | 0
vegetation attached to the pacemaker lead | 0
intracardiac echocardiography | 0
RV lead vegetations | 0
aspiration catheter | 0
vacuum pump | 0
aspiration | 0
smaller vegetation | -0.33
larger vegetation | -0.33
laser lead extraction | 0.33
RA and RV leads extraction | 0.33
pocket inspection | 0.33
suture closure | 0.33
hemostasis | 0.33
72 minutes | 0.33
200 mL blood loss | 0.33
tissue necrosis of the distal upper and lower extremities | 72
lactic acidosis | 72
worsening renal failure | 72
withdrawal of care | 72
death | 72