46-year-old man | 0
Ulcerative colitis | 0
Malaise, fever, loss of appetite | -72
Arrival at emergency department | 0
Blood pressure, heart rate, SpO2, respiratory rate, body temperature | 0
Cardiac arrest | 0
Ventricular fibrillation (VF) | 0
Defibrillation and adrenaline administration | 0
Diagnosis of Brugada syndrome (BS) | 0
Coved-type ST elevation in ECG | 0
Improvement with acetaminophen | 0
Hypercalcemia (HC) level of 14.8 mg/dL | 0
Hypotension and suspected septic shock | 0
Initiation of tazobactam-piperacillin and vasopressors | 0
Extubation on day 2 | 48
Reoccurrence of fever and liver abscess diagnosis | 120
Change of antibiotics to meropenem and vancomycin | 120
Puncture drainage | 120
Positive pilsicainide test result | 720
Implantation of ICD | 720
Discharge | 720
Family history of sudden death | 0
High parathyroid hormone levels and Tc scintigraphy | 0
Tumor resection after discharge | 0
Pathological diagnosis of ectopic parathyroid adenoma | 0
CT and MRI revealing nonfunctional pituitary and adrenal tumors | 0
Diagnosis of multiple endocrine neoplasia type 1 (MEN1) | 0