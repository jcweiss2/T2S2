64 years old | 0
white | 0
male | 0
admitted to the hospital | 0
ground-level fall | -1
dizziness | -1
lightheadedness | -1
hypoglycemia | -1
hemodynamically stable | 0
alert | 0
oriented | 0
bilateral lower extremity pitting edema | 0
superficial forehead abrasion | 0
stage 2 sacral decubitus ulcer | 0
ruptured skin blister | 0
leukocytosis | 0
white blood cell count of 14.7 × 103 cells/μl | 0
neutrophil count of 12.2 × 103 cells/μl | 0
serum creatinine concentration of 1.33 mg/dl | 0
evolving sepsis | 0
septic shock | 24
exacerbation of congestive heart failure | 24
admission to the intensive care unit | 24
bacteremia with methicillin-sensitive Staphylococcus aureus (MSSA) infection | 0
skin infection | 0
acute tubular necrosis | 48
dialysis | 48
infective endocarditis | 0
echocardiography | 0
heart failure with preserved ejection fraction | -720
symptomatic bradycardia | -720
pacemaker placement | -720
hypertension | -720
hyperlipidemia | -720
controlled type 2 diabetes mellitus | -720
dental procedure | -144
computed tomography of the chest | 0
large bilateral pleural effusions | 0
pulmonary vascular congestion | 0
thoracentesis | 24
transudative effusions | 24
blood cultures | 0
MSSA bacteremia | 0
urine cultures | 24
sputum cultures | 24
bronchial washings | 24
transthoracic echocardiogram | 48
moderate pulmonic valve regurgitation | 48
transesophageal echocardiogram (TEE) | 264
mobile mass on the ventricular surface of the pulmonic valve | 264
moderate regurgitation | 264
papillary fibroelastoma | 264
bacterial vegetation | 264
AngioVac procedure | 384
mass debulking | 384
ultrasonography-guided approach | 384
therapeutic anticoagulation | 384
heparin | 384
serial dilation | 384
cardiopulmonary bypass | 384
pigtail catheter | 384
Amplatz Super Stiff guidewire | 384
fluoroscopic guidance | 384
TEE guidance | 384
right heart bypass | 384
mass extraction | 384
pathology | 384
cardiac papillary fibroelastoma (PFE) | 384
Streptococcus salivarius | 384
Rothia spp | 384
linezolid | 384
meropenem | 384
follow-up blood cultures | 408
no bacterial growth | 408
discharged to hospice | 504