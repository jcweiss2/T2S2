48 years old | 0
male | 0
admitted to the hospital | 0
fever | -96
cough | -96
shortness of breath | -96
sputum | -96
amoxicillin | -96
deteriorated | -72
dyspnea | -72
non-invasive mechanical ventilation | -72
Ceftriaxone | -72
bacterial pneumonia | -72
computed tomography | -72
bilateral diffuse consolidation | -72
diabetes mellitus | 0
chronic gout | 0
long-term use of corticosteroids | 0
body temperature | 0
blood pressure | 0
arterial blood gas analysis | 0
PaO2/FiO2 | 0
lung compliance | 0
intubated | 6
mechanical ventilation | 6
prone position | 6
volume-controlled ventilation | 6
transferred to ICU | 24
Mycobacterium tuberculosis | 24
acid-fast bacilli | 24
Human immunodeficiency virus | 24
TB-induced ARDS | 24
VV-ECMO | 24
internal jugular vein cannulation | 24
femoral access vein cannulation | 24
Seldinger technique | 24
blood flow | 24
gas flow | 24
mechanical ventilator setting | 24
tidal volume | 24
end inspiratory plateau pressure | 24
respiratory rate | 24
positive end-expiratory pressure | 24
FiO2 | 24
anti-TB regimens | 24
ethambutol | 24
pyrazinamide | 24
rifampicin/isoniazid | 24
Levofloxacin | 24
meropenem | 24
amikacin | 24
corticosteroids | 24
heparin | 24
anticoagulation regimen | 24
Activated Partial Thromboplastin Time | 24
hypoxemia | 48
lung compliance | 48
improved | 48
chest radiography | 96
improved | 96
weaned from ECMO | 120
extubated | 192
respiratory muscle weakness | 240
corticosteroid-induced myopathy | 240
cerebrospinal fluid examination | 240
normal | 240
tracheostomy | 360
weaned from mechanical ventilation | 840
discharged | 1128