63 years old | 0  
    male | 0  
    admitted to the emergency room | 0  
    weakness | 0  
    nausea | 0  
    vomiting | 0  
    diarrhea | 0  
    ingesting several wild mushrooms | -36  
    severe nausea | -29  
    vomiting | -29  
    diarrhea | -29  
    hypertension | -1464  
    colon carcinoma | -1464  
    surgery | -1464  
    chemotherapy | -1464  
    no metastasis in the liver | -1464  
    did not consume alcohol | -1464  
    did not use any medication | -1464  
    awake | 0  
    fully oriented | 0  
    normal vital signs | 0  
    dehydration | 0  
    normal arterial blood gas analysis | 0  
    nonreactive hepatitis B surface antigen | 0  
    nonreactive hepatitis B core antibody | 0  
    nonreactive immunoglobulin M | 0  
    nonreactive antihepatitis C antibody | 0  
    negative hepatitis B virus DNA analysis | 0  
    admitted to the internal medicine intensive care unit | 0  
    gastric lavage | 0  
    activated charcoal | 0  
    rehydration with 0.9% sodium chloride | 0  
    rehydration with 5% dextrose | 0  
    silibinin bolus dose | 0  
    silibinin continuous infusion | 0  
    acetylcysteine infusion | 0  
    penicillin G infusion | 0  
    multivitamin | 0  
    alpha lipoic acid | 0  
    complete blood count | 0  
    biochemistry measurements | 0  
    blood gas monitoring | 0  
    aspartate aminotransferase 880 U/L | 6  
    alanine aminotransferase 665 U/L | 6  
    lactate dehydrogenase 1,028 U/L | 6  
    total bilirubin 4.9 mg/dL | 6  
    direct bilirubin 1.9 mg/dL | 6  
    prothrombine time 36.5 seconds | 6  
    international normalized ratio 3.11 | 6  
    normal lactate level | 6  
    vitamin K | 6  
    metilprednisolone | 6  
    aspartate aminotransferase 1,836 U/L | 12  
    alanine aminotransferase 1,232 U/L | 12  
    lactate dehydrogenase 1,471 U/L | 12  
    total bilirubin 7.2 mg/dL | 12  
    direct bilirubin 3.1 mg/dL | 12  
    prothrombine time 73.1 seconds | 12  
    international normalized ratio 6.86 | 12  
    metabolic acidosis | 12  
    respiratory alkalosis | 12  
    fresh frozen plasma | 12  
    hemodialysis | 12  
    worsening general condition | 30  
    somnolent | 30  
    mildly tachypneic | 30  
    aspartate aminotransferase 1,900 U/L | 30  
    alanine aminotransferase 1,473 U/L | 30  
    lactate dehydrogenase 2,582 U/L | 30  
    prothrombine time 76.5 seconds | 30  
    international normalized ratio 7.22 | 30  
    hemoglobin 12.5 g/dL | 30  
    platelets 123,000/mm3 | 30  
    consultation for liver transplantation | 30  
    continued therapies | 30  
    hemodialysis | 30  
    fresh frozen plasma | 30  
    aspartate aminotransferase 1,843 U/L | 30  
    alanine aminotransferase 984 U/L | 30  
    lactate dehydrogenase 3,826 U/L | 30  
    prothrombine time 42.6 seconds | 30  
    international normalized ratio 3.71 | 30  
    aspartate aminotransferase 1,207 U/L | 48  
    alanine aminotransferase 1,797 U/L | 48  
    lactate dehydrogenase 4,318 U/L | 48  
    total bilirubin 9.8 mg/dL | 48  
    direct bilirubin 3.3 mg/dL | 48  
    prothrombine time 47.7 seconds | 48  
    international normalized ratio 4.21 | 48  
    hemoglobin 11.8 g/dL | 48  
    platelets 33,000/mm3 | 48  
    high anion gap metabolic acidosis | 48  
    respiratory alkalosis | 48  
    normal fibrinogen level | 48  
    elevated D-dimer concentration | 48  
    no schistocytes | 48  
    flapping tremor | 48  
    blood ammonia level 281 μg/dL | 48  
    hepatic encephalopathy treatment | 48  
    branched chain amino acid solution | 48  
    ornithine-aspartate infusion | 48  
    lactulose | 48  
    aspartate aminotransferase 3,570 U/L | 54  
    alanine aminotransferase 3,282 U/L | 54  
    lactate dehydrogenase 4,379 U/L | 54  
    total bilirubin 12.4 mg/dL | 54  
    prothrombine time 111 seconds | 54  
    international normalized ratio 11.05 | 54  
    platelets 29,000/mm3 | 54  
    hemodialysis | 54  
    fresh frozen plasma | 54  
    prothrombine time 34.6 seconds | 60  
    international normalized ratio 2.92 | 60  
    hemoglobin 8.6 g/dL | 60  
    platelets 12,000/mm3 | 60  
    erythrocyte suspension | 60  
    lost consciousness | 72  
    body temperature 38.2°C | 72  
    pulse rate 112 beats per minute | 72  
    respiratory rate 32 breaths per minute | 72  
    blood pressure 89/57 mmHg | 72  
    meropenem | 72  
    aspartate aminotransferase 1,096 U/L | 78  
    alanine aminotransferase 2,004 U/L | 78  
    lactate dehydrogenase 1,615 U/L | 78  
    prothrombine time 100.6 seconds | 78  
    international normalized ratio 9.87 | 78  
    platelets 7,000/mm3 | 78  
    hemodialysis | 78  
    fresh frozen plasma | 78  
    platelet infusion | 78  
    pure respiratory alkalosis | 78  
    serum lactate 16.59 mg/dL | 84  
    ammonia 415 μg/dL | 84  
    serum creatinine 2.6 mg/dL | 84  
    hepatorenal syndrome | 84  
    arterial blood gas acidosis | 84  
    sedation | 84  
    intubation | 84  
    cardiac arrest | 90  
    resuscitation | 90  
    arterial blood gas acidosis | 90  
    sodium bicarbonate | 90  
    aspartate aminotransferase 329 U/L | 96  
    alanine aminotransferase 855 U/L | 96  
    prothrombine time 77.3 seconds | 96  
    international normalized ratio 7.31 | 96  
    platelets 13,000/mm3 | 96  
    hemoglobin 8.3 g/dL | 96  
    serum creatinine 3.3 mg/dL | 96  
    serum lactate 112 mg/dL | 96  
    arterial blood gas acidosis | 96  
    cardiac arrest | 98  
    death | 98  
    