28 years old | 0
female | 0
admitted to the hospital | 0
right hypochondriac pain | -840
jaundice | -336
passing tea-coloured urine | -336
no known medical illness | 0
no history of surgery | 0
stable | 0
blood pressure of 145/94 mm Hg | 0
pulse rate of 80 bpm | 0
afebrile | 0
mild hyperbilirubinaemia | 0
alanine aminotranferanse (ALT) within the normal range | 0
aspartate aminotranferanse (AST) within the normal range | 0
alkaline phosphatase (ALP) within the normal range | 0
total white cell count was 8.6×10^9/L | 0
full blood count normal | 0
renal profile normal | 0
coagulation profile normal | 0
serum amylase normal | 0
gallstone | 0
no dilated biliary ducts | 0
total bilirubin 57.6 μmol/L | -48
direct 40.2 μmol/L | -48
indirect 17.4 μmol/L | -48
ALP 237 units/L | -48
ALT 251 units/L | -48
AST 266 units/L | -48
total bilirubin 126.4 μmol/L | 0
direct 82.4 μmol/L | 0
indirect 44 μmol/L | 0
ALP 357 units/L | 0
ALT 523 units/L | 0
AST 288 units/L | 0
no recorded fever | 0
dilated intrahepatic and extrahepatic biliary dilatation | 0
lesion in the distal bile duct | 0
impacted soft stone in the common bile duct | 0
CT scan | 0
informed consent | 0
screened for COVID-19 symptoms | -24
denied having travelled abroad | -24
denied having recent mass activity | -24
denied contact with COVID-19 positive person | -24
denied fever | -24
denied sore throat | -24
denied cough | -24
denied difficulty in breathing | -24
denied diarrhoea | -24
signed health declaration document | -24
healthcare staffs screened | -24
donning of PPE | -10
endoscopy system ready | -10
image intensifier ready | -10
patient sent to OT airlock bay | -5
patient wore long sleeve waterproof gown | -5
patient wore cap | -5
patient wore glove | -5
checklist for patient undergoing conscious sedation | -5
intravenous antibiotic | -5
ERCP procedure | 0
aerosol protective barrier | 0
oxygen therapy | 0
vital signs checked | 0
intravenous sedative medication | 0
protective barrier placed | 0
ampulla floppy | 0
bile not present | 0
pus seen on partial sphincterotomy | 0
limited contrast injection | 0
guide wire in bile duct | 0
10-French 9 cm plastic stent deployed | 0
bile flow good | 0
reversal medication | 0
patient fully awake | 0
doffing of PPE | 15
endoscopy equipment disinfected | 30
patient sent to recovery bay | 30
total bilirubin 50 μmol/L | 48
direct 23 μmol/L | 48
indirect 27 μmol/L | 48
total leucocyte count 9.98×10^9/L | 48
ALP 354 units/L | 48
ALT 359 units/L | 48
AST 100 units/L | 48
discharged | 120
oral antibiotics | 120
follow-up | 336
total bilirubin 21.8 μmol/L | 336
direct 15 μmol/L | 336
indirect 6.8 μmol/L | 336
ALP 134 units/L | 336
ALT 21 units/L | 336
AST 20 units/L | 336
scheduled for ERCP and stone clearance | 336