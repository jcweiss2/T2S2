77 years old | 0
male | 0
admitted to the hospital | 0
history of tuberculosis | -87600
chronic obstructive pulmonary disease (COPD) | -87600
hyperthyroidism | -87600
diabetes mellitus (DM) | -87600
confusion | 0
shortness of breath | 0
tachycardia | 0
hypothermia | 0
hypotension | 0
acute respiratory failure | 0
systemic inflammatory response syndrome (SIRS) | 0
intubated | 0
connected to ventilator | 0
decrease in respiratory sounds | 0
right lung marked decrease | 0
coarse rales | 0
prolongation of expirium | 0
bilateral biphasic expiratory ronchi | 0
obstructive pattern on pulmonary function test | 0
Glascow Coma Score 6 | 0
APACHE II 34 | 0
multiple organ dysfunction syndrome (MODS) 8 | 0
pulse 122/min | 0
arterial blood pressure 82/41 mmHg | 0
respiratory rate 30/min | 0
temperature 35°C | 0
leukocyte 27600/mm3 | 0
C-reactive protein (CRP) 52 mg/L | 0
thyrotoxicosis | 0
FT4 8.5 ng/dL | 0
TSH < 0.05 μIU/mL | 0
TRAb 0.9 IU/mL | 0
thyroid ultrasonography hyperechoic nodule 8.5 mm | 0
hyperthyroidism associated with Graves' thyrotoxicosis | 0
propranolol treatment | 0
methimazole treatment | 0
pneumonic infiltration on chest X-ray | 0
ground glass density increase on chest X-ray | 0
no cardiac ischemia on ECG | 0
diastolic dysfunction in echocardiography | 0
temperature 38.4°C at day 2 | 48
no growth on cultures | 48
ampicillin-sulbactam | 48
levofloxacin | 48
acid resistance bacteria (ARB) negative three times | 48
no response to treatment | 48
substituted therapy with piperacillin/tazobactam | 168
trimetoprim/sulfametaxazol | 168
clarithromycin | 168
no temperature decrease | 168
more severe clinical course | 168
no regression of pneumonic infiltration | 168
bronchoscopy performed | 168
fungus ball on thoracic CT | 168
narrow trachea and bronchi lumens | 168
diffuse white-colored plaques | 168
thin-walled necrotic lesion | 168
tuberculosis cavity middle lobe right lung | 168
infiltration around lesion | 168
crescent sign on CT | 168
histopathological examination biopsy specimens | 168
active inflammation | 168
fibrous scarring | 168
microscopic abscess cavity | 168
central bronchiectasis | 168
dense peribronchial inflammation | 168
fibrosis | 168
fungus ball | 168
septate hyphae Aspergillus fumigatus | 168
Aspergillus fumigatus on BAL culture | 168
voriconazole loading dose 400 mg i.v. | 168
voriconazole maintenance dose 200 mg i.v. | 168
disease more severe on day 18 | 432
multiple organ failure (MOF) | 432
death | 432
