32 years old | 0
female | 0
cystic fibrosis | -8760
bronchiectasis | -8760
recurrent hemoptysis | -8760
pancreatic insufficiency | -8760
malnutrition | -8760
admitted to the hospital | 0
massive hemoptysis | 0
broad-spectrum antibiotics | 0
computed tomography angiogram | 0
centrilobular ground-glass opacities | 0
pulmonary hemorrhage | 0
referred to interventional radiology | 0
right common femoral artery access | 0
bronchial artery embolization | 0
left bronchial arteriogram | 0
microcatheter | 0
embolization | 0
post-embolization arteriogram | 0
stasis | 0
preserved patency | 0
discharged | 24
recurrent massive hemoptysis | 3
inhaled tranexamic acid | 3
admitted to the medical intensive care unit | 3
elective intubation | 3
diagnostic bronchoscopy | 3
pulmonary and systemic arterial angiography | 3
embolization | 3
thyrocervical trunk-pulmonary artery fistula | 3
systemic to pulmonary arterial fistulae | 3
embolization of the supreme intercostal artery | 3
embolization of the thyrocervical trunk | 3
post-embolization angiogram | 3
septic shock | 24
Burkholderia cepacian complex | 24
sputum cultures | 24
weaned off vasopressors | 48
transferred out of the MICU | 48
hemoptysis-free | 264
isolated hemoptysis recurrence | 264
repeat CTA | 264
active extravasation | 264
continued enhancement of the pseudoaneurysm | 264
goals of care discussion | 264
repeat embolization | 336
intubation | 336
repeat CTA | 336
pseudoaneurysm | 336
embolization | 336
coil embolization | 336
post-embolization angiogram | 336
stasis | 336
transition to comfort measures | 408
expired | 408
acute respiratory failure | 408
Burkholderia cepacian infection | 408
complication of cystic fibrosis | 408