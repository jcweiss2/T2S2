slipping on wet grass and falling on his left side | -1
presented to the Emergency department | 0
glasgow coma score was 15/15 | 0
vital signs were within normal limits | 0
left hip tenderness | 0
no ecchymosis to the abdomen, flank or thigh | 0
radiograph of his pelvis revealed an undisplaced fracture of his left acetabulum | 0
initial blood tests confirmed his liver dysfunction | 0
pH 7.271 | 0
base excess minus 7.3 | 0
PT 18.2 | 0
INR-1.5 | 0
APTT ratio 1.42 | 0
platelets 73 | 0
bilirubin 63 mmol/l | 0
Hb was unremarkable at 124 g/l | 0
18 g intravenous cannula was inserted | 0
warmed Hartmanns one litre infusion was commenced | 0
referred to the Orthopaedic on call team | 1
blood pressure dropped to 75/51 mm Hg | 2
tachycardic | 2
serum lactate was 9 mmol/l | 2
FAST examination revealed intraabdominal fluid | 2
treated for sepsis in the Emergency department | 2
intensive care, orthopaedic and general registrar attended the patient | 3
pH was 7.227 | 3
base excess of −17.9 | 3
serum lactate of 16.3 mmol/l | 3
Hb was now 75 g/l | 3
arterial blood pressure was 90/60 mm Hg | 3
pulse rate 90/min | 3
left lower abdominal quadrant and upper thigh were now swollen with ecchymosis | 3
diagnosis of haemorrhagic shock was made | 3
massive transfusion pathway was activated | 3
Four units of Blood, 4 units of FFP, 2 adult therapeutic doses of platelets and 10 units of cryoprecipitate were rapidly transfused | 4
noradrenaline infusion to maintain MAP > 65 mm Hg | 4
pelvic binder was in place | 4
CT scan was deemed necessary | 5
CT abdomen confirmed the fracture of the left acetabulum | 6
significant haematoma on left pelvic sidewall adjacent to the fracture | 6
8 mm enhancing nodule suggestive of an internal iliac artery pseudoaneurysm | 6
ill-defined blush of contrast within the haematoma | 6
extra-peritoneal haematoma inseparable from the bladder | 6
cirrhotic liver | 6
incidental 6.7 cm infra-renal aortic aneurysm | 6
transferred to the intensive care unit | 7
CT Angiogram which demonstrated no arterial bleed | 24
prophylactic embolization was recommended | 24
gelfoam embolization of anterior and posterior division segmental branches of the left internal iliac artery | 48
10 lb skeletal traction was applied | 48
developed uncontrollable bleeding from his pin site | 120
skeletal traction was removed | 120
continuous pressure applied to the wound | 120
died on 30 January 2017 | 1224