58 years old | 0
man | 0
schizophrenia | 0
substance abuse | 0
diabetes mellitus | 0
hypertension | 0
headache | -96
chest pain | -96
afebrile | -96
hypertensive | -96
tachycardic | -96
confused | -96
intubated | -96
hyperglycemia | -96
acute kidney injury | -96
admission to emergency department | 0
blood cultures on admission | 0
blood cultures showed no growth | 0
extubated | 24
altered mental status | 24
synthetic cannabinoid intoxication | 24
agitated | 96
tachycardic | 96
hypertensive | 96
abdominal distension | 96
hypotensive | 144
intravenous fluid resuscitation | 144
febrile | 192
respiratory distress | 192
re-intubated | 192
arterial lactate peak | 192
treated with piperacillin-tazobactam | 192
blood cultures from central line | 192
blood cultures from periphery | 192
Lactobacillus species in aerobic bottles | 192
Lactobacillus species in anaerobic bottles | 192
persistent febrile | 192
persistent bandemia | 192
worsening diarrhea | 192
treated with metronidazole | 192
noncontrast CT chest | 192
noncontrast CT abdomen | 192
noncontrast CT pelvis | 192
wall thickening of ascending colon | 192
surrounding inflammatory changes | 192
ileus | 192
C. difficile toxin in stool | 192
C. difficile toxin negative | 192
colonoscopy | 192
diffuse edema from hepatic flexure to cecum | 192
intermittent areas of sparing | 192
severe ulceration | 192
necrotic mucosa | 192
no bleeding on biopsy | 192
ischemic colitis | 192
transesophageal echocardiogram | 192
no vegetation | 192
improved clinically | 240
extubated | 240
discharged | 240
piperacillin-tazobactam course | 240
metronidazole course | 240
- Headache | -24
