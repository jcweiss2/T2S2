48 years old | 0
male | 0
referred to our hospital | 0
right testicular seminoma | 0
pT4 | 0
multiple liver metastases | 0
bulky RPLN metastasis invaded the third portion of the duodenum | 0
human chorionic gonadotropin level of 24 IU/L | 0
LDH at 1060 IU/L | 0
normal alfa-fetoprotein | 0
four cycles of bleomycin | -672
etoposide | -672
cisplatin | -672
cisplatin dose reduced to 90% | -672
start of the fourth cycle of BEP delayed by 1 week | -672
completion of the BEP regimen | -336
hCG normalized | -336
LDH normalized | -336
contrast-enhanced CT | -336
PET-CT at 1 month after the completion of the BEP | -336
disappearance of liver metastases | -336
4-cm RPLN mass remained | -336
positive 18F-FDG uptake | -336
referred to our hospital for further management | -168
tumor markers in the normal range | -168
repeat PET-CT performed | -168
increasing 18F-FDG uptake in RPLN metastases | -168
new uptake in the right iliac lymph node metastases | -168
decided to perform salvage chemotherapy with paclitaxel | 0
ifosfamide | 0
cisplatin | 0
no severe adverse effects during TIP treatment | 168
CT after two courses of TIP demonstrated RPLN metastasis did not respond to chemotherapy | 168
two additional courses of TIP | 336
developed sudden-onset hematochezia | 480
hypovolemic shock | 480
hemoglobin 4.7 g/dL | 480
neutrophil count 4.8 × 109/L | 480
platelet count 4.9 × 109/L | 480
CT depicted dilated bowel loop with massive clot | 480
direct extravasation of contrast from the aorta into the third portion of the duodenum | 480
RPLN mass remained without decrease in size | 480
endoscopic therapy considered impossible | 480
hemodynamically unstable | 480
decision to attempt angioembolization | 480
emergent angiography confirmed presence of PADF | 480
deployed endovascular stent graft in the aorta | 480
control angiography showed minimal residual hemorrhage | 480
extensive fluid infusion | 480
blood transfusion | 480
developed sepsis | 648
disseminated intravascular coagulation | 648
multiple organ failure | 648
massive bleeding recurred | 792
died | 792
septic shock due to graft infection | 792
uncontrolled bleeding | 792
