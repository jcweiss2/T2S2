45 years old | 0
female | 0
accidental flame burns | -120
burns of the chest | -120
burns of the upper limbs | -120
high fever | -120
breathlessness | -120
admitted to the hospital | 0
right internal jugular vein catheter inserted | -120
administration of drugs | -120
administration of volume | -120
high fever | -96
breathing difficulty | -89
sepsis | -89
growth of methicillin-resistant Staphylococcus aureus (MRSA) | -89
antibiotics administered | -89
no clinical improvement | -72
persistent high temperatures | -72
breathlessness | -72
referred to hospital | -72
put on respirator | -72
poor blood gas values | -72
transthoracic echocardiogram | -72
large vegetation on the anterior tricuspid leaflet | -72
no tricuspid regurgitation | -72
trans-oesophageal echocardiogram | -72
ventilated for respiratory decompensation | -24
showering of the pulmonary circuit | -24
tiny vegetations on the ATL | -24
taken for surgery | 0
cardiopulmonary bypass | 0
tricuspid valve approached | 0
cardioplegic arrest | 0
large vegetation on the anterior tricuspid leaflet | 0
vegetation on the chordal apparatus | 0
total vegetectomy | 0
curettage of the anterior tricuspid leaflet | 0
repair of the ATL | 0
native pericardium used | 0
weaned off cardiopulmonary bypass | 0
afebrile | 24
discharged from the hospital | 168
vegetation grew MRSA | 168