68 years old | 0
male | 0
type 1 diabetic | 0
hypertensive | 0
amlodipine | 0
operated for treatment of right inguinal hernia | -175200
admitted to the emergency room | 0
abdominal pain | 0
ketoacidosis decompensation | 0
uremic syndrome | 0
conscious | 0
hemodynamically stable | 0
dyspneic | 0
febrile at 39.6°C | 0
right lumbar tenderness | 0
oliguric | 0
diuresis at 300 ml/24h | 0
altered renal function | 0
creatinine at 92 mg/l | 0
urea at 3.1 g/l | 0
K+ at 6.9 mmol/l | 0
Na+ at 123 mmol/l | 0
blood sugar at 6.5 g/l |,0
alkaline reserves at 8 mEq/l | 0
infectious syndrome | 0
CRP at 418 mg/l | 0
white blood cells at 26000/ml | 0
hemoglobin at 12.3 g/dl | 0
ECBU | 0
leucocyturia 320,000 | 0
hematuria at 120,000 | 0
abdominopelvic CT | 0
single anatomical right kidney | 0
emphysematous pyelonephritis | 0
renal abscess ruptured in the intraperitoneal cavity | 0
moderate abundance of pneumoperitoneum | 0
admitted to intensive care | 0
3 dialysis sessions | 0
insulin therapy | 0
antibiotic therapy | 0
ceftriaxone | 0
metronidazole | 0
ECBU culture | 0
urinary tract infection due to Pseudomonas Aeruginosa | 0
surgical drainage of abscesses | 0
right double J stent | 0
decrease of the infectious syndrome | 48
apyrexia | 48
chronic renal failure | 48
resumption of normal diuresis | 48
creatinine plateau of 20 mg/l | 48
discharged | 240
oral antibiotics | 240
abdominopelvic CT showed clear regression of air bubbles | 672
double J catheter removed | 1008
