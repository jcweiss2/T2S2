61 years old | 0
    male | 0
    visited another hospital | 0
    acute abdominal pain | 0
    fever | 0
    perforated duodenal ulcer | 0
    sepsis | 0
    primary surgical closure | 0
    right internal jugular vein catheterization | 0
    intensive care unit treatment | -120
    stabilized | -120
    transferred to general ward | -144
    CVC removed | -144
    physician assistant | -144
    sitting position | -144
    abruptly complained of shortness of breath | -144
    chest discomfort | -144
    became unconscious | -144
    immediate cardiopulmonary resuscitation | -144
    return of spontaneous circulation | -144
    transthoracic echocardiogram | -144
    multiple air bubbles in right ventricle | -144
    multiple air bubbles in left ventricle | -144
    ostium secundum atrial septal defect | -144
    right-to-left shunt | -144
    air embolism suspected | -144
    brain CT | -144
    chest CT | -144
    gas within centrum semiovale | -144
    gas within cerebral sulci | -144
    gas within cavernous sinuses | -144
    free air in neck | -144
    free air in jugular vein | -144
    free air in left ventricle | -144
    transferred to our hospital | 0
    vital signs on arrival | 0
    blood pressure 107/75 mmHg | 0
    heart rate 134 beats/min | 0
    respiratory rate 30 breaths/min | 0
    temperature 35.8°C | 0
    Glasgow coma scale 3/15 | 0
    chest X-ray | 0
    extensive bilateral infiltrates | 0
    pulmonary edema | 0
    arterial blood gas analysis | 0
    pH 7.141 | 0
    PaCO2 52.3 mmHg | 0
    PaO2 53.6 mmHg | 0
    HCO–3 14.8 mEq/L | 0
    SaO2 74% | 0
    venovenous ECMO support | 0
    stabilized | 168
    pulmonary edema ameliorated | 168
    lung injury ameliorated | 168
    weaned off ECMO | 168
    follow-up echocardiography | 72
    ejection fraction preserved | 72
    no regional wall motion abnormalities | 72
    apical left ventricle thrombus | 72
    anticoagulation therapy | 72
    acute renal failure | 72
    renal failure improved | 72
    no hemodialysis | 72
    Glasgow coma scale score 9 | 168
    diffuse cerebral ischemia | 168
    brain MRI | 168
    tracheostomy | 168
    transferred to general ward | 168
    
    61 years old|0
    male|0
    visited another hospital|0
    acute abdominal pain|0
    fever|0
    perforated duodenal ulcer|0
    sepsis|0
    primary surgical closure|0
    right internal jugular vein catheterization|0
    intensive care unit treatment|-120
    stabilized|-120
    transferred to general ward|-144
    CVC removed|-144
    physician assistant|-144
    sitting position|-144
    abruptly complained of shortness of breath|-144
    chest discomfort|-144
    became unconscious|-144
    immediate cardiopulmonary resuscitation|-144
    return of spontaneous circulation|-144
    transthoracic echocardiogram|-144
    multiple air bubbles in right ventricle|-144
    multiple air bubbles in left ventricle|-144
    ostium secundum atrial septal defect|-144
    right-to-left shunt|-144
    air embolism suspected|-144
    brain CT|-144
    chest CT|-144
    gas within centrum semiovale|-144
    gas within cerebral sulci|-144
    gas within cavernous sinuses|-144
    free air in neck|-144
    free air in jugular vein|-144
    free air in left ventricle|-144
    transferred to our hospital|0
    vital signs on arrival|0
    blood pressure 107/75 mmHg|0
    heart rate 134 beats/min|0
    respiratory rate 30 breaths/min|0
    temperature 35.8°C|0
    Glasgow coma scale 3/15|0
    chest X-ray|0
    extensive bilateral infiltrates|0
    pulmonary edema|0
    arterial blood gas analysis|0
    pH 7.141|0
    PaCO2 52.3 mmHg|0
    PaO2 53.6 mmHg|0
    HCO–3 14.8 mEq/L|0
    SaO2 74%|0
    venovenous ECMO support|0
    stabilized|168
    pulmonary edema ameliorated|168
    lung injury ameliorated|168
    weaned off ECMO|168
    follow-up echocardiography|72
    ejection fraction preserved|72
    no regional wall motion abnormalities|72
    apical left ventricle thrombus|72
    anticoagulation therapy|72
    acute renal failure|72
    renal failure improved|72
    no hemodialysis|72
    Glasgow coma scale score 9|168
    diffuse cerebral ischemia|168
    brain MRI|168
    tracheostomy|168
    transferred to general ward|168