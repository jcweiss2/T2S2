64 years old|0
    male|0
    hospitalized due to remittent high fever| -336
    no gastrointestinal symptoms| -336
    mild back pain over mid back area| -336
    able to walk independently| -336
    blood culture showed Salmonella enterica infection| -336
    meropenem 1g daily for 7 days| -336
    past history of coronary artery bypass grafting surgery due to atherosclerosis| -26208
    steroid-induced diabetes mellitus for 10 years| -87648
    chronic kidney disease| -87648
    readmitted to emergency ward|0
    hypotension|0
    persistently high fever (39.4°C)|0
    severe back pain| -168
    paraplegia| -168
    pain centered in upper back radiating to chest wall| -168
    Visual Analogue Scale (VAS) 7| -168
    weakness of both lower extremities| -168
    sensory loss below chest| -168
    no history of recent trauma| -168
    lost 1 kg weight in past month| -720
    blood sample for hematology|0
    coagulation profile|0
    blood culture|0
    urinary sample to rule out infection source|0
    no leukocytosis|0
    increased neutrophils|0
    decreased lymphocytes|0
    C-Reactive Protein high (111.08 mg/L)|0
    procalcitonin 0.27 ng/mL|0
    blood culture negative|0
    Mantoux test negative|0
    IGRA for tuberculosis negative|0
    HIV testing negative|0
    CD4 cell count 504 cells/mm3|0
    referred to intensive care unit due to septic shock|0
    high dose meropenem injection 1g every 8 hours|0
    renal function normal (upper limit)|0
    maximum urea level 37 mg/dL|0
    maximum creatinine level 1.23 mg/dL|0
    critical condition subsided five days after admission|120
    re-assessed for neurological deficit|120
    consulted orthopedic spine surgeon|120
    midline tenderness over upper thoracic spine region|120
    suspected spinal cord compression|120
    upper motor neuron involvement|120
    decreased sensation from Th5 dermatome|120
    Medical Research Council Scale 0/5 from L2-S1 on both lower extremities|120
    ASIA impairment scale B|120
    MRI revealed wedging on 5th and 6th thoracal vertebrae|120
    intrathecal infiltration of hyperintensity mass in T2 weighted images|120
    suspected granulomatous infection from Mycobacterium tuberculosis|120
    metastatic bone disease as differential diagnosis|120
    posterior stabilization with pedicle screws and rods system on 4th, 5th, 7th, 8th thoracic spines|168
    transpedicular biopsy on 6th vertebra|168
    3 cc purulent discharge oozing from 6th thoracal body|168
    tissue samples obtained for culture|168
    pathological exam|168
    macroscopically similar to granulation tissue from tuberculous infection|168
    debridement attempted|168
    decompression by laminectomy and flavectomy on 5th and 6th thoracal level|168
    similar granulation tissue found underneath laminae and yellow ligament|168
    postoperative ICU admission|168
    pathological exam revealed chronic inflammation|168
    no tuberculoma|168
    no caseous necrotic formation|168
    no malignant cells|168
    tissue culture revealed Salmonella enterica infection|168
    changed antibiotic regimen to ciprofloxacin 400 mg IV twice daily for two weeks|168
    oral ciprofloxacin 500 mg twice daily for 6 weeks|168
    total 8 weeks therapeutic antibiotic|168
    significant improvement of neurological condition|504
    excellent motoric strength (ASIA E)|504
    free of fever|504
    slight discomfort over surgical scar|504
    pain significantly subsided|504
    independently ambulated with spinal brace|504
    discharged three weeks after surgery|504
    symptom-free at 3 month follow-up|2184
    began exercises to strengthen back|2184
    
    <|eot_id|>
    