70 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
farmer | 0 | 0 | Factual
high-grade fever | -120 | 0 | Factual
generalized body ache | -120 | 0 | Factual
headache | -120 | 0 | Factual
altered sensorium | -24 | 0 | Factual
joint pains | -120 | 0 | Factual
epigastric pain | -120 | 0 | Factual
no drug addiction | 0 | 0 | Negated
no intoxication | 0 | 0 | Negated
inguinal lymphadenopathy | 0 | 0 | Factual
mild generalized rash | 0 | 0 | Factual
no eschar | 0 | 0 | Negated
hemodynamically stable | 0 | 0 | Factual
disoriented | 0 | 0 | Factual
no focal neurological deficit | 0 | 0 | Negated
no neck rigidity | 0 | 0 | Negated
acute febrile illness | 0 | 0 | Factual
undifferentiated fever | 0 | 0 | Factual
malaria | 0 | 0 | Negated
dengue | 0 | 0 | Negated
typhoid | 0 | 0 | Negated
leptospira | 0 | 0 | Negated
scrub typhus antigen card | 0 | 0 | Factual
scrub immunoglobulin M | 0 | 0 | Factual
blood and other body fluid cultures | 0 | 0 | Negated
leukocytosis | 0 | 0 | Factual
mild hyperbilirubinemia | 0 | 0 | Factual
transaminitis | 0 | 0 | Factual
slightly raised international normalized ratio | 0 | 0 | Factual
hepatitis B antigen | 0 | 0 | Negated
hepatitis C antibody | 0 | 0 | Negated
mild fatty infiltration of the liver | 0 | 0 | Factual
tablet doxycycline | 0 | 48 | Factual
defervescence | 48 | 48 | Factual
improved orientation | 48 | 48 | Factual
weakness of both lower limbs | 96 | 96 | Factual
weakness of upper limbs | 96 | 96 | Factual
absent deep tendon reflexes | 96 | 96 | Factual
flexor plantar responses | 96 | 96 | Factual
bladder incontinence | 96 | 96 | Factual
no bowel incontinence | 96 | 96 | Negated
breathing difficulty | 96 | 96 | Factual
respiratory distress | 96 | 96 | Factual
intubated | 96 | 96 | Factual
mechanical ventilation | 96 | 240 | Factual
MRI of the brain | 96 | 96 | Factual
MRI of the cervical spine | 96 | 96 | Factual
nerve conduction velocity | 96 | 96 | Factual
motor sensory demyelinating polyneuropathy | 96 | 96 | Factual
cerebrospinal fluid analysis | 96 | 96 | Factual
intravenous immunoglobulin therapy | 96 | 240 | Factual
tablet rifampicin | 96 | 240 | Factual
improvement in weakness | 240 | 240 | Factual
improvement in respiratory parameters | 240 | 240 | Factual
weaned off ventilator | 240 | 240 | Factual
extubated | 240 | 240 | Factual
oral feeding | 240 | 240 | Factual
limb and chest physiotherapy | 240 | 672 | Factual
discharged | 672 | 672 | Factual
full neurological recovery | 672 | 672 | Factual