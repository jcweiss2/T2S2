61 years old | 0
    male | 0
    admitted to the emergency treatment unit | 0
    abdominal pain | -72
    distension | -72
    vomiting | -72
    constipation | -72
    type 2 diabetes mellitus | -131400
    hypertension | -131400
    febrile | 0
    confused | 0
    low volume pulse | 0
    thready pulse | 0
    pulse rate 130 per min | 0
    blood pressure 70/40 mmHg | 0
    rapid breathing 25 per min | 0
    peripheral oxygen saturation 88% | 0
    distended abdomen | 0
    gas in abdomen | 0
    flank dullness | 0
    diffuse tenderness | 0
    guarding | 0
    rigidity | 0
    absent bowel sounds | 0
    septic shock | 0
    intra-abdominal focus | 0
    admitted to intensive care | 0
    arterial blood gas analysis | 0
    septic screening | 0
    broad-spectrum antibiotics | 0
    30 mL/kg intravenous fluid bolus | 0
    subclavian central venous line insertion | 0
    noradrenaline infusion | 0
    adrenaline infusion | 0
    mean arterial pressure 50 mmHg | 0
    lactate level 15 mmol/L | 0
    invasive arterial pressure monitoring | 0
    increased vasopressor requirement | 0
    elective intubation | 0
    hypovolaemia | 0
    moderately impaired cardiac contractility | 0
    1 L crystalloid administered | 0
    dobutamine infusion | 0
    left lateral decubitus X-ray abdomen | 0
    distended small bowel loops | 0
    no air under diaphragm | 0
    ultrasound abdomen | 0
    moderate ascites | 0
    acute kidney injury | 0
    nasogastric tube insertion | 0
    bilious drainage 500 mL | 0
    random blood sugar 250 mg/dL | 0
    absent urine ketone body | 0
    subcutaneous soluble insulin 6 units | 0
    capillary blood sugar 190 mg/dL | 0
    variable-rate intravenous insulin infusion | 0
    blood urea 8.4 mmol/L | 0
    serum creatinine 2 mg/dL | 0
    normal liver profile | 0
    normal clotting profile | 0
    emergency exploratory laparotomy | 0
    midline laparotomy | 0
    faecal peritonitis | 0
    distended small bowel | 0
    fishbone in distal ileum | 0
    sealed 5 mm perforation | 0
    purulent exudate | 0
    resection of 10 cm distal ileum | 0
    end stomas creation | 0
    peritoneal lavage | 0
    pelvic drainage insertion | 0
    increased vasopressor requirement during surgery | 0
    no urine output | 0
    serum lactate 20 mmol/L | 0
    severe metabolic acidosis | 0
    sodium bicarbonate infusion 20 meq/L | 0
    intravenous sedation | 0
    intravenous analgesia | 0
    cardiac arrest | 8
    passed away | 8
    <|eot_id|>
    