58 years old | 0
African American | 0
alcohol abuse | 0
hepatitis C | 0
transferred to university hospital intensive care unit | 0
sepsis | 0
left hand swelling | -72
left hand pain | -72
malaise | -72
catfish bone injury | -72
nausea | -72
edema of dorsum of the hand | 0
edema of thenar eminence | 0
edema extending to wrist | 0
mild pain on active motion | 0
no erythema | 0
no warmth | 0
no crepitus | 0
normal hand x-ray | 0
compartment pressures measured in thenar space | 4
compartment pressures measured in interossei | 4
compartment pressure recorded at 17 mm Hg | 4
duplex of left upper extremity unremarkable | 0
antibiotics initiated | 0
blood cultures obtained | 0
hand swelling increased moderately | 4-6
digit flexion limited | 4-6
digit extension limited | 4-6
progressive hypotension | 4-6
intubation | 4-6
high-dose vasopressor support | 4-6
blood cultures revealed Edwardsiella tarda | 0
infectious disease consultation requested | 0
multiorgan failure | 36
swelling of entire upper extremity | 36
bullae formation | 36
epidermolysis | 36
ischemia to fingertips | 36
Doppler signals within radial artery | 36
Doppler signals within ulnar artery | 36
bullae over remaining extremities | 36
concern for necrotizing fasciitis | 48
concern for myonecrosis | 48
plastic surgery consultation | 48
taken to operating room | 48
dorsal hand incised | 48
flexor compartments of forearm incised | 48
extensor compartments of forearm incised | 48
evaluation revealed serous fluid | 48
normal muscle appearance | 48
normal soft tissue appearance | 48
skin biopsies revealed no necrosis | 48
muscle biopsies revealed no necrosis | 48
intraoperative cultures negative | 48
multiorgan failure progressed | 120
severe acidosis | 120
hemodynamic instability | 120
patient expired | 120
