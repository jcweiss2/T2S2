69 years old | 0
male | 0
high-grade B-cell non-Hodgkin lymphoma | 0
severe chronic ischemic heart disease | 0
arterial hypertension | 0
chronic bronchitis | 0
type 2 diabetes mellitus | 0
admitted to the hospital | 0
fever | -48
weakness | -48
diarrhoea | -48
dyspnoea | -48
septic shock | 0
hypotension | 0
tachycardia | 0
neutropenia | 0
WBC count 0.68 × 10^9/L | 0
ANC 0.6 × 10^9/L | 0
CRP concentration 120 mg/L | 0
kidney injury | 0
lactate acidosis | 0
electrolyte imbalance | 0
hyponatremia | 0
hypokalemia | 0
bilateral opacities at the bases of the lungs | 0
oral candidiasis | 0
herpes labialis | 0
E. coli | 0
C. difficile | 0
meropenem | 0
linezolid | 0
norepinephrine | 0
fluid resuscitation | 0
CRP peaked 286 mg/L | 48
kidney injury progressed | 48
oligoanuric acute kidney insufficiency | 48
continuous diuretic support | 48
fever returned | 312
diarrhoea returned | 312
E. coli | 312
C. difficile | 312
piperacillin | 312
tazobactam | 312
amikacin | 312
fidaxomicin | 312
peripherally inserted central catheter extracted | 312
catheter tip culture negative | 312
recovered | 648
discharged | 648
enrolled in telemedicine project | 648
rituximab | 0
gemcitabine | 0
oxaliplatin | 0
fever | 0
diarrhoea | 0
vomiting | 0
hypertension | 0
tachycardia | 0
ventricular extrasystoles | 0
WBC 3.16 × 10^9/L | 0
ANC 2.95 × 10^9/L | 0
CRP 32 mg/L | 0
intravenous hydration | 0
cefepime | 0
amikacin | 0
granulocyte colony-stimulating factor | 0
E. coli | 0
recovered | 240
discharged | 240