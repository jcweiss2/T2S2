72 years old | 0
female | 0
admitted to the hospital | 0
cough | -168
shortness of breath | -168
weakness | -168
hypoxic | -168
oxygen saturation of 80% | -168
COVID-19 pneumonia | -168
bacterial pneumonia | -168
sepsis | -168
hypertension | 0
hypothyroidism | 0
obesity | 0
dexamethasone | 0
albuterol | 0
nasal cannula oxygen | 0
enoxaparin | 0
vancomycin | 0
meropenem | 0
doxycycline | 0
intravenous piggyback set to gravity containing doxycycline 100 mg in 100 mL of normal saline infiltrated | -48
mild swelling | -48
pain | -48
worsening respiratory failure | -96
endotracheal intubation | -96
transfer to the intensive care unit | -96
norepinephrine | -96
proned periodically | -96
improvement of respiratory status | -96
left hand displayed considerably worsened swelling | -384
large dorsal purplish bulla | -384
pain in her hand and distal forearm | -384
unable to flex her fingers | -384
denies numbness | -384
vascular surgery consulted | -384
no signs of arterial insufficiency on arterial duplex ultrasound and Doppler examination | -384
computed tomography demonstrated a hematoma of the dorsal wrist | -384
venous duplex ultrasound did not find any evidence of venous thrombosis | -384
nonsurgical management and local wound care recommended | -384
hand surgery consulted | -408
hematoma evacuation | -408
faint ulnar and radial Doppler signals | -408
cool fingers | -408
considerable blistering | -408
mottling | -408
intrinsic minus posturing | -408
worsened pain with the passive extension of the interphalangeal and metacarpophalangeal joints of the digits and thumb | -408
limited active range of motion | -408
compartment pressures of 52 and 54 mm Hg in the hypothenar eminence | -408
compartment pressures of 40 and 42 mm Hg in the thenar eminence | -408
delta pressures ranged between -2 and 30 mm Hg | -408
compartment syndrome | -408
emergent decompressive fasciotomy of the left hand | -408
thenar and hypothenar muscle groups were severely edematous | -408
herniated through the volar incisions | -408
two radial incisions on the dorsal surface over the second and fourth metacarpals were made | -408
releasing the interosseous and adductor compartments | -408
evacuating the dorsal hematoma | -408
all compartments were released | -408
dorsal fasciotomies were closed loosely | -408
extubated | -24
reported improved pain | -24
range of motion of all digits was limited | -24
improved from prior to surgery | -24
flexion and extension at the MCP and IP joints to <10° of all digits | -24
improvement in swelling | -24
improved flexion and extension of all digits to >10° at the MCP and IP joints | 0
oppose her thumb as far as her middle finger | 0
discharged | 168
continued to recover function through physical therapy | 168
progressing to form a composite fist | 168
fully extend fingers | 168
necrotic eschar on the dorsal hand was debrided serially | 168
wound was fully healed | 504
mild scar contracture | 504
some limitation of wrist flexion to 60° | 504
full wrist extension | 504
full range of motion in the digit IP and MCP joints | 504
forearm supination and pronation | 504
wrist radial and ulnar deviation | 504
Disabilities of the Arm, Shoulder, and Hand score was 60 of 100 | 504
very satisfied with her outcome | 504
range of motion | 504
ability to perform activities of daily living | 504
resolution of neuropathic pain symptoms | 504