28 years old | 0
female | 0
SLE | -8760
ESKD | -8760
lupus nephritis Grade VI | -8760
maintenance hemodialysis | -8760
hydroxychloroquine | -8760
mycophenolic acid | -8760
fever | -216
cough | -216
fatigue | -216
dyspnea | -216
contact with sister | -168
sister had flu-like illness | -168
admitted to emergency department | 0
fever 38.8°C | 0
persistent cough | 0
fatigue | 0
progressive dyspnea | 0
decreased breath sounds | 0
crepitations at lung bases | 0
SpO2 88% | 0
minor respiratory distress | 0
received 5 L oxygen | 0
desaturated | 0
SpO2 75% | 0
septic shock | 0
intubated | 0
resuscitated with normal saline | 0
noradrenaline | 0
electrocardiogram normal | 0
cardiac enzymes normal | 0
echocardiography normal | 0
lymphocytopenia | 0
increased C-reactive protein | 0
increased d-dimer | 0
increased lactate dehydrogenase | 0
increased ferritin | 0
elevated blood urea nitrogen | 0
elevated creatinine | 0
emergency contrast chest CT scan | 0
bilateral ground-glass opacities | 0
COVID-19 confirmed by RT-PCR | 0
admitted to ICU | 0
full diagnostic work-up | 0
evaluation for SLE flare | 0
elevated anti-dsDNA | 0
decreased serum complement levels | 0
no anti-cardiolipin antibodies | 0
no anti-β2GP1 antibodies | 0
no lupus anticoagulant | 0
no thrombocytopenia | 0
empiric therapy for COVID-19 | 0
lopinavir/ritonavir | 0
ribavirin | 0
piperacillin/tazobactam | 0
prophylactic anticoagulation | 0
hemodialysis every 48 hours | 0
supportive ICU care | 0
double lumen central line inserted | 0
SpO2/FiO2 ratio 150 | 72
prone positioning ventilation | 72
initiation of steroid treatment | 72
pulse methylprednisolone therapy | 72
SpO2/FiO2 ratio 300 | 96
vasopressors discontinued | 96
extubated | 144
high flow nasal cannula | 144
lymphocytes increased | 144
inflammatory biomarkers decreased | 144
oxygen supportive care discontinued | 240
methylprednisolone tapered down | 240
RT-PCR test for COVID-19 negative | 408
repeated microbiology tests negative | 408
discharged to home isolation | 456
maintenance oral steroid therapy | 456