50 years old | 0
female | 0
pruritic urticarial rash | -24
allergic reaction | -24
hypertension | 0
hepatitis C | 0
diabetes mellitus | 0
amlodipine | -24
metoprolol succinate | -24
hydrocortisone | -2
antihistamines | -2
chest pressure | 2
heart palpitations | 2
diaphoresis | 2
respiratory distress | 2
afebrile | 2
respiratory rate 23 breaths per minute | 2
heart rate 155 bpm | 2
blood pressure 220/100 mmHg | 2
diffuse crackles at bilateral lung fields | 2
anion gap metabolic acidosis | 2
respiratory acidosis | 2
lactic acid 14.9 mmol/L | 2
pulmonary edema | 2
bilateral lobe infiltrates | 2
nitroglycerin | 2
enalaprilat | 2
noriepinephrine | 4
vasopressin | 4
bilateral lower lobe consolidation | 4
liver hemangioma | 4
left adrenal gland enlargement | 4
sinus tachycardia | 4
nonspecific ST changes | 4
global dysfunction | 4
decreased ejection fraction | 4
life flighted to cardiac intensive care unit | 4
cardiogenic shock | 4
myocarditis | 4
sepsis | 4
pneumonia | 4
WBC 12.3 × 103/μL | 4
Haemoglobin 13.2 g/dL | 4
Platelets 248 × 103/μL | 4
Sodium 140 mEq/L | 4
Potassium 3 mEq/L | 4
Chloride 98 mEq/L | 4
HCO 12 mEq/L | 4
BUN 17 mg/dL | 4
Creatinine 1.8 mg/dL | 4
Glucose 734 mg/dL | 4
Anion gap 30 mEq/L | 4
Albumin 4 g/dL | 4
AST 50 U/L | 4
ALT 67 U/L | 4
Total bilirubin 0.3 mg/dL | 4
Alkaline phosphatase 107 U/L | 4
pH, arterial 7.00 | 4
pCO2, arterial 45 mmHg | 4
pO2, arterial 66 mmHg | 4
Lactic acid 134 mg/dL | 4
Serum ketones Negative | 4
CK 1637 U/L | 4
MB 126 ng/mL | 4
Troponin T 0.35 ng/mL | 4
nonsmoker | 0
socially drank alcohol | 0
never used recreational drugs | 0
metoprolol succinate 25 mg twice a day | 0
amlodipine 5 mg daily | 0
unremarkable surgical history | 0
unremarkable family history | 0
vasopressors | 4
intra-aortic balloon pump | 4
broad spectrum antibiotics | 4
cortisol stimulation test | 4
normal | 4
nephrology consultation | 4
nonoliguric acute kidney injury | 4
ischemic acute tubular necrosis | 4
contrast-induced nephropathy | 4
renal replacement therapy | 4
hemodynamics improved | 120
intra-aortic balloon pump discontinued | 120
vasopressors discontinued | 120
sodium nitropruside drip | 120
four drug oral blood pressure regimen | 120
weaned off ventilator support | 120
extubated | 120
creatinine plateaued at 1.2 mg/dL | 120
workup for functional adrenal mass | 120
diagnosis of pheochromocytoma | 120
free plasma metanephrine 1877 pg/mL | 120
free plasma normetanephrine 4560 pg/mL | 120
plasma epinephrine 3081 pg/mL | 120
plasma noriepinephrine 8968 pg/mL | 120
24-h urine metanephrine 4462 μg/24 h | 120
24-h urine normetanephrine 2912 μg/24 h | 120
24-h total urine metanephrine 7374 μg/24 h | 120
abdominal CT scan | 120
MIBG scan | 120
doxazosin | 168
metoprolol succinate 50 mg | 168
amlodipine 10 mg | 168
left adrenalectomy | 168
final pathology | 168
well encapsulated minimally fibroadipose tissue | 168
pheochromocytoma | 168
screened for multiple endocrine neoplasm 2 | 168
negative | 168
discharged home | 240
follow-up | 4320
good blood pressure control | 4320
metoprolol 25 mg twice a day | 4320
amlodipine 5 mg daily | 4320