46 years old | 0
female | 0
intracerebral bleeding | -720
intracerebral hemorrhage at the right basal ganglia region | -720
hospitalized in a neurosurgery center | -720
tracheotomy | -60
pneumonia | -60
conservative treatment | -60
transferred to a rehabilitation center | -60
massive hemorrhage | 0
cyanosis | 0
respiratory failure | 0
shocks | 0
cuff air in tracheotomy tube maximally expanded | 0
bleeding did not stop | 0
tracheotomy tube removed | 0
cuffed endotracheal intubation attempted | 0
cuffed endotracheal tube inserted | 0
bleeding stopped | 0
transferred to an intensive care center | 0
blood test | 0
hemoglobin level decreased | 0
cervical CT | 0
bronchoscopy | 0
conservative treatment continued | 0
transfemoral angiography | 168
diagnosis of TIAF | 168
innominate artery made small luminal outpouching to trachea | 168
transferred to the thoracic surgery unit | 168
operation for TIAF | 168
tracheoplasty with bypass graft | 168
rupture area observed | 168
innominate artery rebuilt | 168
tracheoplasty done | 168
tracheostenosis | 744
inflammation | 744
bronchoscopy | 744
endotracheal balloon dilatation | 744
replacement of Montgomery T-tube | 744
continuation of rehabilitation | 744
survives without further complications | 1056
tracheo-innominate artery fistula reported | -131040
tracheotomy | -131040
diphtheria patient | -131040
incidence of tracheo-innominate artery fistula | 0
mechanism of tracheo-innominate artery fistula | 0
pressure necrosis | 0
mechanical erosion | 0
necrosis | 0
invasion into innominate artery | 0
sepsis | 0
radiation therapy | 0
stoma infection | 0
steroid therapy | 0
malnutrition | 0
tracheal mucosal injury | 0
fistulas may occur | 0
common carotid artery | 0
innominate vein | 0
inferior thyroid artery | 0
internal mammary artery | 0
aortic arch | 0
risk factors | 0
long-term mechanical ventilation | 0
high ventilator peak pressures | 0
low-lying tracheostomy sites | 0
previous tracheal resections | 0
high cuff pressures | 0
preventive measures | 0
appropriate humidity | 0
clean maintenance | 0
infection management | 0
smooth tracheal suction | 0
excessive extension of neck | 0
special attention | 0
short neck | 0
children | 0
appropriate size of the tracheotomy tube | 0
excessive movements | 0
head injuries | 0
early detachment of the artificial respirator | 0
appropriate treatment | 0
tracheal granuloma | 0
serious bleeding | 0
tracheo-innominate artery fistula | 0
massive hemorrhage | 0
controlling the hemorrhage | 0
securing the airway | 0
respiratory tract obstruction | 0
respiratory failure | 0
hypovolemic shock | 0
homeostasis | 0
applying pressure | 0
overinflation of the tube cuff | 0
tracheostomy tube removed | 0
oropharyngeal intubation | 0
cuffed oral endotracheal tube | 0
balloon cuff expanded | 0
stomal hemorrhage controlled | 0
digit compression | 0
innominate artery compressed | 0
manubrium | 0
pretracheal fascial plane | 0
tracheostomy wound | 0
index finger | 0
distal compression | 0
pressure continued | 0
transfer of the patient | 0
operating room | 0
homeostasis does not work | 0
overinflation of the balloon cuff | 0
repeatedly carried out | 0
position of oral endotracheal tube | 0
up and down | 0
patient transported | 0
operation room | 0
rigid bronchoscopic examination | 0
trachea | 0
re-bleeding | 0
surgery prepared | 0
evidence of hemorrhage | 0
necrosis | 0
ulcer | 0
indication for surgery | 0
angiography | 0
diagnostic option | 0
lack of time | 0
result may be normal | 0
bleeding at the time of test | 0
ceased already | 0
full median sternotomy | 0
approach for the repair of TIAF | 0
ligation of the innominate artery | 0
resection of a segment of the innominate artery | 0
oversewing of the ends | 0
better survival rate | 0
interposition grafting | 0
direct vascular repair | 0
suturing | 0
innominate artery rebuilt | 0
artificial blood vessel | 0
right subclavian artery | 0
right aorta | 0
tracheoplasty | 0
fifth costal cartilage | 0
domestic research | 0
tracheo-innominate artery fistula after stroke | 0
damage to trachea | 0
repetitive opisthotonos | 0
head trauma | 0
evidence of ulceration | 0
epileptic convulsion | 0
neurological spasticity | 0
abnormal arching of the neck | 0
formation of the TIAF | 0
increased pressure | 0
cannula against the anterior tracheal wall | 0
experience with an unknown case | 0
preventive measures | 0
patients with tracheotomy | 0
frequent observation | 0
rehabilitation unit | 0
appropriate posture | 0
restriction of excessive movements | 0
continuous management of tracheal tubes | 0
sustained management of erosion | 0
ulceration in the trachea | 0
pressure between the anterior wall of trachea | 0
tracheal tube | 0
hemorrhage occurring after tracheotomy | 0
fatal consequences | 0
thorough knowledge | 0
appropriate treatment | 0
prompt execution of treatment | 0