27 years old | 0
male | 0
admitted to the hospital | 0
gingival bleeding | -144
haematuria | -144
haematochezia | -144
pain in the right lower abdomen | -144
swelling | -144
numbness | -144
weakness of the left lower limb | -144
dizziness | -144
fever | -144
cough | -144
expectoration | -144
chest tightness | -144
palpitation | -144
WBC 23.36 × 109/l | -144
neutrophil percentage 68.1% | -144
haemoglobin 110 g/l | -144
platelet count 276 × 109/l | -144
urinary protein 3+ | -144
urinary occult blood 3+ | -144
occult blood in the stool | -144
APPT 85.4 s | -144
prothrombin time 16.6 s | -144
alanine transaminase 86 U/l | -144
albumin 35 g/l | -144
creatinine 65 µmol/l | -144
blood glucose 7.1 mmol/l | -144
anti-infection treatment | -24
haemostasis treatment | -24
symptomatic treatment | -24
gastrointestinal decompression | -24
enema | -24
crystal and colloidal liquid replenishment | -24
volume expansion | -24
blood transfusion | -24
admitted to the intensive care unit | -24
abdominal CT | -24
liver morphology irregular | -24
liver cirrhosis not excluded | -24
WBC 34.24 × 109/l | 0
Hb 66 g/l | 0
APTT 130 s | 0
transferred to Qilu Hospital | 0
past medical history of HBV | 0
no history of drug or food allergy | 0
no history of trauma | 0
no history of surgery | 0
no history of blood transfusion | 0
smoking history | 0
family history of diabetes mellitus | 0
family history of hypertension | 0
no family history of genetic diseases | 0
no family history of infections | 0
body temperature 36.8°C | 0
heart rate 146 beats/min | 0
respiration rate 22 breaths/min | 0
blood pressure 94/66 mmHg | 0
saturation of peripheral oxygen 98% | 0
poor spirit | 0
drowsiness | 0
anaemic appearance | 0
sclera yellow stained | 0
bilateral pupils equal in size | 0
pupils sensitive to light reflection | 0
bleeding at the right subclavian vein catheterization | 0
respiratory sounds thick | 0
no dry and wet rales | 0
heart rate 146 beats/min | 0
rhythm uniform | 0
no pathological murmurs | 0
abdomen bulging | 0
no muscle tension | 0
ecchymosis on both sides of the waist | 0
skin around the umbilicus blue-purple | 0
left lower abdomen tender | 0
right lower abdomen tender | 0
hard mass in the left lower abdomen | 0
liver and spleen not felt | 0
groin circumference of the left lower limb 72 cm | 0
groin circumference of the right lower limb 62 cm | 0
Babinski signs negative | 0
coagulation factor V 54% | 0
coagulation factor VII 28% | 0
coagulation factor VIII 1% | 0
coagulation factor IX 85% | 0
diet prohibition | 0
meropenem anti-infection treatment | 0
vitamin K1 | 0
phenolsulfonamethylamine | 0
aminometrinic acid | 0
batroxobin haemostatic | 0
omeprazole acid suppression | 0
octreotide to inhibit pancreatin secretion | 0
magnesium isoglycyrrhizin | 0
reduced glutathione liver protection | 0
entecavir to inhibit HBV replication | 0
plasma supplements | 0
cold precipitation | 0
infusion of red blood cells | 0
nutrition and symptomatic support treatment | 0
transferred to the Department of Poisoning and Occupational Diseases | 24
black stools | 72
red blood cells and plasma infused | 72
glucose water test | 120
acidified serum haemolysis test | 120
plasma free Hb 41.9 mg/l | 120
direct antiglobulin test | 120
anticoagulant rodenticide not detected | 120
black stools decreased | 168
ecchymosis deepened | 168
blood cultures no anaerobic growth | 168
blood cultures no bacterial growth | 168
coagulation factor V 89% | 168
coagulation factor VII 85% | 168
coagulation factor VIII 1% | 168
coagulation factor IX 92% | 168
tumour markers detected | 288
ferritin 709 ng/ml | 288
carbohydrate antigen (CA) 19-9 294.3 U/ml | 288
CA 125 306.1 U/ml | 288
neuron specific enolase 27.27 ng/ml | 288
immune system examination | 288
systemic lupus erythematosus excluded | 288
bone marrow puncture | 288
abdominal CT showed cholecystitis | 336
swollen lymph nodes in the retroperitoneal area | 336
multiple strip-like low-density shadows in the abdomen and pelvis | 336
peritoneal thickening and soft tissue swelling in the left chest and abdominal wall | 336
laboratory indices improved | 504
blood sent to Haemophilia Diagnosis and Treatment Centre | 504
coagulation factor VIII 5.2% | 504
factor VIII inhibitor 1.5 BU | 504
gene mutation screening | 504
p.Y471H mutation in the PLAT gene | 504
p.Y244Y mutation in the SERPINE1 gene | 504
treatment changed to prednisone | 504
transferred to the Department of Haematology | 504
cryoprecipitate via intravenous drip | 504
symptoms and laboratory examination results improved | 528
discharged | 528
follow-up examinations | 744
follow-up CT of the hip joints | 744
swelling of the left iliopsoas muscle | 744
bleeding cannot be excluded | 744
coagulation factor VIII increased | 744
factor VIII antibody not detected | 744