70 years old | 0
female | 0
admitted to the hospital | 0
hereditary hemorrhagic telangiectasia | -0
severe pulmonary hypertension | -0
diastolic heart failure | -0
mild obstructive sleep apnea | -0
hyperlipidemia | -0
gastroesophageal reflux | -0
hypertension | -0
scheduled for open radical nephrectomy | 0
mass localized to the lower pole | -0
concerning for malignancy | -0
exertional dyspnea | -1092
left and right heart catheterization | -1092
angiographically normal-appearing coronary arteries | -1092
right coronary artery fistula | -1092
severe precapillary pulmonary hypertension | -1092
mean pulmonary artery pressure 45 mmHG | -1092
pulmonary capillary wedge pressure 8 mmHG | -1092
pulmonary vascular resistance 7.8 WU | -1092
cardiac index 3.0 L/min/m2 | -1092
started on sildenafil | -1092
WHO class III symptoms improved to class I or II | -1092
RV enlargement with decreased function | -0
moderate-to-severe eccentric TR | -0
moderately-to-severely dilated right atrium | -0
Doppler-derived estimated systolic pulmonary artery pressure >100 mmHg | -0
low normal left ventricular function | -0
frequent epistaxis | -0
episodes of gastrointestinal bleeding | -0
arterial venous malformations | -0
nasal and upper-gastrointestinal endoscopy | -0
mild OSA treated with CPAP | -0
heart failure with preserved ejection fraction | -0
anemia | -0
30-pound weight loss | -0
synthetic liver dysfunction | -0
elevated PT INR | -0
low albumin | -0
multidisciplinary perioperative consultation | 0
risks, benefits and alternatives discussed | 0
increased risk due to severe pulmonary hypertension | 0
patient consented to proceed with surgery | 0
ASA physical status IV | 0
preoperative transthoracic echocardiography | 0
similar findings to previous echocardiogram | 0
chest x-ray | 0
cardiovascular silhouette at the upper limits of normal | 0
prominent pulmonary arteries | 0
recommended to continue sildenafil | 0
exercise tolerance greater than 4 METS | 0
partial vs. radical nephrectomy discussed | 0
patient elected to have removal of entire left kidney | 0
minimal dyspnea with daily activities | 0
occasionally experiencing lightheadedness during exertion | 0
no angina | 0
no significant orthopnea | 0
no paroxysmal nocturnal dyspnea | 0
no significant edema | 0
no hepatosplenomegaly | 0
frequent epistaxis episodes | 0
elevated PT/INR 1.3 | 0
oral vitamin K ordered | 0
outpatient workup | 0
no evidence of decompensated liver disease | 0
low-grade fibrosis on fibroscan | 0
continued medications | 0
admitted on the day of surgery | 0
no significant changes to medical condition | 0
vitals | 0
temperature 36.6 C | 0
blood pressure 138/77 mmHG | 0
respiratory rate 18/min | 0
pulse oximetry 96% on room air | 0
pain 0/10 | 0
airway exam reassuring | 0
no bleeding episodes | 0
denied new or worsening shortness of breath | 0
denied chest discomfort | 0
ECG | 0
normal sinus rhythm | 0
rate 95 | 0
premature ventricular complexes | 0
inferior and anterolateral T-wave changes | 0
laboratory data | 0
hemoglobin 11.2 g/dl | 0
hematocrit 35.4% | 0
large-bore IV access | 0
radial arterial line | 0
induction of general anesthesia | 0
IV fentanyl | 0
etomidate | 0
lidocaine | 0
rocuronium | 0
intubated with 7.0-mm endotracheal tube | 0
MAC 3 blade | 0
Cormack-Lehane grade I view | 0
no telangiectasias observed | 0
endotracheal tube position confirmed | 0
pulse oximetry, heart rate, and arterial blood pressure stable | 0
Swan-Ganz catheter placed | 0
severe tricuspid regurgitation | 0
right internal jugular venous 9 fr introducer | 0
initial pulmonary artery pressure 96/46 mmHG | 0
mean pulmonary artery pressure 65 mmHG | 0
systemic arterial pressure 125/74 mmHG | 0
initial arterial blood gas | 0
pH 7.33 | 0
pCO2 43 mmHG | 0
pO2 145 mmHG | 0
HCO3 22.7 mEq/L | 0
correction of hypercarbia and mild acidosis | 0
inhaled nitric oxide 20 ppm initiated | 0
improvement in pulmonary artery pressures | 0
fluid balance maintained | 0
adequate urine output | 0
replacement of blood loss | 0
transversus abdominal plane block | 0
real-time ultrasound guidance | 0
1:1 mixture of 0.25% bupivacaine and 1.3% liposomal bupivacaine | 0
general anesthesia maintained with sevoflurane | 0
total surgical time less than 60 min | 0
open technique with flank incision | 0
patient remained hemodynamically stable | 0
final arterial blood gas analysis | 0
pH 7.38 | 0
pCO2 38 mmHG | 0
pO2 182 mmHG | 0
transferred to surgical intensive care unit | 0
inhaled nitric oxide weened over 3 h | 0
cardiac output and pulmonary artery pressures reached baseline values | 0
no evidence of pulmonary arterial crisis | 0
extubated on postoperative day 0 | 24
noninvasive positive pressure ventilation | 24
weened to nasal cannula | 24
pulse oximetry saturation 93-96% | 24
pain adequately controlled | 24
numerical rating scale <4 | 24
multimodal regimen | 24
PO and IV acetaminophen | 24
Ultram | 24
incremental doses of fentanyl | 24
expected return of bowel function | 24
no placement of nasogastric tube | 24
able to tolerate oral diet | 48
transferred to step-down unit | 48
able to ambulate with assistance | 48
discharged to home on postoperative day 3 | 72
pathologic specimens returned as renal cell carcinoma | 72
clear cell type | 72
high-grade histologic pathology | 72
classification pT1bG4 | 72
clear margins | 72
continued to progress as expected | 72
able to resume normal daily activities | 72
turned 71 years old during hospitalization | -0