21 years old | 0
male | 0
obese | 0
admitted to the hospital | 0
cough | -72
fevers | -72
shortness of breath | -72
pleuritic chest pain | -72
light-headedness | -72
near syncope | -72
dyspnoea | -72
COVID-19 | 0
sub-massive PE | 0
unfractionated heparin | 0
hypotensive | 12
massive PE | 12
catheter-directed thrombolysis | 12
improved clinically | 24
discharge planned | 24
acute respiratory failure | 96
hypotension | 96
intubated | 96
cardiac arrest | 96
return of spontaneous circulation | 96
vasopressors | 96
extracorporeal membrane oxygenation | 96
recurrent massive PE | 96
repeat catheter-directed thrombolysis | 96
ventilation parameters improved | 144
vasopressors discontinued | 144
weaning of ECMO | 144
deep venous thrombus | 144
inferior vena cava filter | 144
low-molecular-weight heparin | 144
septic shock | 240
right thigh haematoma | 240
compartment syndrome | 240
surgical debridement | 240
rivaroxaban | 240
discharged | 1248
home | 1608
anticoagulated | 1608
no major adverse events | 1936