72 years old | 0
female | 0
bilateral breast cancers | -6720
occipital neck mass | -12960
shortness of breath | 0
haemoglobin of 4.2 g/dl | 0
cyst | -19680
minor trauma | -19680
mass growth | -720
mass drainage | -720
mass bleeding | -720
portion of the mass fell out | -120
severe diffuse swelling | -240
afebrile | 0
haemodynamically stable | 0
hypertensive to 170/70 mmHg | 0
oxygen saturation of 100% | 0
clear lung sounds | 0
severe upper and lower extremity pitting oedema | 0
baseball-sized malodorous occipital mass | 0
thick oozing purulent drainage | 0
white blood cell count of 8.3*103/μl | 0
haemoglobin of 4.7 g/dl | 0
albumin of 2.9 g/dl | 0
INR of 1.6 | 0
B-type natriuretic peptide (BNP) level of 666 pg/ml | 0
mild interstitial oedema | 0
transfused three units of packed red blood cells | 12
febrile to 101.2 °F | 12
tachycardic to 110 bpm | 12
acetaminophen | 12
temperature increased to 102 °F | 24
heart rate increased to 120 bpm | 24
tachypnoeic to 30 breaths per minute | 24
hypertensive to 200/60 mmHg | 24
lactate level of 2.7 mEq/l | 24
white blood cell count of 24.3*103/μl | 24
E. coli in blood cultures | 24
vancomycin | 24
piperacillin–tazobactam | 24
creatinine doubled | 36
INR of 2.4 | 36
platelet count fell | 36
fibrinogen of 224 mg/dl | 36
d-dimer level of 4668 ng/ml | 36
bilevel non-invasive positive pressure ventilation | 36
transferred to the medical intensive care unit (MICU) | 36
hypotensive to 80/40 mmHg | 36
vasopressors initiated | 36
pyuria with greater than 180 white blood cells per hpf | 36
intubated | 36
sedated | 36
pan-CT scan | 48
obstructing left distal ureteric stone | 48
proximal dilation and hydronephrosis | 48
operating room for extraction and stenting | 60
weaned from vasopressors | 72
extubated | 84
chest X-ray showed increasing pulmonary oedema | 84
oliguric | 84
creatinine elevated to 6.4 mg/dl | 84
urgently dialyzed | 84
transferred back to the general medicine service | 240
discharged from the hospital | 672
haemodialysis | 672
neck mass excised | 672
pathology showed a benign haemangioma | 672
infected haematoma and abscess formation | 672