58 years old | 0
    woman | 0
    hypertension | -175200
    generalized anxiety disorder | -175200
    depression | -175200
    hepatitis C | -175200
    retroperitoneal leiomyosarcoma | -175200
    radical resection | -175200
    segmental duodenectomy | -175200
    inferior vena cava closure | -175200
    nausea | -48
    vomiting | -48
    right upper quadrant abdominal pain | -48
    recurrent disease | -48
    chemotherapy | -48
    neutropenic fever | -48
    neutropenic fever | -48
    ifosfamide dose reduction | -48
    acute altered mental status | -24
    thiamine prophylaxis | -24
    bisacodyl | -24
    docusate-senna | -24
    clonidine | -24
    losartan | -24
    nifedipine ER | -24
    ondansetron | -24
    dexamethasone | -24
    metoclopramide | -24
    oxycodone ER | -24
    fluconazole | -24
    paroxetine | -24
    confusion | -24
    memory impairment | -24
    inability to follow commands | -24
    incoherent speech | -24
    delirium | -24
    thiamine dose increased | -24
    IV thiamine | -24
    neurological decline | -24
    methylene blue | -24
    paroxetine discontinued | -24
    confusion worsened | 0
    delirium worsened | 0
    sinus tachycardia | 0
    hypertension | 0
    diaphoresis | 0
    fever | 0
    combativeness | 0
    hyperreflexia | 0
    ocular clonus | 0
    spontaneous muscular clonus | 0
    facial tremors | 0
    serotonin syndrome concern | 0
    methylene blue discontinued | 0
    ondansetron discontinued | 0
    lorazepam | 0
    metoprolol | 0
    acetaminophen | 0
    hydromorphone | 0
    transfer to critical care unit | 0
    intubation | 0
    normal laboratory tests | 0
    unremarkable sepsis workup | 0
    normal head imaging | 0
    IV thiamine continued | 0
    supportive care | 0
    mentation improvement | 144
    extubation | 144
    normal memory | 144
    fluent speech | 144
    discharged | 360
    follow-up appointment | 720
    ifosfamide unsafe | 720
    alternative therapy options | 720
    surgical resection | 4320
    no evidence of disease | 4320
    
    
    58 years old|0
    woman|0
    hypertension|-175200
    generalized anxiety disorder|-175200
    depression|-175200
    hepatitis C|-175200
    retroperitoneal leiomyosarcoma|-175200
    radical resection|-175200
    segmental duodenectomy|-175200
    inferior vena cava closure|-175200
    nausea|-48
    vomiting|-48
    right upper quadrant abdominal pain|-48
    recurrent disease|-48
    chemotherapy|-48
    neutropenic fever|-48
    neutropenic fever|-48
    ifosfamide dose reduction|-48
    acute altered mental status|-24
    thiamine prophylaxis|-24
    bisacodyl|-24
    docusate-senna|-24
    clonidine|-24
    losartan|-24
    nifedipine ER|-24
    ondansetron|-24
    dexamethasone|-24
    metoclopramide|-24
    oxycodone ER|-24
    fluconazole|-24
    paroxetine|-24
    confusion|-24
    memory impairment|-24
    inability to follow commands|-24
    incoherent speech|-24
    delirium|-24
    thiamine dose increased|-24
    IV thiamine|-24
    neurological decline|-24
    methylene blue|-24
    paroxetine discontinued|-24
    confusion worsened|0
    delirium worsened|0
    sinus tachycardia|0
    hypertension|0
    diaphoresis|0
    fever|0
    combativeness|0
    hyperreflexia|0
    ocular clonus|0
    spontaneous muscular clonus|0
    facial tremors|0
    serotonin syndrome concern|0
    methylene blue discontinued|0
    ondansetron discontinued|0
    lorazepam|0
    metoprolol|0
    acetaminophen|0
    hydromorphone|0
    transfer to critical care unit|0
    intubation|0
    normal laboratory tests|0
    unremarkable sepsis workup|0
    normal head imaging|0
    IV thiamine continued|0
    supportive care|0
    mentation improvement|144
    extubation|144
    normal memory|144
    fluent speech|144
    discharged|360
    follow-up appointment|720
    ifosfamide unsafe|720
    alternative therapy options|720
    surgical resection|4320
    no evidence of disease|4320

    58 years old | 0
    woman | 0
    hypertension | -175200
    generalized anxiety disorder | -175200
    depression | -175200
    hepatitis C | -175200
    retroperitoneal leiomyosarcoma | -175200
    radical resection | -175200
    segmental duodenectomy | -175200
    inferior vena cava closure | -175200
    nausea | -48
    vomiting | -48
    right upper quadrant abdominal pain | -48
    recurrent disease | -48
    chemotherapy | -48
    neutropenic fever | -48
    neutropenic fever | -48
    ifosfamide dose reduction | -48
    acute altered mental status | -24
    thiamine prophylaxis | -24
    bisacodyl | -24
    docusate-senna | -24
    clonidine | -24
    losartan | -24
    nifedipine ER | -24
    ondansetron | -24
    dexamethasone | -24
    metoclopramide | -24
    oxycodone ER | -24
    fluconazole | -24
    paroxetine | -24
    confusion | -24
    memory impairment | -24
    inability to follow commands | -24
    incoherent speech | -24
    delirium | -24
    thiamine dose increased | -24
    IV thiamine | -24
    neurological decline | -24
    methylene blue | -24
    paroxetine discontinued | -24
    confusion worsened | 0
    delirium worsened | 0
    sinus tachycardia | 0
    hypertension | 0
    diaphoresis | 0
    fever | 0
    combativeness | 0
    hyperreflexia | 0
    ocular clonus |A|0
    spontaneous muscular clonus | 0
    facial tremors | 0
    serotonin syndrome concern | 0
    methylene blue discontinued | 0
    ondansetron discontinued | 0
    lorazepam | 0
    metoprolol | 0
    acetaminophen | 0
    hydromorphone | 0
    transfer to critical care unit | 0
    intubation | 0
    normal laboratory tests | 0
    unremarkable sepsis workup | 0
    normal head imaging | 0
    IV thiamine continued | 0
    supportive care | 0
    mentation improvement | 144
    extubation | 144
    normal memory | 144
    fluent speech | 144
    discharged | 360
    follow-up appointment | 720
    ifosfamide unsafe | 720
    alternative therapy options | 720
    surgical resection | 4320
    no evidence of disease | 4320