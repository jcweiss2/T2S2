56 years old | 0
male | 0
admitted to the hospital | 0
intermittent chest tightness | -168
shortness of breath | -168
worsening of symptoms | -24
tremor of the hands | -24
loss of appetite | -24
general malaise | -24
loss of consciousness | -24
no history of alcohol consumption | 0
no history of drug abuse | 0
no history of hypertension | 0
no history of diabetes | 0
no history of heart diseases | 0
no family history of hypertension | 0
no family history of diabetes | 0
no family history of heart diseases | 0
abdomen was soft | 0
right upper quadrant tenderness | 0
no rebound pain | 0
no muscle tension | 0
body temperature 39.2 °C | 0
blood pressure 98/56 mmHg | 0
heart rate 84 beats per min | 0
respiratory rate 26 breaths per min | 0
white blood cell count was 22.22×10^9/L | 0
neutrophil percentage was 91.7% | 0
platelet count was 26 × 10^9/L | 0
pH was 7.28 | 0
PCO2 was 27 mmHg | 0
PO2 was 64 mmHg | 0
HCO3- was 12.7 mmol/L | 0
BE was -12.5 mmol/L | 0
C-reactive protein level was > 90 mg/L | 0
interleukin 6 was > 5000 pg/mL | 0
procalcitonin was > 100 ng/mL | 0
myoglobin was > 2000 ug/L | 0
cranial computed tomography showed soft tissue of the posterior top of the nasopharynx was slightly thicker | 0
thoracic CT showed bilateral pneumonia | 0
thoracic CT showed lung air sac in the right lung apex | 0
thoracic CT showed multiple nodules in bilateral lungs | 0
thoracic CT showed bilateral pleural effusion | 0
abdominal and pelvic CT showed foci with a slightly lower density in the right lobe of the liver | 0
abdominal and pelvic CT showed mixed density in segment IV of the liver near the first porta hepatis | 0
needle-like high-density shadow in the liver | 0
drainage from the indwelling gastric tube was brown | 0
purulent infection | 0
history of eating fish a few days before the onset of disease | -72
fishbone puncture through the stomach wall and into the liver | 0
PLA caused by fishbone puncture | 0
severe pneumonia | 0
acute respiratory failure | 0
septic shock | 0
anti-inflammatory rescue therapy | 0
electrolyte correction | 0
nutritional support | 0
recurrent fever | 192
inflammatory index did not decrease | 192
repeat abdominal CT showed combined density | 192
PLA was considered | 192
laparoscopic exploration | 216
inspection hole was made above the navel | 216
introduction of the laparoscope | 216
three trocars were introduced | 216
dense adhesions between the pylorus and hepatic hilum | 216
liver was obviously swollen at the root of the ligamentum teres | 216
incision | 216
white foreign body about 2 cm long was found | 216
fishbone was confirmed after removal | 216
abscess cavity was found | 216
abscess cavity was incised | 216
white pus was drained | 216
abscess cavity was expanded | 216
drainage tube was placed | 216
patient recovered smoothly | 240
small amount of reddish drainage fluid was observed | 240
inflammatory indexes decreased | 264
symptoms and discomfort disappeared | 264
drainage tube was removed | 264
patient was discharged | 288
follow-up at 2 wk after discharge was unremarkable | 432
follow-up at 2 mo after discharge was unremarkable | 864