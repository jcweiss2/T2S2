53 years old | 0
male | 0
admitted to the hospital | 0
exertional dyspnea | -168
productive cough | -960
thymectomy | -1200
adjuvant radiotherapy | -1200
diagnosed with sarcoidosis | -60
transbronchial lung biopsy | -60
anti-tuberculosis chemotherapeutic regimen | -10
cavitary lesion detected | -10
blood pressure 90/60 mmHg | 0
body temperature 39.3 | 0
pulse rate 152 beats per minute | 0
respiration rate 32 breaths per minute | 0
inspiratory crackles in both lower lung fields | 0
haziness and disseminated nodules in both lung fields | 0
conglomerated cavities in the right upper lobe | 0
multiple micronodular densities and multiple cavitary nodules | 0
ground glass opacity (GGO) in both lower lobes | 0
white blood cell count 3500 cells/mm3 | 0
hemoglobin 15.2 g/dL | 0
platelet cell count 253,000 cells/mm3 | 0
erythrocyte sedimentation rate 36 mm/h | 0
C-reactive protein level 17.29 mg/dL | 0
mildly elevated aspartate aminotransferase (AST) level | 0
normal renal function | 0
HIV test negative | 0
arterial blood gas analysis | 0
pH 7.44 | 0
PaCO2 34.0 mmHg | 0
PaO2 60.5 mmHg | 0
bicarbonate (HCO3) level 22.8 mmol/L | 0
SaO2 91.9% | 0
admitted to the intensive care unit | 0
bronchoalveolar lavage (BAL) | 0
cell count from the BAL fluid 119/µL | 0
cell differential showed 30% macrophages | 0
cell differential showed 60% lymphocytes | 0
cell differential showed 10% neutrophils | 0
polymerase chain reaction (PCR) positive for Pneumocystis jirovecii | 0
direct florescent antibody (DFA) positive for Pneumocystis jirovecii | 0
culture for cytomegalovirus (CMV) negative | 0
trimethoprim/sulfamethoxazole administered | 0
methylprednisolone administered | 0
neutrophil dihydrorhodamine test normal | 0
T lymphocytes (CD3) 290/µL | 0
B lymphocytes (CD19) 0/µL | 0
CD4 148/µL | 0
CD8 132/µL | 0
immunoglobulin levels low | 0
IgG 507 mg/dL | 0
IgA 31 mg/dL | 0
IgM <3 mg/dL | 0
video-assisted thoracoscopic biopsy | 0
biopsy specimens revealed diffuse thickening of the alveolar wall | 0
fibrosis and lymphocyte infiltration | 0
analysis of a smear of the specimen for acid-fast bacilli negative | 0
immunohistochemical analysis for CMV, HSV, and adenovirus antigens negative | 0
diagnosed with Good's syndrome | 0
supportive ventilatory care | 0
antibiotic treatment for acute respiratory distress syndrome | 0
intravenous immunoglobulin (IVIG) infusions | 0
pneumonia and diarrhea did not improve | 2160
infection worsened | 2160
culture of the pleural fluid and material from the catheter tip showed Candida albicans | 2160
died of septic shock and multi-organ failure | 2160