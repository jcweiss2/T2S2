6 years old | 0
female | 0
right wrist swelling | -48
right wrist pain | -48
stepped on right wrist | -48
moderate pain | -48
pain worsened | -24
redness | -24
swelling of the joint | -24
subjective fever | -24
febrile at 39.4°C | 0
tachycardic with heart rate of 140 bpm | 0
wrist swollen | 0
erythematous | 0
tender to palpation | 0
exquisite pain elicited by motion | 0
limited range of motion of the joint | 0
elevated erythrocyte sedimentation rate (ESR) at 40 mm/h | 0
elevated C-reactive protein (CRP) at 13.5 mg/dL | 0
blood cultures drawn | 0
Orthopedic Surgery consultation | 0
joint aspiration | 0
extraction of frankly purulent fluid | 0
Gram stain demonstrated gram-positive cocci with numerous neutrophils | 0
fluid sent for culture | 0
admitted to the hospital | 0
treatment with intravenous (IV) clindamycin | 0
arthrotomy | 24
incision of the joint capsule | 24
seropurulent fluid expressed | 24
joint space copiously irrigated | 24
continued IV clindamycin | 24
repeat ESR at 85 mm/h | 48
repeat CRP at 11 mg/dL | 48
afebrile | 48
pain well controlled by acetaminophen | 48
joint aspiration fluid culture positive for Streptococcus pyogenes | 72
blood culture positive for Streptococcus pyogenes | 72
Infectious Disease consultation | 72
antibiotic regimen switched to IV cefazolin | 72
repeat arthrotomy | 96
no return of fluid on joint entry | 96
joint irrigated and closed | 96
continued IV cefazolin | 96
serial ESR and CRP trending downward | 96
repeat blood culture | 48
no growth after 48 hours | 48
discharged | 144
oral cephalexin course | 144
ESR normalized | 168
CRP normalized | 168
completion of oral antibiotic course | 168
