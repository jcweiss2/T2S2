24 years old | 0
lady | 0
admitted to ICU | 0
refractory status epilepticus | 0
history of repeated hospital admission for seizure attacks | -672
difficult peripheral intravenous access | 0
central vein catheterized | 0
seizure controlled on four anti-epileptic medications | 0
intravenous levetiracetam | 0
sodium valproate | 0
phenytoin | 0
septic shock | 0
ventilator associated pneumonia (VAP) | 0
coagulopathic | 0
platelet count of 48,000/cu mm | 0
prothrombin time of 21 s | 0
international normalized ratio of 1.75 | 0
intravenous nor-adrenaline support | 0
intravenous Colistin | 0
intravenous tigecycline | 0
mechanical ventilatory support | 0
volume assist control mode of ventilation | 0
fraction of inspired oxygen of 0.5 | 0
positive end-expiratory pressure of 10 cm of H2O | 0
intravenous midazolam 2 mg as required | 0
Richmond Agitation Sedation Scale (RASS) of zero | 0
delirious | 0
agitated off sedation | 0
accidental catheter removal (ACR) | 0
progressively agitated | 2
RASS +3 to +4 | 2
MAP decreased to 50 mmHg | 2
attempts to establish peripheral intravenous access was unsuccessful | 2
intranasal midazolam 10 mg | 2
RASS dropped to one | 10
MAP did not drop further | 10
peripheral intravenous access established | 10
intermittent Phenylephrine boluses | 10
further sedation administered as required | 10
central venous access reestablished | 12
septic shock progressively improved | 24
weaned off the ventilator | 120
extubated | 120