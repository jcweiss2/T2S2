32 years old | 0
male | 0
admitted to the hospital | 0
painful right lower limb swelling | -120
difficulty to walk | -120
generalized weakness | -120
fever | -120
history of hepatitis C | 0
history of intravenous drug abuse | 0
focal tenderness | 0
ecchymosis | 0
marked edema of knee joint | 0
turbid yellowish synovial fluid | 0
cellulitis | 0
septic arthritis of the knee | 0
piperacillin | 0
metronidazole | 0
abnormal vital signs | 0
blood pressure of 98/54 mmHg | 0
heart rate of 123 b/min | 0
respiratory rate of 22/min | 0
oxygen saturation of 92% | 0
temperature of 38.1°C | 0
nonsteroidal anti-inflammatory drugs | 0
white blood cells 11,060/μL | 0
C-reactive protein: 36.8 mg/dL | 0
hematocrit: 40.7% | 0
hemoglobin:14.3 g/dL | 0
platelets of 184,000/μL | 0
D-dimers: 127,5 μg/L | 0
urea: 100 mg/dL | 0
creatinine: 0.81 mg/dL | 0
erythrocyte sedimentation rate: 108 mm/h | 0
Na: 145 mmol/L | 0
K: 4.6 mmol/L | 0
creatine kinase: 1210 IU/L | 0
lactate dehydrogenase: 355 IU/L | 0
cutaneous ecchymosis | 0
necrosis in rectus femoris | 0
necrosis in vastus lateralis | 0
knee arthrotomy | 12
synovectomy | 12
irrigation with 9 L of saline | 12
debridement of all infected soft tissues | 12
fasciotomy | 12
necrosis of the fascia | 12
S. aureus infection | 12
vancomycin | 12
intensive care unit | 12
daily evaluation of the open wound | 12
irrigation | 12
aggressive surgical debridement | 12
foul-smelling necrotic materials | 84
surgical exploration | 84
extensive necrosis of the fascia | 84
popliteal and peroneal artery thrombosed aneurysm | 84
hematoma/thrombus evacuation | 84
stent insertion | 84
reconstructive and plastic surgeries | 240
septic shock | 336
above-the-knee amputation | 336
metabolic and hemodynamic support | 336
discharged | 4176