68 years old | 0
male | 0
admitted to hospital | 0
elective laparoscopy | 0
excisional lymph node biopsy | 0
intra-abdominal lymphadenopathy | 0
enlarged lymph node in the small bowel mesentery | 0
diathermy | 0
placement of Surgicel | 0
uncomplicated post-operative stay | 0
discharged home | 24
histopathology of the lymph node | 24
diffuse large B-cell lymphoma | 24
commenced on rituximab, cyclophosphamide, doxorubicin, vincristine and prednisolone | 24
R-CHOP chemotherapy regiment | 24
good clinical response | 576
abdominal pain | -576
fever | -576
presented to the emergency department | -576
computed tomography scan of the abdomen and pelvis | -576
high-grade mechanical bowel obstruction | -576
transition point in the mid abdomen | -576
mesenteric soft tissue mass | -576
interloop free fluid | -576
mesenteric congestion | -576
gas locules adjacent to the soft tissue mass | -576
mesenteric venous gas | -576
bowel ischemia | -576
diagnostic laparotomy | -552
thick fibrous band | -552
epiploic appendage of the transverse colon | -552
mass at the root of the small bowel mesentery | -552
closed-loop small bowel obstruction | -552
Surgicel used at the site of the previous mesenteric lymph node excisional biopsy | -552
complete adhesiolysis | -552
sepsis | -528
inotropic support | -528
acute renal failure | -528
hemofiltration | -528
ischemic hepatitis | -528
coagulopathy | -528
intensive care | -528
total acute inpatient stay | -504
transferred to subacute care | -504
rehabilitation | -504
discharged home | 0
hematology follow-up | 0