81 years old|0
male|0
hypertension|0
hyperlipidemia|0
remote smoking|0
chronic obstructive pulmonary disease|0
peptic ulcer disease|0
maroon stools|-72
bright red blood per rectum|-72
lightheadedness|-72
daily intake of baby aspirin|0
previous melena episode|0
no recent melena|0
no abdominal pain|0
no nausea|0
no vomiting|0
no fevers|0
no chills|0
orthostatic|0
intravenous fluids|0
emergency colonoscopy|0
3 colonic polyps removed|0
diverticuli as bleeding source|0
re-hospitalized for COPD|1440
massive painless hematochezia|1440
IV steroids|1440
hypovolemic shock|1440
intubation|1440
ICU care|1440
extubation|1440
another massive painless hematochezia|1440
initial bleeding scan negative|1440
large transfusion requirement|1440
stabilized|1440
another episode of massive hematochezia|1440
2nd bleeding scan positive in splenic flexure and sigmoid colon|1440
increased uptake in distal abdominal aorta|1440
increased uptake in right common iliac|1440
radiologically read as physiological blood pooling|1440
angiography negative|1440
active hematochezia|1440
hypotension|1440
received 9 units of blood|1440
differential diagnoses of diverticular bleed|1440
differential diagnoses of peptic ulcer disease|1440
differential diagnoses of arteriovenous malformations|1440
differential diagnoses of severe hemorrhoids|1440
repeat urgent colonoscopy|1440
transverse colon diverticular disease|1440
descending colon diverticular disease|1440
left hemicolectomy|1440
exploratory laparotomy|1440
total abdominal colectomy|1440
excision of AE fistula|1440
previous abdominal aortic aneurysm|1440
aortoenteric fistula secondary to stent|1440
AAA repair 14 years prior|1440
massive lower GI bleed|1440
hematochezia|1440
melena history|1440
right iliac artery aneurysm|1440
one-year follow-up|1440
good health at follow-up|1440
