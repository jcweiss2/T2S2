66 years old | 0
male | 0
white | 0
admitted to the hospital | 0
intense abdominal pain | 0
acute renal failure | 0
urea 178 mg/dL | 0
serum creatinin 7.92 mg/dL | 0
amphotericin B deoxycholate | -24
nasal leishmaniasis | -24
HIV infection | -8760
gastroesophageal reflux disease | -8760
former smoker | -8760
HIV viral load 92,494 copies/ml | 0
CD4 count 5 cells/mm3 | 0
CD4/CD8 ratio 0.08 | 0
pancytopaenic | 0
haemoglobin 6.0 g/dL | 0
leucocytes 1,620 cells/μL | 0
lymphocytes 142 cells/μL | 0
platelets 64,000 cells/μL | 0
afebrile | 0
emaciated | 0
severe nasal lesion | 0
ulcer in the hard palate | 0
extensive necrotic lesion | 0
dysphonic | 0
consolidative lesions in both lungs | 0
small bilateral pleural effusions | 0
haemodialysis | 0
amphotericin B treatment | 0
amphotericin B lipid complex | 3
L-AmB 4 mg/kg/day | 3
acute respiratory distress | 384
pulmonary sepsis by P. aeruginosa | 384
admission to the intensive care unit | 384
melena | 384
severe blood dyscrasia | 384
testicular mass | 384
local swelling | 384
hyperemia | 384
multiseptate fluid collection | 384
diagnostic orchiectomy | 384
swollen testicle | 384
areas of necrosis | 384
fluid accumulation | 384
unfavourable clinical outcome | 600
death | 600
genitourinary histoplasmosis | 648
histology and culture of testicular sample analysis | 648
disseminated histoplasmosis | 648
nasal lesions | -24
mucocutaneous leishmaniasis | -24
nasal biopsy | -24
antigen detection | 0
serology | 0
culture | 0
amastigotes | 0
yeast structures | 0
Giemsa stain | 0
testicular lesion | 384
epididymo-orchitis | 384
histoplasmosis | 384
AIDS | -8760
testicular tuberculosis | 0
granulomatous diseases | 0
differential diagnosis | 0