60 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
fever | -48 | 0 | Factual
abdominal pain | -48 | 0 | Factual
edema of the scrotum | -48 | 0 | Factual
edema of the penis | -48 | 0 | Factual
edema of the perineum | -48 | 0 | Factual
edema of the right gluteal region | -48 | 0 | Factual
hypertension | 0 | 0 | Factual
osteoporosis | 0 | 0 | Factual
hemorrhoids | 0 | 0 | Factual
blood pressure 103/62 mmHg | 0 | 0 | Factual
heart rate 135/min | 0 | 0 | Factual
oxygen saturation 88% | 0 | 0 | Factual
white blood cell count 13.11/μL | 0 | 0 | Factual
C-reactive protein level 61.4 mg/dL | 0 | 0 | Factual
serum creatinine 4.3 mg/dL | 0 | 0 | Factual
blood urea 157 mg/dL | 0 | 0 | Factual
blood sugar 142 mg/dL | 0 | 0 | Factual
procalcitonin 8.53 ng/mL | 0 | 0 | Factual
SARS-CoV-2 infection suspected | 0 | 0 | Possible
RT-PCR test for SARS-CoV-2 | 0 | 0 | Factual
RT-PCR test result negative | 0 | 0 | Factual
CT of the abdomen and pelvis | 0 | 0 | Factual
inflammatory infiltration of the subcutaneous tissues | 0 | 0 | Factual
liquefaction and gas in the subcutaneous tissues | 0 | 0 | Factual
necrosis of scrotum and penis | 0 | 0 | Factual
edema of the subcutaneous tissues | 0 | 0 | Factual
Fournier's gangrene diagnosed | 0 | 0 | Factual
surgery | 0 | 0 | Factual
resection of the necrotic tissues | 0 | 0 | Factual
bilateral orchiectomy | 0 | 0 | Factual
excision of the penile and scrotal skin | 0 | 0 | Factual
antibiotic therapy | 0 | 432 | Factual
meropenem | 0 | 432 | Factual
metronidazole | 0 | 432 | Factual
linezolid | 0 | 432 | Factual
intensive care unit | 0 | 0 | Factual
mechanical ventilation | 0 | 0 | Factual
broad-spectrum antibiotics | 0 | 0 | Factual
supportive and nutritional therapies | 0 | 0 | Factual
colostomy | 0 | 0 | Factual
wound debridement | 0 | 0 | Factual
negative pressure wound therapy | 0 | 0 | Factual
sedation discontinued | 0 | 0 | Factual
extubated | 0 | 0 | Factual
oxygen on low flow | 0 | 0 | Factual
hemodynamically stable | 0 | 0 | Factual
diuresis stimulated | 0 | 0 | Factual
inflammatory markers decreased | 0 | 0 | Factual
culture of the pus material | 0 | 0 | Factual
Escherichia coli | 0 | 0 | Factual
Pseudomonas aeruginosa | 0 | 0 | Factual
antibiotic therapy modified | 0 | 576 | Factual
cephazolin | 0 | 576 | Factual
NPWT discontinued | 0 | 0 | Factual
free-skin grafts | 0 | 0 | Factual
discharged | 1104 | 1104 | Factual
nursing home | 1104 | 0 | Factual
continous nursing care | 1104 | 0 | Factual
free-skin graft care | 1104 | 0 | Factual
regular dressing changes | 1104 | 0 | Factual
physiotherapy | 1104 | 0 | Factual
testosterone supplementation | 1104 | 0 | Factual
colostomy reversal | 0 | 0 | Possible