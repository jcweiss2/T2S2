28 years old | 0
male | 0
white | 0
admitted to the hospital | 0
found unresponsive | -1
EMS performed 12-lead electrocardiogram | -1
ECG interpreted as acute anterior myocardial infarction | -1
brought to a Chest Pain-Accredited facility | 0
arrival to the ED | 0
consciousness was waxing and waning | 0
Kussmaul breathing | 0
hypothermic | 0
hypoxic | 0
required 3 L of supplemental oxygen | 0
blood pressure was 116/42 mmHg | 0
heart rate 90 beats per minute | 0
pupils were equal and reactive to light | 0
oral mucous membranes were dry | 0
heart had regular rate and rhythm | 0
no murmurs | 0
no jugular venous distension | 0
no edema of the lower extremities | 0
radial and dorsal pedal pulses were intact | 0
demonstrated Kussmaul breathing | 0
clear to auscultation bilaterally | 0
abdomen was soft and nontender | 0
skin had multiple tattoos | 0
no rashes or lesions | 0
obtunded | 0
arousable | 0
able to follow commands | 0
initial arterial blood gas showed pH 6.85 | 0
carbon dioxide 14.0 kPa | 0
oxygen 164.0 kPa | 0
bicarbonate 2.3 mmol/L | 0
base excess −29.6 mmol/L | 0
potassium of 9.0 mmol/L | 0
Cardiology was consulted | 0
initial arrival ECG demonstrated an irregular rhythm | 0
rSR’ with down-sloping S-wave and inverted T-waves | 0
Cardiology agreed these findings were likely secondary to hyperkalemia | 0
empiric treatment was started with calcium carbonate and insulin therapy | 0
ED repeat ECG showed improvement | 1
reduction in rSR’ in V1 and V2 | 1
initial laboratory data showed sodium 115 mmol/L | 0
potassium 9.0 mmol/L | 0
chloride 76 mmol/L | 0
blood urea nitrogen 88 mmol/L | 0
creatinine 4.8 mmol/dL | 0
glucose 1375 mmol/L | 0
calcium 7.9 mmol/L | 0
alkaline phosphatase 112 μkat/L | 0
bicarbonate <5.0 mmol/L | 0
alanine aminotransferase 40 μkat/L | 0
aspartate aminotransferase 26 μkat/L | 0
albumin 3.5 g/L | 0
total bilirubin 0.5 μmol/L | 0
osmolality 330 mmol/kg | 0
creatinine phosphokinase 176 units/L | 0
troponin-I 0.596 μg/L | 0
c-reactive protein 0.1 mg/L | 0
glomerular filtration rate (GFR) 15 mL/s | 0
creatinine kinase-MB 5.3 μg/L | 0
myoglobin 551 nmol/L | 0
white blood cell count 29.4×10^9/L | 0
hemoglobin 8.1 g/L | 0
hematocrit 25% | 0
mean corpuscular volume 86.8 fL | 0
platelet count 301×10^9/L | 0
intubated | 0
central venous access and dialysis catheter were placed | 0
covered with a Bair Hugger and multiple heated blankets | 0
intravenous access was started | 0
aggressive volume resuscitation was started | 0
admitted to the Intensive Care Unit (ICU) | 0
diabetic ketoacidosis | 0
hyperosmolar coma | 0
type I diabetes mellitus | 0
non-compliance with insulin therapies | 0
alcohol use | 0
severe dehydration | 0
severe electrolyte and metabolic derangements | 0
acute renal failure | 0
sepsis | 0
type-II myocardial infarction | 0
Nephrology was consulted | 1
life-threatening electrolyte abnormalities | 1
potential need for emergent dialysis | 1
empiric antibiotic therapy with vancomycin and meropenem | 1
Chest radiography confirmed a left lower-lobe aspiration pneumonia | 2
lactic acidosis | 2
cardiac troponin-I level was 0.596 μg/L | 0
subsequent 19.1 μg/L | 12
peaking at 20.452 μg/L | 24
trending downwards | 48
weight-based heparin infusion and antiplatelet therapy | 12
Cardiology consultation concluded that this was likely a representation of a WHO fourth universal definition type-II myocardial infarction | 12
no significant cardiac history | 0
presentation of DKA and profound hypovolemia | 0
sixth day of his hospital course | 120
biochemically and clinically improved | 120
eager for discharge | 120
no documented seizures or agonal nocturnal respirations | 120
medical therapies were optimized | 120
discharged home | 120
atorvastatin 80 mg P.O. QHS | 120
aspirin 81 mg p.o. daily | 120
metoprolol tartrate 12.5 mg p.o. BID | 120
amlodipine 5 mg p.o. daily | 120
Levemir 25 units subcutaneous qam | 120
10 units subcutaneous qpm | 120
nov-Log subcutaneous carb count | 120
Cardiology follow-up | 168
non-ST-elevation myocardial infarction | 168
history of syncope | 168
continued isolated dizzy spells | 168
prior Brugada-like ECG findings | 168
high-risk diabetes | 168
left heart catheterization | 168
selective coronary angiogram | 168
left ventriculo-gram | 168
normal epicardial coronary arteries | 168
ejection fraction of 65% | 168
referred for electrophysiology consultation | 168
no family history suggestive of sudden cardiac death | 0
no proband-positive Brugada syndrome family history | 0