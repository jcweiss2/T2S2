55 years old | 0
male | 0
admitted to the hospital | 0
ingested sodium chlorite | -2
ingested whiskey | -2
ingested ibuprofen | -2
attempted to hang himself | -2
found lying on the floor | -1
cyanotic | -1
lowered consciousness | -1
vomited | -1
transported to the hospital | -1
Glasgow Coma Scale score 13 | 0
body temperature 33.6°C | 0
heart rate 110/min | 0
blood pressure 150/80 mm Hg | 0
respiratory rate 28/min | 0
pulse oximetry 65% | 0
generalized skin cyanosis | 0
neck markings after strangulation | 0
silent abdomen | 0
incontinence for urine and feces | 0
blood samples from the arterial line rendered chocolate-brown serum | 0
depression | 0
previous suicide attempt | 0
alcohol abuse | 0
sedated | 0
intubated | 0
mechanically ventilated | 0
hemoglobin 179 g/L | 0
erythrocytes 5.45 × 10^12/L | 0
hematocrit 0.54 | 0
leukocytes 28.5 × 10^9/L | 0
platelet count 279 × 10^9/L | 0
body urea nitrogen 5.5 mg/dL | 0
creatinine 142 μmol/L | 0
potassium 7.5 mM | 0
osmolality 351 mosm/L | 0
arterial lactate 6.5 mM | 0
myoglobin 433 ng/mL | 0
bilirubin elevated to 28 mM | 0
arterial blood gas analysis | 0
pH 7.25 | 0
PaCO2 4.45 kPa | 0
PaO2 52.45 kPa | 0
BE -12.2 mmol/L | 0
HCO3 14.1 mmol/L | 0
SaO2 99% | 0
lactate 6.48 mmol/L | 0
methemoglobinemia 40.1% | 0
methylene blue administration | 2
continuous venovenous hemodiafiltration | 4.5
anuria | 4.5
hyperkalemia | 4.5
metabolic acidosis | 4.5
hemodialysis | 8.5
lactate level dropped to 2.55 mmol/L | 14
methemoglobinemia decreased to 15.2% | 14
methemoglobinemia decreased to 10.2% | 29
hemolytic anemia | 24
disseminated intravascular coagulation | 24
norepinephrine drip | 20
hypotension | 20
bronchopneumonia | 192
sepsis | 192
gastric and esophageal ulceration improved | 240
weaned from mechanical ventilation | 312
intermittent hemodialysis | 408
urine output 2500 mL/24 h | 528
blood urea 12 mg/dL | 528
creatinine 428 μmol/L | 528
estimated GFR 15.6 mL/min | 528
transferred to a medium care facility | 528
transferred to a psychiatric ward | 1008
discharged from hospital | 1536