82 years old | 0
female | 0
admitted to emergency department | 0
cognitive regression | -168
deterioration | -168
decreased oral intake | -168
fever | -168
hypertension | -6720
chronic atrial fibrillation | -6720
bilateral salpingo-oophorectomy | -6720
total abdominal hysterectomy | -6720
clavicle fracture | -2880
bed-dependent state | -1092
GCS was 8 | 0
SaO2 was 92–95% | 0
ABP was 90/60 mmHg | 0
pulse was 120–136 bpm | 0
respiratory rate was 25–35/min | 0
ED transthoracic echocardiogram | 0
contrast-enhanced thoracoabdominal computed tomography | 0
intubated | 0
vasopressor support | 0
transferred to ICU | 0
perianal abscess | 0
perianal fistula | 0
abscess drained | 0
sedation with dexmedetomidine/propofol | 0
analgesia with fentanyl/morphine | 0
ventilatory weaning | 0
tracheostomy | 672
short thyromental distance | 672
short neck | 672
limited neck extension | 672
open surgical tracheostomy | 672
enteral feeding solution remnants in tracheostomy aspirations | 48
pulsative air filling in nasogastric drainage bag | 48
bedside bronchoscopy | 48
trachea and esophagus joined | 48
contrast-enhanced cervical and thorax CT | 48
mini laparotomy | 72
tube jejunostomy | 72
Sengstaken–Blakemore tube insertion | 96
gastric balloon inflated | 96
esophagus balloon inflated | 96
SBt placement | 96
patient adaptation to mechanical ventilation improved | 96
air leak into GIS prevented | 96
reflux of GIS content into tracheobronchial tree prevented | 96
discharged | unknown