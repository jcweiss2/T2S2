65 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
recurrent fever | -744 | 0 | Factual
nausea | -168 | 0 | Factual
vomiting | -168 | 0 | Factual
highest body temperature 38 ℃ | -744 | 0 | Factual
neutrophil count 6.96×10^9/L ↑ | 0 | 0 | Factual
monocyte count 0.86×10^9/L ↑ | 0 | 0 | Factual
lymphocyte percentage 14.9% ↓ | 0 | 0 | Factual
red blood cell count 3.17×10^12/L ↓ | 0 | 0 | Factual
hemoglobin content 87 g/L ↓ | 0 | 0 | Factual
hematocrit 0.28 L/L ↓ | 0 | 0 | Factual
average red blood cell hemoglobin concentration 312 g/L ↓ | 0 | 0 | Factual
platelet count 363×10^9/L ↑ | 0 | 0 | Factual
platelet distribution width 8.3 fl ↓ | 0 | 0 | Factual
C-reactive protein (CRP) 52.01 mg/L ↑ | 0 | 0 | Factual
Klebsiella pneumoniae sepsis | -744 | 0 | Factual
secondary infectious thrombocytopenia | 0 | 0 | Factual
liver abscess | 0 | 0 | Factual
bilateral lung inflammation | 0 | 0 | Factual
type 2 diabetes | 0 | 0 | Factual
hypertension grade 3 | 0 | 0 | Factual
vancomycin | 0 | 24 | Factual
caspofungin | 0 | 24 | Factual
dexamethasone | 0 | 24 | Factual
posaconazole oral suspension | 0 | 24 | Factual
liver abscess puncture and drainage | 24 | 24 | Factual
endogenous endophthalmitis (left) | 48 | 48 | Factual
orbital cellulitis (left) | 48 | 48 | Factual
rubeosis iridis (left) | 48 | 48 | Factual
exudative retinal detachment (left) | 48 | 48 | Factual
diabetic retinopathy (right) | 48 | 48 | Factual
intravitreal injection with vancomycin and ceftazidime | 48 | 72 | Factual
left eyeball enucleation | 168 | 168 | Factual
moxifloxacin | 168 | 192 | Factual
sulperazon | 168 | 192 | Factual
fever again | 192 | 192 | Factual
computed tomography (CT) examination | 216 | 216 | Factual
inflammation of both lungs | 216 | 216 | Factual
pericardial effusion | 216 | 216 | Factual
bilateral pleural thickening and effusion | 216 | 216 | Factual
atelectasis in right inferior lobe | 216 | 216 | Factual
liver cyst | 216 | 216 | Factual
liver abscess | 216 | 216 | Factual
right renal cyst | 216 | 216 | Factual
myoma of the uterus | 216 | 216 | Factual
convulsion with unconsciousness | 360 | 360 | Factual
transferred to the respiratory intensive care unit | 360 | 360 | Factual
lacunar infarction | 360 | 360 | Factual
encephalomalacia | 360 | 360 | Factual
bilateral pleural effusion | 360 | 360 | Factual
lower lobe of the right lung insufficiently inflated | 360 | 360 | Factual
intracranial infection | 360 | 360 | Factual
lumbar puncture | 360 | 360 | Factual
cerebrospinal fluid (CSF) analysis | 360 | 360 | Factual
microbial metagenomic next-generation sequencing (mNGS) | 360 | 360 | Factual
Klebsiella pneumoniae with drug-resistant gene blaSHV | 360 | 360 | Factual
meropenem | 360 | 720 | Factual
body temperature improved | 360 | 720 | Factual
blood routine improved | 360 | 720 | Factual
CRP improved | 360 | 720 | Factual
CT examination | 720 | 720 | Factual
pulmonary edema and pleural effusion dissipated | 720 | 720 | Factual
CSF analysis | 720 | 720 | Factual
discharged from the hospital | 744 | 744 | Factual