48 years old | 0
male | 0
mason | 0
admitted to the hospital | 0
fever | -72
cough | -72
breathlessness | -72
type 2 diabetes mellitus | -8760
poor glycemic control | -8760
body temperature 39.7°C | 0
respiratory rate 28 breaths/min | 0
heart rate 128 bpm | 0
blood pressure 100/60 mm Hg | 0
mucopurulent sputum | 0
decreased breath sounds on the left lung base | 0
no bilateral crackles | 0
total leukocyte count 15.9 G/L | 0
Neutrophil predominance | 0
platelet 78 G/L | 0
C-reactive protein (CRP) 324.6 mg/l | 0
hemoglobin A1c (HbA1c) 9.09% | 0
small pleural effusion | 0
consolidated lung base | 0
Ziehl-Neelsen stain negative | 0
sputum culture | 0
blood culture | 0
pleural fluid culture | 0
Gram-negative bacilli | 0
abundant white blood cells | 0
turbidity in blood culture bottle | 96
smooth white non-hemolytic colonies | 96
non-fermenting colonies | 96
catalase-positive | 96
oxidase-positive | 96
identified as Aeromonas salmonicida | 96
treated with cefoperazone-sulbactam | 0
treated with azithromycin | 0
treated with gentamicin | 0
antibiotics changed to piperacillin-tazobactam | 96
antibiotics changed to fosfomycin | 96
antibiotics changed to meropenem | 96
antibiotics changed to ciprofloxacin | 96
high fever | 24
tachypnea | 24
thick mucopurulent sputum | 24
16S rRNA gene sequencing | 120
identified as B. pseudomallei | 120
immunochromatographic assay positive | 120
sensitive to amoxicillin/clavulanic acid | 120
sensitive to ceftazidime | 120
sensitive to meropenem | 120
sensitive to sulfamethoxazole/trimethoprim | 120
sensitive to piperacillin/tazobactam | 120
transferred to Hue Central hospital | 168