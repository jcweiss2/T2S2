68 years old | 0
    woman | 0
    presented with dyspnea | -72
    presented with wheezing | -72
    presented with productive cough | -72
    albuterol use at home | -72
    completed corticosteroid regimen | -168
    weight gain of 30 pounds | -168
    COPD exacerbations history | -87600
    treated with antibiotics | -87600
    treated with beta 2 agonists | -87600
    treated with long-acting muscarinic antagonist | -87600
    treated with systemic corticosteroids | -87600
    last hospitalization | -5760
    no intubation history | 0
    no stridor history | 0
    no reflux symptoms history | 0
    mMRC symptom score 3 | 0
    150 pack-year smoking history | 0
    quit smoking 1 month prior | -720
    sleeps in seated position | 0
    dyspnea when lying flat | 0
    chairbound due to dyspnea | 0
    hypertension | 0
    depression | 0
    obstructive sleep apnea | 0
    end-stage renal disease | 0
    hemodialysis | 0
    medications: fluticasone/salmeterol | 0
    medications: tiotropium | 0
    medications: albuterol as needed | 0
    medications: prednisone | 0
    medications: 3L oxygen by nasal cannula | 0
    medications: CPAP at night | 0
    medications: simvastatin | 0
    medications: diltiazem SR | 0
    medications: sertraline | 0
    completed pulmonary rehabilitation 2 years prior | -17520
    physical exam: alert | 0
    physical exam: moderate respiratory distress | 0
    temperature 98.6 F | 0
    blood pressure 150/72 | 0
    pulse rate 90/min | 0
    respiratory rate 26/min | 0
    BMI 36 kg/m² | 0
    oxygen saturation 96% on 6L/min oxygen | 0
    Cushingoid facies | 0
    centripetal obesity | 0
    rapid regular cardiac rhythm | 0
    no cardiac murmur | 0
    bilateral expiratory wheezing | 0
    no pedal edema | 0
    chest radiograph no infiltrates | 0
    chest radiograph no congestion | 0
    sinus tachycardia on ECG | 0
    non-specific ST changes on ECG | 0
    hemoglobin 11 g/dL | 0
    glucose 147 mg/dL | 0
    potassium 4.7 mEq/L | 0
    creatinine 9.1 mg/dL |!0
    admitted with COPD exacerbation | 0
    received intravenous glucocorticoids | 0
    received albuterol nebulizer treatments | 0
    received BiPAP | 0
    received broad-spectrum antibiotics | 0
    continued hemodialysis | 0
    improved oxygenation | 24
    improved symptoms | 24
    PFT FEV1/FVC 62% | 0
    PFT FEV1 41% predicted | 0
    GOLD 3 classification | 0
    alternative diagnosis pursued | 24
    transthoracic echocardiogram LVEF 70% | 24
    normal RV function | 24
    Grade 1 diastolic dysfunction | 24
    normal valves | 24
    negative thrombophilia workup | 24
    CT neck unremarkable | 24
    dynamic expiratory CT: emphysema | 24
    dynamic expiratory CT: 11mm pulmonary nodule | 24
    dynamic expiratory CT: tracheobronchial collapse | 24
    dynamic expiratory CT: bronchus intermedius collapse | 24
    TM diagnosis | 24
    declined lung biopsy | 24
    agreed on silicone stent | 24
    bronchoscopy performed | 24
    Y stent placed | 24
    discharged next day | 24
    arterial blood gases pH 7.35 | 24
    pCO2 47 | 24
    PO2 85 | 24
    oxygen 3L/min on discharge | 24
    good inhaler technique | 24
    found hypotensive | 48
    found unresponsive | 48
    acute hypoxic respiratory failure | 48
    admitted to ICU | 48
    endotracheal intubation | 48
    intravenous vasopressors | 48
    systemic corticosteroids | 48
    broad-spectrum antibiotics | 48
    nebulized bronchodilators | 48
    mucolytic agents | 48
    chest radiograph no infiltrates | 48
    chest radiograph no edema | 48
    chest radiograph no pneumothorax | 48
    normal stent position | 48
    sepsis ruled out | 48
    myocardial ischemia ruled out | 48
    COPD exacerbation improved | 48
    placed on home hospice | 72
    discharged | 72