63 years old | 0
    man | 0
    admitted to his local general hospital | 0
    feeling unwell for a fortnight | -336
    blood culture confirmed the presence of vancomycin resistant enterococcal (VRE) | 0
    transthoracic esophageal echocardiogram confirmed dehiscence of the aortic valve | 0
    aortic valve replacement for aortic stenosis | -2880
    aortic root abscess | 0
    mitral valve vegetations | 0
    patent foramen ovale (PFO) | 0
    inferior vena cava Eustachian valve | 0
    transfer to our institution | 0
    liver failure | 0
    renal failure | 0
    bilirubin 54 mg/dL | 0
    alkaline phosphatase 222 IU/L | 0
    alanine aminotransferase 1211 IU/L | 0
    continuous veno-venous hemofiltration (CVVHF) | 0
    heparin as the anticoagulant | 0
    initial blood tests revealed a platelet count of 179 × 10³ per mm³ | 0
    significant drop in platelet count to 35 × 10³ per mm³ | 72
    heparin induced thrombocytopenia (HIT) | 72
    enzyme-linked immunosorbent assay serotonin release assay | 72
    heparin stopped | 72
    Danaparoid as hemofiltration anticoagulation | 72
    platelet counts dropped to 16 × 10³ per mm³ | 168
    off heparin for over a week | 168
    redo-aortic valve replacement | 0
    mitral valve repair | 0
    closure of the PFO | 0
    repair of the aortic root abscess | 0
    excision of the Eustachian valve | 0
    ventilator dependence | 0
    tracheostomy | 0
    renal failure needing renal replacement therapy | 0
    cardiovascular support for 22 days | 528
    milrinone 10 ml/h | 528
    noradrenaline 20 ml/h | 528
    vasopressin 2 IU/h | 528
    appropriate weaning | 4320
    discharged | 4320
    SDF device used to examine sub-lingual microvasculature | 48
    sepsis signs | 48
    pyrexia | 48
    low systemic vascular resistance | 48
    increased inflammatory markers | 48
    increased inotropic-vasoconstrictor support | 48
    HIT present | 48
    sepsis well-controlled | 1128
    platelet count recovered | 1128
    SDF data not recorded between 90 h and 47 days | 90
    clinically stable | 90
    CI: 3.7 L/min/m² | 48
    MAP: 66 mmHg | 48
    SVRI: 1038 dynes×s/cm⁵/m² | 48
    pH: 7.42 | 48
    lactate: 4.9 mmol/L | 48
    NA: 0.3 mcg/kg/min | 48
    VA: 1 IU/h | 48
    CI: 2.9 L/min/m² | 60
    MAP: 55 mmHg | 60
    SVRI: 1178 dynes×s/cm⁵/m² | 60
    pH: 7.36 | 60
    lactate: 6.9 mmol/L | 60
    NA: 0.2 mcg/kg/min | 60
    VA: 1 IU/h | 60
    CI: 2.8 L/min/m² | 90
    MAP: 74 mmHg | 90
    SVRI: 1885 dynes×s/cm⁵/m² | 90
    pH: 7.2 | 90
    lactate: 6.6 mmol/L | 90
    NA: 0.26 mcg/kg/min | 90
    VA: 4 IU/h | 90
    CI: 2.8 L/min/m² | 1128
    MAP: 52 mmHg | 1128
    SVRI: 1715 dynes×s/cm⁵/m² | 1128
    pH: 7.45 | 1128
    lactate: 1.1 mmol/L | 1128
    NA: 0.06 mcg/kg/min | 1128
    VA: None | 1128
    
    63 years old | 0
    man | 0
    admitted to his local general hospital | 0
    feeling unwell for a fortnight | -336
    blood culture confirmed the presence of vancomycin resistant enterococcal (VRE) | 0
    transthoracic esophageal echocardiogram confirmed dehiscence of the aortic valve | 0
    aortic valve replacement for aortic stenosis | -2880
    aortic root abscess | 0
    mitral valve vegetations | 0
    patent foramen ovale (PFO) | 0
    inferior vena cava Eustachian valve | 0
    transfer to our institution | 0
    liver failure | 0
    renal failure | 0
    bilirubin 54 mg/dL | 0
    alkaline phosphatase 222 IU/L | 0
    alanine aminotransferase 1211 IU/L | 0
    continuous veno-venous hemofiltration (CVVHF) | 0
    heparin as the anticoagulant | 0
    initial blood tests revealed a platelet count of 179 × 10³ per mm³ | 0
    significant drop in platelet count to 35 × 10³ per mm³ | 72
    heparin induced thrombocytopenia (HIT) | 72
    enzyme-linked immunosorbent assay serotonin release assay | 72
    heparin stopped | 72
    Danaparoid as hemofiltration anticoagulation | 72
    platelet counts dropped to 16 × 10³ per mm³ | 168
    off heparin for over a week | 168
    redo-aortic valve replacement | 0
    mitral valve repair | 0
    closure of the PFO | 0
    repair of the aortic root abscess | 0
    excision of the Eustachian valve | 0
    ventilator dependence | 0
    tracheostomy | 0
    renal failure needing renal replacement therapy | 0
    cardiovascular support for 22 days | 528
    milrinone 10 ml/h | 528
    noradrenaline 20 ml/h | 528
    vasopressin 2 IU/h | 528
    appropriate weaning | 4320
    discharged | 4320
    SDF device used to examine sub-lingual microvasculature | 48
    sepsis signs | 48
    pyrexia | 48
    low systemic vascular resistance | 48
    increased inflammatory markers | 48
    increased inotropic-vasoconstrictor support | 48
    HIT present | 48
    sepsis well-controlled | 1128
    platelet count recovered | 1128
    SDF data not recorded between 90 h and 47 days | 90
    clinically stable | 90
    CI: 3.7 L/min/m² | 48
    MAP: 66 mmHg | 48
    SVRI: 1038 dynes×s/cm⁵/m² | 48
    pH: 7.42 | 48
    lactate: 4.9 mmol/L | 48
    NA: 0.3 mcg/kg/min | 48
    VA: 1 IU/h | 48
    CI: 2.9 L/min/m² | 60
    MAP: 55 mmHg | 60
    SVRI: 1178 dynes×s/cm⁵/m² | 60
    pH: 7.36 | 60
    lactate: 6.9 mmol/L | 60
    NA: 0.2 mcg/kg/min | 60
    VA: 1 IU/h | 60
    CI: 2.8 L/min/m² | 90
    MAP: 74 mmHg | 90
    SVRI: 1885 dynes×s/cm⁵/m² | 90
    pH: 7.2 | 90
    lactate: 6.6 mmol/L | 90
    NA: 0.26 mcg/kg/min | 90
    VA: 4 IU/h | 90
    CI: 2.8 L/min/m² | 1128
    MAP: 52 mmHg | 1128
    SVRI: 1715 dynes×s/cm⁵/m² | 1128
    pH: 7.45 | 1128
    lactate: 1.1 mmol/L | 1128
    NA: 0.06 mcg/kg/min | 1128
    VA: None | 1128

    63 years old | 0
    man | 0
    admitted to his local general hospital | 0
    feeling unwell for a fortnight | -336
    blood culture confirmed the presence of vancomycin resistant enterococcal (VRE) | 0
    transthoracic esophageal echocardiogram confirmed dehiscence of the aortic valve | 0
    aortic valve replacement for aortic stenosis | -2880
    aortic root abscess | 0
    mitral valve vegetations | 0
    patent foramen ovale (PFO) | 0
    inferior vena cava Eustachian valve | 0
    transfer to our institution | 0
    liver failure | 0
    renal failure | 0
    bilirubin 54 mg/dL | 0
    alkaline phosphatase 222 IU/L | 0
    alanine aminotransferase 1211 IU/L | 0
    continuous veno-venous hemofiltration (CVVHF) | 0
    heparin as the anticoagulant | 0
    initial blood tests revealed a platelet count of 179 × 10³ per mm³ | 0
    significant drop in platelet count to 35 × 10³ per mm³ | 72
    heparin induced thrombocytopenia (HIT) | 72
    enzyme-linked immunosorbent assay serotonin release assay | 72
    heparin stopped | 72
    Danaparoid as hemofiltration anticoagulation | 72
    platelet counts dropped to 16 × 10³ per mm³ | 168
    off heparin for over a week | 168
    redo-aortic valve replacement | 0
    mitral valve repair | 0
    closure of the PFO | 0
    repair of the aortic root abscess | 0
    excision of the Eustachian valve | 0
    ventilator dependence | 0
    tracheostomy | 0
    renal failure needing renal replacement therapy | 0
    cardiovascular support for 22 days | 528
    milrinone 10 ml/h | 528
    noradrenaline 20 ml/h | 528
    vasopressin 2 IU/h | 528
    appropriate weaning | 4320
    discharged | 4320
    SDF device used to examine sub-lingual microvasculature | 48
    sepsis signs | 48
    pyrexia | 48
    low systemic vascular resistance | 48
    increased inflammatory markers | 48
    increased inotropic-vasoconstrictor support | 48
    HIT present | 48
    sepsis well-controlled | 1128
    platelet count recovered | 1128
    SDF data not recorded between 90 h and 47 days | 90
    clinically stable | 90
    CI: 3.7 L/min/m² | 48
    MAP: 66 mmHg | 48
    SVRI: 1038 dynes×s/cm⁵/m² | 48
    pH: 7.42 | 48
    lactate: 4.9 mmol/L | 48
    NA: 0.3 mcg/kg/min | 48
    VA: 1 IU/h | 48
    CI: 2.9 L/min/m² | 60
    MAP: 55 mmHg | 60
    SVRI: 1178 dynes×s/cm⁵/m² | 60
    pH: 7.36 | 60
    lactate: 6.9 mmol/L | 60
    NA: 0.2 mcg/kg/min | 60
    VA: 1 IU/h | 60
    CI: 2.8 L/min/m² | 90
    MAP: 74 mmHg | 90
    SVRI: 1885 dynes×s/cm⁵/m² | 90
    pH: 7.2 | 90
    lactate: 6.6 mmol/L | 90
    NA: 0.26 mcg/kg/min | 90
    VA: 4 IU/h | 90
    CI: 2.8 L/min/m² | 1128
    MAP: 52 mmHg | 1128
    SVRI: 1715 dynes×s/cm⁵/m² | 1128
    pH: 7.45 | 1128
    lactate: 1.1 mmol/L | 1128
    NA: 0.06 mcg/kg/min | 1128
    VA: None | 1128