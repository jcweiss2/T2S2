38-week gestational age | 0
    female | 0
    3.2 kg birth weight | 0
    born via cesarean section for breech presentation | 0
    respiratory distress | -216
    tachypnea | -216
    fever | -216
    feeding refusal | -216
    admitted to peripheral hospital neonatal ICU | -192
    pneumonia | -192
    septicemia | -192
    left lung consolidation | -192
    right lung cysts | -192
    oxygen therapy | -192
    intravenous antibiotics | -192
    chest X-ray on day 7 of admission | -168
    aggravating cystic lesions in right lung | -168
    referred to our hospital | -72
    admitted to our neonatal ICU | 0
    mild respiratory distress | 0
    family members COVID-19-positive | -672
    nasopharyngeal swab for SARS-CoV-2 RNA | 0
    SARS-CoV-2 PCR positive | 24
    tachypnea | 0
    respiratory rate 72 breaths/min | 0
    subcostal retractions | 0
    intercostal retractions | 0
    absent breath sounds on right chest | 0
    heart sounds better audible on right side | 0
    normal white blood cell count | 0
    Hb 13 gm/dL | 0
    blood gas pH 7.25 | 0
    pO2 55 | 0
    bicarbonate 18 | 0
    base deficit 4 | 0
    pCO2 55 | 0
    O2 saturation 90-95% | 0
    chest X-ray | 0
    chest tomography | 0
    left lung opacities | 0
    left lung consolidation | 0
    right cystic lesions | 0
    chest CT suggested CPAM | 0
    echocardiogram normal | 0
    blood culture sterile | 0
    multidisciplinary team discussion | 0
    decision to monitor closely | 0
    surgical resection indication if no improvement | 0
    respiratory distress treatment with oxygen | 0
    FiO2 50% | 0
    intravenous antibiotics | 0
    clinical improvement after 7 days | 168
    off oxygen | 168
    respiratory distress signs disappeared | 168
    normal feeding resumed | 168
    discharged | 168
    out-patient follow-up after 8 weeks | 168
    control chest CT after 8 weeks | 168
    complete resolution of cystic lesions | 168
    post-pneumonia healing changes | 168
    
    <|eot_id|>
    38-week gestational age | 0
    female | 0
    3.2 kg birth weight | 0
    born via cesarean section for breech presentation | 0
    respiratory distress | -216
    tachypnea | -216
    fever | -216
    feeding refusal | -216
    admitted to peripheral hospital neonatal ICU | -192
    pneumonia | -192
    septicemia | -192
    left lung consolidation | -192
    right lung cysts | -192
    oxygen therapy | -192
    intravenous antibiotics | -192
    chest X-ray on day 7 of admission | -168
    aggravating cystic lesions in right lung | -168
    referred to our hospital | -72
    admitted to our neonatal ICU | 0
    mild respiratory distress | 0
    family members COVID-19-positive | -672
    nasopharyngeal swab for SARS-CoV-2 RNA | 0
    SARS-CoV-2 PCR positive | 24
    tachypnea | 0
    respiratory rate 72 breaths/min | 0
    subcostal retractions | 0
    intercostal retractions | 0
    absent breath sounds on right chest | 0
    heart sounds better audible on right side | 0
    normal white blood cell count | 0
    Hb 13 gm/dL | 0
    blood gas pH 7.25 | 0
    pO2 55 | 0
    bicarbonate 18 | 0
    base deficit 4 | 0
    pCO2 55 | 0
    O2 saturation 90-95% | 0
    chest X-ray | 0
    chest tomography | 0
    left lung opacities | 0
    left lung consolidation | 0
    right cystic lesions | 0
    chest CT suggested CPAM | 0
    echocardiogram normal | 0
    blood culture sterile | 0
    multidisciplinary team discussion | 0
    decision to monitor closely | 0
    surgical resection indication if no improvement | 0
    respiratory distress treatment with oxygen | 0
    FiO2 50% | 0
    intravenous antibiotics | 0
    clinical improvement after 7 days | 168
    off oxygen | 168
    respiratory distress signs disappeared | 168
    normal feeding resumed | 168
    discharged | 168
    out-patient follow-up after 8 weeks | 168
    control chest CT after 8 weeks | 168
    complete resolution of cystic lesions | 168
    post-pneumonia healing changes | 168