9 years old | 0
    male | 0
    admitted to the hospital | 0
    painful skin eruption | -720
    skin eruption started on the abdomen | -720
    skin eruption progressed to cover almost the entire body | -720
    fever (39°C) | -720
    generalized malaise | -720
    erythematous macules | 0
    papules | 0
    necrotic plaques | 0
    hemorrhagic crusts | 0
    flexural accentuation of the lesions in the axillae | 0
    flexural accentuation of the lesions in the groin | 0
    flexural accentuation of the lesions in the neck | 0
    oral mucosa involvement | 0
    small painful ulcers on the tongue | 0
    small painful ulcers on the inner lip | 0
    mild leukocytosis | 0
    elevated erythrocyte sedimentation rate | 0
    elevated C-reactive protein | 0
    anemia | 0
    skin biopsy from necrotic plaque | 0
    focal full-thickness epidermal necrosis | 0
    exocytosis | 0
    vacuolar interface dermatitis | 0
    superficial perivascular lymphocytic infiltrate | 0
    deep perivascular lymphocytic infiltrate | 0
    focal hemorrhage | 0
    diagnosis of FUMHD | 0
    systemic antibiotics (azithromycin, 250 mg/d) | 0
    systemic steroids (30 mg/d) | 0
    left the hospital | 240
    returned to the hospital | 720
    treated with intravenous immunoglobulins (IVIG) | 720
    treated with cyclosporine | 720
    worsening skin lesions | 720
    impaired renal function | 720
    ulceronecrotic papules increased in number and size | 720
    ulceronecrotic plaques increased in number and size | 720
    ulceronecrotic papules became confluent | 720
    ulceronecrotic plaques became confluent | 720
    ulcerative lesions secondarily infected with Pseudomonas aeruginosa | 720
    Pseudomonas aeruginosa cultured from the skin | 720
    Pseudomonas aeruginosa cultured from the blood | 720
    development of gangrenous ulcers | 720
    central black eschars | 720
    erythematous borders | 720
    ecthyma gangrenosum | 720
    transferred to the intensive care unit | 720
    systemic vancomycin | 720
    systemic gentamycin | 720
    deterioration | 720
    tachypnea | 720
    tachycardia | 720
    hypothermia | 720
    systemic inflammatory response syndrome | 720
    supportive measures | 720
    intravenous fluids | 720
    refractory hypotension | 720
    myocardial dysfunction | 720
    generalized edema | 720
    fulminant sepsis | 720
    multiple organ failure | 720
    death | 720
    
    
    9 years old | 0
    male | 0
    admitted to the hospital | 0
    painful skin eruption | -720
    skin eruption started on the abdomen | -720
    skin eruption progressed to cover almost the entire body | -720
    fever (39°C) | -720
    generalized malaise | -720
    erythematous macules | 0
    papules |Cozzio et al, 200410 72 Male Monoclonal T cell MI: NegativeSI: Sepsis, pancytopenia MTX, IVIG Cozzio et al, 200410 26 Female Monoclonal T cell MI: NegativeSI: Sepsis, pancytopenia SS, MTX, PUVA Aytekin et al, 200511 27 Female Unknown MI: NegativeSI: Sepsis SS, ATB, IVIG, acyclovir Malnar et al, 200612 60 Male Unknown MI: PositiveSI: Sepsis, pulmonary thromboembolism, thrombosis of superior mesenteric artery SS, ATB ABS, Antibiotics; DDS, diamino-diphenyl sulphone; MI, mucosal involvement; MTX, methotrexate; SI, systemic involvement; SS, systemic steroids.∗ Fever and severe generalized, progressive ulceronecrotic papules and plaques were constant clinical features in all patients.Adapted from Nofal A, Assaf M, Alakad R, Amer H, Nofal E, Yosef A. Febrile ulceronecrotic Mucha-Habermann disease: proposed diagnostic criteria and therapeutic evaluation. Int J Dermatol. http://dx.doi.org/10.1111/ijd.13195. Published online December 23, 2015.
    <|eot_id|><|start_header_id|>assistant<|end_header_id|>
    9 years old | 0
    male | 0
    admitted to the hospital | 0
    painful skin eruption | -720
    skin eruption started on the abdomen | -720
    skin eruption progressed to cover almost the entire body | -720
    fever (39°C) | -720
    generalized malaise | -720
    erythematous macules | 0
    papules | 0
    necrotic plaques | 0
    hemorrhagic crusts | 0
    flexural accentuation of the lesions in the axillae | 0
    flexural accentuation of the lesions in the groin | 0
    flexural accentuation of the lesions in the neck | 0
    oral mucosa involvement | 0
    small painful ulcers on the tongue | 0
    small painful ulcers on the inner lip | 0
    mild leukocytosis | 0
    elevated erythrocyte sedimentation rate | 0
    elevated C-reactive protein | 0
    anemia | 0
    skin biopsy from necrotic plaque | 0
    focal full-thickness epidermal necrosis | 0
    exocytosis | 0
    vacuolar interface dermatitis | 0
    superficial perivascular lymphocytic infiltrate | 0
    deep perivascular lymphocytic infiltrate | 0
    focal hemorrhage | 0
    diagnosis of FUMHD | 0
    systemic antibiotics (azithromycin, 250 mg/d) | 0
    systemic steroids (30 mg/d) | 0
    left the hospital | 240
    returned to the hospital | 720
    treated with intravenous immunoglobulins (IVIG) | 720
    treated with cyclosporine | 720
    worsening skin lesions | 720
    impaired renal function | 720
    ulceronecrotic papules increased in number and size | 720
    ulceronecrotic plaques increased in number and size | 720
    ulceronecrotic papules became confluent | 720
    ulceronecrotic plaques became confluent | 720
    ulcerative lesions secondarily infected with Pseudomonas aeruginosa | 720
    Pseudomonas aeruginosa cultured from the skin | 720
    Pseudomonas aeruginosa cultured from the blood | 720
    development of gangrenous ulcers | 720
    central black eschars | 720
    erythematous borders | 720
    ecthyma gangrenosum | 720
    transferred to the intensive care unit | 720
    systemic vancomycin | 720
    systemic gentamycin | 720
    deterioration | 720
    tachypnea | 720
    tachycardia | 720
    hypothermia | 720
    systemic inflammatory response syndrome | 720
    supportive measures | 720
    intravenous fluids | 720
    refractory hypotension | 720
    myocardial dysfunction | 720
    generalized edema | 720
    fulminant sepsis | 720
    multiple organ failure | 720
    death | 720
    