76 years old | 0
male | 0
admitted to the hospital | 0
bladder cancer | -672
regional lymph node involvement | -672
Clostridium difficile infection (CDI) | -672
vomiting | -72
watery diarrhea | -72
anorexia | -72
mild odynophagia | -72
oral vancomycin | -72
acute renal dysfunction | 0
lactic acidosis | 0
leukocytosis with bandemia | 0
basilar atelectasis | 0
diffuse colonic wall-thickening | 0
peri-colonic fat-stranding | 0
normal saline | 0
lactated ringers | 0
norepinephrine | 0
broad-spectrum intravenous antibiotics | 0
septic shock | 0
mental status excellent | 4
urine output in excess of 0.5 mL/kg/hr | 4
resolving lactic acidosis | 4
unexplained back pain | 6
worsening shock | 6
multi-organ failure | 6
emergent endotracheal intubation | 6
orogastric tube placement | 6
bilateral hydropneumothorax | 6
pneumomediastinum | 6
placement of bilateral chest tubes | 6
dark fluid from each pleural space | 6
esophageal perforation suspected | 6
pleural fluid analysis | 6
elevated amylase level | 6
Gram stain revealed Gram-positive cocci and rods | 6
pleural cultures grew multiple species of aerobic Gram-positive organisms | 6
mixed refractory acidemia | 12
continuous veno-venous hemodiafiltration | 12
mechanical ventilation | 12
vasopressor support | 12
CT of the chest | 24
esophageal perforation confirmed | 24
locules of air communicating from the pleural spaces to the distal esophagus | 24
orogastric tube penetrating across the perforation into the lesser sac of the stomach | 24
endoscopic intervention | 72
extensive esophageal necrosis | 72
complete separation of the lower esophagus from the stomach | 72
unsutured fully-covered self-expanding metal stent deployed | 72
parental nutrition | 72
chest tubes maintained | 72
vasopressors titrated off | 168
dialysis discontinued | 168
extubated | 168
mediastinitis | 216
recurrent respiratory failure | 216
comfort-focused approach | 216
passed away | 216