73 years old | 0
male | 0
inoperable adenocarcinoma of the right lung | -8760
concurrent chemoradiotherapy | -8760
Salmonella Group D necrotising pneumonia | -8760
extra-thoracic extension | -8760
empyema necessitans | -8760
haemoptysis | 0
purulent discharge | 0
invasive pulmonary aspergillosis | 0
voriconazole | 0
acetaminophen | 0
cefoperazone-sulbactam | 0
metronidazole | 0
vancomycin | 0
piperacillin-tazobactam | 0
meropenem | 0
acidotic breathing | 960
severe metabolic acidosis | 960
raised anion gap | 960
no lactic acidosis | 960
normal serum osmolal gap | 960
no exposure to salicylate | 960
no exposure to toxic alcohols | 960
no exposure to glycols | 960
elevated creatinine | 960
elevated beta-hydroxybutyrate | 960
elevated urine anion gap | 960
discontinuation of acetaminophen | 960
N-acetylcysteine infusion | 960
transfer to intensive care unit | 960
improvement of acid-base imbalance | 1008
discharge from ICU | 1032
massive haemoptysis | 1464
death | 1464
pyroglutamic acidosis | 960
chronic acetaminophen ingestion | -960
glutathione depletion | -960
cysteine depletion | -960
renal impairment | -960
voriconazole treatment | 0