Mayer-Rokitansky-Küster-Hauser syndrome | 0 | 0 | Factual
27 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
sigmoid neovaginoplasty | -7560 | -7560 | Factual
lower abdominal pain | -336 | 0 | Factual
bilateral pelvic pain | -336 | 0 | Factual
no routinely irrigating or dilating her neovagina | -7560 | 0 | Factual
penetrative sexual intercourse | -7560 | -168 | Factual
life stressors | -168 | 0 | Factual
no intercourse | -168 | 0 | Factual
CT imaging of the abdomen | 0 | 0 | Factual
tubular, heterogenous, fluid-filled structure | 0 | 0 | Factual
outpatient referral to the gynecologist | 0 | 0 | Factual
abdominal pain acutely worsened | 24 | 24 | Factual
diaphoresis | 24 | 24 | Factual
significant distress due to pain | 24 | 24 | Factual
vitals were unremarkable | 24 | 24 | Factual
leukocytosis | 24 | 24 | Factual
absolute neutrophils | 24 | 24 | Factual
repeat abdominal CT | 24 | 24 | Factual
increasing inflammatory process | 24 | 24 | Factual
empiric intravenous piperacillin-tazobactam | 24 | 24 | Factual
transferred emergently to hospital | 24 | 24 | Factual
hypotensive | 48 | 48 | Factual
tachycardic | 48 | 48 | Factual
afebrile | 48 | 48 | Factual
tachypneic | 48 | 48 | Factual
oxygen saturation | 48 | 48 | Factual
IV fluid boluses | 48 | 48 | Factual
antimicrobials changed | 48 | 48 | Factual
exploratory laparotomy | 48 | 48 | Factual
cystoscopy | 48 | 48 | Factual
vaginoscopy | 48 | 48 | Factual
normal bladder | 48 | 48 | Factual
normal urethra | 48 | 48 | Factual
obliterated introitus | 48 | 48 | Factual
diffuse intra-abdominal spillage | 48 | 48 | Factual
perforated sigmoid neovagina | 48 | 48 | Factual
purulent fluid drained | 48 | 48 | Factual
intrabdominal drains placed | 48 | 48 | Factual
intubated | 48 | 168 | Factual
mechanical ventilation | 48 | 168 | Factual
septic shock | 48 | 168 | Factual
vasopressor agents | 48 | 168 | Factual
antimicrobials transitioned | 168 | 168 | Factual
peritoneal culture | 168 | 168 | Factual
blood cultures remained negative | 168 | 168 | Factual
weaned off vasopressors | 192 | 192 | Factual
extubated | 192 | 192 | Factual
transferred to general floor | 288 | 288 | Factual
Infectious Diseases team consulted | 288 | 288 | Factual
antimicrobial management | 288 | 288 | Factual
discharged home | 360 | 360 | Factual
abdominal wound vacuum | 360 | 360 | Factual
IV piperacillin-tazobactam | 360 | 504 | Factual
follow-up with primary care doctor | 360 | 504 | Factual
follow-up with urologist | 360 | 504 | Factual
follow-up with infectious diseases physician | 360 | 504 | Factual
readmitted with sepsis | 504 | 504 | Factual
generalized malaise | 504 | 504 | Factual
diffuse abdominal pain | 504 | 504 | Factual
white blood count | 504 | 504 | Factual
absolute neutrophil count | 504 | 504 | Factual
d-dimer | 504 | 504 | Factual
lactate | 504 | 504 | Factual
CT of chest, abdomen and pelvis | 504 | 504 | Factual
bilateral pleural effusions | 504 | 504 | Factual
loculated left pleural effusion | 504 | 504 | Factual
multiple new abdominal abscesses | 504 | 504 | Factual
transcutaneous drainage catheter | 504 | 504 | Factual
open anterior midline wound | 504 | 504 | Factual
wound vacuum | 504 | 504 | Factual
hypoxemia | 504 | 504 | Factual
transferred to ICU | 504 | 504 | Factual
IV piperacillin-tazobactam continued | 504 | 504 | Factual
placement of right perihepatic drain | 504 | 504 | Factual
aspiration of purulence | 504 | 504 | Factual
unsuccessful drainage of peri-splenic collection | 504 | 504 | Factual
blood cultures remained negative | 504 | 504 | Factual
Interventional radiology reconsulted | 504 | 504 | Factual
drained fluid from abscesses | 504 | 504 | Factual
broad-spectrum PCR | 504 | 504 | Factual
improved clinically | 672 | 672 | Factual
antimicrobials narrowed | 672 | 672 | Factual
discharged | 672 | 672 | Factual
broad-spectrum PCR results | 672 | 672 | Factual
Gleimia europaea | 672 | 672 | Factual
Alistipes onderdonkil | 672 | 672 | Factual
Varibaculum timonense | 672 | 672 | Factual
Jonquetella anthropi | 672 | 672 | Factual
follow-up at adult infectious diseases clinic | 1008 | 1008 | Factual
improved clinically | 1008 | 1008 | Factual
repeat CT abdomen | 1008 | 1008 | Factual
decreased size of abscesses | 1008 | 1008 | Factual
transitioned to oral amoxicillin-clavulanate | 1008 | 1008 | Factual
complete resolution of abscesses | 1008 | 1008 | Factual