38 years old | 0
male | 0
accidental traumatic forearm amputation | 0
steel rope hit arm | 0
amputated distal forearm | 0
wrapped in saline-saturated gauze | 0
cooled on ice | 0
applied tourniquet | 0
replantation decision | 0
broad spectrum antibiotic treatment | 0
replantation surgery | 0
arterial inflow | 0
venous outflow | 0
microbiological testing samples | 0
arterial anastomosis | 48
venous anastomosis | 48
saphenous vein grafts | 48
Coldex skin substitute | 48
swelling | 168
increasing skin necrosis | 168
venous congestion | 168
re-exploration | 168
thrombosis of blood vessels | 168
avital extensor muscles | 168
avital flexor muscles | 168
superficial fungal contamination | 168
amputation at proximal forearm | 168
Amphotericin B | 168
surgical debridement | 168
Bacillus cereus complex | 168
Yersinia enterocolitica | 168
Staphylococcus capitis | 168
Pseudomonas putida | 168
Aspergillus fumigatus | 168
Mucor circinelloides | 168
uncertainty about Mucor invasiveness | 168
Isavuconazol | 384
Tienam | 384
acute renal failure | 432
multi-organ failure | 432
intensive care unit transfer | 432
histologic confirmation of colonization | 360
no angioinvasive infection | 360
preserved ulna length | 360
fasciocutaneous hatchet flap | 840
meshed skin graft | 840
ulnar stump length of 7 centimeters | 840
graft healed well | 1512
transferred to rehabilitation center | 1512
no further complications | 1512
