9 years old | 0
male | 0
admitted to the hospital | 0
periumbilical abdominal pain | -96
watery diarrhea | -96
vomiting | -96
fever | -96
discharged home with analgesics | -48
hospitalized due to worsening of previous symptoms | -24
antibiotics started | -24
transferred to service for diagnostic procedures and surgical evaluation | -24
dysuria | -24
oliguria | -24
abdominal pain | 0
signs of peritonitis | 0
prescribed fasting, antibiotics and maintenance fluid | 0
ultrasound examination | 0
hypothesis of MIS-C | 0
serology requested | 0
RT-PCR nasopharynx/oropharynx swab requested | 0
persistent abdominal pain | 0
diarrhea episodes | 0
persistent tachycardia | 0
abdominal CT | 12
perforated appendix | 12
pelvic abscess | 12
appendectomy and exploratory laparotomy | 12
abscess formation in the pelvis | 12
drain placed in the cavity | 12
anatomopathological examination of the appendix | 12
inflammatory infiltrate with neutrophils and mononuclear cells | 12
hemorrhage | 12
extensive areas of wall necrosis with loss of mucosa | 12
IHC positive for SARS-CoV-2 | 12
RT-PCR positive for SARS-CoV-2 | 12
admitted to the pediatric intensive care unit | 12
fluid resuscitation | 12
oxygen support through nasal cannula | 12
laboratory tests | 12
echocardiogram | 12
normal echocardiogram results | 12
hemodynamically stable | 12
clinical improvement | 12
discharged home | 216
elevated C-reactive protein | 0
elevated fibrinogen | 0
elevated d-dimer | 0
elevated ferritin | 0
leukocytosis | 0
lymphopenia | 0
elevated INR | 0
elevated troponin | 0
elevated creatine kinase | 0
COVID-19 infection confirmed | 0
MIS-C suspected | 0
SARS-CoV-2 infection confirmed | 0
appendicitis | -96
acute inflammatory abdomen | 0
gastrointestinal symptoms | 0
systemic inflammation | 0
coagulation dysfunction | 0
positive RT-PCR | 0
positive serology | 0
asymptomatic previous infection | 0
IgG positive | 0
IgM inconclusive | 0
RT-PCR nasopharynx/oropharynx swab positive | 0
SARS-CoV-2 detected in appendix tissue | 12
viral infection in appendix | 12
MIS-C diagnosed | 216
SARS-CoV-2 infection diagnosed | 0
appendicitis as a complication of SARS-CoV-2 | 12
acute abdomen as a presentation of COVID-19 | 0
GI symptoms in COVID-19 patients | 0
inflammatory profile | 0
coagulation dysfunction | 0
MIS-C as a post-infectious hyperinflammatory complication of SARS-CoV-2 | 216
direct viral effect on tissues | 216
viral entry through ACE 2 | 0
terminal ileitis | 0
appendicitis as a complication of SARS-CoV-2 | 12
inflammation associated with viral entry | 12
reactive lymphoid hyperplasia | 12
luminal obstruction | 12
appendicolith formation | 12
mesenteric adenopathy | 12
malhotra et al | 0
acute appendicitis as a post-infectious hyperinflammatory complication of SARS-CoV-2 | 216
acute GI infection and inflammation trigger the development of appendicitis | 216
cause of appendicitis remains poorly understood | 216
family clusters | 0
seasonal pattern | 0
viral trigger | 0
acute abdominal pain in COVID-19 patients | 0
diagnostic dilemma | 0
delaying management of surgical abdomen | 0
performing unnecessary surgery | 0
iatrogenic morbidity and mortality | 0
strain on healthcare resources | 0
high-risk exposure for healthcare workers | 0
optimum clinical and surgical management | 0
pediatric surgeons and clinicians awareness of GI manifestation of MIS-C | 0
differentiation of MIS-C from other surgical pathologies | 0
broad clinical spectrum of COVID-19 in pediatric population | 0
different phenotypes | 0
latest reports in literature | 0
viral infection in IHC and RT-PCR analysis of appendix | 12
consideration of MIS-C and SARS-CoV-2 infection in diagnostic hypotheses | 0
children with acute abdomen | 0