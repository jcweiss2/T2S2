52 years old | 0
male | 0
admitted to the hospital | 0
high grade fever | 0
shortness of breath | 0
hypotension | 0
urosepsis | 0
poor oral intake | -168
significant weight loss | -168
no history of cough | 0
no history of expectoration | 0
no history of nausea | 0
no history of vomiting | 0
no history of dysuria | 0
no history of bleeding | 0
no history of loose bowel movements | 0
no alteration of higher mental functions | 0
drinking unpasteurized camel milk | -168
hypertension | 0
diabetes | 0
single | 0
denies sexual activities | 0
served in the military | 0
no past history of sexual transmitted diseases | 0
no past history of blood transfusion | 0
no past history of homosexuality | 0
no travel outside the country | 0
moderate distress | 0
febrile | 0
decreased breath sounds | 0
blood pressure 100/50 mmHg | 0
carotid pulsations visible | 0
no bruits | 0
non-elevated jugular venous pressure | 0
normal heart sounds | 0
abdomen soft | 0
abdomen non-tender | 0
no hepatospleenomegaly | 0
no pain on deep palpation | 0
hemoglobin 85 g/liter | 0
total leucocyte count 6200/mm3 | 0
normal platelet count | 0
C reactive protein 222 mg/L | 0
no malaria parasites | 0
internal hemorrhoids | 0
gastritis | 0
gastric biopsy for Helicobacter pylori stain negative | 0
no mediastinal lymphadenopathy | 0
no hilar lymphadenopathy | 0
no axillary lymphadenopathy | 0
pleural effusion | 0
pericardial effusion | 0
no focal changes in liver | 0
no focal changes in pancreas | 0
no focal changes in spleen | 0
no focal changes in kidneys | 0
no focal changes in adrenals | 0
no retroperitoneal lymphadenopathy | 0
no intraperitoneal lymphadenopathy | 0
free abdominal fluid | 0
non-typhoidal Salmonella Group D | 0
sensitive to piperacillin/tazobactam | 0
sensitive to ciprofloxacin | 0
sensitive to ampicillin | 0
resistant to cefuroxime | 0
resistant to gentamicin | 0
resistant to trimethoprim/sulfamethoxazole | 0
positive ELISA result | 0
positive Western blot test | 0
HIV infection | 0
cytology report negative for malignancy | 0
sputum smears negative | 0
sputum cultures negative | 0
ciprofloxacin 200 mg IV twice daily | 0
switched to piperacillin/tazobactam | 72
total duration of treatment 7 days | 168
urine culture negative | 168
discharged | 168