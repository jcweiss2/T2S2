57 years old | 0
male | 0
admitted to the hospital | 0
cough | -504
hemoptysis | -504
pleuritic chest pain | -504
dyspnea on exertion | -504
general malaise | -504
kidney transplantation | -1512
end-stage renal disease | -1512
chronic hemodialysis treatment | -1512
family history of proteinuria | -1512
hypertension | -1512
hypercholesterolemia | -1512
asthma bronchiale | -1512
corticosteroids | -672
Pneumocystis jirovecii prophylaxis | -672
trimethoprim-sulfamethoxazole | -672
mycophenolate mofetil | 0
tacrolimus | 0
methylprednisolone | 0
increased leukocyte count | 0
eosinophilia | 0
systemic involvement | 0
diffuse erythematous or maculopapular eruption | 0
pruritis | 0
DRESS syndrome | 0
fever persisted | 0
rash persisted | 0
discharged | 24
low blood pressure | 168
dizziness | 168
nausea | 168
atypical chest pain | 168
elevated CRP level | 168
elevated troponin I levels | 168
non-ST elevation myocardial infarction | 168
reduced dose of low molecular weight heparin | 168
blood cultures positive for R. equi | 192
R. equi sepsis | 192
meropenem | 192
vancomycin | 192
tapering of immunosuppression | 192
voriconazole stopped | 192
levofloxacin | 216
hypoxic respiratory failure | 240
intensive care unit | 240
CRP level | 240
lactate dehydrogenase level | 240
P. jirovecii pneumonia | 240
trimethoprim-sulfamethoxazole | 240
methylprednisolon | 240
primaquine | 264
clindamycine | 264
moxifloxacin | 672
rifampicin | 672
oral antibiotic regimen | 672
discharged home | 1008
follow-up | 1008
clinical and radiological evolution | 1008
resolution of lung lesion | 1008