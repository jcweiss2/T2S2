39 years old | 0
woman | 0
virgo intacta | 0
heavy menstrual bleeding | -720
submucous leiomyoma | -720
office hysteroscopy | -672
active bleeding | -672
decision to postpone procedure | -672
administration of GnRH agonists | -672
second-look office diagnostic hysteroscopy | -432
difficult entry into uterine cavity | -432
leiomyoma dimensions incompatible with resection | -432
procedure stopped | -432
discharged home | -432
administration of GnRH agonist (goserelin) | -432
admitted to emergency department | -24
mild pelvic pain | -24
vomiting | -24
no fever | -24
no bleeding | -24
ultrasound revealed leiomyoma | -24
no free pelvic fluid | -24
blood analysis no leukocytosis | -24
normal C-reactive protein | -24
prescribed paracetamol | -24
discharged | -24
presented to emergency department | 0
4-day history of intermittent fever | -96
abdominal pain | 0
abdominal distension | 0
multiple episodes of vomiting | -48
limited oral intake | -48
normotensive | 0
normal heartrate | 0
tympanic temperature 37.3 °C | 0
facial flushing | 0
cold extremities | 0
mottled skin | 0
immediate care | 0
large-bore venous catheters | 0
IV fluid infusion | 0
administration of large-spectrum antibiotics | 0
blood samples collected | 0
urine samples collected | 0
vaginal ultrasound performed | 0
normal-sized uterus | 0
leiomyoma | 0
no signs of perforation | 0
virtual uterine cavity | 0
adnexa in retro8-uterine position | 0
limited mobility | 0
previously undiagnosed endometriosis | 0
13-centimeter fluid-filled cystic mass | 0
dilated right fallopian tube | 0
left ovary normal | 0
left fallopian tube normal | 0
no free fluid in pelvic cavity | 0
mildly painful ultrasound | 0
transferred to intermediate care unit | 0
blood analysis no anemia | 0
leukocytosis 16.630/mL | 0
neutrophilia 91% | 0
C-reactive protein 291 mg/dL | 0
acute renal lesion | 0
anuric status | 0
high-volume crystalloid infusion | 0
blood creatinine 4.54 mg/dL | 0
arterial blood gasometry metabolic alkalosis | 0
pH 7.57 | 0
pCO2 43.4 mmHg | 0
HCO3– 39.9 mEq/L | 0
lactate 31 mmol/L | 0
abdominal X-ray | 0
distension of stomach | 0
distension of small bowel | 0
no pneumoperitoneum | 0
CT scan ordered | 0
marked distension of gastric chamber | 0
distension of proximal small bowel | 0
no apparent extrinsic compression | 0
fluid collection in pelvis | 0
possibly cystic | 0
normal liver | 0
normal biliary ducts | 0
normal pancreas | 0
normal kidneys | 0
no hydronephrosis | 0
emergency exploratory laparotomy | 0
ruptured right fallopian tube | 0
hemoperitoneum | 0
generalized pelvic infection | 0
microbial analysis | 0
ampicillin-sensitive E. coli | 0
sub-total hysterectomy | 0
bilateral adnexectomy | 0
transferred to intensive care unit | 0
stage 4 multiple organ failure | 0
mechanical ventilation | 0
administration of vasopressors (dopamine) | 0
hypoperfusion acute kidney injury (KDIGO 3) | 0
responded to fluid resuscitation | 0
aminergic support | 0
full recovery of kidney function | 120
discharged home | 288
oral antibiotics | 288
post-operative evaluation | 288
histological findings acute salpingitis | 288
peritonitis | 288
endometriotic cysts | 288
uterine leiomyomas | 288
no uterine perforation | 288
counseled hormone replacement therapy | 288
