78 years old | 0
female | 0
shortness of breath | -240
dyspnea | -240
acute non-ST segment elevation myocardial infarction | -240
chest pain | -240
tracheal intubation | -240
ventilator-assisted ventilation | -240
vasodilation | -240
hypertension | -13140
coronary heart disease | -13140
cerebral infarction | -4380
anterior wall myocardial infarction | -4380
decreased blood pressure | 0
increased heart rate | 0
fever | 0
septic shock | 0
cardiogenic shock | 0
blood oxygen saturation (SpO2) fluctuations | 0
thick breath sounds | 0
moist rale | 0
heart rate 100 bpm | 0
low and blunt heart sound | 0
no noise in each valve area | 0
dry necrosis of the right lower foot | 0
scattered ecchymoses | 0
serum creatine kinase-MB concentration 25.8 ng/mL | 0
white blood cell count 24.25 × 10^9/L | 0
double lung infection | 0
moderate mitral regurgitation | 0
mild aortic regurgitation | 0
imipenem and cilastatin sodium | -72
anti-infection | -72
dopamine | -72
norepinephrine | -72
anti-shock treatment | -72
percutaneous coronary intervention (PCI) | -72
coronary angiography | -72
right coronary artery stent implantation | -72
stent implantation | -72
vascular opening | -72
body temperature increased | -48
white blood cell count 33.74 × 10^9/L | -48
right lower extremity dry skin necrosis | -48
scattered ecchymoses | -48
right middle iliac artery occlusion | -48
endotracheal tube | -48
fever | -48
SpO2 over 97% | -48
medium flow oxygen inhalation | -48
mid-thigh amputation | 0
tracheal catheter | 0
dopamine 5 µg/kg per min | 0
norepinephrine 0.06 µg/kg per min | 0
non-invasive blood pressure 95/45 mmHg | 0
heart rate 98 bpm | 0
SpO2 99% | 0
left radial artery puncture catheter | 0
arterial blood pressure monitoring | 0
anesthesia system | 0
tracheal catheter | 0
ventilation | 0
ultrasound-guided right-side improved fascia iliaca compartment block | 0
local anesthetics (0.33% ropivacaine hydrochloride 30 mL) | 0
in-plane technique | 0
needle implantation | 0
deep surface of the fascia iliaca | 0
anesthetic plane testing | 5
acupuncture | 5
acupuncture | 10
midazolam 2 mg | 0
sufentanil 10 µg | 0
cisatracurium 6 mg | 0
etomidate 6 mg | 0
general anesthesia induction | 0
1% sevoflurane inhalation anesthesia | 0
anesthesia maintenance | 0
operation duration 65 min | 0
bispectral index 45-60 | 0
vasoactive drugs | 0
blood pressure regulation | 0
heart rate regulation | 0
vital signs stable | 0
CPOT score 2 | 6
Ramsay sedation score 3 | 6
postoperative analgesia satisfactory | 6
inflammatory indicators improved | 48
tracheal intubation removed | 48
discharged | 168