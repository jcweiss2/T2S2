66 years old | 0
female | 0
admitted to the hospital | 0
complaining of cough | 0
tachypnoea | 0
chills | 0
weakness | 0
reduced oxygen saturation | 0
diabetes mellitus | -672
hypertension | -672
dyslipidemia | -672
hypothyroidism | -672
deteriorated to hypoxic respiratory failure | 0
intubated and ventilated | 0
septic shock | 0
acute kidney injury | 0
haemodialysis | 0
high white blood cell count | 0
low platelets | 0
high activated partial thromboplastin time | 0
normal international normalised ratio | 0
normal prothrombin time | 0
high fibrinogen | 0
high D-dimer | 0
high C-reactive protein | 0
high creatinine | 0
high alanine aminotransferase | 0
high aspartate aminotransferase | 0
high alkaline phosphatase | 0
recent travel | -168
tested positive for COVID-19 | 0
computed tomography scan of the head | 504
focal left parietal centrum semiovale vasogenic oedema | 504
magnetic resonance imaging head | 504
widespread susceptibility weighted imaging blooming hypointense foci | 504
microbleeds | 504
juxtacortical white matter | 504
perilesional oedema | 504
no evidence of abscess formation | 504
tiny foci of microbleeds in the internal capsules | 504
critical illness-associated cerebral microbleeds | 504
discharged | -1 
Note: The time stamp for "discharged" is not explicitly mentioned in the text, so it is assumed to be at the end of the hospital stay, which is not specified. Therefore, a timestamp of -1 is assigned, indicating that the discharge time is unknown.