4 years old | 0
female | 0
Mexican | 0
relapsed refractory pre-B cell ALL | -199 
diagnosis of standard risk pre-B ALL | -199 
blasts that coexpressed CD19, CD22, CD58, CD10, CD38 | -199 
cytogenetics that revealed p53 deletion, t(1;19) with a complex karyotype | -199 
no CNS disease | -199 
treated with the National Mexican Protocol | -199 
no evidence of morphologic or minimal residual disease via flow cytometry | -199 
relapsed | -199 
failed reinduction chemotherapy | -199 
failed two cycles of blinatumomab | -199 
treated with reinduction therapy per ALL R3 | -199 
did not achieve remission | -199 
high burden of extramedullary disease in the liver, spleen, kidneys, lymph nodes | -199 
chloroma to left orbit causing a significant cranial nerve II palsy | -199 
renal insufficiency requiring long-term electrolyte replacement | -199 
bridging oral chemotherapy with 6-mercaptopurine and methotrexate | -14 
Staphylococcal epidermidis central catheter infection | -336 
septic shock | -336 
treated with a 10-day course of vancomycin | -336 
lymphoid depleting chemotherapy | -14 
fludarabine | -14 
cyclophosphamide | -14 
fever | -168 
nausea | -168 
headache | -168 
fatigue | -168 
admitted to the emergency department | -168 
initial resuscitation | -168 
work-up | -168 
initiation of broad-spectrum antibiotics | -168 
admitted to the hematology/oncology team | -168 
transferred to the PICU | -132 
septic shock with hypotension | -132 
afebrile | -132 
blood pressure was 69/31 | -132 
heart rate 165 beats per minute | -132 
respiratory rate 56 breaths per minute | -132 
oxygen saturation was 100% on room air | -132 
poor perfusion | -132 
capillary refill time of 5 seconds | -132 
pulses were 3+ in bilateral radial arteries | -132 
intubation | -131 
persistent shock | -131 
contacted the patient’s oncology team | -131 
discuss expected prognosis | -131 
ECMO candidacy | -131 
consent for venoarterial ECMO | -96 
cannulated in the PICU for venoarterial ECMO | -96 
indwelling central catheter was removed | -96 
anticoagulation was managed with systemic heparin | -96 
CRRT via Prismaflex | -96 
therapeutic plasma exchange (TPE) | -96 
broad-spectrum antimicrobial therapy | -96 
meropenem | -96 
ceftazidime/avibactam | -96 
gentamicin | -96 
micafungin | -96 
rapidly weaned off vasoactive and inotropic support | -72 
initiated on milrinone | -72 
afterload reduction | -72 
improvement in systemic vascular resistance | -72 
good antegrade flow across the aortic valve | -72 
no left atrial decompression | -72 
bacteremia cleared | -72 
cardiac dysfunction quickly improved | -72 
repeat echo demonstrating low normal biventricular systolic function | -72 
EF of 51% | -72 
ECMO clamp trial | -72 
decannulated | 120 
extubated | 240 
CAR T-cell infusion (tisagenlecleucel) | 408 
transferred to the hematology/oncology service | 408 
developed cytokine release syndrome | 408 
tocilizumab | 408 
brief PICU readmission | 408 
identified to be in remission | 720 
discharged from the hospital | 720