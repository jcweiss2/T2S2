2260-g male infant | 0
born at 34 weeks | 0
central placenta previa | 0
hemorrhage | 0
hyperthyroidism | 0
full dose of dexamethasone | 0
Apgar score 8 at 1 minute | 0
Apgar score 9 at 5 minutes | 0
admitted to the neonatal intensive care unit | 0
intubated | 0
respiratory distress | -30
pulmonary hemorrhage | 0
high-frequency oscillatory ventilation | 0
inhalational nitric oxide | 3
PPHN | 3
surfactant | 0
umbilical venous catheter | 0
umbilical artery catheter | 0
hypotension | 0
substantial fluid administration | 0
intensive inotropic support | 0
hydrocortisone 2 mg/kg q8h | 0
epinephrine | 0
dopamine | 0
mean arterial pressure increased to 92 mmHg | 168
hyperbilirubinemia | 0
greatest indirect bilirubin 434 μmol/L | 0
blood exchange | 0
albumin 2 g | 0
acute hypokalemia | 336
serum potassium 2.1 mmol/L | 336
potassium replacement 0.3 mmol/kg/h | 336
oral repletion 4 mmol/kg/d | 336
serum potassium 2.8-3.3 mmol/L | 336
fetal echocardiography at 24 weeks | -1344
structurally normal heart | -1344
pediatric cardiology consultation | 0
transthoracic echocardiogram | 0
right-to-left shunting across foramen ovale | 0
large patent ductal arteriosus | 0
second transthoracic echocardiogram | 72
mean pulmonary artery pressure 35 mmHg | 72
LVEF 67% | 72
atrial left-right shunt | 72
patent ductal shunt | 72
PPHN persistent | 72
third transthoracic echocardiogram | 264
PPHN ameliorated | 264
mean pulmonary artery pressure 23 mmHg | 264
normal IVS thickness | 264
profound cardiomegaly | 720
grade III/IV harsh systolic ejection murmur | 720
transthoracic echocardiogram at day 30 | 720
IVS thickening 13.8 mm | 720
LVPW thickening 6 mm | 720
IVS/LVPW 2.3 | 720
hypertrophic cardiomyopathy | 720
outflow tract obstruction not observed | 720
peak velocity 0.85 m/s | 720
aortic coarctation ruled out | 720
negative maternal risk factors | 720
negative familial history | 720
normal maternal oral glucose tolerance test | 720
normal glycated hemoglobin | 720
propranolol 0.2 mg q8h | 720
captopril 0.02 mg q8h | 720
no arrhythmia | 720
transesophageal echocardiograms | 720
IVS thickness decreased to 3 mm | 1440
asymptomatic | 720
supplemental oxygen discontinued | 720
normal tandem mass spectroscopy | 720
normal exome sequencing | 720
discharged | 1080
MAP 65 mmHg | 1440
normal cardiologic evaluation | 1440
hypotension responsive to fluid and inotropic support | 0
hydrocortisone weaned over 5 days | 0
MAP remained at 85 ± 7.4 mmHg | 0
serum potassium normalized | 336
serial echocardiograms showing IVS decrease | 720
spontaneous reversal of hypertrophy | 720
hypertension | 720
hyperglycemia | 720
GI hemorrhage | 720
perforation | 720
cerebral palsy | 720
increased MAP | 720
normal LVOT flow | 720
remission of left ventricular hypertrophy | 1440
improvement of septal configuration | 1440
discharge follow-up | 1440
HCM associated with HC | 0
genetic HCM ruled out | 720
metabolic causes ruled out | 720
prenatal causes ruled out | 720
maternal causes ruled out | 720
HC suppresses inflammatory response | 0
HC induces adrenergic receptors | 0
HC inhibits catecholamine metabolism | 0
HC increases intracellular calcium | 0
HC enhances adrenergic response | 0
HC-related myocardial thickening | 0
HC acts through IGF1 | 0
HC induces LV hypertrophy | 0
thickened IVS blocking blood flow | 720
arrhythmias risk | 720
beta blockers | 720
calcium channel blockers | 720
septal myectomy | 720
ablation | 720
implantable cardioverter-defibrillator | 720
HC-induced HCM benign | 720
HCM resolution post HC discontinuation | 720
hypertension related to HCM | 720
increased hypertrophy with HC dose/duration | 0
insulin with HC may increase hypertrophy | 0
risk/benefit HC in septic shock | 0
HCM monitoring recommendations | 0
novel therapeutic approaches | 0
