40 years old | 0
male | 0
admitted to the hospital | 0
hematemesis | 0
catheter ablation of the left atrium | -672
medically refractory rapid AF | -672
pleuritic chest pain | -504
odynophagia | -504
malaise | -504
headache | -504
fevers | -504
sepsis | 0
temperature of 100.8°F | 0
heart rate 96 bpm | 0
blood pressure 89/50 mm Hg | 0
responsive to fluid resuscitation | 0
thoracic CT with intravenous contrast | 0
small locules of gas along the esophageal wall | 0
abutting the left atrium | 0
no definite esophageal perforation or AEF | 0
transferred to cardiothoracic intensive care unit | 0
gated thoracic CT with intravenous contrast | 24
punctate foci of gas between the left atrium and the esophagus | 24
concerning esophageal leak | 24
no clear AEF | 24
Gastroenterology consultation | 24
upper endoscopy without CO2 insufflation | 24
esophagus could not be adequately examined | 24
minimal insufflation with CO2 | 24
large amount of fresh blood in the mid esophagus | 24
confirmation of AEF | 24
new-onset left hemiplegia | 29
left gaze deviation | 29
lethargy | 29
emergent surgery | 29
3 × 5 mm defect in the posterior wall of the left atrium | 29
visibility of esophageal fibers through a perforation | 29
postoperative cranial CT without contrast | 53
new right middle cerebral artery territory ischemic stroke | 53
cranial CT angiography | 53
normal vasculature | 53
Streptococcus mitis bacteremia | 120
no evidence of infective endocarditis on transthoracic echocardiogram | 120
discharged home on intravenous antibiotics | 480
six-week treatment | 480
outpatient rehabilitation | 480
significant clinical improvement | 2160
mild left-sided neurological deficits | 2160