54 years old | 0
man | 0
admitted to the hospital | 0
insulin dependent diabetes mellitus | 0
hepatitis C chronic infection | 0
liver cirrhosis child B | 0
esophageal varices | 0
right sided facial weakness | -168
right sided headache | -168
blocked right nostril | -168
fever of 7 days | -168
treatment for presumed bell's palsy | -168
short course of steroids | -168
BP 140/70 mmHg | 0
pulse of 92 beat per minute | 0
oxygen saturation of 99% | 0
temperature of 38.2 Celsius | 0
swelling of the right side of the face | 0
right eye complete ptosis | 0
chemosis | 0
injection | 0
mid dilated fixed pupil | 0
right frozen globe | 0
multiple cranial nerves palsies | 0
II | 0
III | 0
IV | 0
V1 | 0
VI |0
VII |0
no other focal neurological deficits |0
right central retinal artery occlusion |0
edematous retina |0
right side black discoloration |0
pale mucosa |0
high WBC count |0
hyperglycemia |0
abnormal kidney function |0
pansinusitis |0
IV fluids |0
insulin |0
IV liposomal amphotericin |0
linezolid |0
ceftazidime |0
complicated fungal infection |0
right radical endoscopic sinus surgery |24
extubated |24
pansinusitis |24
inflammatory changes |24
bony defect |24
nasal swab positive for Mucor species |24
invasive mucormycosis |96
afebrile |24
blood sugar improved |24
kidney function improved |24
serum creatinine 260 µmol/L |96
amphotericin toxicity |96
contrast induced nephropathy |96
IV fluids support continued |96
IV amphotericin continued |96
deteriorated |192
decreased level of consciousness |192
confusion |192
GCS drop to 9/15 |192
vital signs stable |192
non contrast head CT showed no new changes |192
presumed hepatic encephalopathy |192
lactulose |192
broad spectrum antibacterial agents |192
monitoring of mental status |192
level of consciousness not improved |360
brain MRI |360
total occlusion of the right internal carotid artery |360
right anterior cerebral artery occlusion |360
right middle cerebral artery occlusion |360
edema effect |360
compression of the right posterior cerebral artery |360
secondary massive infarction |360
hemorrhagic change |360
secondary mass effect |360
significant midline shift |360
declared brain dead |408
apnea test positive |408
withdraw of care discussed |408
family objected |408
passed away |504
refractory septic shock |504
