69 years old | 0
male | 0
Caucasian | 0
admitted to the hospital | 0
abdominal pain | -48
nausea | -48
atrial fibrillation | 0
diabetes | 0
chronic kidney disease | 0
left thoracotomy for lung cancer resection | 0
micropenis | -336
microhematuria | -336
urinalysis | -336
cystoscopy | -336
CT scan | -336
left perinephric mass | -336
enlarged peri-renal and para-aortic lymph nodes | -336
retroperitoneal streaky changes | -336
CT-guided peri-renal lesion biopsy | -336
atypical cellular proliferation | -336
surveillance | -336
increasing abdominal pain | -336
tachycardia | 0
abdomen distended | 0
abdomen tender | 0
positive fluid wave | 0
leukocytosis | 0
ultrasound-guided paracentesis | 0
bloody fluid | 0
repeat CT imaging | 0
concern for urine extravasation | 0
fluid analysis | 0
serum-ascites albumin gradient (SAAG) <1.1 g/dL | 0
paracentesis | 72
bloody fluid | 72
urology consultation | 72
retrograde pyelogram | 72
urine extravasation | 72
left ureteral stent | 72
left nephrostomy tube | 72
urinary diversion | 72
discharged home | 96
readmitted | 120
syncopal event | 120
painful abdominal distention | 120
frequent paracenteses | 120
hemorrhagic ascites | 120
surgical oncology consultation | 192
tumor markers | 192
AFP | 192
CEA | 192
CA 19-9 | 192
diagnostic laparoscopy | 192
purplish discoloration | 192
thickening of omentum | 192
inflammatory reaction | 192
biopsy of omentum | 192
frozen section analysis | 192
atypical cellular proliferation | 192
necrosis | 192
bloody peritoneal fluid | 192
systemic inflammatory response | 216
intensive care unit admission | 216
exploratory laparotomy | 240
omentectomy | 240
sepsis | 240
tissue necrosis | 240
normal liver | 240
normal gallbladder | 240
normal pancreas | 240
serositis | 240
necrotic greater omentum | 240
peri-renal mass | 240
Gerota’s fascia | 240
lower lobe of left kidney | 240
bloody ascites fluid | 240
high-grade angiosarcoma | 240
palliative chemotherapy | 240
clinical status decline | 288
death | 312