53 years old | 0
female | 0
admitted to the hospital | 0
intermittent abdominal pain | -43800
fever | -43800
cholecystectomy | -28800
abdominal pain worsened | -72
hyperpyrexia | -72
chills | -72
jaundice | -72
dyspnea | -72
decreased oxygen saturation | -72
elevated total bilirubin | -72
liver-protective therapy | 0
anti-infective treatment | 0
hepatectomy | 0
cholangioplasty | 0
left hepaticolithotomy | 0
second biliary duct exploration | 0
choledocholithotomy | 0
T-tube drainage | 0
accretion lysis | 0
liver showed nodular and atrophic changes | 0
cirrhosis | 0
splenomegaly | 0
splenic varices | 0
elevated total bilirubin | 144
worsened coagulation function | 144
respiratory failure | 192
septicemia | 192
Pseudomonas aeruginosa | 192
bilateral pulmonary infection | 192
bilateral pleural effusion | 192
tracheal intubation | 192
ventilator support | 192
packed red blood cell transfusion | 192
fresh frozen plasma transfusion | 192
noradrenaline bitartrate | 192
artificial liver support therapy | 336
plasmapheresis | 336
reintubation | 360
disturbance of consciousness | 360
decreased oxygen saturation | 360
discontinuation of treatment | 480
liver failure | 480
respiratory failure | 480
septicemia | 480
death | 480
DRESS syndrome | -672 
diffuse erythematous or maculopapular eruption | -672 
pruritis | -672 
fever persisted | 0
rash persisted | 0 
discharged | 24