68 years old | 0
male | 0
heavy smoker | 0
no previous medical history | 0
no known history of allergy | 0
no known history of asthma | 0
admitted to the hospital | 0
near cardiac arrest | -1
persistent severe hypotension | -1
made spicy pork kidneys for dinner | -3
gasping on the armchair | -1
telephone-assisted cardiopulmonary resuscitation (CPR) | -1
spontaneous circulation restored | -0.25
severely hypotensive | 0
norepinephrine administration | 0
afebrile | 0
tachycardic | 0
tachypneic | 0
oxygen saturation of 85% | 0
drowsy yet awake | 0
Glasgow coma scale of 4-5-6 | 0
auscultation of the heart failed to reveal any murmurs | 0
lung sounds were clear | 0
abdomen was soft with no tenderness or guarding | 0
skin examination did not reveal any efflorescence | 0
tick embedded in the skin extracted | 0
mechanical ventilation initiated | 0
electrocardiogram showed sinus tachycardia | 0
white cell count of 14,700 per cubic millimetre | 0
C-reactive protein elevated to 64 mg/l | 0
procalcitonin (0.1 ng/ml) | 0
renal functions normal | 0
hepatic enzymes normal | 0
lactate markedly elevated (6.3 mmol/l) | 0
bed-side echocardiography failed to reveal hypovolemia | 0
high left ventricle ejection fraction | 0
whole-body CT showed consolidation of the lower lobe in the left lung | 0
suspected pneumonia | 0
treated empirically for pneumonia and septic shock | 0
itchy skin | -2
postprandial timing | -2
serum tryptase sample obtained | 2
serum tryptase significantly higher than normal | 2
total IgE levels elevated | 2
investigation of potential trigger | 2
specific IgE against alpha-gal highly positive | 4
allergologist consultation requested | 4
diagnosed with alpha-gal syndrome | 4
vasoplegic shock | 0
cardiac arrest | -1
alpha-gal syndrome as a causative factor | 4
rapid progression to cardiac arrest | -1
galactose-alpha-1,3-galactose expressed on glycoproteins and glycolipids of mammals | 0
specific IgE antibodies formation | 0
tick saliva contains immunologically active substances | 0
IL-4 causes isotype switching to IgE antibodies production | 0
majority of patients sensitised to alpha-gal will never develop the alpha-gal syndrome | 0
typical case of alpha-gal syndrome has an adult-life onset | 0
clinical symptoms usually delayed and start 3–6 hours after ingestion | 0
symptomatology includes typical allergic reactions | 0
abdominal pain without skin involvement | 0
anaphylaxis or anaphylactic shock | 0
diagnosis mainly based on history of eating red meat | 0
detecting specific IgE antibodies | 0
prick tests with extracts of beef or pork unreliable | 0
red meat a source of alpha-gal | 0
milk and milk-based products contain alpha-gal | 0
butter contains alpha-gal | 0
sweets containing gelatine contain alpha-gal | 0
some medicaments contain alpha-gal | 0
treatment of acute allergic reaction does not differ from standard practice | 0
patients should know that any further tick bite can increase the titres of alpha-gal antibodies | 0
patients advised to avoid mammalian meat products | 0
avoidance of dairy products and other mediators of alpha-gal not routinely advised | 0
life-threatening protracted delayed vasoplegic shock | 0
animal organ consumption | -3
tick bite | -3
initially mistaken for sepsis | 0
tick-borne anaphylaxis due to alpha-gal syndrome | 4
severe protracted anaphylaxis in this type of allergy | 0
alpha-gal syndrome a potentially life-threatening syndrome | 0
primary source of this IgE–binding epitope are mammalian products | 0
sensitisation to this antigen requires a tick bite | 0
typical cases present as a delayed anaphylaxis after red meat consumption | 0
atypical clinical manifestation without common allergic symptomatology and trigger may occur | 0
diagnostic errors may occur | 0
importance of avoiding mental shortcuts in the diagnostic process | 0
tick-borne diseases tend to rise in incidence and prevalence | 0
alpha-gal syndrome yet rare | 0