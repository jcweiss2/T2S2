29 years old | 0  
    male | 0  
    admitted to the hospital | 0  
    cardiogenic shock | -432  
    biventricular failure | -432  
    ejection fraction 5-10% | -432  
    myopericarditis | -432  
    constrictive physiology | -432  
    peripherally inserted central catheter (PICC) line placed | -432  
    discharged on milrinone | -432  
    presented to Emergency Department | -432  
    septic shock | -432  
    PICC line removed | -432  
    started on IV vancomycin | -432  
    started on piperacillin/tazobactam | -432  
    transferred to intensive care unit | -432  
    vasopressor support | -432  
    Chryseobacterium indologenes grew from admission PICC line | 0  
    Chryseobacterium indologenes grew from peripheral blood cultures | 0  
    PICC line dressing contaminated with tap water during bathing | 0  
    antibiotics changed to ciprofloxacin | 0  
    antibiotics continued on piperacillin/tazobactam | 0  
    weaned off vasopressor support | 0  
    underwent pericardiectomy | 264  
    completed 14 days of antibiotics | 408  
    discharged from the hospital | 504  
    stable vital signs | 504  
    labs | 504  
    seen in outpatient cardiology clinic | 8760  
    remains in good health | 8760  
    no evidence of recurrent infection | 8760  
    fevers | 0  
    chills | 0  
    progressive fatigue | -432  
    dyspnoea on exertion | -432  
    non"ischemic cardiomyopathy | -432  
    viral myopericarditis | -432  
    computed tomography angiography | -432  
    cardiomegaly | -432  
    dilated right atrium | -432  
    passive hepatic congestion | -432  
    right ventricular failure | -432  
    pericardial calcification | -432  
    no evidence of constrictive pericarditis | -432  
    echocardiogram showed biventricular failure | -432  
    features of constrictive pericarditis | -432  
    cardiac magnetic resonance imaging | -432  
    left ventricular ejection fraction 23% | -432  
    right ventricular ejection fraction 36% | -432  
    delayed gadolinium enhancement | -432  
    scarring/fibrosis | -432  
    non"coronary artery disease hyperenhancement pattern | -432  
    no evidence of infiltrative process | -432  
    prior myocarditis | -432  
    diastolic septal bounce | -432  
    concentrically thickened pericardium | -432  
    atrial flutter | -432  
    rapid ventricular response | -432  
    radiofrequency ablation | -432  
    cardiogenic shock | -432  
    stabilized on inotrope therapy | -432  
    discharged on home milrinone infusion | -432  
    seen by cardiothoracic surgery | -432  
    plans for elective pericardiectomy | -432  
    symptom burden | -432  
    fever 38.7°C | 0  
    chills for 1 day | 0  
    no other complaints | 0  
    home medications | 0  
    furosemide 40 mg once daily | 0  
    losartan 12.5 mg once daily | 0  
    metoprolol succinate 12.5 mg once daily | 0  
    milrinone 0.25 µg/kg/min | 0  
    spironolactone 12.5 mg once daily | 0  
    initial vitals | 0  
    fever 38.7°C | 0  
    tachycardia | 0  
    heart rate 110 | 0  
    blood pressure 96/57 mmHg | 0  
    exam | 0  
    tachycardic heart | 0  
    normal rhythm | 0  
    no murmurs | 0  
    no rubs | 0  
    no gallops | 0  
    no signs of elevated jugular venous pressure | 0  
    no lower extremity edema | 0  
    bilateral radial pulses 2+ | 0  
    dorsalis pedis pulses 2+ | 0  
    lungs clear | 0  
    normal work of breathing | 0  
    no redness around PICC line | 0  
    no drainage around PICC line | 0  
    chest X-ray showed no abnormalities | 0  
    electrocardiogram | 0  
    sinus tachycardia | 0  
    normal axis | 0  
    RSR' pattern in V1 | 0  
    QRS duration 90 ms | 0  
    non"specific T wave flattening | 0  
    removal of PICC line | 0  
    fever 39.5°C | 0  
    severe rigours | 0  
    hypotension | 0  
    blood pressure 70/40 mmHg | 0  
    elevated lactate 5.5 mmol/L | 0  
    blood cultures drawn peripherally | 0  
    blood cultures drawn from PICC line | 0  
    started on empiric vancomycin | 0  
    started on empiric piperacillin/tazobactam | 0  
    transferred to cardiac intensive care unit | 0  
    vasopressor support | 0  
    septic shock | 0  
    catheter"related bloodstream infection | 0  
    advanced heart failure service consulted | 0  
    plans for pericardiectomy | 0  
    preliminary report of blood cultures | 0  
    Gram"negative rods | 0  
    speciated as Chryseobacterium indologenes | 0  
    cultures from PICC line positive | 0  
    peripheral blood cultures positive | 0  
    infectious disease team consulted | 0  
    started on ciprofloxacin | 0  
    continued on piperacillin/tazobactam | 0  
    susceptibility testing | 0  
    sensitive to ciprofloxacin | 0  
    sensitive to piperacillin | 0  
    sensitive to trimethoprim/sulfamethoxazole | 0  
    resistant to meropenem | 0  
    improved clinically | 0  
    remained afebrile | 0  
    weaned off vasopressor support | 0  
    follow"up blood cultures negative | 0  
    interval echocardiogram | 0  
    dilated left ventricle | 0  
    hypertrophied left ventricle | 0  
    diastolic septal bounce | 0  
    constrictive pericarditis | 0  
    ejection fraction 30"35% | 0  
    dilated right ventricle | 0  
    reduced systolic function | 0  
    no valvular stenosis | 0  
    no regurgitation | 0  
    no vegetations | 0  
    right heart catheterization | 0  
    left heart catheterization | 0  
    discordance of ventricular pressures | 0  
    diastolic equalization of pressures | 0  
    optimal timing of pericardiectomy discussed | 0  
    repeat blood cultures negative | 0  
    pericardiectomy on hospital day 11 | 264  
    intraoperative findings | 264  
    dense adhesions | 264  
    calcium deposits | 264  
    adhesions taken down | 264  
    complete pericardium removal | 264  
    follow"up transthoracic echocardiogram | 264  
    left ventricular ejection fraction 50"55% | 264  
    right ventricular systolic function improved | 264  
    continued on piperacillin/tazobactam | 264  
    continued on ciprofloxacin | 264  
    discharged after antibiotic completion | 504  
    inotrope independent | 504  
    guideline"directed medical therapy | 504  
    furosemide 40 mg once daily | 504  
    metoprolol succinate 12.5 mg once daily | 504  
    sacubitril"valsartan 24"26 mg every 12 h | 504  
    followed by outpatient cardiologist | 504  
    seen in October 2019 | 8760  
    great improvement in functional status | 8760  
    denied heart failure symptoms | 8760  
    NYHA Class I | 8760  
    no evidence of recurrent infection | 8760  
    Gram"negative bacilli | 0  
    non"motile | 0  
    indole"positive | 0  
    environmental sources | 0  
    systemic illness | 0  
    congestive heart failure | 0  
    constrictive myopericarditis | 0  
    indwelling PICC line | 0  
    tap water contamination hypothesis | 0  
    sleeve failure | 0  
    water seepage | 0  
    contamination of PICC line dressing | 0  
    appropriate antibiotics | 0  
    line removal | 0  
    fluoroquinolone treatment | 0  
<|eot_id|>
    