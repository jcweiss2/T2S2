26 6/7 weeks gestational age | -672
normal spontaneous vaginal delivery | -672
40-year-old mother | -672
G3P1011 | -672
history of sickle trait | -672
admitted to the Neonatal Intensive Care Unit | 0
prematurity | 0
respiratory distress syndrome | 0
chronic lung disease | 0
suspected sepsis | 0
metabolic acidosis | 0
anemia | 0
suspected necrotizing enterocolitis | 0
cow’s milk protein allergy | 0
newborn screening | -240
diagnosis of SCD | -240
repeat hemoglobin electrophoresis | -150
SCD-SS type | -150
irritable | -589
swelling of the left thigh | -589
tenderness | -589
minimal active movement | -589
non-displaced fracture of the left femoral shaft | -589
periosteal reaction | -589
splint | -579
healing fracture | -579
calcium normal | -579
phosphorus normal | -579
vitamin D normal | -579
alkaline phosphatase level 599 units/L | -593
alkaline phosphatase level 699 units/L | -672
bluish sclera | -579
OI type 1 | -579
genetic testing | -579
13th percentile for length | 540
below the third percentile for weight | 540
no further fractures | 540
hospitalized for sickle cell pain crisis | 8760
irritability | 8760
inability to bear weight on right lower extremity | 8760
no new fractures | 8760
hospitalized for sickle cell pain crisis | 14520
irritability | 14520
inability to bear weight on right lower extremity | 14520
no new fractures | 14520
folic acid | 540
prophylactic penicillin | 540
vitamin D supplementation | 540
referred to a comprehensive center for OI | 540