60 years old | 0
female | 0
nausea | -2
vomiting | -2
steroid treatment | -672
malignant lymphoma | -672
abdominal pain | -2
abdominal mass | -2
increased inflammation | -2
acidosis | -2
abdominal CT | -2
thickness of the descending colon | -2
swelling of surrounding lymph nodes | -2
ascites | -2
decreased blood pressure | -1
decreased level of consciousness | -1
sepsis | -1
colectomy | 0
stoma creation | 0
admitted to ICU | 0
early rehabilitation | 0
multiple organ failure | 1
tracheotomy | 288
GCS 4 | 288
anisocoria | 288
abnormal light reflex | 288
disorder of eye movement | 288
facial muscle paralysis | 288
severe flaccid weakness | 288
diminished deep tendon reflexes | 288
MRC sum score 0 | 288
head CT | 288
ICUAW | 288
active rehabilitation | 288
nutritional support | 288
glycemic control | 288
MRC score improved to 50 | 4320
discharged | 4320