46 years old | 0
male | 0
Caribbean-Black | 0
admitted to the hospital | 0
fever | -48
cough | -48
shortness of breath | -48
systolic blood pressures of 140 mm Hg | 0
heart rate of 142 beats per minute | 0
respiratory rate of 28 breaths per minute | 0
oxygen saturation of 88% on room air | 0
hypertension | 0
tachycardia | 0
tachypnea | 0
normal jugular venous pulse | 0
scattered bilateral crackles | 0
no peripheral edema | 0
atrial flutter (AFL) | 0
2 to 1 atrioventricular block | 0
rate-related ST-T segment changes | 0
chest radiograph did not reveal any acute cardiopulmonary disease | 0
preserved left ventricular ejection fraction | 0
no regional wall motion abnormalities | 0
D-dimer 357 ng/dL | 0
pro-brain natriuretic peptide 413 pg/mL | 0
cardiac biomarkers | 0
CK-MB 15 U/L | 0
troponin I 0.12 ng/mL | 0
mild hypoxia on 24% fractional inspiration of oxygen | 0
estimated alveolar-arterial gradient of 17 mm Hg | 0
amiodarone and digoxin bolus | 0
moderate-intensity beta-blockade | 0
initiated on an amiodarone infusion | 0
atenolol | 0
cardioversion with 100 J | 12
transitioned to atrial fibrillation with rapid ventricular response | 12
COVID-19 test returned positive | 12
transferred to another quarantine facility | 24
intensive care unit (ICU) capabilities | 24
discharged to home quarantine | 72
oral low dose, twice daily amiodarone | 72
follow-up visit | 168
1-week Holter monitor | 168
reverted to normal sinus rhythm | 48
anticoagulation was deferred | 48
CHADS-VASc score of 0 | 48
HAS-BLED score of 0 | 48
anemia | 0
mild rhabdomyolysis | 0
hypokalemia | 0
hypomagnesemia | 0
hypophosphatemia | 0
electrolyte abnormalities | 0
aggressively repleted | 24
tachycardia | 0
adequate volume resuscitation | 24
judicious intravenous crystalloid hydration | 24