23 years old | 0
female | 0
learning disability | -175200 (assuming childhood onset, approximately 20 years prior)
meningitis | -175200
generalized abdominal pain | -48
peritonitis | 0
abdominal ultrasonography | 0
periappendicular fat infiltration | 0
intraperitoneal effusion | 0
septic shock | 0
median laparotomy | 0
appendicular perforation | 0
purulent effusion | 0
perforation of cecal tumoral mass | 0
tumor fixation posteriorly | 0
invasion of adjacent structures | 0
liver palpation | 0
right annexe palpation | 0
adenomegaly in right mesocolon | 0
tumor adhesion to second duodenum | 0
right hemicolectomy R2 | 0
ileostomy | 0
postoperative septic shock | 0
transfer to university hospital | 0
12 days ICU stay | 288
pathological examination | 0
mesenchymal tumor | 0
immunohistochemical diagnosis of schwannoma | 0
thoracoabdominopelvic CT scan | 720
tumoral residue in right iliac fossa | 720
multidisciplinary meeting discussion | 720
decision for complementary resection | 720
restore digestive continuity | 2160
tumoral residue invading right annexe | 2160
right iliac vessels invasion | 2160
right ureter invasion | 2160
outpatient follow-up | 0
CT scan control at 2 years | 17520
mesenteric recurrence | 17520
stability of tumoral residue | 17520
exploratory laparotomy | 17520
unresectable mesenteric mass | 17520
parietal nodules | 17520
surgical biopsies of nodules | 17520
neurofibromatous nature confirmed | 17520
multidisciplinary meeting decision on adjuvant treatment | 17520
suspected neurofibromatosis | 17520
lack of oncogenetic investigation | 17520
4-year follow-up | 35040
right nephrostomy | 35040
ureter compression | 35040
learning disability | -175200
transfer to university hospital |DONE
