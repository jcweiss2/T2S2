27 years old | 0
male | 0
admitted to our emergency department | 0
recurrent fever | -1008
fatigue | -1008
unconsciousness | -24
bilateral lung infection | -1008
high WBC count | -1008
low RBC count | -1008
low hemoglobin | -1008
low platelet count | -1008
high CRP concentration | -1008
prescribed moxifloxacin | -1008
refused admission | -1008
temperature 38.5°C | 0
pulse rate 129 beats/min | 0
respiratory rate 42 beats/min | 0
transcutaneous saturation of oxygen 65% | 0
blood pressure 85/55 mmHg | 0
infusion of norepinephrine | 0
intubated | 0
mechanical ventilation | 0
moist crackles | 0
anoxia | 0
hyperventilation | 0
low partial pressures of oxygen | 0
low partial pressures of carbon dioxide | 0
pH 7.516 | 0
higher WBC count (34.45 × 10⁹/L) | 0
higher CRP concentration (80.78 mg/L) | 0
lower hemoglobin (90.00 g/L) | 0
lower platelet count (80.78 × 10⁹/L) | 0
RBC count 3.36 × 10¹²/L | 0
mean corpuscular volume 120.1 fL | 0
mean corpuscular hemoglobin 40.8 pg | 0
elevated erythrocyte sedimentation rate | 0
elevated ferritin | 0
severe multiple patchy shadows in both lungs | 0
consolidation | 0
worsened pneumonia | 0
initial diagnosis of severe pneumonia | 0
sputum samples for mNGS | 0
detected Epstein–Barr virus | 0
detected Mycobacterium kansasii | 0
chromosomal copy number analysis duplication on chromosome 8 | 0
alveolar lavage fluid for mNGS | 48
detected Cordyceps portugal | 48
confirmed M. kansasii | 48
confirmed chromosome 8 duplication | 48
bone marrow aspiration | 48
evidence of infection in bone marrow | 48
karyotype analysis trisomy 8 | 48
immunophenotypic analysis ruled out leukemia | 48
blood cultures detected Candida Portugal | 48
diagnosis of severe pneumonia | 0
respiratory failure | 0
septic shock | 0
anemia | 0
thrombocytopenia | 0
trisomy 8 | 0
treatment with moxifloxacin | -1008
treatment with imipenem | 0
treatment with vancomycin | 0
ambroxol | 0
omeprazole | 0
enteral nutrition | 0
discontinuation of vancomycin | 72
addition of fluconazole | 120
administration of methylprednisolone 500 mg daily | 168
discontinuation of imipenem | 240
substitution with piperacillin–tazobactam | 240
reduction of methylprednisolone to 250 mg daily | 240
extubation | 288
reduction of methylprednisolone to 120 mg daily | 312
reduction of methylprednisolone to 60 mg daily | 384
transfer to Department of Respiratory Medicine | 408
discharged | 456
no notable history of past illness | 0
no notable personal or family history | 0
no abnormalities on physical examination other than respiratory | 0
no obvious abnormalities on liver and spleen ultrasonography | 0
no gastrointestinal involvement | 0
no progression to hematological malignancy | 0
no MDS | 0
