58 years old | 0
male | 0
admitted to the hospital | 0
fever | -72
perineal erythema | -72
pain | -72
mild seasonal allergies | 0
ingual herniorrhaphy | -2628
fexofenadine | 0
pseudoephedrine | 0
perineal cellulitis | 0
subcutaneous air | 0
Fournier's gangrene | 0
normotensive | 0
tachycardic | 0
increased heart rate | 0
no cardiac murmurs | 0
no ST, T-wave changes | 0
no third heart sound | 0
no peripheral edema | 0
no jugular venous distention | 0
clear lungs | 0
SpO2 98% | 0
hemoglobin 14.9 g/dL | 0
hematocrit 44% | 0
white blood cell count 12.7 × 10^3 / mL | 0
platelet count 146,000 / mL | 0
sodium 135 mmol / L | 0
potassium 4.3 mmol / L | 0
chloride 99 mmol / L | 0
HCO3 26 mmol / L | 0
blood urea nitrogen 16 mg / dL | 0
creatinine 1.14 mg / dL | 0
midazolam 2 mg | -1
propofol 200 mg | -1
fentanyl 100 mcg | -1
sevoflurane 2-3% | -1
fentanyl 500 mcg | -1
dilaudid 1 mg | -1
LMA placement | -1
surgical debridement | 0
tachypnea | 0
respiratory rate 35 breaths / minute | 0
surgical blood loss 200 mL | 0
LMA removal | 1
laryngospasm | 1
tachycardia | 1
hypertension | 1
positive pressure ventilation | 1
propofol | 1
succinylcholine | 1
orotracheal intubation | 1
bilateral rales | 1
pink frothy secretions | 1
tachycardia | 2
hypertension | 2
SpO2 85-88% | 2
FiO2 100% | 2
pH 7.27 | 2
PaCO2 59 mmHg | 2
PaO2 46 mmHg | 2
HCO3 16 mmol / L | 2
base excess -1.9 | 2
oxygen saturation 75% | 2
lactate 1.27 mmol / L | 2
SIMV | 2
tidal volume 750 mL | 2
pressure support 10 cm H2O | 2
PEEP 10 cm H2O | 2
PEEP increased to 12 cm H2O | 4
SpO2 > 90% | 4
ICU admission | 4
SIMV | 4
tidal volume 580 mL | 4
FiO2 100% | 4
pressure support 15 cm H2O | 4
PEEP 12 cm H2O | 4
pH 7.6 | 4
PaCO2 25 mmHg | 4
PaO2 165 mmHg | 4
HCO3 27 mmol / L | 4
SpO2 99% | 4
FiO2 weaned to 40% | 12
pH 7.45 | 12
PCO2 41 mmHg | 12
PaO2 78 mmHg | 12
HCO3 28 mmol / L | 12
base excess 3.8 | 12
oxygen saturation 96% | 12
re-debridement | 48
extubation | 72
shortness of breath | 72
pH 7.49 | 72
PCO2 39 mmHg | 72
PaO2 62 mmHg | 72
HCO3 29 mmol / L | 72
SpO2 93% | 72
CPAP 10 cm H2O | 72
furosemide 40 mg | 72
oxygenation improved | 72
furosemide 20 mg | 96
oxygen weaned off | 144
discharged | 168
follow-up at 3 months | 2160
skin grafting | 2160
no general anesthesia-related complications | 2160