72 years old | 0
    woman | 0
    decreased consciousness level | 0
    stupor status | 0
    elective left internal carotid artery stenting | -72
    transient ischemic attack | -72
    diabetes mellitus | 0
    hypertension | 0
    ischemic heart disease | 0
    aspirin | 0
    clopidogrel | 0
    statins | 0
    amlodipine | 0
    valsartan | 0
    antidiabetics | 0
    sudden fall in consciousness level | -72
    right hemiplegia (1/5–2/5) | 0
    brain computed tomography scan without contrast | 0
    ruled out hemorrhagic stroke | 0
    Doppler sonography on carotid arteries | 0
    totally occluded left internal carotid artery | 0
    emergent left internal carotid artery catheterization | 0
    unfractionated heparin (5000 units) injection | 0
    carotid artery wired through thrombosis | 0
    thrombosuction | 0
    alteplase (30 mg) injection | 0
    carotid stent thrombosis reoccurrence | 0
    second thrombosuction | 0
    carotid filtering for distal protection | 0
    second carotid stenting procedure | 0
    edge dissection | 0
    stent malposition | 0
    iatrogenic edge dissection | 0
    third left internal carotid artery stenting | 0
    postdilation with noncompliant balloon | 0
    patency of left internal carotid artery flow | 0
    M2 branch occlusion | 0
    transfer to intensive care unit | 0
    intravenous nitroglycerin | 0
    systolic blood pressure maintained between 120 mmHg and 130 mmHg | 0
    control brain computed tomography scan | 48
    massive infarction in middle cerebral artery area | 48
    sepsis | 96
    ventilator-associated pneumonia | 96
    disseminated intravascular coagulation | 96
    expired | 96
    no previous coronary stenting | 0
    resided in rural area | 0
    considerable distance from nearest hospital | 0
    no vascular surgeon available | 0
    high glucose levels at admission | 0
    suspected hypercoagulable state | 0
    resistance to clopidogrel | 0
    noncompliance | 0
    under-expansion stent use | 0
    oversized stent use | 0
    unavailability of appropriate carotid stent | 0
    lack of proximal protection | 0
    no thrombectomy facilities for cerebral arteries | 0
    consultation with neuro-intervention expert by phone | 0
    transferred to catheterization laboratory | 0
    angiography view confirmed carotid stent thrombosis | 0
    total cut off in left internal carotid artery | 0
    blood flow became normal | 0
    edge dissection at distal border of second stent | 0
    stent deployment on overlapping site | 0
    M1 and M3 branches normal | 0
    discharge after first procedure | 24
    complications at home | -72
    no history of previous coronary stenting | 0
    emergent procedure | 0
    dual antiplatelet therapy | 0
    long lesion development in artery | 0
    hypercoagulable state | 0
    dual-layer stent use | 0
    multiple stent use | 0
    bailout procedures | 0
    stent thrombosis | 0
    acute carotid stent thrombosis | 0
    subacute carotid stent thrombosis | 0
    early stent thrombosis | 0
    repeated early stent thrombosis | 0
    carotid stent thrombosis classification | 0
    stent thrombosis risk factors | 0
    patient-related risk factors | 0
    technical risk factors | 0
    early diagnosis | 0
    prompt revascularization | 0
    thromboaspiration | 0
    thrombectomy | 0
    thrombolytic therapy | 0
    mechanical thrombectomy | 0
    intravenous abciximab | 0
    recombinant tissue plasminogen activator | 0
    percutaneous approach | 0
    facilitated thrombolysis | 0
    aspiration thrombectomy | 0
    angioplasty | 0
    adjuvant therapy | 0
    blood sugar control | 0
    clopidogrel (150 mg) administration | 0
    information about compliance | 0
    well-equipped intensive care unit | 0
    prolonged hospital stay | 0
    P2Y12 platelet function tests | 0
    high-risk patients | 0
    hypercoagulable state evaluation | 0
    elective procedures postponed | 0
    carotid artery stent thrombosis prevention | 0
    carotid artery stenting complications | 0
    carotid endarterectomy complications | 0
    carotid stent thrombosis management | 0
    carotid stent thrombosis treatment strategies | 0
    carotid stent thrombosis incidence | 0
    carotid stent thrombosis mortality rate | 0
    carotid stent thrombosis long-term follow-up | 0
    carotid stent thrombosis differential diagnosis | 0
    carotid stent thrombosis causes | 0
    carotid stent thrombosis risk factors | 0
    carotid stent thrombosis recurrence | 0
    carotid stent thrombosis classification | 0
    carotid stent thrombosis timing | 0
    carotid stent thrombosis prevention measures | 0
    carotid stent thrombosis case presentation | 0
    carotid stent thrombosis experience sharing | 0
    carotid stent thrombosis adjuvant therapy | 0
    carotid stent thrombosis endovascular approach | 0
    carotid stent thrombosis complications | 0
    carotid stent thrombosis resolution | 0
    carotid stent thrombosis outcome | 0
    carotid stent thrombosis follow-up | 0
    carotid stent thrombosis patient care | 0
    carotid stent thrombosis ICU management | 0
    carotid stent thrombosis reperfusion-induced brain edema | 0
    carotid stent thrombosis blood pressure control | 0
    carotid stent thrombosis mortality causes | 0
    carotid stent thrombosis patient death | 0
    carotid stent thrombosis case report | 0
    carotid stent thrombosis discussion | 0
    carotid stent thrombosis recommendations | 0
    carotid stent thrombosis conclusion | 0
    