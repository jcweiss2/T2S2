43 years old | 0
male | 0
shortness of breath | -336
non-productive cough | -672
subjective fevers | -672
chills | -672
weakness | -672
malaise | -672
denied autoimmune conditions | 0
denied systemic conditions | 0
denied immune-compromising conditions | 0
denied sick contacts | 0
denied recent travel | 0
denied tuberculosis exposure | 0
denied chemical exposure | 0
denied nausea | 0
denied vomiting | 0
denied diarrhea | 0
denied muscular weakness | 0
denied neurological symptoms | 0
denied orthopnea | 0
denied paroxysmal nocturnal dyspnea | 0
able to walk five blocks without dyspnea | 0
no known drug allergies | 0
20 pack year smoking history | 0
desk job | 0
no occupational exposure to environmental pollutants | 0
admission to emergency room | 0
afebrile | 0
respiratory rate 26 breaths/min | 0
heart rate 115 beats/min | 0
room air saturation 75% | 0
blood pressure 90/60 mm Hg | 0
hyperkeratosis over index fingers | 0
thickening over metacarpophalangeal joints | 0
thickening over proximal interphalangeal joints | 0
treated with 6 L oxygen via nasal cannula | 0
received 30 cc/kg normal saline | 0
white blood cell count 25,000 units/L | 0
hemoglobin 13.5 g/dL | 0
platelet count 385 × 109/L | 0
sodium 133 mg/dL | 0
BUN 13 mg/dL | 0
creatinine 0.69 mg/dL | 0
troponin 0.09 μg/L | 0
B-type natriuretic peptide 79 pg/mL | 0
normal alkaline phosphatase | 0
normal bilirubin | 0
aspartate transaminase 259 units/L | 0
alanine transaminase 266 units/L | 0
CPK 7,500 International Units/L | 0
albumin 2.4 g/dL | 0
globulin 4.2 g/dL | 0
arterial blood gas 7.37/43/52 on 6 L oxygen | 0
lactic acid 2.4 mg/dL | 0
ESR 35 mm/h | 0
CRP 24 mg/L | 0
procalcitonin 34 ng/mL | 0
ANA speckled pattern 1:320 | 0
anti-Jo-1 antibody positive | 0
anti-CCP antibody positive 153 | 0
CT chest showing pericardial effusion 1.3 cm | 0
non-confluent ill-defined opacities in both lungs | 0
consolidations with air bronchograms in right middle lobe | 0
consolidations with air bronchograms in lower lobes | 0
atelectasis | 0
chest X-ray showing small right pleural effusion | 0
chest X-ray showing patchy right opacity | 0
ECHO showing moderate to large pericardial effusion | 0
intensive care unit transfer | 48
worsening hypoxia | 48
worsening hypotension | 48
treated with non-invasive positive pressure ventilation | 48
mechanical ventilation | 48
maximal ventilator support | 48
pulmonary artery catheterization | 48
continued decline | 48
decision for VV ECMO | 96
diagnosis of severe ARDS | 96
radiographic findings suspicious for acute interstitial pneumonia | 0
negative bronchoscopic serology | 0
negative viral serology | 0
negative fungal serology | 0
negative bacterial serology | 0
negative mycobacterial serology | 0
treated with vancomycin | 0
treated with zosyn | 0
treated with azithromycin | 0
mechanic's hands | 0
non-specific interstitial pneumonia | 0
ILD | 0
elevated CK | 0
positive anti-Jo-1 | 0
suspicion of AS | 0
treated with methylprednisolone 1 g daily for 3 days | 0
treated with methylprednisolone 125 mg four times daily for 4 days | 0
treated with methylprednisolone 60 mg four times daily for 4 days | 0
prednisone 40 mg daily at discharge | 0
minimal vasopressor requirements | 0
follow-up ECHO showing worsening pericardial effusion | 0
pericardial window | 0
fluid analysis negative for infection | 0
discharge surveillance ECHO showing no fluid re-accumulation | 0
non-oliguric renal failure | 0
acute tubular necrosis | 0
hypotension contributing to renal failure | 0
sepsis contributing to renal failure | 0
rhabdomyolysis not contributing | 0
CPK peak 7,500 International Units/L | 0
upper gastrointestinal bleed | 0
erosive gastritis | 0
managed with proton pump inhibitors | 0
improvement in respiratory status | 0
improvement in cardiovascular status | 0
improvement in renal status | 0
decannulated from ECMO | 96
transition to mechanical ventilation | 96
extubated | 96
improved clinical dyspnea | 96
discharged home | 96
instructed to wean steroids | 96
follow-up with rheumatology | 96
20 pack year smoking history |,0
