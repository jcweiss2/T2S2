70 years old | 0
female | 0
admitted to the hospital | 0
increasing abdominal pain | -72
chronic obstructive pulmonary disease (COPD) | 0
smoking | 0
hypertension | 0
dyslipidemia | 0
osteoporosis | 0
appendectomy | -0 (assuming it happened long before admission)
left partial mastectomy for breast cancer | -0 (assuming it happened 13 years prior)
right femoral hernia repair | -8760 (assuming it happened 1 year prior)
ruptured abdominal aortic aneurysm (AAA) | 0
infra-renal aortic prosthesis | 0
ligation of inferior mesenteric artery | 0
bilateral iliac thrombosis | 2
aorto-bifemoral bypass | 2
NSTEMI | 24
coronary angiography | 24
non-revascularizable occluded circumflex artery | 24
medical treatment | 24
right brachial artery thrombosis | 48
right brachial embolectomy | 48
post-operative ileus | 48
diffuse abdominal pain | 576
leukocytosis | 576
CT of abdomen | 576
air in the left retroperitoneum | 576
possible free air above the bladder | 576
descending colon wall thickening | 576
contrast extravasation | 576
left colic perforation | 576
ischemic colitis | 576
exploratory laparotomy | 600
ischemia of small bowel | 600
ischemia of descending and sigmoid colon | 600
ischemia of rectum | 600
resection of small bowel | 600
primary anastomosis | 600
left colectomy | 600
sigmoidectomy | 600
proctectomy | 600
transverse terminal colostomy | 600
Jackson-Pratt (JP) drains | 600
exacerbated COPD | 744
volume overload | 744
failed extubations | 744
infarction of inferior pole of spleen | 888
left renal artery thrombosis | 888
non-enhancing left kidney | 888
possible air bubbles in peri-renal tissue | 888
intra-abdominal fluid collections | 888
laparotomy | 912
necrosis of inferior pole of spleen | 912
necrosis of left kidney | 912
splenectomy | 912
left nephrectomy | 912
terminal transverse colostomy | 912
percutaneous feeding tube | 912
Pseudomonas aeruginosa | 912
piperacillin-tazobactam | 912
fungal infection | 936
voriconazole | 936
sepsis | 960
respiratory failure | 960
acute kidney injury | 960
diffuse non-peritonitic abdominal pain | 960
enteric feeding formula | 960
perforated small bowel | 960
anastomotic leak | 960
Mucor sp. | 984
liposomal amphotericin B | 984
comfort measures | 1008
death | 1012