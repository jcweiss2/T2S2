61 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
non-smoking | 0 | 0 | Factual
hypertension | -672 | 0 | Factual
chronic cough | -168 | 0 | Factual
dyspnea | -168 | 0 | Factual
weight loss | -168 | 0 | Factual
nausea | -72 | 0 | Factual
vomiting | -72 | 0 | Factual
cachexia | 0 | 0 | Factual
scleral icterus | 0 | 0 | Factual
jaundice | 0 | 0 | Factual
dry mucous membranes | 0 | 0 | Factual
normal bowel sounds | 0 | 0 | Factual
no pain | 0 | 0 | Factual
no distension | 0 | 0 | Factual
no organomegaly | 0 | 0 | Factual
decreased breath sounds | 0 | 0 | Factual
tachycardia | 0 | 0 | Factual
hypotension | 0 | 0 | Factual
hyponatremia | 0 | 0 | Factual
elevated alkaline phosphatase | 0 | 0 | Factual
elevated total bilirubin | 0 | 0 | Factual
elevated aspartate aminotransferase | 0 | 0 | Factual
elevated alanine aminotransferase | 0 | 0 | Factual
pulmonary parenchymal nodules | 0 | 0 | Factual
lung mass | 0 | 0 | Factual
pleural effusion | 0 | 0 | Factual
dilated common bile duct | 0 | 0 | Factual
distended gall bladder | 0 | 0 | Factual
pancreatic head mass | 0 | 0 | Factual
biliary obstruction | 0 | 0 | Factual
biopsy of lung mass | 24 | 24 | Factual
biliary stenting | 24 | 24 | Factual
lung adenocarcinoma | 0 | 0 | Factual
metastases to brain | 0 | 0 | Factual
radiation therapy | 48 | 168 | Factual
adjunctive chemotherapy | 48 | 168 | Factual
carboplatin | 48 | 168 | Factual
pemetrexed | 48 | 168 | Factual
pembrolizumab | 48 | 168 | Factual
whole brain radiation | 72 | 168 | Factual
severe pneumonia | 168 | 168 | Factual
sepsis | 168 | 168 | Factual
death | 168 | 168 | Factual