15-month-old male | 0
Wiskott–Aldrich syndrome | 0
thrombocytopenia | 0
eczema | 0
immunodeficiency | 0
mutations in the WAS gene | 0
no protein expression of WAS | 0
four-base-pair deletion in intron-8 | 0
diagnosis of WAS | 0
admitted to the hospital for HSCT | 0
thrombocytopenic after birth | -10920
genetic studies | -10920
human leukocyte antigen (HLA) unmatched sister | -10920
required unrelated donor | -10920
platelets transfusions (two) | -8760
worsening petechiae | -8760
intermittent hematochezia | -8760
intravenous immunoglobulin therapy monthly | -10920
prophylactic trimethoprim-sulfamethoxazole | -10920
no significant history of infection before transplantation | -10920
admitted at 13 months of age | -240
preconditioning therapy for HSCT | -240
fludarabine | -240
melphalan | -240
thiotepa | -240
antithymocyte globulin | -240
bone marrow completely ablated | -240
Escherichia coli sepsis | -240
started on antibiotics | -240
hemodynamic instability | -192
admitted to the Pediatric Intensive Care Unit on HD#8 | -192
refractory septic shock | -192
intubation | -192
volume resuscitation | -192
inotropic support | -192
venoarterial ECMO on HD#9 | -168
cannulated with 14-French arterial cannula in right carotid artery | -168
cannulated with 14-French venous cannula in right internal jugular vein | -168
echocardiogram after cannulation | -168
severely diminished left ventricular function | -168
left atrial hypertension | -168
balloon atrial septostomy | -168
inotropic support weaned off within 72 hours | -168
continuous renal replacement therapy (CRRT) on HD#10 | -144
fluid overload | -144
unrelated HLA donor stem cell transplant through ECMO circuit on HD#10 | -144
received ABO-mismatched cord blood transplant | -144
CD34+ count of 4.7 × 10^5/kg | -144
total nucleated cell count of 1.12 × 10^8/kg | -144
cord blood infused on arterial side | -144
left-sided paralysis on HD#13 | -120
emergent head computed tomography | -120
acute intraparenchymal hemorrhages in right posterior temporal lobe | -120
acute intraparenchymal hemorrhages in left occipital lobe | -120
4 mm right to left midline shift | -120
decannulated from ECMO | -120
brain magnetic resonance on HD#16 | -96
stable right greater than left occipital lobe hematomas | -96
watershed infarction along right parasagittal centrum semiovale | -96
signs of engraftment on HD#22 (day +12) | 288
extubated on HD#36 | 432
fluorescence in situ hybridization XY showed 100% donor cells on HD#40 (day +30) | 720
transitioned to peritoneal dialysis on HD#57 | 1248
discharged to the floor on HD#69 | 1656
neurologic examination improvement | 1656
renal function improvement | 1656
discharged home on HD#94 | 2256
peritoneal catheter removed 10 days after discharge | 2256 + 240 = 2496
recovered from neurologic injury with no sequelae | 8760
remained asymptomatic from WAS standpoint | 8760
complete donor engraftment | 8760
no evidence of mixed chimerism | 8760
no signs of chronic graft versus host disease | 8760
white blood count and absolute neutrophil count monitored during hospital course | various
eczema |+0
peritoneal catheter removed 10 days after discharge | 2496
