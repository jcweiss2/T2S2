87 years old | 0
female | 0
TAVI performed | -2160
severe symptomatic aortic stenosis | -2160
non-insulin dependent diabetes mellitus | 0
chronic hypertension | 0
coronary artery disease | 0
gastro-oesophageal reflux disease | 0
osteoarthritis | 0
right total knee replacement | 0
cervical spine fixation | 0
fever | -720
convulsive seizure | -720
acute ischaemic stroke | -720
decreased level of consciousness | -720
dysarthria | -720
admitted to ICU | -720
TTE negative for vegetations | -720
CT head showed acute right cerebellar infarction | -720
blood cultures negative | -720
empiric antibiotics | -720
fever curve reduced | -720
transferred to tertiary hospital | 0
blood pressure 105/49 mmHg | 0
sinus tachycardia | 0
pulse 108 | 0
temperature 38°C | 0
oxygen saturation 96% | 0
soft systolic murmur | 0
crackles in dependent lung regions | 0
GCS 9/15 | 0
pseudobulbar signs | 0
inability to swallow | 0
dysarthria | 0
bilateral motor weakness | 0
right upper extremity MRC 1/5 | 0
left upper extremity MRC 3/5 | 0
decreased lower extremity tone | 0
bilateral extensor plantar reflexes | 0
no peripheral stigmata of endocarditis | 0
respiratory distress | 0
intubated | 0
hypoxaemia | 0
bilateral lower lobe opacities | 0
aspiration pneumonia | 0
normochromic normocytic anaemia | 0
haemoglobin 10 g/dL | 0
normal leucocyte count | 0
thrombocytopenia | 0
platelet count 71 × 10³/µL |=
CRP 104 mg/L | 0
low albumin 21.1 g/L | 0
normal liver function | 0
normal renal function | 0
blood cultures grew Corynebacterium | 0
TTE repeated | 0
no vegetations | 0
no para-valvular leak | 0
LVEF 60% | 0
subacute right cerebellar infarct | 0
TOE performed | 24
large vegetation 1.3×0.6 cm | 24
aortic root pseudoaneurysm | 24
aortic root abscess | 24
CT angiography | 48
pseudoaneurysm 2.5×2.0 cm | 48
suspected infection | 48
infective endocarditis diagnosed | 24
prosthetic valve endocarditis | 24
hospital acquired pneumonia | 0
meropenem/levofloxacin | 0
vancomycin | 0
CRP decreased | 144
fever persisted | 0
transferred to France | 192
blood cultures grew Corynebacterium amycolatum | 192
aortic root and valve replacement | 312
homograft implanted | 312
vegetations cultures grew Corynebacterium | 312
post-operative chylothorax | 312
septic shock | 312
ventilator associated pneumonia | 312
prolonged mechanical ventilation | 312
tracheostomy | 312
daptomycin | 312
rifampin | 312
transferred back to ICU | 432
GCS 6/15 | 432
lumbar puncture | 432
slight protein elevation | 432
MRI head confirmed previous findings | 432
cervical MRI showed degenerative disease | 432
EEG no seizures | 432
axonal neuropathy | 432
muscle weakness | 432
critical illness polyneuropathy | 432
critical illness myopathy | 432
intermittent consciousness changes | 432
recurrent CVAs | 432
sepsis | 432
improved consciousness | 432
rifampin discontinued | 432
drug rash | 432
elevated liver enzymes | 432
meropenem | 432
daptomycin continued | 432
ventilator associated pneumonia | 432
catheter-related infection | 432
urinary tract infection | 432
PEG placement | 432
nutrition optimized | 432
physiotherapy | 432
infection control | 432
weaned off ventilator | 432
tracheostomy in situ | 432
tolerated pureed diet | 432
TTE showed mild aortic regurgitation | 432
preserved LVEF | 432
CRP 4.64 mg/L | 432
discharged home | 1080
home health nurse | 1080
afebrile | 1080
able to follow commands | 1080
interacts with family | 1080
