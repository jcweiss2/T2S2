74 years old | 0
    woman | 0
    schizophrenia | 0
    referred to hospital with high-grade fever | 0
    high-grade fever | 0
    unaware of febrile status prior to admission | -72
    no chest pain | 0
    no cough | 0
    no dyspnea | 0
    no palpitation | 0
    no urinary complaints | 0
    no bowel complaints | 0
    no history of tuberculosis | 0
    no history of malignancy | 0
    no previous hospital admissions | 0
    denied smoking | 0
    denied drinking alcohol | 0
    denied illicit drug use | 0
    no recent travel history | 0
    temperature 39.1°C | 0
    pulse rate 110 beats/min | 0
    blood pressure 100/60 mmHg | 0
    respiratory rate 24/min | 0
    oxygen saturation 99% | 0
    Glasgow Coma Scale E4V4M6 | 0
    non-tender mass in lower right back | -720
    cardiovascular examination unremarkable | 0
    abdominal examination unremarkable |* 0
    leukocytosis 23,300 cells/mm3 | 0
    polymorphic neutrophil predominance 93.8% | 0
    hemoglobin 8.6 g/dL | 0
    platelet count 339,000/mm3 | 0
    CPK 125 IU/L | 0
    blood urea nitrogen 23.3 mg/dl | 0
    creatinine 0.97 mg/dl | 0
    CRP 15.26 mg/dl | 0
    blood sugar 116 mg/dl | 0
    HbA1c 5.4% | 0
    HIV test negative | 0
    urine protein +/- | 0
    urine nitrite 1+ | 0
    urine leukocyte 2+ | 0
    urine glucose negative | 0
    urine occult blood negative | 0
    urine ketones negative | 0
    subcutaneous abscess suspected | 0
    ultrasound examination | 0
    low echoic mass reaching right kidney | 0
    CT large mass right retroperitoneum | 0
    abscess extended into subcutaneous space | 0
    staghorn calculus | 0
    surgical drainage | 0
    admitted to intensive care unit | 0
    septic shock | 0
    M. morganii detected in abscess fluid | 0
    M. morganii detected in urine culture | 0
    blood cultures negative | 0
    repeat CT with contrast | 0
    right renal abscess | 0
    staghorn calculus | 0
    retroperitoneum abscess improvement | 0
    iliopsoas abscess from renal abscess | 0
    urinary tract infection uncontrolled | 0
    M. morganii sensitive to piperacillin/tazobactam | 0
    M. morganii sensitive to meropenem | 0
    M. morganii sensitive to cefmetazole | 0
    M. morganii sensitive to gentamycin | 0
    M. morganii sensitive to amikacin | 0
    M. morganii sensitive to levofloxacin | 0
    M. morganii resistant to cephalosporins | 0
    M. morganii resistant to ampicillin | 0
    meropenem administered | 0
    salvage nephrectomy | 0
    post-operative recovery exceptional | 0
    intravenous meropenem 0.5g every 8h for 2 weeks | 0
    responded well to initial treatment | 0
    oral levofloxacin 250mg for 4 weeks | 0
    discharged to nursing home | 672
    <|eot_id|>
    