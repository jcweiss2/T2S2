28 years old | 0
female | 0
8 weeks pregnant | 0
acute severe asthma | -10
short non-infective prodrome | -10
hypoxic cardiac arrest | -10
ventricular fibrillation | -10
resuscitation to sinus tachycardia | -10
endotracheal intubation | -10
therapeutic cooling to 33°C | 0
salbutamol | 0
ipratropium | 0
aminophylline | 0
hydrocortisone | 0
magnesium | 0
ketamine | 0
inhalation anesthesia with 1 MAC isoflurane | 0
severe hypercapnic acidosis | 0
neuromuscular blockade | 0
inadequate minute ventilation | 0
generalised status myoclonus | 48
absent motor response to painful stimulus | 96
preserved pupillary reflexes | 96
preserved corneal reflexes | 96
preserved cough reflexes | 96
preserved gag reflexes | 96
spontaneously breathing | 96
severe GSM | 96
refractory to three antiepileptic medications | 96
generalised periodic discharges | 96
no discernable background rhythm | 96
reversible causes of coma eliminated | 96
no agreement about neurological outcome | 192
plasma neuron-specific enolase | 240
somatosensory-evoked potential | 240
brain magnetic resonance imaging | 240
bilateral basal ganglia and frontoparietal cortex infarction | 240
medical consensus regarding poor prognosis | 240
extubated | 264
died | 288