40 days old | 0
    male | 0
    neonate | 0
    twin | 0
    born of normal vaginal delivery | 0
    gestation 36 weeks | 0
    referred for management of tricuspid valve mass | 0
    admitted to neonatal intensive care unit | -480
    neonatal seizures | -480
    necrotizing enterocolitis | -480
    blood cultures | -480
    negative blood cultures | -480
    anti-convulsants | -480
    intravenous antibiotics | -480
    piperacillin tazobactam | -480
    amikacin | -480
    peripheral venous access | -480
    no invasive procedures | -480
    echocardiography | -480
    no structural heart disease | -480
    tricuspid mass | -480
    referred to our center | 0
    admission | 0
    not febrile | 0
    deeply icteric | 0
    no focal neurologic deficits | 0
    no clinical heart failure | 0
    normal cardiovascular examination | 0
    small cephalhematoma | 0
    computed tomography brain scan | 0
    petechial hemorrhages | 0
    no space occupying lesions | 0
    echocardiography | 0
    vegetation attached to tricuspid valve | 0
    Doppler examination | 0
    mean tricuspid inflow gradient 5 mmHg | 0
    blood cultures collected | 0
    blood cultures positive | 0
    fungal cultures | 0
    white yeast-like colonies | 0
    K. ohmeri identified | 0
    Gram staining | 0
    oval budding yeast cells | 0
    antifungal susceptibility test | 0
    Amphotericin <0.25 mcg/L | 0
    Fluconazole 2 mcg/L | 0
    Voriconazole <0.12 mcg/L | 0
    Flucytosine <1 mcg/L | 0
    intravenous amphotericin B | 0
    packed cell transfusion | 0
    planned surgical removal | 0
    hemodynamic compromise | 48
    fungal septicemia | 48
    death | 48

    40 days old | 0
    male | 0
    neonate | 0
    twin | 0
    born of normal vaginal delivery | 0
    gestation 36 weeks | 0
    referred for management of tricuspid valve mass | 0
    admitted to neonatal intensive care unit | -480
    neonatal seizures | -480
    necrotizing enterocolitis | -480
    blood cultures | -480
    negative blood cultures | -480
    anti-convulsants | -480
    intravenous antibiotics | -480
    piperacillin tazobactam | -480
    amikacin | -480
    peripheral venous access | -480
    no invasive procedures | -480
    echocardiography | -480
    no structural heart disease | -480
    tricuspid mass | -480
    referred to our center | 0
    admission | 0
    not febrile | 0
    deeply icteric | 0
    no focal neurologic deficits | 0
    no clinical heart failure | 0
    normal cardiovascular examination | 0
    small cephalhematoma | 0
    computed tomography brain scan | 0
    petechial hemorrhages | 0
    no space occupying lesions | 0
    echocardiography | 0
    vegetation attached to tricuspid valve | 0
    Doppler examination | 0
    mean tricuspid inflow gradient 5 mmHg | 0
    blood cultures collected | 0
    blood cultures positive | 0
    fungal cultures | 0
    white yeast-like colonies | 0
    K. ohmeri identified | 0
    Gram staining | 0
    oval budding yeast cells | 0
    antifungal susceptibility test |;