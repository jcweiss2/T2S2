83 years old | 0
female | 0
admitted to the emergency department | 0
fever | 0
vomiting | 0
diffuse abdominal pain | 0
abdominal pain in the right upper quadrant | 0
rheumatoid arthritis | -6720
atrial fibrillation | -6720
asthma | -6720
cerebrovascular disease | -6720
hysterectomy | -6720
intestinal obstruction | -6720
oral steroids | -6720
methotrexate | -6720
clopidogrel | -6720
omeprazole | -6720
paracetamol | -6720
hormone replacement therapy | -6720
nonsteroidal anti-inflammatory drug | -6720
tenderness in the right upper quadrant | 0
guarding in the right upper quadrant | 0
temperature 37.6°C | 0
leukocytosis | 0
C-reactive protein 306 mg/L | 0
abnormal liver enzymes | 0
ALT 137 U/L | 0
AST 97 U/L | 0
GGT 220 U/L | 0
total blood bilirubin level 30.5 mmol/L | 0
plain abdominal radiography | 0
circular gas pattern in the area of the gallbladder | 0
emphysematous cholecystitis | 0
computed tomography | 0
gas in the gallbladder wall | 0
gas-fluid level within the organ | 0
emergency laparoscopic cholecystectomy | 0
extensive inflammation and necrosis of the gallbladder | 0
gallbladder punctured | 0
intraoperative cholangiography | 0
biliary obstruction excluded | 0
cholecystectomy | 0
bubbling from the gallbladder wall | 0
resection of the gallbladder completed | 0
extensive laparoscopic abdominal lavage | 0
drainage | 0
intravenous antibiotic therapy | 0
discharged | 264
pathological analysis of the resected gallbladder | 264
full-thickness infarctive necrosis | 264
abscess | 264
single small calculus at the gallbladder neck | 264
microbiological analysis of the pus | 264
Clostridium perfringens | 264