18 years old | 0
male | 0
admitted to the hospital | 0
new-onset headache | -72
blurred vision | -72
kidney transplant | -672
end-stage kidney disease | -672
immunousuppression | -672
mycofenolate sodium | -672
methylprednisolone | -672
estimated glomerular filtration rate (eGFR) | -672
proteinuria | -672
chronic kidney transplant disease stage 3bA1 | -672
status post vascular rejection | -672
chronic calcineurin-inhibitor toxicity | -672
contrast-enhancing intracerebral lesions | -672
perifocal edema | -672
methylprednisolone therapy | -672
dexamethasone | -672
brain biopsy | -672
cerebral PTLD | -672
diffuse large B-cell lymphoma | -672
positive for Ebstein-Barr virus | -672
CT scan of the thorax | -672
abdomen sonography | -672
bone marrow biopsy | -672
high-dose cytarabin | -672
Rituximab | -672
MRI scan | -672
complete remission of PTLD | -672
impairment of the transplant function | -672
eGFR 25.4 mL/min/1.73 qm | -672
CKD-EPI equation | -672
cytomegalovirus (CMV) reactivated | -672
pneumocystis jirovecii pneumonia | -672
Rituximab only | -672
antiviral and antibiotic therapy | -672
mycofenolate sodium tapered | -672
leukopenia | -672
infections | -672
generalized seizure | -672
cerebral MRI scan | -672
recurrence of PTLD | -672
intravenous HDMTX | -672
Leukovorine | -672
Rituximab | -672
vigorous hydration | -672
high-flux hemodialysis (HFHD) | -672
MTX-level in serum | -672
leucocytes | -672
acute kidney failure | -672
sepsis | -672
intensive care unit | -672
invasive ventilation | -672
CMV- and E.coli pneumonia | -672
acute kidney transplant failure | -672
follow up cerebral MRI scan | -672
small regredience of PTXLD | -672
cerebral radiation | -672
no relevant response of the disease | -672
elected radiotherapy | -672
dialysis parameters | -672
MTX-level measurements | -672
MTX administration | -672
Gambro machine AK 200 | -672
high-flux dialyser (Polyflux 170H) | -672
dialysate SelectBag One AX 450 G | -672
potassium 4 mmol/L | -672
calcium 1.50 mmol/L | -672
glucose 1.0 g/L | -672
dialysate flow | -672
blood flow | -672
unfractionated heparin | -672
dialysis sessions | -672
MTX clearance | -672
fluorescence polarization immunoassay | -672
TDx analyser | -672
MTX toxicity | -672
renal impairment | -672
kidney function | -672
acute kidney failure | -672
bone marrow toxicity | -672
severe CMV- and E.coli pneumonia | -672
sepsis | -672
acute kidney transplant failure | -672
MTX elimination | -672
HFHD | -672
vigorous hydration | -672
alkalinization of the urine | -672
leucovorin rescue | -672
MTX clearance | -672
renal replacement therapy | -672
hemodialysis | -672
hemodiafiltration | -672
Charcoal hemoperfusion/hemofiltration | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDMTX | -672
MTX clearance | -672
HFHD | -672
MTX elimination | -672
renal function | -672
kidney function | -672
acute kidney failure | -672
nephrotoxicity | -672
hematological toxicities | -672
leucopenia | -672
anemia | -672
thrombocytes | -672
infection | -672
CMV-colonization | -672
CMV-activation | -672
posttransplant immunosuppressive therapy | -672
impaired kidney function | -672
rituximab | -672
HDM