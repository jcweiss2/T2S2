68 years old | 0
male | 0
admitted to the hospital | 0
abdominal pain | -168
clear breath sounds | 0
no dry and wet rales | 0
abdomen soft and flat | 0
no tenderness | 0
no rebound tenderness | 0
old surgical scar | 0
no swelling of the liver | 0
no swelling of the spleen | 0
chronic inflammation of the lungs | 0
thickening of the lower esophageal wall | 0
enlarged mediastinal lymph nodes | 0
no other organ metastases | 0
malignant tumor of the esophageal mucosa | 0
squamous cell carcinoma | 0
ulceration | 0
radical surgery for esophageal carcinoma | 264
postoperative histopathology | 264
pathological mitosis | 264
tumor infiltration | 264
cancer metastasis | 264
no nerve invasion | 264
immunohistochemistry | 264
positive expression of p40 | 264
positive expression of CK5/6 | 264
positive expression of EGFR | 264
positive expression of p53 | 264
negative expression of CK7 | 264
negative expression of p16 | 264
negative expression of CD34 | 264
negative expression of S-100 | 264
stage IIIa moderately differentiated ulcerative esophageal squamous cell carcinoma | 264
high fever | 288
dyspnea | 288
blood pressure 80/50 mmHg | 288
neck wound clean and dry | 288
white blood cells 34.38 × 10^9/L | 288
neutrophils 95.7% | 288
C-reactive protein 207.26 mg/L | 288
procalcitonin >100 ng/mL | 288
urinary leukocytes 62.20/µL | 288
leukocytes per high-power field 11.20 | 288
increased exudative lesions in both lungs | 288
postoperative changes in the esophagus | 288
sepsis | 288
meropenem administration | 288
blood cultures suggested growth of E. fergusonii | 336
E. fergusonii identified | 336
drug sensitivity testing | 336
E. fergusonii sensitive to cefuroxime | 336
E. fergusonii sensitive to cefuroxime axetil | 336
E. fergusonii sensitive to ceftazidime | 336
E. fergusonii sensitive to ceftriaxone | 336
E. fergusonii sensitive to cefepime | 336
E. fergusonii sensitive to cefoxitin | 336
E. fergusonii sensitive to amoxicillin–clavulanic acid | 336
E. fergusonii sensitive to piperacillin–tazobactam | 336
E. fergusonii sensitive to cefoperazone–sulbactam | 336
E. fergusonii sensitive to imipenem | 336
E. fergusonii sensitive to ertapenem | 336
E. fergusonii sensitive to amikacin | 336
E. fergusonii sensitive to tigecycline | 336
E. fergusonii sensitive to cotrimoxazole | 336
fever subsided | 432
clinical indicators improved | 432
repeat blood culture negative | 648
patient recovered | 720
discharged from the hospital | 720
follow-up | 1440
no specific discomfort | 1440
postoperative adjuvant radiation therapy | 1440