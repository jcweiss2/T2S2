49 years old | 0
male | 0
admitted to the hospital | 0
fever | -96
pyrexia | -96
cough | -96
shortness of breath | -96
Covid-19 positive | -96
diabetes | -8760
sliding-scale insulin | -8760
HbA1c 12.3% | 0
fasting blood sugar 250 mg/dL | 0
post prandial blood sugar 350 mg/dL | 0
interleukin 637.93 pg/mL | 0
C-reactive protein 17.84 mg/L | 0
D-Dimer 460 ng/mL | 0
creatinine 0.8 mg/dl | 0
lymphocyte 9.5% | 0
neutrophil 84% | 0
injection Remdesivir IV | 0
methylprednisolone IV | 0
intensive care unit | 0
recovered from Covid | 240
bilateral pneumonia | 240
swelling and discomfort in the left eye | 240
malaise | 240
proptosis | 240
chemosis | 240
periorbital cellulitis | 240
partial ophthalmoplegia | 240
visual acuity 6/6 | 240
magnetic resonance imaging | 240
mucormycosis of the rhino-orbital-cerebral extension | 240
bone erosion | 240
surgery scheduled for FESS and debridement | 240
general anesthesia | 240
glycopyrrolate 0.2 mg | 240
fentanyl 150 mg | 240
preoxygenation with 100% oxygen | 240
propofol 100 mg | 240
rapid sequence induction | 240
scoline 2 mg/kg | 240
intubation | 240
xylocard 1.5 mg/kg | 240
thoracic pack | 240
postintubation pulse oximetry | 240
five-lead ECG | 240
NIBP | 240
end-tidal carbon dioxide | 240
temperature | 240
urine output monitoring | 240
oxygen | 240
nitrous | 240
sevoflurane 1% | 240
vecuronium 0.1 mg/kg | 240
elective ventilation | 240
discharged | 720