51 year old | 0
male | 0
admitted to ICU | 0
bilateral nephrectomy | 0
invasive urothelial cancer | 0
hemodynamic monitoring | 0
uneventful first 24 hours | 0
high fever | 48
distributive shock pattern | 48
elevated C-reactive protein | 48
septic shock consideration | 48
cultures realized | 48
CT scan abdomen | 48
no abscess | 48
septic shock patient | 48
no problematic source | 48
antibiotics started | 48
Tazocin 4 g TDS | 48
amikacin 25 mg/kg | 48
resuscitated | 48
adequate volume loading | 48
noradrenaline infusion | 48
0.1 mcg/kg/min | 48
continuous veno-venous hemofiltration | 48
deteriorated after 72 hours | 72
increased noradrenaline infusion | 72
1.9 mcg/kg/min | 72
received 5 L fluids | 72
high fever 39.5°C | 72
enlarging antimicrobial coverage consideration | 72
drug-resistant gram-negative bacteria coverage | 72
fungal infections coverage | 72
cultures negative | 72
senior nephrologist-intensivist consulted | 72
bilateral adrenal glands resection consideration | 72
Addison’s disease diagnosis | 72
hydrocortisone 100 mg bolus | 72
hydrocortisone 300 mg infusion | 72
condition normalized | 72
antimicrobials stopped | 72
