54 years old|0
    African-American woman|0
    past medical history of deep vein thrombosis|-672
    past medical history of remote provoked pulmonary embolism|-672
    presented to the Emergency Department|0
    fevers|-336
    progressive shortness of breath|-336
    cough|-336
    >2 weeks duration of fevers|-336
    >2 weeks duration of progressive shortness of breath|-336
    >2 weeks duration of cough|-336
    history of provoked pulmonary embolism in 2012|-40320
    anticoagulated with warfarin for 3 months after 2012|-40320
    initial presentation to the Emergency Department|0
    oxygen saturation 99% on room air|0
    blood pressure 100/70 mmHg|0
    heart rate 75 b.p.m.|0
    respiratory rate 30 breaths/min|0
    elevated D-dimer 2.86 mg/L|0
    elevated ferritin 683.2 ng/mL|0
    elevated lactate dehydrogenase 929 U/L|0
    elevated aspartate aminotransferase 190 U/L|0
    elevated alanine aminotransferase 131 U/L|0
    decreased platelet count 98|0
    decreased white blood cell count 3.9|0
    decreased absolute lymphocyte count 0.59|0
    elevated probrain natriuretic peptide 2016 pg/mL|0
    initial troponin elevation 0.100 ng/mL|0
    troponin trended down|0
    electrocardiogram showed right ventricular strain|0
    transthoracic echocardiogram revealed dilated right ventricle with McConnell’s sign|0
    computed tomography angiography of the chest|0
    large pulmonary embolism in the right main pulmonary artery|0
    additional smaller pulmonary emboli in the left upper and lower lobe|0
    computed tomography chest evidence of right heart strain|0
    scattered ground-glass opacities with rounded morphology|0
    oxygen saturation 84% on 4.5 L nasal cannula in ICU|0
    cardiovascular exam normal|0
    lungs clear to auscultation bilaterally|0
    mild respiratory distress with accessory muscle use|0
    increased oxygen supplementation|0
    hypoxic on 10 L non-rebreather|0
    intubated|0
    intubated for 14 days|0
    managed with volume control without ARDS protocol|0
    required norepinephrine intermittently|0
    transthoracic echocardiogram confirmed severe right ventricular dilatation|24
    transthoracic echocardiogram confirmed moderate pulmonary hypertension|24
    right ventricular thrombus 1.3 cm × 1.3 cm|24
    thrombus on anterior tricuspid leaflet|24
    thrombus in dilated inferior vena cava 1.4 cm × 1.9 cm|24
    positive COVID-19 PCR on day 4|96
    started on azithromycin 500 mg for 1 day|0
    transitioned to doxycycline on day 1|24
    started on hydroxychloroquine on day 1|24
    hydroxychloroquine loading dose 400 mg twice a day on day 1|24
    hydroxychloroquine 200 mg twice a day for 4 days|24
    doxycycline 100 mg twice a day for 5 days|24
    treated with intravenous heparin on day 1|24
    transitioned to enoxaparin 80 mg twice a day on day 14|336
    catheter-directed thrombolysis discussed|24
    intravenous anticoagulation not pursued|24
    screened for thrombosis using Doppler imaging|336
    right popliteal deep vein thrombosis|336
    weaned down to room air|336
    evaluated by physical medicine and rehabilitation|336
    inpatient rehabilitation therapy|336
    hoarse voice|336
    D-dimer remained elevated at 2.35 mg/L on discharge|456
    discharged on therapeutic enoxaparin|456
    discharged to inpatient rehabilitation unit|456
    instructed to report to primary care physician and cardiologist|456
    no follow-up to date|456
    <|eot_id|>
    