60 years old | 0
female | 0
admitted to the hospital | 0
seizure-like activity | -120
unwitnessed fall | -120
laceration on the forehead | -120
nausea | -96
vomiting | -96
diarrhea | -96
generalized weakness | -96
severe fatigue | -96
non-specific headaches | -168
low back pain | -168
neck pain | -168
hearing loss | -168
hallucinations | -72
epilepsy | 0
chronic obstructive pulmonary disease | 0
hypertension | 0
hyperlipidemia | 0
depression | 0
anxiety | 0
migraines | 0
multiple sclerosis | 0
fever | 0
tachycardia | 0
hypertension | 0
bilateral periorbital ecchymosis | 0
forehead laceration | 0
tachycardia with regular rhythm | 0
no murmurs | 0
no rubs | 0
no gallops | 0
clear lungs | 0
fluent speech | 0
no aphasia | 0
cranial nerves II-XII intact | 0
5/5 muscle strength | 0
intact sensation | 0
normal reflexes | 0
negative Babinski sign | 0
no dysmetria | 0
no nuchal rigidity | 0
negative Kernig and Brudzinski maneuvers | 0
elevated white blood cell count | 0
elevated lactic acid | 0
low potassium | 0
low sodium | 0
elevated glucose | 0
elevated troponin | 24
ECG with sinus tachycardia | 0
ECG with non-specific ST-segment depression | 0
CT scan with small frontal scalp hematoma | 0
MRI with progressive periventricular white matter lesions | 0
blood cultures positive for yeast | 48
lumbar puncture | 48
started on amphotericin | 48
cerebrospinal fluid with low glucose | 48
cerebrospinal fluid with elevated protein | 48
cerebrospinal fluid with positive Cryptococcus antigen | 48
added flucytosine to treatment | 48
became unresponsive | 96
became hypoxic | 96
required endotracheal intubation | 96
became bradycardic | 96
cardiac arrest | 96
advance cardiac life support | 96
return of spontaneous circulation | 96
elevated troponin | 96
ECG with Q waves | 96
ECG with poor R wave progression | 96
ECG with ST-segment elevations | 96
echocardiogram with hypokinesis | 96
echocardiogram with basal hyperkinesis | 96
diagnosed with Takotsubo cardiomyopathy | 96
deteriorated clinically | 120
required increasing vasopressor support | 120
required significant ventilator support | 120
no cough reflex | 120
no corneal reflex | 120
no pharyngeal reflex | 120
transitioned to comfort care | 144
passed away | 144