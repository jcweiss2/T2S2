44 years old | 0
male | 0
Darier6White disease | -8760
symptom onset during infancy | -43800
first diagnosed in 1995 | -216576
mild acne | -43800
seborrheic distribution | -43800
summertime exacerbations | -43800
treated with systemic retinoids | -216576
multiple complications from 1995 to 2014 | -216576
sepsis episodes | -216576
Kaposi varicelliform eruption | -216576
frequent local infections | -216576
Staphylococcus aureus infections | -216576
Morganella morganii infections | -216576
atypical Mycobacterium cutaneous infection in 2005 | -131040
infections treated with antibiotics | -216576
disease peak during 2013 | -17520
widespread erythema | -17520
hypertrophic warty keratotic papules | -17520
plaques | -17520
cysts | -17520
nodules | -17520
giant comedones | -17520
severe macerations | -17520
severe fetor | -17520
leonine-like facies | -17520
diffuse palmo-plantar keratoderma | -17520
extreme cachexia | -17520
tachycardia | -17520
normal neuropsychiatric evaluation | -17520
skin biopsy findings | -17520
keratotic plugs | -17520
dyskeratosis | -17520
corps ronds | -17520
grains | -17520
suprabasal clefts | -17520
Periodic acid-Schiff staining negative | -17520
anemia | -17520
leukocytosis | -17520
hypoalbuminemia | -17520
Staphylococcus aureus skin culture | -17520
Morganella morganii skin culture | -17520
Streptococcus group G skin culture | -17520
S aureus blood culture | -17520
negative fungal infection tests | -17520
negative HIV serology | -17520
negative herpes simplex PCR | -17520
negative varicella zoster PCR | -17520
low blood iron | -17520
low folic acid | -17520
low transferrin | -17520
low vitamin D | -17520
normal immune function tests | -17520
negative genetic test for 3-base deletion | -17520
treated with broad-spectrum antibiotics | -17520
high-dose oral isotretinoin | -17520
topical keratolytic therapy | -17520
infections responded well | -17520
partial response of cutaneous disease | -17520
discharged | -17520
presented to ICU 10 months later | -240
severe sepsis | -240
severe hypoglycemia | -240
widespread erythema | -240
died 2 days after admission | 48
| Header 1 | Header 2 |
|----------|----------|
| Item 1   | Item 2   |
| Item 3   | Item 4   |
