54 years old | 0\
male | 0\
admitted to the hospital | 0\
pre-syncope | -2\
syncope | -2\
left-sided chest tightness | -2\
generalized fatigue | -672\
weight loss | -672\
diffuse erythematous rash | 0\
weight 41 kg | 0\
blood pressure 96/60 mm Hg | 0\
unremarkable cardiac examination | 0\
unremarkable respiratory examination | 0\
normal sinus rhythm | 0\
raised troponin concentration | 0\
eosinophil count 7.6 × 10^9/l | 0\
referred to cardiology | 0\
diagnosis of myocarditis | 0\
cardiac magnetic resonance imaging | 24\
eosinophilic myocarditis | 24\
coronary angiography | 24\
no evidence of coronary artery disease | 24\
skin biopsy | 24\
cardiac biopsy | 24\
edoxaban | 24\
prednisolone | 24\
discharged | 48\
missed appointment | 336\
neck swelling | 336\
admitted to hospital | 336\
eosinophil count 19.7 × 10^9 cells/l | 336\
increase dose of prednisolone | 336\
computed tomography of neck | 336\
lymphadenopathy | 336\
T-cell lymphoma | 336\
cyclophosphamide | 336\
sepsis | 360\
cholecystitis | 360\
new onset of seizures | 360\
reduction in consciousness | 360\
Glasgow Coma Scale 9/15 | 360\
head computed tomography | 360\
multiple bilateral acute infarctions | 360\
transferred to intensive care unit | 360\
history of hepatitis B | -8760\
history of asthma | -8760\
history of intravenous drug use | -8760\
history of excessive use of alcohol | -8760\
diffuse subendocardial late gadolinium enhancement | 360\
mild left ventricular systolic impairment | 360\
eczematous changes | 360\
bone marrow biopsy | 360\
no increase in eosinophils | 360\
axillary lymph node biopsy | 360\
T-cell lymphoma | 360\
infarcts involving frontal, parietal, and left temporo-occipital regions | 360\
apical tear | 360\
intramural myocardial tear | 360\
small apical cavity | 360\
mobile structures attached to dissected myocardium | 360\
diastolic flow in the apical cavity | 360\
systolic flow out of the apical cavity | 360\
cyclophosphamide therapy | 360\
partial response | 360\
reduction of eosinophil count | 360\
palliation | 432