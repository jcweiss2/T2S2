65 years old | 0\
female | 0\
liver cirrhosis | -672\
chronic hepatitis B | -672\
hepatocellular carcinoma | 0\
scheduled for left lobe hepatectomy | 0\
glycopyrrolate | 0\
propofol | 0\
rocuronium | 0\
remifentanil | 0\
sevoflurane | 0\
intubated | 0\
mechanical ventilation | 0\
electrocardiography | 0\
arterial blood pressure | 0\
central venous pressure | 0\
SpO2 | 0\
stable vital signs | 0\
sudden decrease in arterial blood pressure | 1\
tachycardia | 1\
ST elevation on EKG | 1\
resuscitation with colloid and catecholamines | 1\
intraoperative ultrasonography | 1\
massive air emboli in both heart | 1\
diagnosis of VAE and PAE | 1\
arterial blood gas analysis | 1\
catecholamine administration | 1\
systolic blood pressure and heart rate maintained | 10\
central venous pressure maintained | 10\
end-tidal carbon dioxide restored | 10\
arterial blood gas analysis | 30\
norepinephrine infusion | 30\
fluid resuscitation | 30\
air emboli in left heart disappeared | 70\
hepatectomy restarted | 70\
completion of hepatectomy | 70\
total anesthesia time | 300\
total fluid administered | 300\
total urinary output | 300\
blood loss | 300\
intensive care unit | 300\
intubated and ventilated mechanically | 300\
response to intense pain | 300\
systolic pressure maintained | 300\
norepinephrine infusion | 300\
postoperative laboratory findings | 300\
abnormal PT/PTT | 300\
fibrinogen | 300\
d-dimer | 300\
antithrombin III | 300\
CK-MB | 300\
troponin-T | 300\
postoperative EKG | 300\
ST elevation | 300\
trans-thoracic echocardiogram | 24\
normal EKG findings | 24\
no patent foramen ovale | 24\
stable vital signs | 24\
norepinephrine infusion tapered out | 24\
unchanged mental status | 120\
brain CT and MRI | 120\
multiple acute cerebral infarctions | 120\
weaned to spontaneous ventilation | 264\
extubated | 264\
unstable vital signs | 360\
intravenous administration of catecholamines | 360\
panperitonitis | 360\
expired due to cardiac arrest | 744\
septic shock | 744