79 years old | 0
male | 0
admitted to the hospital | 0
severe COVID-19 | 0
coronary atherosclerotic heart disease | 0
cerebral infarction | 0
fever | -168
fatigue | -168
anorexia | -168
body temperature 38.5 °C | -168
body temperature fluctuated between 36.5 °C and 38 °C | -168
pulmonary bacterial infection | 0
respiratory failure | 0
co-morbid diseases | 0
poor nutrition | 0
nasogastric tube insertion | 0
physical examination | 0
nasal septum deviation assessment | 0
nasal inflammation assessment | 0
obstruction assessment | 0
cerebrospinal fluid rhinorrhea assessment | 0
laboratory examinations | 0
anti-infection treatment | 0
antiviral treatment | 0
cardiac function improvement treatment | 0
blood transfusions | 0
symptomatic treatments | 0
brain computed tomography (CT) scan | 0
multiple small punctate hypodense foci next to the lateral ventricles bilaterally | 0
ischemic changes | 0
acute ischemic stroke | 0
chest CT | 0
scattered patches and cloudy fuzzy shadows in both lungs | 0
COVID-19 infection | 0
gastric juice extraction | 0
ultrasound examination | 0
nasogastric tube positioning | 0
circular nasogastric tube and comet tail sign | 0
nutrient solution injection | 0
patient stable without adverse reactions | 0
discharge | unknown