52 years old | 0
    male | 0
    hepatitis C virus infection | -4320
    liver cirrhosis | -4320
    portal hypertension | -4320
    grade 1 esophageal varices | -4320
    HIV infection | -4320
    Tenvir-EM (tenofovir 300 mg/emtricitabine 200 mg) | -672
    efavirenz 600 mg | -672
    follow up | -336
    severe epigastric pain | -264
    breathlessness | -264
    nausea | -264
    vomiting | -264
    denied fever | -264
    denied cough | -264
    denied diarrhea | -264
    denied chest pain | -264
    conscious | 0
    Glasgow coma scale 14/15 | 0
    lethargic | 0
    dehydrated | 0
    blood pressure 90/42 mmHg | 0
    pulse rate 133 beats per minute | 0
    temperature 36° Celsius | 0
    tachypneic | 0
    respiratory rate 36 per minute | 0
    oxygen saturation 92% | 0
    mildly icteric | 0
    no flapping tremor | 0
    minimal crepitations | 0
    reduced vocal resonance | 0
    soft abdomen | 0
    moderate ascites | 0
    pitting edema up to the knees | 0
    insignificant cardiovascular examination | 0
    severe metabolic acidosis | 0
    arterial blood gas pH 7.08 | 0
    HCO3- 12 mmol/L | 0
    base excess -16.9 mmol/L | 0
    pCO2 32 mmHg | 0
    lactate level 12.4 mmol/L | 0
    serum ammonia 116 mmol/L | 0
    ALT 55 mmol/L | 0
    bilirubin 37 mmol/L | 0
    elevated WBC 21 × 10^9 | 0
    elevated C-reactive protein 4.0 mmol/L | 0
    unremarkable amylase | 0
    chest radiograph minimal interstitial opacities | 0
    ECG normal sinus rhythm | 0
    ECG no ischemic changes | 0
    intubated | 0
    managed in ICU | 0
    intravenous amoxicillin/clavulanic acid 1.2 g twice daily | 0
    intravenous metronidazole 500 mg twice daily | 0
    continuous veno2venous hemofiltration (CVVH) | 0
    persistent lactic acidosis | 0
    discontinued antiretroviral therapy | 0
    peritoneal fluid analysis unremarkable | 0
    abdominal CT scan unremarkable | 0
    CD4 36 cells/uL | 0
    CD8 27 cells/uL | 0
    gram-negative rod Escherichia coli in blood cultures | 0
    septicemic shock | 0
    E. coli bacteremia | 0
    multiorgan dysfunction | 0
    lactic acid level remained high | 0
    deterioration in liver function | 0
    succumbed to illness | 72
    