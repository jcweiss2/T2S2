36 years old| 0
female | 0
labial pain | -72
swelling | -72
fevers | -72
hypertension | 0
BMI 56 kg/m² | 0
polysubstance abuse | 0
intravenous drug use | 0
opioid abuse | 0
tobacco use | 0
asthma | 0
bipolar disorder | 0
obsessive-compulsive disorder | 0
chronic pain syndrome | 0
homelessness | 0
cesarean section | 0
temperature 38.4°C | 0
blood pressure 135/69 | 0
heart rate 121 bpm | 0
respiratory rate 18 | 0
right labial abscess | 0
mons abscess | 0
opened wound | 0
drainage | 0
leukocytosis 16.5 | 0
lactic acid 0.6 mmol/L | 0
hemoglobin A1C 5.6 | 0
Streptococcus viridians | 0
Staphylococcus aureus | 0
Enterococcus faecalis | 0
Actinomyces species | 0
Corynebacterium species | 0
soft-tissue inflammatory stranding | 0
subcutaneous gas | 0
necrotizing infection | 0
sepsis protocol | 0
IV fluids | 0
vancomycin | 0
piperacillin-tazobactam | 0
clindamycin | 0
left against medical advice | 0
psychiatric assignment officer assessment | 0
four-point restraints | 0
combative behavior | 0
security involvement | 0
police department involvement | 0
surgical debridement | 17
skin-sparing debridement | 17
vulvar NSTI | 17
mons NSTI | 17
second-stage debridement | 41
wound dressings changed daily | 0
Veraflow™ wound vacuum placed | 240
delayed-primary closure | 672
mons pubis panniculectomy | 672
Blake drain placed | 672
Blake drain removed | 1344
broad-spectrum antibiotics transitioned to Augmentin | 0
severe agitation | 0
maladaptive personality | 0
emotional dysregulation | 0
four-point restraints utilized | 0
IV access lost | 0
attempts to leave hospital | 0
intentional wound disruptions | 0
vacuum changes 2-3× per day | 0
pain exacerbations | 0
IV narcotics | 0
psychiatry consultation | 0
palliative care consultation | 0
haloperidol | 0
lorazepam | 0
olanzapine | 0
quetiapine | 0
trazadone | 0
hydroxyzine | 0
scheduled acetaminophen | 0
NSAIDs | 0
gabapentin | 0
oral narcotics | 0
IV opiates discontinued | 0
suboxone regimen initiated | 0
multidisciplinary meetings | 0
discharge planning | 0
women's shelter referral | 0
outpatient chemical dependency referral | 0
gynecology follow-up | 0
transferred to jail | 0
loss to follow-up | 0
