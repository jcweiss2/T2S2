56 years old | 0
    female | 0
    anemia | 0
    high sedimentation rate | 0
    referred to investigate probable malignancy | 0
    diabetes mellitus | 0
    hypertension | 0
    hyperthyroidism | 0
    body temperature 38.0°C | 0
    pulse rate 75 beats/min | 0
    blood pressure 91/55 mm Hg | 0
    tenderness on the left iliac fossa | 0
    bilateral chest radiography showed pleural effusions | 0
    bilateral chest radiography showed minimal infiltration | 0
    blood samples taken for culture | 0
    urine samples taken for culture | 0
    levofloxacin IV 0.5 g antibiotic treatment | 0
    cultures showed Escherichia coli | 24
    antibiotic regimen changed to piperacillin/tazobactam | 24
    antibiotic regimen changed to linezolid | 24
    constipation | 72
    abdominal examination revealed diffuse distension | 72
    abdominal examination revealed tenderness | 72
    abdominal examination revealed sluggish bowel sounds | 72
    abdominal radiography detected air-fluid levels | 72
    abdominal ultrasonography showed free peritoneal fluid | 72
    contrast-enhanced chest MDCT scan performed | 72
    chest MDCT showed bilateral pleural effusion | 72
    chest MDCT showed compression atelectasis | 72
    chest MDCT showed hypodense mass at right breast | 72
    chest MDCT showed calcifications at right breast | 72
    chest MDCT showed enlarged thyroid gland | 72
    chest MDCT showed filling defect secondary to free-floating thrombus | 72
    free-floating thrombus at descending aorta | 72
    thrombus causing partial obstruction of aortic lumen | 72
    sagittal images showed thrombus clinging to aortic wall via peduncle | 72
    coronal images showed thrombus clinging to aortic wall via peduncle | 72
    no signs of aneurysm | 72
    no signs of dissection | 72
    no signs of cardiac thrombus | 72
    abdominal CT revealed massive ascites | 72
    abdominal CT revealed wedge-shaped renal infarction | 72
    echocardiography showed mild mitral regurgitation | 72
    intravenous fluids | 72
    broad spectrum antibiotics | 72
    enoxaparin sodium | 72
    total parenteral nutrition | 72
    surgery not viable | 72
    clinical course worsened with respiratory distress | 144
    clinical course worsened with sepsis | 144
    clinical course worsened with visceral ischemia | 144
    transferred to ICU | 144
    unconscious | 168
    intubated | 168
    leukocyte count 12.3×10^9/L | 168
    hemoglobin 10.5 g/dL | 168
    thrombophilia workup normal | 168
    potassium 3.31 mmol/L | 168
    creatinine 2.14 mg/dL | 168
    lactate dehydrogenase 439 U/L | 168
    albumin 2.79 g/dL | 168
    emergency hemodialysis | 168
    albumin replacement | 168
    decrease in blood pressure | 168
    treated with positive inotropic agents | 168
    cardiac arrest | 216
    full organ support | 216
    cardiovascular resuscitation | 216
    death | 216
  