69 years old | 0
male | 0
hypertension | 0
CKD stage 5 | 0
hemodialysis | 0
consumed 6 bilimbi fruits | -48
uncontrollable hiccups | -45
malaise | -45
abdominal discomfort | -45
macroscopic hematuria | -45
nausea | -28
vomiting | -28
decrease in the level of consciousness | -24
dysarthria | -24
myoclonus of the upper limbs | -24
seizures | -24
admitted to the hospital | 0
mechanical ventilation | 0
orotracheal intubation | 0
Richmond Agitation Sedation Scale score of −3 | 0
hemodynamically stable | 0
blood pressure of 110/60 mm Hg | 0
heart rate of 68 bpm | 0
diffuse ecchymoses on the trunk and extremities | 0
hemoglobin of 13.1 g/dL | 0
hematocrit of 39.3% | 0
white blood cells of 13,600/mL | 0
band form count of 3% | 0
179,000 platelets/mL | 0
urea blood levels of 86.8 mg/dL | 0
serum creatinine of 7.11 mg/dL | 0
serum sodium of 139 mEq/L | 0
serum potassium of 3.93 mEq/L | 0
hypoattenuation in the periventricular deep white matter and centrum semiovale | 0
lumbar puncture | 0
transparent, colorless cerebrospinal fluid | 0
22 red blood cells | 0
normal concentrations of glucose, white blood cells, and proteins | 0
negative results from the bacterial test, China ink test, analysis for fungi, and acid-fast staining | 0
phenytoin | 0
midazolam | 0
sustained low-efficiency daily dialysis (SLEDD) | 0
severe hypotension | 6
norepinephrine | 72
hemodynamic worsening | 72
infectious process | 72
hemoglobin of 12.5 g/dL | 72
hematocrit of 38.8% | 72
white blood cells of 16,700/mL | 72
band form count of 8% | 72
180,000 platelets/mL | 72
C-reactive protein (CRP) levels to 320 mg/dL | 72
antibiotic therapy | 72
piperacillin-tazobactam | 72
septic shock secondary to ventilator-associated tracheobronchitis | 72
seizures during attempts to reduce the dose of the sedative medications | 96
further tests | 96
immunosuppression with intravenous methylprednisolone | 96
search for rheumatic diseases | 96
electroencephalogram (EEG) | 120
epileptogenic activity | 120
thiopental | 120
family confirmed that the patient had consumed bilimbi fruit | 120
EEG detected a decrease in paroxysmal activity | 192
therapy with thiopental, midazolam, and valproic acid | 192
attempt to intensify hemodialysis | 192
EEG suggested improvement of the seizure disorder | 240
thiopental and midazolam were gradually decreased | 240
valproic acid increased | 240
dose of noradrenaline had to be increased | 288
fever (38.5°C) | 288
lactate of 3.9 mmol/L | 288
white blood cells of 21,500/mL | 288
band form count of 9% | 288
CRP of 107 mg/dL | 288
septic shock of unknown origin | 288
meropenem, vancomycin, and gentamicin | 288
blood, tracheal aspirate, and catheter samples were collected | 288
isolates of multidrug-resistant Klebsiella pneumoniae | 288
tigecycline | 288
conscious and responsive, with no sedatives | 336
persistent myoclonus in the lower limbs | 336
no new episodes of generalized tonic-clonic seizures | 336
SLEDD was maintained with low clinical tolerability | 336
worsening of the clinical status | 552
progressive increase in vasoactive drug doses | 552
fever | 552
leukocytosis | 552
increased CRP levels | 552
died of circulatory failure | 648