7-year-old | 0  
    girl | 0  
    admitted to the hospital | 0  
    periodic fever of over 38℃ | -144  
    headache | -144  
    abdominal pain | -144  
    watery diarrhea | -144  
    projectile vomiting | -144  
    severe headache | -144  
    lethargy | -144  
    conjugated pneumococcal vaccines | 0  
    Haemophilus influenzae type b vaccines | 0  
    neck stiffness | 0  
    Bruzinski sign positive | 0  
    Kernig sign positive | 0  
    no abnormality in motor function | 0  
    muscle strength intact | 0  
    sensation intact | 0  
    deep tendon reflexes hyper-reactive | 0  
    white blood cell counts 21,150/µL | 0  
    segmented neutrophils 89% | 0  
    lymphocytes 6.3% | 0  
    ESR 57 mm/hr | 0  
    CRP 9.52 mg/dL | 0  
    fasting blood sugar 169 mg/dL | 0  
    CSF white blood cells 1,500/µL | 0  
    CSF segmented neutrophils 30% | 0  
    CSF red blood cells 250/µL | 0  
    CSF sugar 25 mg/dL | 0  
    CSF protein 117 mg/dL | 0  
    no bacteria on gram staining | 0  
    PCR for tuberculosis negative | 0  
    herpes simplex virus antibody test negative | 0  
    co-agglutination test negative | 0  
    cryptococcus antigen test negative | 0  
    ceftriaxone | 0  
    amikacin | 0  
    steroid injections | 0  
    vancomycin | 48  
    fever over 39℃ | 48  
    severe headache | 48  
    vomiting | 48  
    altered mental status | 48  
    stuporous | 48  
    delirious | 48  
    suspected increased intracranial pressure | 48  
    diplopia | 48  
    brain MRI performed | 48  
    no brain edema | 48  
    fever continued | 72  
    headache continued | 72  
    pain in both legs | 72  
    worsening mental status | 72  
    repeated CSF examination | 72  
    repeated blood tests | 72  
    white blood cells 37,860/µL | 72  
    segmented neutrophils 88.2% | 72  
    lymphocytes 5.3% | 72  
    ESR 50 mm/hr | 72  
    CRP 17.19 mg/dL | 72  
    fasting blood sugar 142 mg/dL | 72  
    CSF white blood cells 2,000/µL | 72  
    CSF segmented neutrophils 35% | 72  
    CSF red blood cells 250/µL | 72  
    CSF sugar 73 mg/dL | 72  
    CSF protein 319 mg/dL | 72  
    gram-positive rods confirmed | 72  
    L. monocytogenes identified | 72  
    ampicillin | 72  
    antimicrobial susceptibility test | 72  
    IgG 872 mg/dL | 72  
    IgA 208 mg/dL | 72  
    IgM 257 mg/dL | 72  
    IgE 960 IU/mL | 72  
    C3 113 mg/dL | 72  
    C4 28.2 mg/dL | 72  
    CH50 51.1 U/mL | 72  
    CD3 61.3% | 72  
    CD4 32.7% | 72  
    CD8 35.2% | 72  
    CD19 17% | 72  
    ultrasound of thymus normal | 72  
    responded to pain stimulation | 96  
    confused conversation | 96  
    no voluntary movement | 96  
    pupillary reflexes slow | 96  
    nystagmus | 96  
    muscle strength decreased to grade 2 | 96  
    respiratory difficulty | 96  
    semicoma level | 96  
    transferred to intensive care unit | 96  
    ventilator support initiated | 96  
    brain CT | 96  
    hydrocephalus | 96  
    parenchymal edema | 96  
    brain stem extrusion | 96  
    increased third and fourth cerebral ventricles | 96  
    increased lateral ventricles | 96  
    extraventricular drainage performed | 96  
    additional extraventricular drainage on sixth day | 144  
    additional extraventricular drainage on fourteenth day | 336  
    CSF white blood cells 32/µL | 408  
    CSF red blood cells 3,100/µL | 408  
    CSF sugar 99 mg/dL | 408  
    CSF protein 169 mg/dL | 408  
    no bacteria detected | 408  
    no bacteria on blood culture | 408  
    no bacteria on CSF culture | 408  
    worsening hydrocephalus | 528  
    consciousness not improving | 528  
    ventriculoperitoneal shunt performed | 528  
    off ventilator support | 600  
    appropriate response | 600  
    language no longer confused | 600  
    vital signs stable | 744  
    transferred to general ward | 744  
    brain CT on 38th day | 912  
    communicating hydrocephalus | 912  
    ventriculostomy | 912  
    parenchymal edema | 912  
    recovered consciousness | 1464  
    recovered motor functions | 1464  
    discharged | 1464  

