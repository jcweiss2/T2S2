72 years old | 0
male | 0
admitted to the emergency room | 0
fever | 0
penile pain | 0
vomiting | 0
diarrhea | 0
history of hemodialysis | -6120
history of diabetic nephropathy | -6120
history of percutaneous transluminal angioplasty | -unknown
lanthanum carbonate hydrate | -unknown
calcium carbonate | -unknown
cilostazol | -unknown
lansoprazole | -unknown
cinacalcet | -unknown
amlodipine | -unknown
enalapril maleate | -unknown
carvedilol | -unknown
non-smoker | 0
does not consume alcohol regularly | 0
good general condition | 0
physical examination | 0
penile pain worsened | 9
lost consciousness | 9
Glasgow Coma Scale score of 3 | 0
blood pressure of 84/58 mmHg | 0
respiratory rate of 28 breaths per minute | 0
heart rate of 102 beats per minute | 0
temperature of 37.6°C | 0
oxygen saturation of 100% | 0
cold sweat | 0
swelling and dark brownish changes at the glans | 0
white blood cell count of 5,600 /μL | 0
hemoglobin of 10.2 g/dL | 0
platelets of 81,000 /μL | 0
sodium of 141 mmol/L | 0
potassium of 5.3 mmol/L | 0
chloride of 103 mmol/L | 0
creatinine of 9.71 mg/dL | 0
blood urea nitrogen of 47.7 mg/dL | 0
albumin of 3.3 g/dL | 0
calcium of 9.4 mg/dL | 0
phosphorus of 5.8 mg/dL | 0
parathyroid hormone of 280 pg/mL | 0
C-reactive protein of 129.8 mg/L | 0
total bilirubin of 1.5 mg/dL | 0
aspartate aminotransferase of 34 IU/L | 0
alanine aminotransferase of 10 IU/L | 0
atrial blood gas with oxygen flow rate of 15 L/min | 0
pH of 7.031 | 0
PaCO2 of 62.4 Torr | 0
PaO2 of 80.6 Torr | 0
HCO3 of 15.7 mEq/L | 0
anion gap of 25.0 mmol/L | 0
respiratory condition deteriorated | 3
intubated | 3
admitted to the intensive care unit | 3
blackish changes on the entire penis and scrotum | 3
test incision in the perineum, penis, and scrotum | 3
no evidence of effusion | 3
contrast-enhanced computed tomography of the pelvic region | 3
poor contrast enhancement of the penis | 3
no intestinal necrosis | 3
no evidence of abscess or gas in the penis | 3
treated with antibiotics | 3
treated with vasoactive agents | 3
treated with hydrocortisone | 3
treated with continuous hemodiafiltration dialysis | 3
metabolic acidosis and hyperkalemia progressed | 12
died | 12
postmortem blood culture showed Streptococcus dysgalactiae subsp. equisimilis | 12
diagnosis of STSS | 12
antimicrobial susceptibility results of SDSE | 12
pathological autopsy | 12
calcification of the aorta | 12
ischemic necrosis of the stomach | 12
ischemic necrosis of the lower gastrointestinal tract | 12
calcified lesions and numerous infected thrombi | 12
septic emboli associated with Gram-positive Streptococcus | 12
calcium deposition in small arteries | 12