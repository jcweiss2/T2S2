65 years old | 0\
male | 0\
multiple blisters and erosions all over his body including oral mucosa, scalp with superadded maggot infection | -432\
previous episodes of such lesions | -720\
treated with steroids and some unknown generic medications | -720\
lesions all over the body | -180\
febrile | 0\
numerous flaccid blisters and erosions covering more than 85% of body surface area with some of them covered with slough and maggots | 0\
Nikolsky sign was strongly positive | 0\
diagnosis of PV was confirmed by a skin biopsy | 0\
tzanck smear | 0\
intravenous (IV) dexamethasone pulse (120 mg) | 0\
supportive care such as fluids, fresh frozen plasma (FFP) and dressings | 0\
intravenous antibiotics (Piperacillin/Tazobactam and Teicoplanin) | 0\
oozing from skin ulcerations and hemorrhagic excoriation with peeling of skin | 0\
maintained on 1 mg/kg of oral methyl prednisolone | 72\
no improvement in the skin lesions and general condition of the patient worsened further with hypoproteinemia | 168\
developed pleural effusion | 168\
blood culture showed enterobacter | 168\
pus culture from erosions show Staphylococcus aureus and Proteus mirabilis | 168\
intravenous Tigecycline and vancomycin | 168\
erosions still persisted and did not show any sign of re-epithelialization | 168\
perilesional Nikolsky sign was still positive | 168\
developed new blisters | 168\
sepsis with persistent high grade fever | 168\
albumin levels fell to 2.1 mg | 168\
hold the “Pulse therapy” of IV methyl prednisolone and cyclophosphamide | 168\
plan for one TPE cycle | 168\
TPE was performed | 216\
Nikolsky sign became negative | 240\
no new lesions appeared | 240\
exudation from the lesions reduced drastically | 240\
dressings also started to remain dry | 240\
lesions showed 60-70% re-epithelization | 288\
lesions showed 90% healing | 312\
oral lesions also healed completely | 312\
little erosions on back, anterior aspect of thigh and buttocks persisted | 312\
given “Pulse therapy” of IV methyl prednisolone (1 gm/day) and cyclophosphamide (500 mg/day) | 312\
further improvement in the lesions | 336\
patient was clinically stable | 336\
plan was to given one more TPE cycles for three sessions | 336\
discharged on maintained dose of monthly IV dexamethosone pulse along with daily oral prednisolone (60 mg/day) | 360