77 years old | 0
female | 0
breast cancer | 0
chemotherapy | 0
radiation to the chest | 0
severe aortic stenosis | 0
coronary artery disease | 0
90% occlusion of the left anterior descending artery | 0
tissue aortic valve replacement | 0
saphenous vein graft bypass | 0
midline sternotomy | 0
induction of anesthesia | 0
intubation | 0
left internal mammary artery dissection | 0
atretic left internal mammary artery | 0
unusable left internal mammary artery | 0
use of greater saphenous vein | 0
small greater saphenous vein | 0
discontinuation of cardiopulmonary bypass | 0
decline in cerebral head saturations | 0
reduced mean arterial perfusion | 0
reduced cerebral artery perfusion | 0
vasopressor use | 0
intensive care unit admission | 0
extubated 2 h postoperatively | 2
persistent lactic acidosis | 15
high-dose vasopressor support | 15
mean arterial perfusion pressure goal >65 mm Hg | 15
mixed cardiogenic and vasoplegic shock | 15
lethargic | 15
leftward gaze | 15
right upper extremity weakness | 15
symptoms resolved over 15 minutes | 15
bilateral tongue ecchymoses | 15
tongue numbness | 15
dysgeusia | 15
CT scan negative for acute hemorrhage | 15
CT angiogram negative for large vessel occlusion | 15
transient ischemic attack | 15
mild calcification at bifurcation of right common carotid artery | 15
50% focal stenosis of distal left common carotid artery | 15
completely occluded right lingual artery | 15
mild distal collateral flow | 15
multifocal irregularities in left lingual artery | 15
normal platelet count | 15
normal prothrombin time | 15
normal INR | 15
normal fibrinogen | 15
no prior vasculitic disease | 15
normal ADAMTS13 inhibitor screen | 15
volume resuscitation with crystalloid | 15
volume resuscitation with colloid | 15
low-dose epinephrine | 15
high-dose norepinephrine | 15
high-dose vasopressin | 15
systemic vascular resistance improvement over 2 days | 15
otolaryngology consultation | 15
serial tongue examinations | 15
flexible bronchoscopes for disease monitoring | 15
persistent tongue numbness | 15
persistent dysgeusia | 15
supportive therapy | 15
symptom improvement with shock treatment | 15
no surgical intervention | 15
tongue sensation return to baseline at 2 months | 1440
taste return to baseline at 2 months | 1440
bilateral lingual artery involvement confirmed | 15
atretic vessels systemically | 0
small internal mammary arteries | 0
small saphenous veins | 0
reduced cerebral perfusion intraoperatively | 0
transient ischemic attack postoperatively | 15
atherosclerotic emboli possibility | 15
shower emboli during aortic cross clamp | 0
short duration of endotracheal intubation | 2
multifactorial etiology | 15
bilateral tongue ischemia | 15
lingual artery disease confirmed by imaging | 15
improved symptoms without surgery | 15
high mortality associated with tongue ischemia | 0
possible surgical debridement in severe cases | 0
conservative management | 0
self-amputation possibility | 0
self-resolution possibility | 0
speech and language alterations | 0
swallowing difficulties | 0
prompt diagnosis | 0
management strategies | 0
