16 years old | 0
female | 0
admitted to the hospital | 0
fever | -336
generalized weakness | -336
joint pain | -336
auricular perichondritis | -336
arthritis | -336
no skin rash | -336
no abdominal pain | -336
no headaches | -336
no visual disturbances | -336
no changes in urinary or bowel habits | -336
no change in weight | -336
no ill contacts | -336
red and swollen ears | 0
joint line tenderness | 0
no limitations of active or passive range of motion | 0
no joint swelling or redness | 0
normal chest shape and contour | 0
no murmurs | 0
no added sounds | 0
no wheeze or crackles | 0
splenomegaly | 0
temperature 39°C | 0
pulse rate 102 BPM | 0
blood pressure 102/80 mmHg | 0
respiratory rate 18 respirations per minute | 0
oxygen saturation 98% | 0
hemoglobin 11.9 g/dL | 0
mean corpuscular volume 79.2 mm3 | 0
platelets 308,000/mm3 | 0
white blood cell count 14,600/mm3 | 0
C-reactive protein 369 mg/L | 0
erythrocyte sedimentation rate 110 mm/hr | 0
lactate dehydrogenase 561 U/L | 0
broad spectrum antibiotics | 0
intravenous fluids | 0
paracetamol | 0
Brucella antibodies negative | 24
cytomegalovirus negative | 24
Epstein-Barr virus negative | 24
rheumatoid factor negative | 24
antinuclear antibodies negative | 24
hepatitis A immunoglobulin antibodies negative | 24
bone marrow aspirate showed increased numbers of cytologically normal monocytes | 24
blasts not increased | 24
lymphocytes and plasma cells normal | 24
Leishmania testing negative | 24
abdominal ultrasound showed enlarged spleen | 48
whole-body computed tomography scan showed enlarged spleen and mesenteric lymph node enlargement | 48
echocardiography showed significant apical hypokinesia | 48
pulmonary hypertension 50 mmHg | 48
tricuspid regurgitation | 48
mobile echo-dense structure on the pulmonic valve | 48
blood film showed microcytic hypochromic red blood cells | 72
Rouleaux formation | 72
leukocytosis with segmented neutrophils and occasional monoblasts | 72
transferred to hematology/oncology facility | 72
fever | 96
tachycardia 110 bpm | 96
hypotension 90/58 mmHg | 96
leukocytosis 51,000/mm3 | 96
absolute neutrophil count 36,000/mm3 | 96
HBG 7.5 g/dL | 96
CRP 240 mg/L | 96
ESR 145 mm/hr | 96
broad spectrum antibiotics | 96
urine and blood cultures negative | 120
transferred to ICU | 120
ferritin 3200 ng/mL | 144
fibrinogen 1.43 mg/dL | 144
total serum bilirubin 2.7 mg/dL | 144
direct serum bilirubin 1.2 mg/dL | 144
LDH 583 U/L | 144
cytoplasmic anti-neutrophil cytoplasmic antibodies negative | 144
perinuclear ANCA negative | 144
antinuclear antibodies negative | 144
RF negative | 144
Anti-Jo negative | 144
anti-Sjögren’s-syndrome-related antigen A and B antibodies negative | 144
anti-double-stranded DNA negative | 144
anti-smith negative | 144
anti-scl-70 antibodies negative | 144
palpable purpuric and bullous skin lesions | 168
skin biopsy showed epidermal edema | 168
diffuse interstitial neutrophilic infiltration | 168
no evidence of vasculitis | 168
diagnosis of RP with HLH | 168
treated with paracetamol | 168
IV fluids | 168
2 units of packed RBCs | 168
prednisolone 60 mg | 168
IVIG | 168
hydroxyurea | 168
warfarin 5 mg per day | 168
furosemide 40 mg per day | 168
cyclosporine 100 mg twice daily | 168
prednisone 60 mg | 168
remission | 336
relapse | 504
bone marrow examination showed AML | 504
cytarabine 100 mg/m2 | 504
allopurinol | 504
heart failure | 504
incomplete treatment protocol for AML | 504
died due to Enterococcus fecium sepsis and multiorgan failure | 720