64 years old | 0
male | 0
obesity | 0
olfactory groove meningioma | 0
left-sided optic neuropathy | 0
bifrontal craniotomy | -24
endoscopic resection | -24
intra- and postoperative empiric antibiotics | -24
steroids | -24
pneumcephalus | -24
non-contrast computed tomography (NCCT) scan | -24
palpable collection below the scalp | -120
worsening pneumocephalus | -120
large scalp collection | -120
disorientation | -144
unsteady gait | -144
worsening of intracranial and extracranial air | -168
decline of mental status | -168
decline of respiratory status | -168
bradycardia | -168
tachypnea | -168
hypoxia | -168
endotracheal intubation | -168
emergent bedside needle decompression | -168
endoscopic exploration and repair of the anterior cranial fossa defect | -168
profound hypotension | -168
multiple vasopressors | -168
diffuse pulmonary edema | -168
acute respiratory distress syndrome | -168
white blood cell count of 44 | -168
erythrocyte sedimentation rate of 49 mm/h | -168
C-reactive protein of 11.7 mg/dL | -168
procalcitonin of 1.17 ng/mL | -168
platelet count of 521 | -168
lactate of 2.25 mmol/L | -168
creatinine of 2.3 mg/dL | -168
broad-spectrum antibiotics | -168
improved pneumocephalus | -216
normalized laboratory parameters | -240
improved kidney function | -240
weaned off vasopressors | -240
extubation | -264
CSF sampling | -408
white blood cell count of 25 | -408
glucose of 111 mg/dL | -408
protein of 194 mg/dL | -408
lactic acid of 4.1 mmol/L | -408
near-complete resolution of pneumocephalus | -1296
admitted to the hospital | 0 
tension pneumocephalus | -168 
systemic inflammatory response syndrome (SIRS) | -168 
multiorgan dysfunction | -168 
catecholamine surge | -168 
increased intracranial pressure | -168 
central dysregulation | -168 
emergent decompression | -168 
surgical repair of the cranial fossa defect | -168 
critical care support | -168 
reversal of tension pneumocephalus | -216 
reversal of SIRS response | -216 
infection | -168 
postoperative state | -24 
SIRS-like response | -24 
close observation | 0 
timely neurosurgical intervention | 0 
supportive care | 0 
progressive pneumocephalus | -120