55 years old | 0
male | 0
admitted to emergency department | 0
dyspnea | 0
fever | -168
cough | -168
whitish sputum | -168
former smoker | 0
5-pack-year | 0
no alcohol abuse history | 0
no known history of pulmonary diseases | 0
no underlying diseases | 0
no medications or herbal medicines | 0
atypical chest pain | -72
admitted to coronary care unit | -72
normal coronary angiography | -72
normal chest radiography | -72
chest computed tomography | -72
diffuse bronchial wall thickening | -72
no evidence of emphysema | -72
flu-like symptoms | -72
fever | -72
cough | -72
sore throat | -72
myalgia | -72
conservative medication | -72
no antiviral agents | -72
blood pressure 130/90 mm Hg | 0
heart rate 113 beats/min | 0
respiratory rate 26 breaths/min | 0
body temperature 37.8℃ | 0
conscious | 0
acute ill-looking appearance | 0
normal conjunctiva | 0
no palpable lymph nodes | 0
bilateral expiratory wheezes | 0
white blood cells 15,200/mm3 | 0
neutrophils 84.9% | 0
lymphocytes 8.6% | 0
eosinophils 0.5% | 0
hemoglobin 16.0 g/dL | 0
platelets 144,000/mm3 | 0
C-reactive protein 46.5 mg/L | 0
liver function tests normal | 0
renal function tests normal | 0
serologic tests for autoantibodies negative | 0
rheumatoid factor negative | 0
human immunodeficiency virus negative | 0
venereal disease research laboratory test negative | 0
CD4 count normal | 0
arterial blood gas analysis | 0
pH 7.45 | 0
PaO2 81.8 mm Hg | 0
PaCO2 38.5 mm Hg | 0
rapid influenza diagnostic test negative | 0
anti-mycoplasma antibody negative | 0
urinary antigen tests for Legionella negative | 0
urinary antigen tests for pneumococcus negative | 0
sputum and blood cultures negative | 0
special stain for acid-fast bacilli negative | 0
serum galactomannan assay positive | 24
ceftriaxone and clarithromycin | 0
community-acquired pneumonia | 0
acute exacerbation of asthma | 0
methylprednisolone | 24
bilateral wheezes | 24
no history of asthma | 24
no history of pulmonary diseases | 24
piperacillin/tazobactam plus levofloxacin | 96
worsening leukocytosis | 96
hypoxemia | 96
respiratory failure | 96
mechanically ventilated | 96
intensive care unit | 96
fever subsided | 192
C-reactive protein level declined | 192
chest radiographic findings improved | 192
high fever | 216
worsening chest radiographic findings | 216
bronchoscopy | 216
extensive yellow-whitish exudative pseudomembranes | 216
trachea and both main bronchi | 216
airway narrowing | 216
acute-angle branching hyphal elements | 216
bronchoalveolar lavage fluid | 216
Aspergillus species colonies | 216
repeat serum GM assays positive | 216
polymerase chain reaction of BAL fluid positive for influenza B | 216
probable IPA | 216
voriconazole | 216
progressively worsened | 240
no documented bacterial infection | 240
died | 336