33 years old |
