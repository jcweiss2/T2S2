40 years old|0
male|0
motorcycle collision|0
hypotensive|0
alert|0
left needle thoracostomy|0
decreased breath sounds|0
hypotensive upon arrival|0
blood pressure 60 mmHg systolic|0
intubated|0
massive transfusion protocol activated|0
left chest deformity|0
left chest tube placed|0
initial return of >2000 cc blood|0
taken to operating room emergently for left thoracotomy|0
multiple comminuted rib fractures|0
multiple large pulmonary lacerations|0
left diaphragm injury|0
bilateral hemothoraces|0
fragment of bone abutting pericardium|0
thoracotomy converted to clamshell thoracotomy|0
pericardium incised|0
heart intact|0
tractotomy required to control pulmonary hemorrhage|0
left chest packed|0
exploratory laparotomy performed|0
superficial splenic lacerations|0
left humerus fracture|0
left scapula fracture|0
postoperative hypotension|0
systolic blood pressures in low 80s mmHg|0
hypoxic|0
massive transfusion including 38 packed red blood cells|0
massive transfusion including 36 plasma|0
massive transfusion including 4 units of platelets|0
hospital's blood supply exhausted|0
poor prognosis|0
started on vasopressors|0
resuscitation continued|0
failed to respond to additional fluid resuscitation|0
hemorrhage controlled|0
empiric hydrocortisone 100 mg dose|0
empiric hydrocortisone continued every 8 h|0
patient stabilized with systolic blood pressures into 150s mmHg|0
vasopressors weaned|0
fluids decreased|0
family contacted|24
history of hypopituitarism from previous head trauma|24
taking levothyroxine for several years|24
taking hydrocortisone for several years|24
returned to operating room 2 days later for washout|48
rib fixation|48
closure of left chest|48
extubated on posttrauma day 6|144
left bronchopulmonary fistula|144
pulmonary embolism|144
heparin-induced thrombocytopenia|144
discharged on 47th day of hospitalization|1128
returned to work|8760
no respiratory difficulty|8760
