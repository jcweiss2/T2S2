67 years old | 0
male | 0
admitted to the hospital | 0
fever | -336
cough | -336
shortness of breath | -336
renal transplant | -6720
end-stage renal disease | -6720
diabetic nephropathy | -6720
hypertension | 0
diabetes mellitus | 0
antihypertensive therapy | 0
insulin use | 0
immunosuppressive therapy | 0
mycophenolate mofetil | -672
tacrolimus | -672
prednisone | -672
dyspnea | 0
body temperature of 38.0°C | 0
respiratory rate of 28 breaths/minute | 0
oxygen saturation of 98% | 0
blood pressure of 134/71 mmHg | 0
heart rate of 101 beats/minute | 0
pulmonary moist rale | 0
pitting edema in the lower extremities | 0
white blood cell count of 8.2×10^9 cells/L | 0
neutrophils of 89.5% | 0
hemoglobin level of 114 g/L | 0
platelet count of 187×10^9 cells/L | 0
potassium ion of 6.59 mmol/L | 0
creatinine of 193 μmol/L | 0
C reactive protein of 199 g/L | 0
HIV test negative | 0
pleural effusion | 0
bilateral airspace opacities | 0
pneumonia | 0
methylprednisolone | 0
imipenem/cilastatin | 0
trimethoprim–sulfamethoxazole | 0
continuous venovenous hemodialysis | 0
mechanical ventilation | 72
respiratory failure | 72
heart failure | 72
Chest CT scan | 72
discrete scattered patchy consolidation in both lungs | 72
sputum culture | 72
Candida albicans | 72
blood culture | 72
negative results | 72
teicoplanin | 120
caspofungin | 120
T. asahii fungemia | 216
sepsis | 240
multiple organ failure | 240
death | 240
Vitek 2 YST yeast identification kit | 240
antifungal susceptibility test | 240
amphotericin B | 240
itraconazole | 240
fluconazole | 240
voriconazole | 240
5-fluorocytosine | 240