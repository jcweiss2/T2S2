30 years old| 0
woman | 0
abnormal liver function (2-year history) | 0
admitted to the hospital | 0
persistent jaundice | 0
abdominal distension | 0
intermittent mild fever | -720
serologic antibodies negative for hepatitis virus A | 0
serologic antibodies negative for hepatitis virus B | 0
serologic antibodies negative for hepatitis virus C | 0
serologic antibodies negative for hepatitis virus E | 0
serologic antibodies negative for Epstein-Barr virus | 0
serologic antibodies negative for cytomegalovirus | 0
serologic antibodies negative for rubella virus | 0
antibodies of autoimmune diseases negative | 0
alpha fetoprotein (AFP) negative | 0
no alcohol abuse | 0
no hepatotoxic prescriptions | 0
no gastrointestinal hemorrhage | 0
no surgery in the last few months | 0
abdominal contrast-enhanced CT showing liver cirrhosis with moderate ascites | -168
no space occupying lesions in the liver | -168
temperature 38.1°C | 0
heart rate 98 bpm | 0
normal breathing | 0
normal blood pressure | 0
fully conscious | 0
thyroid non-tender | 0
no thyromegaly | 0
bulging abdomen | 0
positive ascites sign | 0
pitting edema | 0
ecchymosis on both lower limbs | 0
total leukocyte count 3.19×10^9/L | 0
neutrophil percentage 63.3% | 0
red blood cell count 3.46×10^12/L | 0
hemoglobin 10.7 g/L | 0
platelets 80×10^9/L | 0
bone marrow biopsy normal | 0
no infection found | 0
liver function persistently worsened | 0
increasing bilirubin | 0
coagulopathy | 0
low serum ceruloplasmin 0.108 g/L | 0
higher urinary copper 5.5 μmol/L | 0
normal blood copper 9.7 μmol/L | 0
Kayser Fleischer ring detected by slit lamp | 0
positive ATP-7B gene detection (Wilson disease) | 0
New Wilson index score 13 | 0
thyroid-stimulating hormone <0.005 mU/L | 0
free thyroxine 50.67 pmol/L | 0
thyrotrophin receptor antibody 4.52 IU/L | 0
thyroid Doppler ultrasound showing non-uniform density with rich blood flow | 0
apparent abnormal liver function | 0
anti-thyroid drugs contraindicated | 0
radioactive iodine therapy considered | 0
iodine level in 24-h thyroid uptake 4.1% | 0
anti-copper treatment not effective | 0
liver transplantation considered as only solution | 0
polyene phosphatidyl choline used | 0
ademetionine 1,4-butanedisulfonate used | 0
diuretics used | 0
infusion of albumin | 0
infusion of plasma | 0
persistent mild fever | 0
liver function deteriorated | 0
no suitable liver donation | 0
hepatic encephalopathy developed | 384
progressed to coma | 432
plasma exchange | 432
mechanical ventilation | 432
supportive treatments in ICU | 432
persistently comatose condition | 432
increasing serum bilirubin level | 432
bleeding in gastrointestinal tract | 432
bleeding in respiratory tract | 432
bleeding in urinary tract | 432
family members stopped treatment | 432
died | 432
