41 years old | 0
male | 0
admitted to the hospital | 0
pain in the right lower posterior teeth | -168
swelling and pain in the oral and maxillofacial head and neck regions | -168
difficulty in breathing | -48
difficulty in swallowing | -48
placed a cigarette butt dipped in the pesticide "Miehailin" into the "dental cavity" | -168
visited a local community clinic | -144
removed the cigarette butt | -144
received an infusion of anti-inflammatory drugs | -144
odontogenic infections gradually became aggravated | -144
spread bilaterally to the floor of the mouth, submandibular space, neck, chest, waist, back, temporal and other areas | -144
mentally exhausted | -168
poor diet | -168
poor sleep | -168
weight loss of approximately 2.5 kg | -168
acutely painful face | 0
extensive swelling and pneumatosis in the bilateral temporal, oral, maxillofacial, neck, chest, waist and back regions | 0
skin redness and high temperature | 0
submandibular space and neck regions pulsated when touched | 0
puncture revealed purulent fluid which was black, thin, with bubbles and had a foul odor | 0
mouth opening was less than 1 cm | 0
leukocyte count was 13.53 × 10^9/L | 0
neutrophil ratio was 88.40% | 0
hypersensitive C-reactive protein was > 180 mg/L | 0
procalcitonin was 9.8 ng/mL | 0
electrolyte results were abnormal | 0
liver and kidney function test results were abnormal | 0
platelet count was 41.0 × 10^9/L | 0
D-dimer level was 1184 ng/mL | 0
blood culture indicated infection with Streptococcus viridans | 0
drug sensitivity testing indicated that the organism was sensitive to penicillin antibiotics | 0
computed tomography scans showed extensive swelling and pneumatosis in soft tissues bilaterally | 0
upper respiratory tract was narrowed slightly | 0
bilateral lung pneumothorax was observed | 0
small amount of effusion was seen bilaterally in the pleura and pericardium | 0
lung pneumothorax was more serious on the left side | 0
compression ratio was approximately 20%-30% | 0
pulmonary infection was seen in both lungs | 0
transferred to the intensive care unit | 0
oral and maxillofacial surgeons organized consultations and discussion of treatment plans | 0
extensive abscess incision and drainage in the oral and maxillofacial head and neck regions | 0
thoracic and pericardial puncture, catheter drainage and pneumothorax management | 0
management of back and waist infections | 0
anesthesia and respiratory management | 0
platelets and blood transfusion | 0
intensive care, antimicrobial administration, nutritional support, water, electrolytes and acid-base stability | 0
platelets decreased to 22.00 × 10^9/L | 24
liver and kidney function tests were abnormal | 24
electrolytes were abnormal | 24
liver and kidney function continued to deteriorate | 48
septic shock | 72
respiratory and cardiac arrest | 72
cardiopulmonary resuscitation | 72
died | 72
severe multi-space infections bilaterally in the oral and maxillofacial head and neck regions | 0
secondary infections of the thorax, back and waist | 0
mediastinal abscess | 0
bilateral pneumothorax | 0
bilateral pulmonary infection | 0
purulent pleural effusion | 0
pericardial effusion | 0
secondary thrombocytopenia | 0
septic shock | 72
acute hepatic and renal insufficiency | 72
multi-space infections in the oral and maxillofacial head and neck regions | 0
odontogenic infection | -168
toothache | -168
dental pain | -168
use of pesticide "Miehailin" | -168
toxicity of pesticides | 0
secondary thrombocytopenia | 0
spread of odontogenic infection | -144
timely incision and drainage | 0
respiratory obstruction | 0
mortality in multi-space infections | 72