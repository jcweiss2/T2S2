40 years old | 0
    female | 0
    referred | -336
    diagnosed with WOPN | -336
    WOPN size 13 × 9 × 7.4 cm | -336
    acute severe pancreatitis | -504
    initial admission | -336
    acute severe epigastric pain | -336
    leukocytosis 2.73 × 103/µl | -336
    neutrophils 91% | -336
    serum amylase 1,309 U/l | -336
    total bilirubin 1.9 mg/dl | -336
    direct bilirubin 0.5 mg/dl | -336
    AST 126 U/l | -336
    ALT 343 U/l | -336
    alkaline phosphatase 104 U/l | -336
    endoscopic retrograde cholangiopancreatography | -336
    common bile duct sludge | -336
    no intensive care | -336
    high-grade fever | -336
    abdominal pain | -336
    CT scan pancreatic necrosis | -336
    fluid collection at pancreatic body | -336
    high-grade fever persisted | -336
    intravenous antibiotics | -336
    EUS-guided drainage | -336
    10 Fr × 7 cm double pigtail stent | -336
    prophylactic antibiotics | -336
    re-admitted | -240
    severe abdominal pain | -240
    sepsis | -240
    CT scan enlargement of pancreatic collection | -240
    increased enhancement of the rim | -240
    septation | -240
    air inside | -240
    repeat EUS-guided drainage | -240
    infected WOPN | -240
    procedure left lateral decubitus position | -240
    curvilinear echoscope GF UC-140P | -240
    partially clogged stent | -240
    large collection with turbid content | -240
    turbid content | -240
    air inside | -240
    punctured abscess using 19-gauge needle | -240
    aspirated purulent fluid | -240
    fluid sent for culture | -240
    contrast injection | -240
    8.5 Fr tapered tip Teflon catheter | -240
    10 Fr tapered tip Teflon catheter | -240
    10 Fr × 7 cm double pigtail stent inserted | -240
    multiseptated collection | -240
    thick pus | -240
    turbid pus | -240
    placed two additional stents | -240
    different puncture site | -240
    extended course of intravenous antibiotics | -240
    discharged | 792
    hospitalization 33 days | 792
    follow-up MRI 6 weeks later | 1008
    small pancreatic fluid collection | 1008
