53 years old | 0
    female | 0
    admitted to the hospital | 0
    blurred vision | 0
    retinal ischemia | 0
    cotton wool spots | 0
    macular edema | 0
    hypertensive retinopathy | 0
    1.5 g/dL monoclonal protein | 0
    immunoglobulin G (IgG) kappa type | 0
    negative hypercoagulable panel | 0
    normal blood cell counts | 0
    elevated erythrocyte sedimentation rate | 0
    elevated lactate dehydrogenase | 0
    slightly elevated creatinine (1.1 mg/dL) | 0
    total immunoglobulin G 1176 mg/dL | 0
    free light chains (FLC) ratio 28.12 | 0
    high free kappa (274 mg/L) | 0
    no monoclonal protein in 24-hour urine collection | 0
    no significant proteinuria | 0
    skeletal survey showed no lytic lesions | 0
    bone marrow aspiration and biopsy showed 10%–15% plasma cells | 0
    diagnosed with smoldering myeloma | 0
    plasma cell directed therapy recommended | 0
    started triple therapy with bortezomib, lenalidomide, and dexamethasone | -168
    acute renal failure | -168
    creatinine rise from 1.4 to 6.9 mg/dL | -168
    urinalysis showed 1+ protein | -168
    greater than five red blood cells per high power field | -168
    no casts seen | -168
    serum albumin 3.1 g/dL | -168
    negative hepatitis serologies | -168
    normal-sized kidneys | -168
    no evidence of obstruction | -168
    renal biopsy indicated | -168
    renal biopsy showing shrunken glomeruli with bloodless appearance | -168
    diffuse interstitial edema | -168
    focal mild interstitial inflammation | -168
    acute tubular injury | -168
    rare granular casts | -168
    no atypical, fractured crystalline eosinophilic casts | -168
    interstitial fibrosis | -168
    tubular atrophy | -168
    endothelial swelling | -168
    intimal edema | -168
    concentric fibroplasia | -168
    entrapped red blood cells | -168
    luminal obliteration | -168
    no definite thrombi | -168
    no fibrinoid necrosis | -168
    Congo Red stain negative for amyloid | -168
    no light chain restriction | -168
    electron microscopy confirmed absence of amyloid fibrils | -168
    subendothelial lucent widening | -168
    diffusely wrinkled glomerular basement membranes | -168
    intracytoplasmic vacuoles | -168
    loss of microvilli | -168
    acute tubular injury | -168
    no crystals or abnormal lysosomes | -168
    diagnosis of acute thrombotic microangiopathy | -168
    bortezomib discontinued | -168
    no recovery of renal function | -168
    remained dialysis-dependent | -168
    progressive decline of vision | -168
    no response to intravitreal anti-VEGF | -168
    partial response to steroids | -168
    presented with shock | 2160
    recurrent pericardial effusions | 2160
    congestive heart failure | 2160
    ejection fraction 25% | 2160
    severe left ventricular systolic dysfunction | 2160
    moderate pulmonary hypertension | 2160
    pulmonary hypertension detected two days after renal biopsy | -168
    normal ejection fraction | -168
    diagnosis of primary pulmonary hypertension | -168
    cardiac arrest | 2160
    resuscitated | 2160
    transferred to ICU | 2160
    broad antibiotic therapy started | 2160
    no clear infection source identified | 2160
    echocardiogram showed moderate pericardial effusion | 2160
    enlarged right atrium | 2160
    enlarged right ventricle | 2160
    tricuspid regurgitation | 2160
    no tamponade | 2160
    pulmonary artery systolic pressure (PASP) 85.28 mmHg | 2160
    previous PASP 52 mmHg | 2160
    left ventricular ejection fraction 60%–65% | 2160
    pericardiocentesis drained 325 mL | 2160
    negative cytopathology | 2160
    negative fluid cultures | 2160
    serum protein electrophoresis showed 0.66 g/dL monoclonal band | 2160
    IgG 1226 mg/dL | 2160
    serum kappa FLC 340.8 mg/L | 2160
    kappa/lambda FLC ratio 16.15 | 2160
    skeletal survey showed no lytic lesions | 2160
    abdominal fat pad biopsy negative for amyloid | 2160
    low C3 levels (54 mg/dL) | 2160
    normal C4 (19 mg/dL) | 2160
    normal Factor I | 2160
    normal Factor H | 2160
    ADAMTS13 activity 17% | 2160
    negative ADAMTS13 inhibitor screen | 2160
    negative antiphospholipid antibody panel | 2160
    peripheral neuropathy | 2160
    plasma VEGF negative | 2160
    negative anti-myelin associated glycoprotein antibodies | 2160
    multiple episodes of lactic acidosis | 2160
    repeated intubations | 2160
    severe right heart failure | 2160
    initiated on treprostinil | 2160
    cardiac arrest refractory to resuscitative efforts | 2160
    partial autopsy requested | 2160
    ulcer with fat layer exposure on left foot | 2160
    bilateral serous pleural effusions | 2160
    pericardial sac contained 200 mL serous fluid | 2160
    heart weighted 440 g | 2160
    no significant atherosclerosis | 2160
    no thrombi | 2160
    concentric left ventricular hypertrophy | 2160
    dilated right ventricle | 2160
    congested lungs | 2160
    spleen weighted 100 g | 2160
    subcapsular wedge-shaped infarcts | 2160
    no enlarged lymph nodes | 2160
    bilaterally atrophic kidneys | 2160
    liver weighted 1330 g | 2160
    nutmeg appearance | 2160
    severe renal interstitial fibrosis | 2160
    shrunken glomeruli | 2160
    concentric fibrointimal thickening | 2160
    splenic artery changes | 2160
    pulmonary artery changes | 2160
    myocyte hypertrophy | 2160
    minimal fibrosis | 2160
    no amyloid deposition | 2160
    centrolobular congestion and necrosis | 2160
    death | 2160

<|end_header_id|>

