35 years old | 0
female | 0
past medical history acute lymphocytic leukemia | -8784
in remission since 1997 | -8784
diabetes mellitus | 0
bipolar disorder | 0
recurrent urinary tract infections | 0
obesity | 0
status post gastric bypass surgery | 0
altered mental status | -24
bedbound for 3 months | -720
withdrawn | -720
decreased appetite | -720
poor nutrition | -720
afebrile | 0
tachycardic to 150 bpm | 0
tachypneic to 30-40 bpm | 0
hypotensive to 72/52 mm Hg | 0
severe cachexia | 0
mottled bilateral upper extremities | 0
necrotic sacral decubitus ulcer | 0
sluggish bilateral pupils | 0
right-sided downward gaze preference | 0
roving eye movements | 0
pH 7.564 | 0
PCO2 23 mm Hg | 0
PO2 67 mm Hg | 0
lactic acid of 5.3 mmol/L | 0
leukocytosis of 19.2 K/UL | 0
neutrophilic predominance | 0
sodium 137 mmol/L | 0
potassium 3.8 mmol/L | 0
blood urea nitrogen (BUN) 10 mg/dL | 0
creatinine 0.6 mg/dL | 0
albumin 1.5 g/dL | 0
total bilirubin 1.4 mg/dL | 0
direct bilirubin 0.6 mg/dL | 0
aspartate transaminase (AST) 26 IU/L | 0
alkaline phosphatase 109 IU/L | 0
alanine transaminase (ALT) 18 IU/L | 0
total protein 3.4 g/dL | 0
ammonia levels were elevated to 261umol/L | 0
negative urine toxicology | 0
unremarkable noncontract head computed tomography (CT) | 0
septic shock | 0
treated for septic shock with empiric broad-spectrum antibiotics | 0
intravenous fluids | 0
vasopressors | 0
stress-dose hydrocortisone | 0
continuous video electroencephalogram (EEG) | 0
generalized delta-range background slowing | 0
excess beta activity | 0
generalized sharply contoured waveforms with triphasic morphology | 0
Duloxetine XR 30 mg OD | 0
Gabapentin 800 mg BID | 0
Quetiapine XR 800 mg OD | 0
Alprazolam 1 mg OD | 0
Glargine 40 units OD | 0
Lispro 9 units TID | 0
acute hypoxemic respiratory failure | 48
intubation | 48
urine cultures grew ESBL E coli | 48
respiratory cultures grew ESBL E coli | 48
blood cultures were positive for M morganii | 48
stool cultures were positive for P mirablis | 48
high-dose dextrose intravenous solution | 48
lactulose | 48
rifaximin | 48
l-carnitine | 48
broad-spectrum antibiotics | 48
new seizure activity | 72
rhythmic jerking movements of her head, jaw, and tongue | 72
right downward gaze | 72
IV benzodiazepines | 72
levetiracetam | 72
second continuous video EEG | 72
near-continuous approximately 0.5 to 1.5 Hz left hemispheric posteriorly predominant blunted lateralized periodic discharges | 72
focal epilepsy | 72
severe diffuse cerebral dysfunction | 72
brain magnetic resonance imaging (MRI) | 72
diffuse gyriform restricted diffusion throughout the cerebral hemispheres and insula bilaterally | 72
elevated ammonia levels of 551 µmol/L | 72
continuous veno-venous hemodialysis (CVVHD) | 72
urine and plasma amino acids were abnormal | 72
elevated glutamine | 72
elevated glutamic acid | 72
elevated asparagine | 72
elevated urinary ornithine | 72
normal arginine | 72
normal citrulline | 72
zinc levels were not measured | 72
carnitine levels were normal | 72
acylcarnitine/carnitine ratio levels were elevated | 72
tracheostomy | 528
able to track motion with her eyes | 528
minimal responsiveness to painful stimuli | 528
death | 0