46 years old | 0 | 0 
male | 0 | 0 
admitted to the hospital | 0 | 0 
ulcerative colitis | -720 | 0 
malaise | -72 | 0 
fever | -72 | 0 
loss of appetite | -72 | 0 
chills | -72 | 0 
nausea | -72 | 0 
cardiac arrest | 0 | 0 
chest compression | 0 | 0 
tracheal intubation | 0 | 0 
ventricular fibrillation | 0 | 0 
defibrillation | 0 | 0 
adrenaline administration | 0 | 0 
Brugada syndrome | 0 | 0 
coved-type ST elevation | 0 | 0 
hypercalcemia | 0 | 0 
hypotension | 24 | 24 
septic shock | 24 | 24 
tazobactam-piperacillin administration | 24 | 168 
vasopressors administration | 24 | 168 
extubation | 48 | 48 
fever reoccurred | 120 | 120 
liver abscess | 120 | 120 
meropenem administration | 120 | 504 
vancomycin administration | 120 | 504 
puncture drainage | 120 | 504 
infection controlled | 504 | 504 
pilsicainide test | 720 | 720 
implantable cardioverter defibrillator implantation | 720 | 720 
discharged | 720 | 720 
sudden death in family history | -8760 | 0 
ectopic parathyroid adenoma | 720 | 720 
tumor resection | 720 | 720 
multiple endocrine neoplasia type 1 | 720 | 720 
nonfunctional pituitary adenoma | 720 | 720 
nonfunctional adrenal tumor | 720 | 720 
electrocardiogram taken on October 4, 2021 | -360 | -360 
electrocardiogram taken on June 28, 2021 | -420 | -420 
electrocardiogram taken on March 24, 2021 | 0 | 0 
electrocardiogram taken on September 25, 2017 | -1440 | -1440 
early repolarization | -1440 | 0 
J point elevation | -1440 | 0 
high parathyroid hormone levels | 720 | 720 
Tc scintigraphy | 720 | 720 
abnormal uptake in the anterior mediastinum | 720 | 720 
tumor in the pituitary gland | 720 | 720 
tumor in the adrenal gland | 720 | 720 
computed tomography scan | 24 | 24 
blood sample data | 24 | 24 
lactate level increased | 24 | 24 
white blood cell count increased | 24 | 24 
procalcitonin level increased | 24 | 24 
contrast-enhanced CT scan | 120 | 120 
acetaminophen administration | 0 | 0 
body temperature 40.2°C | 0 | 0 
body temperature 38.9°C | 0 | 0 
serum calcium level 14.8 mg/dL | 0 | 0 
serum calcium level 9.7 mg/dL | -360 | -360 
serum calcium level 13.8 mg/dL | -420 | -420