18 years old | 0
female | 0
hypertension | 0
syphilis | 0
type 2 diabetes | 0
mechanical fall | -720
pruritic scalp | -720
purulent drainage from sinuses on the scalp | -720
altered mental status | 0
fever | 0
heart rate of 127 bpm | 0
respiratory rate of 22 breaths/min | 0
blood pressure of 144/80 mmHg | 0
oxygen saturation of 98% on room air | 0
oriented to person and place, but not to time | 0
erythematous and edematous face, scalp and right ear | 0
large fluctuant mass with purulent drainage over the occipital and parietal portions of the scalp | 0
posterior auricular mass without signs of active drainage | 0
hyperglycemia to 700 | 0
anion gap metabolic acidosis with serum bicarbonate of 20 | 0
ketonuria | 0
extensive multifocal scalp swelling along the right temporal, right posterior parietal and left frontal regions | 0
diabetic ketoacidosis | 0
cellulitis of the scalp with concern for underlying abscesses | 0
admitted to the intensive care unit | 0
continuous infusion of insulin | 0
broad-spectrum coverage with intravenous Vancomycin and Cefepime | 0
incision and drainage of scalp lesion | 48
10-cm subgaleal abscess with large amounts of purulence evacuated | 48
initial admission blood cultures grew MRSA | 72
paranasal sinus CT with intravenous contrast did not show involvement | 72
transesophageal echocardiogram without evidence for endocarditis | 72
pulse irrigation of the wounds and sharp debridement | 96
serial bedside debridements | 96
scalp wound measured 20 cm in length, 10 cm in width and 2 cm depth | 120
right posterior auricular wound measured 7 × 7 × 2 cm | 120
wounds of the scalp and post-auricular region were definitively closed with split-thickness skin grafts | 120
100% take of the grafts on postoperative day 7 | 168
discharged on hospital day 32 | 672
intravenous Vancomycin to complete a full 7-week course | 672