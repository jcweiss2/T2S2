23 years old | 0
woman | 0
admitted to Medical Intensive Care Unit | 0
organophosphorus poisoning | 0
mechanical ventilation | 0
ionotropic support | 0
left femoral artery catheter inserted | 0
fever (102°F) | 168
tachycardia | 168
erythematous papules on left lower limb | 216
white blood cell count 16,500/mm3 | 216
neutrophils 84% | 216
lymphocytes 12% | 216
monocytes 3% | 216
eosinophils 1% | 216
blood cultures sent | 216
intra-arterial catheter removed | 216
skin lesions biopsied | 216
histopathology | 216
culture | 216
skin lesions became blackish with necrotic areas | 264
blood culture yielded Pseudomonas aeruginosa | 264
catheter tip culture yielded Pseudomonas aeruginosa | 264
skin lesion culture yielded Pseudomonas aeruginosa | 264
ceftazidime sensitive | 264
biopsy revealed acute neutrophilic infiltration | 264
perivascular area pronounced | 264
necrotic area | 264
treated with ceftazidime | 264
lesions resolved completely | 528
full recovery from organophosphorus poisoning | 528
discharged home | 528
+ Fever (102°F) | 168
+ Tachycardia | 168
+ Erythematous papules on left lower limb | 240
+ White blood cell count 16,500/mm3 | 240
+ Neutrophils 84% | 240
+ Lymphocytes 12% | 240
+ Monocytes 3% | 240
+ Eosinophils 1% | 240
+ Blood cultures sent | 240
