3 years old | 0
female | 0
admitted to the emergency department | 0
fever | 0
diarrhea | 0
abdominal pain | 0
severe dehydration | 0
critically ill | 0
pediatric intensive care unit admission | 0
feverish | 0
tachypneic | 0
rapid shallow breathing | 0
hypotensive | 0
blood pressure 60/40 mmHg | 0
severe dehydration | 0
dry tongue | 0
sunken eyes | 0
poor skin turgor | 0
oliguria | 0
pale | 0
purpuric eruption | 0
no organomegaly | 0
no lymphadenopathy | 0
pancytopenia | 0
absolute neutropenia | 0
renal impairment | 0
electrolyte imbalance | 0
hyperuricemia | 0
coagulopathy | 0
disseminated intravascular coagulation | 0
high inflammatory markers | 0
stool culture positive for Escherichia coli | 0
blood culture positive for Escherichia coli | 0
intravenous fluid therapy | 0
blood components transfusion | 0
correction of electrolyte disturbance | 0
antibiotic therapy | 0
provisional diagnosis of acute infectious gastroenteritis | 0
sepsis | 0
severe dehydration | 0
acute renal failure | 0
disseminated intravascular coagulation | 0
pelvi-abdominal ultrasound normal | 0
bone marrow aspirate | 0
hypocellular bone marrow | 0
no abnormal cells | 0
discharged | 336
follow-up visit | 504
unexplained irritability | 504
abnormal behavior | 504
hallucinations | 504
failure to recognize parents | 504
vital signs stable | 504
hematological indices normal | 504
coagulation parameters normal | 504
renal panel normal | 504
serum electrolytes normal | 504
brain imaging studies | 504
magnetic resonance imaging | 504
magnetic resonance arteriography | 504
magnetic resonance venography | 504
thrombosis in left sigmoid and transverse sinuses | 504
thrombophilia workup | 504
no thrombocytosis | 504
normal coagulation profile | 504
normal protein C and S | 504
normal antithrombin III | 504
genetic testing for thrombophilia mutations panel | 504
pediatric cardiologist assessment | 504
electrocardiogram normal | 504
echocardiography normal | 504
low molecular weight heparin | 504
discharged | 528
follow-up appointment | 528
readmitted | 672
fever | 672
pallor | 672
abdominal enlargement | 672
leukocytosis | 672
anemia | 672
thrombocytopenia | 672
peripheral smear with blast cells | 672
abdominal ultrasonography with hepatosplenomegaly | 672
bone marrow examination | 672
hypercellular bone marrow | 672
blast cells 96% | 672
immunophenotyping | 672
positive CD10 | 672
positive CD20 | 672
positive CD79a | 672
diagnosis of Common ALL | 672
induction therapy | 672
consolidation | 672
thrombophilia mutations panel result | 720
positive factor XIII V34L | 720
positive MTHFR A1298C homozygous | 720
positive factor V Leiden heterozygous | 720
follow-up MRV | 744
complete recanalization of thrombosed sinuses | 744
no new thrombi | 744
complete remission | 1008
regular follow-up | 1008
no thrombotic events | 1008
no leukemia relapses | 1008