56 years old | 0
female | 0
abnormal vaginal discharge | -336
visited a gynecologist | -336
vaginal culture | -336
cervical cytology | -336
endometrial cytology | -336
fever of 40 °C | -336
lower abdominal pain | -336
taken to the emergency room | -336
blood pressure 71/46 mmHg | -336
marked tenderness from right upper quadrant to lower abdomen | -336
fluid resuscitation therapy crystalloids 500 mL/h | -336
high procalcitonin 75.49 ng/mL | -336
abdominal CT no free air or massive ascites | -336
full stomach | -336
edema of the small intestine | -336
intra-peritoneal source of infection not detected preoperatively | -336
severe sepsis | -336
severe pan-peritonitis | -336
exploratory laparotomy | -336
purulent ascites | -336
no injury in the gastrointestinal tract | -336
uterus intact | -336
ovaries and fallopian tubes red and swollen | -336
bilateral salpingitis | -336
preserve uterine adnexa | -336
peritoneal lavage | -336
drainage | -336
administered 4000 mL crystalloid fluid | -336
poor increase in blood pressure | -336
edema of the small intestine worsened | -336
intubated | -336
managed postoperatively due to concern of worsening respiratory status | -336
noradrenaline administered | 0
intensive care | 0
intubation management started | 0
meropenem 1.5 g/day | 0
extubated | 48
noradrenaline tapered | 72
noradrenaline terminated | 72
oral intake started | 96
drainage tube removed | 96
GAS found in vaginal fluid culture | 144
GAS found in ascitic fluid culture | 144
intravenous antibiotics stopped | 144
body temperature rose to 38.1 °C | 144
oral levofloxacin prescribed | 144
discharged | 240
condition good after 2 months | 1440
infection did not recur | 1440
