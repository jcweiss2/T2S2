63 years old | 0
male | 0
admitted to the hospital | 0
history of right median nerve EHE | -72
treated with wide local excision | -72
pain along his right arm | -48
radiograph of the right elbow | -48
radiograph of the chest | -48
diagnosed with a benign muscular pathology | -48
conservative treatments | -48
pain persisted | -48
pain worsened | -24
CT scan of the right upper extremity | -12
post-surgical changes | -12
no evidence of recurrence | -12
PET-CT | -8
abnormal uptake in the right forearm | -8
no abnormal uptake in the area of pain | -8
no evidence of metastatic disease | -8
biopsy of the FDG avid area | -8
traumatic neuroma | -8
continue conservative treatments | -8
radiograph of the right upper extremity | -4
abnormality over the cortical surface | -4
new lytic lesion | -4
repeat PET-CT | 0
FDG avidity of the mid to distal right humeral shaft | 0
periosteal changes | 0
medial soft tissue mass | 0
satellite nodules in the humeral neck area | 0
CT-guided biopsy of the right humeral mass | 0
recurrence of high-grade EHE | 0
soft tissue recurrence | 0
local bone metastasis of EHE | 0
surgical resection of his tumor | 4
dyspnea on exertion | 4
lower extremity swelling | 4
difficult to take a deep breath | 4
CT imaging of the chest with angiography | 4
new interstitial-nodular opacities | 4
edema or infectious-inflammatory etiology | 4
no acute pulmonary embolism | 4
cardiac work-up | 4
unremarkable | 4
discharged home | 4
symptoms improved | 4
no longer huffing | 4
dyspnea when climbing stairs | 4
pre-anesthesia medical evaluation | 4
lungs were clear to auscultation | 4
able to lay flat without dyspnea | 4
resting oxygen saturation was 96% | 4
pre-procedure chest radiograph | 4
bilateral pulmonary opacities | 4
interstitial/septal thickening | 4
upper lung predominant fine reticulation/micronodularity | 4
surgical removal of his tumor | 8
pathology revealed high-grade EHE | 8
nodal involvement | 8
clear margins | 8
successfully extubated | 8
required supplemental oxygen | 8
chest CT angiogram | 8
segmental PE | 8
atelectasis | 8
right diaphragm paralysis | 8
worsening interstitial-nodular opacities | 8
transthoracic echocardiogram | 8
new severe right heart failure | 8
fully anticoagulated with heparin | 8
received diuretics | 8
clinical status continued to decline | 12
respiratory failure | 12
septic shock | 12
transfer to the intensive care unit | 12
intubated | 12
treated with broad spectrum antibiotics | 12
bronchoscopy | 12
bloody secretions | 12
mildly edematous airway | 12
no focal endobronchial abnormality | 12
no area of bleeding | 12
bronchoalveolar lavage | 12
negative for malignancy | 12
chest imaging | 12
diffuse alveolar filling process | 12
suspicious for alveolar hemorrhage | 12
treated empirically with high-dose steroids | 12
no response | 12
succumbed to hypoxia | 16
autopsy | 16
acute bronchopneumonia | 16
organizing fibrinous pneumonia | 16
right pulmonary artery thromboembolism | 16
EHE in a lymphangitic and intraparenchymal distribution | 16