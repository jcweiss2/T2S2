28 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
8 weeks pregnant | 0 | 0 | Factual
acute severe asthma | -10 | 0 | Factual
short non-infective prodrome | -10 | 0 | Factual
hypoxic cardiac arrest | -10 | 0 | Factual
ventricular fibrillation | -10 | 0 | Factual
resuscitation to sinus tachycardia | -10 | -10 | Factual
endotracheal intubation | -10 | -10 | Factual
therapeutically cooled to 33°C | 0 | 24 | Factual
salbutamol | 0 | 48 | Factual
ipratropium | 0 | 48 | Factual
aminophylline | 0 | 48 | Factual
hydrocortisone | 0 | 48 | Factual
magnesium | 0 | 48 | Factual
ketamine | 0 | 48 | Factual
inhalation anesthesia with 1 MAC isoflurane | 0 | 48 | Factual
severe hypercapnic acidosis | 0 | 48 | Factual
inadequate minute ventilation | 0 | 48 | Factual
neuromuscular blockade | 0 | 48 | Factual
generalised status myoclonus | 48 | 240 | Factual
absent motor response to painful stimulus | 96 | 240 | Factual
preserved pupillary reflexes | 96 | 240 | Factual
preserved corneal reflexes | 96 | 240 | Factual
preserved cough reflexes | 96 | 240 | Factual
preserved gag reflexes | 96 | 240 | Factual
spontaneously breathing | 96 | 240 | Factual
severe GSM | 96 | 240 | Factual
refractory to three antiepileptic medications | 96 | 240 | Factual
electroencephalography showed generalised periodic discharges | 96 | 240 | Factual
no discernable background rhythm | 96 | 240 | Factual
reversible causes of coma eliminated | 96 | 240 | Factual
biochemical causes eliminated | 96 | 240 | Factual
metabolic causes eliminated | 96 | 240 | Factual
septic causes eliminated | 96 | 240 | Factual
drug causes eliminated | 96 | 240 | Factual
plasma neuron-specific enolase | 240 | 240 | Factual
NSE 51 mcg/L | 240 | 240 | Factual
somatosensory-evoked potential | 240 | 240 | Factual
myoclonus motion artefacts | 240 | 240 | Factual
brain magnetic resonance imaging | 240 | 240 | Factual
bilateral basal ganglia and frontoparietal cortex infarction | 240 | 240 | Factual
severe hypoxic encephalopathy | 240 | 240 | Factual
medical consensus regarding poor prognosis | 240 | 240 | Factual
extubated | 240 | 240 | Factual
died | 264 | 264 | Factual
comfort measures | 240 | 264 | Factual