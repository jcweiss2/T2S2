severe headache | -24
right periorbital and mid-facial swelling | 0
fever | -336
headache | -336
light pain in the right ear | -336
purulent secretion from the ear | -336
swelling and redness of the skin behind the right ear | -336
tinnitus | -336
hearing disorder | -336
right acute mastoiditis | -336
treated with antibiotics | -336
treated with painkillers | -336
treated with anti-inflammatory drugs | -336
symptoms improved slightly | -192
severe headache | -192
anorexia | -192
high fever | -192
confusion | -192
admitted to hospital | 0
ophthalmological examination | 0
right facial and periorbital swelling | 0
right blepharoptosis | 0
chemosis | 0
proptosis | 0
visual acuity of 7/12 on her right eye | 0
no visual fields abnormalities | 0
intraocular pressures in both eyes were normal | 0
no relative afferent pupillary defect | 0
color vision was normal | 0
no signs of optic disc swelling | 0
febrile | 0
conscious | 0
somnolent | 0
no neurological deficits | 0
blood cultures were taken | 0
inflammatory parameters were significantly elevated | 0
renal and liver functions within normal limits | 0
tests for vasculitis were negative | 0
tests for human immunodeficiency virus (HIV) were negative | 0
tests for diabetes were negative | 0
prothrombin G20210A mutation | 0
coagulation profile was normal | 0
urinalysis was normal | 0
magnetic resonance imaging (MRI) of the brain | 0
non-opacification of the right cavernous sinus | 0
treated with high-dose intravenous Ceftriaxone | 0
treated with anticoagulation with Enoxaparin | 0
did not receive corticosteroids | 0
blood cultures were positive for Streptococcus pneumoniae | 48
continued prior antibiotic treatment | 48
developed shortness of breath | 96
reduced oxygen saturation | 96
chest X-ray revealed unilateral homogeneous opacification | 96
referred to the Intensive Care Unit (ICU) | 96
needed non-invasive mechanical ventilation | 96
antibiotics were changed to Amikacin and Piperacillin–Tazobactam | 96
symptoms resolved | 168
transferred back to our Service | 168
control contrast-enhanced magnetic resonance angiography (CE–MRA) | 168
persistence of the lacunar image in the right cavernous sinus | 168
ophthalmological symptoms improved | 168
periorbital swelling has diminished | 168
discharged | 336
on oral anticoagulant – Acenocoumarol | 336
follow-up CT venogram will indicate resolution of the thromboses | 504
full recovery | 504