47 years old | 0
male | 0
hepatitis C | 0
hemophilia A | 0
ulcerative colitis | 0
prednisone 40 mg | -240
admitted to the medical intensive care unit | 0
temperature 34.4°C | 0
heart rate 96 bpm | 0
blood pressure 107/51 | 0
respiratory rate 14 breaths per minute | 0
oxygen saturation 97% | 0
cachectic | 0
abdomen distended | 0
abdomen diffusely tender | 0
rectal examination positive for gross blood | 0
non-contrast abdomen and pelvis computed tomography scan | 0
pancolitis | 0
antibiotics started | 0
transferred to the surgical intensive care unit | 0
hypotension | 24
vasopressors | 24
respiratory failure | 24
mechanical ventilation | 24
leukocytosis | 24
lactic acidosis | 24
weaned off vasopressors | 48
extubated | 48
Clostridium difficile antigen negative | 48
antibiotics narrowed | 48
sudden onset sharp abdominal pain | 144
peritoneal signs | 144
non-contrast abdominal CT scan | 144
pneumoperitoneum | 144
colitis | 144
ascites | 144
loop ileostomy rescue procedure | 144
small bowel appeared normal | 144
ascites appeared clear | 144
extubated postoperatively | 144
supraventricular tachycardia | 216
respiratory failure | 216
mechanical ventilation | 216
hypotension | 216
vasopressors | 216
large-volume serosanguinous ascites drainage | 216
intraoperative ascites cultures grew Candida | 216
intraoperative ascites cultures grew Methicillin-resistant Staphylococcus aureus | 216
intraoperative ascites cultures grew E. coli | 216
antibiotic therapy initiated | 216
sputum cultures grew 1+ Aspergillus fumigatus | 216
repeat endotracheal aspirate culture negative | 216
non-contrast chest CT scan | 216
intubated | 216
weaned off vasopressors | 264
abdominal examination improved | 264
peritoneal signs | 336
acute hypotension | 336
vasopressors | 336
black ileostomy output | 336
bleeding from the intra-abdominal drain | 336
bright red blood per rectum | 336
emergent exploratory laparotomy | 336
small bowel necrotic | 336
seventy-three centimeters of small bowel resected | 336
primary anastomosis performed | 336
profuse intra-abdominal bleeding | 360
hemodynamically unstable | 360
massive transfusion | 360
aggressive attempts to correct coagulopathy | 360
goals of care changed to comfort measures | 360
died | 372
third ET aspirate culture positive for 2+ A. fumigatus | 372
pathologic evaluation of the resected bowel | 372
hemorrhagic gangrenous bowel | 372
granular friable ulcerated mucosa | 372
transmural bowel necrosis | 372
fungi within the bowel wall | 372
fungi within the artery wall | 372
fungi within the lumen | 372
Gomori Methenamine Silver stain characteristic of Aspergillus species | 372