78 years old | 0
male | 0
chronic obstructive pulmonary disease (COPD) | 0
prostate cancer | 0
status post radical prostatectomy | 0
subsequent radiation therapy | 0
radiation colitis | 0
presented to the emergency department | 0
recent onset shortness of breath | -48
altered mental status | -48
productive cough | -48
subjective fevers | -48
confused | -24
unable to get into bed | -24
rushed to the emergency department | 0
recent hospitalization 2 months prior | -1440
COPD exacerbation | -1440
suspected bowel obstruction | -1440
hypotensive | 0
blood pressure 92/61 | 0
tachycardic | 0
heart rate 130 | 0
tachypneic | 0
respiratory rate 25 | 0
hypoxic | 0
oxygen saturation 71% | 0
afebrile | 0
temperature 99.9°F (37.7°C) | 0
alert | 0
oriented | 0
diminished breath sounds | 0
scattered crackles | 0
noninvasive positive pressure ventilation with BiPAP | 0
leukocytosis | 0
white blood cell 30.6 | 0
12% bands | 0
lactic acidosis | 0
lactic acid 3.6 mmol/l | 0
acute kidney injury | 0
creatinine 1.5 mg/dl | 0
chest X-ray left upper and lower lobe opacity | 0
pneumonia severity index 131 | 0
Class V management strategy | 0
mortality 27%-31.1% | 0
admitted to the intensive care unit | 0
acute on chronic hypoxic hypercapnic respiratory failure | 0
left-sided pneumonia | 0
intubation | 24
mechanical ventilation | 24
broad-spectrum antibiotics vancomycin | 0
piperacillin-tazobactam | 0
azithromycin | 0
healthcare-associated pneumonia (HCAP) | 0
blood cultures positive for P. multocida | 48
ownership over five cats | 0
deep involvement in cat care and grooming | 0
no scratch or bite marks | 0
no signs of skin infection or abscess | 0
antibiotic regimen switched to ampicillin-sulbactam | 48
clinical status improved | 168
successful extubation | 168
discharge | 432
extended care facility | 432
amoxicillin-clavulanic acid | 432
14 days of antibiotic therapy | 432
