Here is the table of events and timestamps:

79 years old | 0
male | 0
hypertension | 0
ischemic heart disease | 0
scheduled for elective TAVR | 0
severe symptomatic aortic stenosis | 0
coronary artery bypass graft surgery | -11
mitral valve repair | -11
transthoracic echocardiography | -11
aortic valve area 0.6 cm2 | -11
transvalvular max and mean gradients 61 and 33 mm Hg | -11
left ventricular ejection fraction 45% | -11
right transcarotid approach | 0
fluoroscopic and transesophageal echocardiographic guidance | 0
TAVR procedure | 0
TAVR procedure duration 1 hour | 1
SAPIEN 3 valve deployed | 1
postprocedural TEE | 1
prosthesis in good position | 1
no visible paravalvular leak | 1
gastric aspiration with orogastric tube | 1
blood-tinged secretions | 1
extubated in the operating room | 1
transferred to the intensive care unit | 1
progressive chest pain | 2
shivering | 2
computed tomography (CT) | 2
pneumomediastinum | 2
right hydropneumothorax | 2
esophageal perforation suspected | 2
right thoracic drain inserted | 2
serosanguinous liquid drained from the pleural space | 2
300 milliliters | 2
esophagogastroscopy | 2
4-cm vertical perforation of the middle third of the esophagus | 2
returned to the operating room | 9
right thoracotomy and repair of an esophageal perforation | 9
lysis of extensive pleural adhesions | 9
esophageal laceration site | 9
large vertebral osteophyte | 9
primary closure of the esophageal wall in two layers | 9
intercostal muscular flap mobilized | 9
three thoracic drains left in place | 9
transferred to the intensive care unit | 9
pneumonia | 9
severe delirium | 9
congestive heart failure with pulmonary edema | 9
withdrawal of care | 30
death | 30