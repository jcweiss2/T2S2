55 years old | 0
African American | 0
male | 0
admitted to the hospital | 0
alcohol withdrawal symptoms | 0
headache | 0
tremors | 0
sweating | 0
chronic pulmonary obstructive disease | -8760
alcohol dependence | -17520
denied history of liver disease | 0
denied sleep disturbances | 0
denied memory changes | 0
denied seizures | 0
stable vital signs | 0
anxious | 0
tremulous | 0
slow and delayed response to questions | 0
unsteady gait | 0
scleral icterus | 0
skin icterus | 0
gynecomastia | 0
bibasilar crackles | 0
liver edge palpable 3cm below costal margin | 0
asterixis | 0
nail clubbing | 0
non-pitting edema of the legs | 0
macrocytic anemia | 0
hemoglobin 11.3 g/dl | 0
Mean Corpuscular Volume (MCV) 101.8 fL | 0
platelet count 83,000/μL | 0
total protein 8.2 g/dL | 0
albumin 2.8 g/dL | 0
total Bilirubin 3.9 mg/dL | 0
Aspartate Aminotransferase (AST) 69 U/L | 0
Alanine Aminotransferase (ALT) 36 U/L | 0
ammonia level 124 mcg/dl | 0
International Normalized Ratio (INR) 1.6 | 0
early cirrhosis | 0
chlordiazepoxide-based alcohol withdrawal protocol | 0
lactulose for hepatic encephalopathy | 0
300 mg of chlordiazepoxide | -72
good control of withdrawal symptoms | -72
mental status deteriorated | 240
upgraded to intensive care unit | 240
urine drug screen positive for benzodiazepines | 240
repeat ammonia level 121 mcg/dl | 240
septic work-up unremarkable | 240
diagnosis of benzodiazepine-induced hepatic encephalopathy | 240
single dose of flumazenil 1mg | 240
improvement of mental status | 240
effect short-lived | 240
repeated single doses of flumazenil | 240
flumazenil drip at 0.25 mg/hour | 240
persistent nausea | 240
treated with ondansetron | 240
flumazenil well tolerated | 240
attempts to decrease infusion rate | 240
deterioration of mental status | 240
repeated urine benzodiazepine testing positive | 240
flumazenil drip for 28 days | 240
tapered off successfully | 672
mental status returned to normal | 672
repeat urine benzodiazepine test negative | 672
discharged home | 672