23 years old|0
    female|0
    admitted to the hospital|0
    labor pains of gradually increasing intensity|0
    denied fever symptoms|0
    denied shortness of breath|0
    denied cough|0
    denied sore throat|0
    initial temperature 37°C|0
    BP 138/89 mm Hg|0
    heart rate 103 beats/min|0
    external OS 2 cm|0
    premature rupture of membrane|0
    meconium-stained liquor|0
    fetal distress|0
    hemoglobin 10.2gm%|0
    COVID Rapid Antigen Test positive|0
    mild cough for the last seven days|0
    not vaccinated with first dose of Covishield|0
    cervix unsuitable for normal vaginal delivery|0
    emergency caesarean section|0
    healthy live born male neonate|0
    baby weighed 2.86 kg|0
    routine RT PCR test not done|0
    baby transferred to nursery|0
    blood sent for matching|0
    1 unit B+ blood transferred to mother|0
    postpartum hemorrhage developed|24
    heavy vaginal bleeding|24
    probable cause atonicity of uterus|24
    Inj carboprost|24
    tranexamic acid|24
    Inj methergine|24
    IV syntocinon|24
    per rectal misoprostol|24
    PPH persisted|24
    BP 106/64 mmHg|24
    respiratory rate 17 per min|24
    heart rate 120 beats per minute|24
    abdomen reopened|24
    uterus flabby|24
    devascularization performed|24
    bilateral uterine and ovarian arteries located|24
    B4lynch suture done|24
    uterus partially contracted|24
    abdomen closed|24
    2 litres of blood lost|24
    3 units B+ blood transfused|24
    sent to COVID HDU ward|24
    oral feeding started|40
    slight respiratory distress|48
    O2 saturation dropped to 92%|48
    blood sent for investigation|48
    managed with IV piperacillin/tazobactam|48
    IV metronidazole|48
    Inj pantoprazole|48
    Tab ivermectin|48
    Tab montelukast|48
    Tab cetirizine|48
    Inj ondansetron|48
    Tab zinc|48
    Tab vitamin C|48
    Capsules vitamin D|48
    Infusion paracetamol|48
    Tab paracetamol|48
    1 unit blood transfused|72
    condition gradually improved|72
    no need for tracheal intubation|72
    O2 saturation maintained 96–98%|72
    abdominal stitches removed|192
    repeat blood report on 10th day|240
    D-Dimer 9.78 mg/L|240
    C-Reactive Protein 129 mg/L|240
    WBC count 16200 /μL|240
    Haemoglobin 8.2 g/dL|240
    Interleukin 49.7 pg/mL|240
    Ferritin 224.1 ng/mL|240
    RT PCR negative|336
    discharged|360
    
    <|eot_id|>
    23 years old|0
    female|0
    admitted to the hospital|0
    labor pains of gradually increasing intensity|0
    denied fever symptoms|0
    denied shortness of breath|0
    denied cough|0
    denied sore throat|0
    initial temperature 37°C|0
    BP 138/89 mm Hg|0
    heart rate 103 beats/min|0
    external OS 2 cm|0
    premature rupture of membrane|0
    meconium-stained liquor|0
    fetal distress|0
    hemoglobin 10.2gm%|0
    COVID Rapid Antigen Test positive|0
    mild cough for the last seven days|0
    not vaccinated with first dose of Covishield|0
    cervix unsuitable for normal vaginal delivery|0
    emergency caesarean section|0
    healthy live born male neonate|0
    baby weighed 2.86 kg|0
    routine RT PCR test not done|0
    baby transferred to nursery|0
    blood sent for matching|0
    1 unit B+ blood transferred to mother|0
    postpartum hemorrhage developed|24
    heavy vaginal bleeding|24
    probable cause atonicity of uterus|24
    Inj carboprost|24
    tranexamic acid|24
    Inj methergine|24
    IV syntocinon|24
    per rectal misoprostol|24
    PPH persisted|24
    BP 106/64 mmHg|24
    respiratory rate 17 per min|24
    heart rate 120 beats per minute|24
    abdomen reopened|24
    uterus flabby|24
    devascularization performed|24
    bilateral uterine and ovarian arteries located|24
    B4lynch suture done|24
    uterus partially contracted|24
    abdomen closed|24
    2 litres of blood lost|24
    3 units B+ blood transfused|24
    sent to COVID HDU ward|24
    oral feeding started|40
    slight respiratory distress|48
    O2 saturation dropped to 92%|48
    blood sent for investigation|48
    managed with IV piperacillin/tazobactam|48
    IV metronidazole|48
    Inj pantoprazole|48
    Tab ivermectin|48
    Tab montelukast|48
    Tab cetirizine|48
    Inj ondansetron|48
    Tab zinc|48
    Tab vitamin C|48
    Capsules vitamin D|48
    Infusion paracetamol|48
    Tab paracetamol|48
    1 unit blood transfused|72
    condition gradually improved|72
    no need for tracheal intubation|72
    O2 saturation maintained 96–98%|72
    abdominal stitches removed|192
    repeat blood report on 10th day|240
    D-Dimer 9.78 mg/L|240
    C-Reactive Protein 129 mg/L|240
    WBC count 16200 /μL|240
    Haemoglobin 8.2 g/dL|240
    Interleukin 49.7 pg/mL|240
    Ferritin 224.1 ng/mL|240
    RT PCR negative|336
    discharged|360