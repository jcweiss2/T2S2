32 years old | 0
female | 0
lymphangioleiomyomatosis | -8760
multiple lymphangioleiomyomas in the retroperitonium | -8760
repeated spontaneous pneumothoraces | -8760
drainage | -8760
low ejection fraction | -720
intubated | -720
ventilated | -720
respiratory failure | -720
bronchopneumonia | -720
multiresistant Pseudomonas aeruginosa | -720
sepsis | -720
disseminated intravascular coagulopathy | -720
severe bleeding from the nose | -720
severe bleeding from the hypopharynx | -720
severe bleeding from the lower respiratory tract | -720
mechanical ventilation | -720
venovenous ECMO (VV-ECMO) | -720
arteriovenous ECMO (AV-ECMO) | -720
cannulation of the vena jugularis interna dextra | -720
cannulae from the VV-ECMO | -720
arterial cannula | -720
ascending aorta | -720
donor lungs | -144
sequential bilateral lung transplant | 0
clamshell incision | 0
severely hypokinetic right and left ventricles | 0
large thrombus in the left atrium | 0
pulmonary veins | 0
diffuse bleeding | 0
coagulopathy | 0
10 L blood loss | 0
AV-ECMO | 0
poor myocardial function | 0
sternotomy | 0
severe pulmonary edema | 6
continuous leakage of edematous fluid | 6
endotracheal tube | 6
tidal volumes | 6
peak pressure | 6
positive end-expiratory pressure | 6
cardiovascular support | 6
high-dose norepinephrine | 6
arterial blood gas | 6
good oxygenation | 6
immunosuppression therapy | 6
tacrolimus | 6
mycophenolate mofetil | 6
corticosteroids | 6
anticoagulation | 6
heparin | 6
activated coagulation time (ACT) | 6
thrombi in both left and right atria | 6
thrombolysis | 6
alteplase | 6
pulmonary artery | 6
rescue procedure | 6
left atrial thrombus | 8
second dose of alteplase | 8
pulmonary edema | 8
resolution | 8
full dose of thrombolytic agent | 24
no further thrombi | 24
lung function | 24
improvement | 24
radiological findings | 24
acute kidney injury | 48
continuous renal replacement therapy | 48
heart function | 48
improvement | 48
ECMO support | 192
stop | 192
sternotomy | 192
closure | 192
P. aeruginosa infection | 192
resolution | 192
weaning | 192
rehabilitation | 192
poor muscle strength | 192
transbronchial biopsy | 192
tissue rejection | 192
A 1–2 | 192
pulses of steroids | 192
loss of consciousness | 192
posterior reversible encephalopathy syndrome | 192
electroencephalograph | 192
epileptic status | 192
antiepileptic medications | 192
stenosis of the right main bronchus | 2160
biodegradable stent | 2160
ELLA-CS s.r.o. | 2160
pulmogenic sepsis | 2160
multiorgan failure | 2160
continuous renal replacement therapy | 2160
extubation | 4320
rehabilitation | 4320
discharge | 5040
good quality of life | 5040
no signs of stenosis | 5040
stationary spirometric values | 5040
FEV1 38% | 5040