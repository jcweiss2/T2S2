21 years old | 0
female | 0
admitted to the hospital | 0
low-grade fever | -72
abdominal pain | -168
conscious | 0
anxious | 0
pale | 0
blood pressure on the lower side of normal | 0
distended abdomen | 0
tuberculosis ruled out | 0
vasculitis ruled out | 0
erect X-ray normal | 0
abdomen ultrasonography normal | 0
septic shock | 72
altered sensorium | 72
intubated | 72
transferred to ICU | 72
magnetic resonance imaging of head normal | 72
cerebrospinal fluid study normal | 72
serum sodium level normal | 72
leukocytosis | 72
anemia | 72
thrombocytopenia | 72
deranged liver function tests | 72
echocardiography showed mild diastolic dysfunction | 72
ejection fraction >60% | 72
noradrenaline infusion started | 72
vasopressin infusion started | 72
broad-spectrum antibiotics started | 72
platelet transfusion | 72
packed cell transfusion | 72
repeat ultrasonography of the abdomen showed thickened and dilated nonobstructed bowel loops | 120
coarse hepatic echo-texture | 120
gastro surgeon refused active management | 120
high nasogastric aspirates | 120
feed intolerance | 120
prokinetics used | 120
started accepting nasogastric feeds | 144
enteral feed started | 144
rapidly rising intraabdominal pressure | 144
deterioration in hemodynamics | 144
increasing metabolic acidemia | 144
hyponatremia | 144
passed large amounts of fresh blood-mixed loose stools | 144
bedside abdominal ultrasonography suspected presence of air shadows within the hepatic portal vein | 144
CT scan abdomen showed pneumatosis intestinalis | 144
gas in portal venous system | 144
exploratory laparotomy | 144
multiple areas of gangrenous patches | 144
dusky discoloration of the jejunum | 144
air bubbles in the subserosa | 144
major mesenteric vessels pulsating | 144
no evidence of thrombus | 144
no atherosclerosis | 144
no visible occlusion | 144
no bowel perforation | 144
surgical incisions in the wall of the jejunum | 144
succumbed | 148
postmortem examination not conducted | 148