22 years old | 0
male | 0
admitted to the hospital | 0
fever | -360
escharotic skin lesions | -360
purpuric skin lesions | -360
ibuprofen administration | -240
diclofenac sodium administration | -240
cephalosporin antibiotics administration | -96
alcoholism history | -1752
severe obesity | 0
black necrotic eschar | 0
subcutaneous nodules | 0
enlarged lymph nodes | 0
purpuric and necrotic crusted lesions | 0
thrombosis in small saphenous vein | 0
thrombosis in bilateral great saphenous vein | 0
thrombosis in cephalic vein | 0
large fresh cerebral infarction | 0
intracranial infection | 0
lung infection | 0
pleurisy | 0
pericardial effusion | 0
elevated WBC count | 0
elevated neutrophils | 0
elevated lymphocytes | 0
elevated monocytes | 0
elevated eosinophils | 0
thrombocytopenia | 0
elevated PT | 0
elevated APTT | 0
elevated D-dimer | 0
decreased fibrinogen | 0
decreased antithrombin III | 0
skin lesion pain | 24
back pain | 24
headache | 24
vertigo | 24
sputum-free cough | 24
diarrhea | 24
stomach ache | 24
abdominal pain | 168
hematemesis | 168
blood in stool | 168
gastrointestinal bleeding | 168
multiple pulmonary emboli | 168
liver damage | 168
hepatic vein thrombosis | 168
portal vein thrombosis | 168
splenic vein thrombosis | 168
superior mesenteric vein thrombosis | 168
inguinal swelling | 168
difficulty breathing | 240
irritability | 240
decreased blood oxygen saturation | 240
respiratory failure | 240
sedative administration | 240
subclavian vein catheterization | 240
hypernutrition administration | 240
liver function damage | 240
renal function damage | 240
hypokalemia | 240
hyperchloremia | 240
hypernatremia | 240
metabolic acidosis | 240
coma | 240
continuous renal replacement therapy | 480
consciousness improvement | 480
tar-like stools | 480
occult blood positive | 480
platelet increase | 480
oxygen mask administration | 480
returned to dermatology | 528
elevated blood chloride | 576
decreased oxygen partial pressure | 576
decreased HGB | 576
femoral artery catheterization | 576
radial artery catheterization | 576
central venous catheterization | 576
active bloody stools | 720
bruise on right upper limb | 720
fever | 864
decreased HGB | 864
red liquid in gastric tube | 984
palpitations | 984
shortness of breath | 984
convulsions | 984
worsened breathing difficulty | 1056
oxygen saturation decrease | 1056
thoracentesis catheter drainage | 1056
tracheal intubation | 1056
mechanical ventilation | 1056
improved condition | 1248
normal body temperature | 1344
returned to dermatology | 1344
varicose veins in stomach | 1368
chronic gastritis | 1368
splenic infarction | 1584
resolved portal vein thrombosis | 1608
resolved hepatic vein thrombosis | 1608
resolved inferior vena cava thrombosis | 1608
reduced thigh skin lesions | 1608
softened skin texture | 1608
resolved purpura lesions | 1608
stable vital signs | 1608
stable laboratory indicators | 1608
weight loss | 1608
discharged | 1608
increased WBC count | 0
increased eosinophils | 0
decreased AT | 0
decreased serum protein | 0
decreased albumin | 0
elevated transaminase | 0
elevated bilirubin | 0
elevated bile acids | 0
elevated muscle enzymes | 0
elevated creatinine | 0
elevated uric acid | 0
elevated fasting glucose | 0
elevated serum iron | 0
proteinuria | 0
fecal occult blood | 0
decreased protein C | 0
negative autoantibodies | 0
decreased complement C3 | 0
elevated C-reactive protein | 0
Klebsiella pneumoniae infection | 0
Stenotrophomonas maltophilia infection | 0
human herpesvirus type 5 infection | 0
oral Candida infection | 0
epidermal serous callus | 0
liquefaction degeneration | 0
vascular stenosis | 0
fibrinoid necrosis | 0
inflammatory thrombosis | 0
collagen necrosis | 0
adipose hyperplasia | 0
fat cell necrosis | 0
inflammatory cell infiltration | 0
continuous renal replacement therapy | 0
mechanical ventilation | 0
plasma infusion | 0
clotting factor infusion | 0
RBC apheresis | 0
platelet apheresis | 0
antibiotics administration | 0
glucocorticoids administration | 0
IVIG administration | 0
hemostatic agents | 0
acid suppression | 0
liver protection | 0
AIPF diagnosis | 0
acute cellulitis | 0
sepsis | 0
DIC | 0
multiple organ failure | 0
acute gastrointestinal bleeding | 0
acute respiratory distress | 0
pulmonary embolism | 0
cerebral infarction | 0
portal vein thrombosis | 0
splenic infarction | 0
deep vein thrombosis | 0
liver damage | 0
no bleeding points found | 168
no special bronchoscopy findings | 240
no Mycobacterium tuberculosis | 0
no mycoplasma/chlamydia | 0
no fungal detection | 0
no parasite detection | 0
no dsDNA pathogens | 0
no ssDNA pathogens | 0
no EBV/CMV DNA | 0
no Gram-positive bacteria in blood | 240
no growth in urine culture | 168
no growth in stool culture | 168
negative fungal microscopy | 168
negative fecal occult blood | 480
negative sputum microscopy | 168
negative G/GM tests | 240
