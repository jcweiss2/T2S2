14 years old | 0
male | 0
admitted to the hospital | 0
fever | -24
pain in the left side of the hip | -24
denies any injuries | 0
denies medical problems | 0
denies intake of any medications | 0
denies previous hospitalizations | 0
denies recent tours | 0
family history unremarkable | 0
temperature 38℃ | 0
blood pressure 110/70 mmHg | 0
heart rate 88/min | 0
respiratory rate 22/min | 0
tenderness over the lateral aspect of the left side of the hip | 0
hemoglobin level 14.6 g/dL | 0
WBC count 6,400/mm3 | 0
neutrophils 79% | 0
platelet count 176,000/mm3 | 0
ESR 12 mm/h | 0
CRP 3.1 mg/dL | 0
hip radiography no abnormal findings | 0
pelvic CT no abnormal findings | 0
transient synovitis considered | 0
antibiotics not prescribed | 0
body temperature risen to 38.9℃ | 72
pain at the sacroiliac joint on the FABERE test | 72
hip MRI scan showed synovitis and capsulitis | 72
empiric administration of vancomycin | 72
empiric administration of ceftriaxone | 72
condition deteriorated | 120
fever 40.4℃ | 120
respiratory rate >40/min | 120
difficulty breathing | 120
ABGA pH 7.399 | 120
ABGA pCO2 32.7 mmHg | 120
ABGA PO2 52.7 mmHg | 120
ABGA O2 Sat 88% | 120
dyspnea | 120
oxygen supply via a nasal cannula | 120
respiratory status worsened | 144
ABGA PaO2/FiO2 137 mmHg | 144
bilateral lower lobe infiltrates on chest radiographs | 144
bilateral and symmetric compartmental consolidation on chest CT | 144
ARDS diagnosed | 144
synchronized intermittent mandatory ventilation | 144
tidal volume 360 mL | 144
FiO2 40% | 144
PEEP 12 cmH2O | 144
WBC count 2,400/mm3 | 144
platelet count 58,000/mm3 | 144
ESR 40 mm/h | 144
CRP 13.8 mg/dL | 144
blood cultures yielded E. cloacae | 144
antibiotic regimen changed to ceftriaxone and amikacin | 144
methylprednisolone administration initiated | 144
defervescence occurred | 120
need for ventilatory support reduced | 120
breathing room air | 168
pain in the left side of the hip lessened | 168
discharged from ICU | 168
follow-up chest radiograph showed improvement | 240
parenteral antimicrobial therapy maintained | 240
methylprednisolone tapered | 240
repeat hip MRI scan showed improvement | 312
repeat blood culture grew no bacteria | 96
discharged from hospital | 1104
serum immunoglobulin normal | 1104
serum complement levels normal | 1104
no further tests for immunologic disorder | 1104