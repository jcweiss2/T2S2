40 years old | 0
    African-American woman | 0
    chronic eczema | 0
    previous alcohol abuse | 0
    gout | 0
    hypothyroidism | 0
    presented with worsening eruption | 0
    presented with intermittent diarrhea | 0
    cutaneous eruption began | -1440
    desquamation of the hands | -1440
    desquamation of the feet | -1440
    desquamation of the perioral skin | -1440
    desquamation of the perineal skin | -1440
    associated pain | -1440
    associated swelling | -1440
    concurrent hair loss | -1440
    increasing weakness | -5760
    fatigue | -5760
    intermittent diarrhea | -5760
    70 pounds unintentional weight loss | -5760
    1 to 2 glasses of wine a day | 0
    smoking | 0
    no significant family history | 0
    not on any medications | 0
    dermatologic examination found erythematous desquamative patches | 0
    erosions | 0
    crusted lesions involving distal fingers of both hands | 0
    left dorsal arm involvement | 0
    sacrum involvement | 0
    perineum involvement | 0
    left medial leg involvement | 0
    bilateral distal feet involvement | 0
    predilection for acral interdigital web spaces | 0
    diffuse nonscarring alopecia of the scalp | 0
    scaling patches on the vermillion lips | 0
    punch biopsy of the left medial thigh | 0
    psoriasiform epidermal spongiosis | 0
    slight superficial perivascular lymphohistiocytic infiltrate | 0
    diffuse hypogranulosis | 0
    broad overlying parakeratosis | 0
    ballooning degeneration of the spinous layer | 0
    nutritional deficiency dermatitis | 0
    methicillin-resistant Staphylococcus aureus sepsis | 0
    Escherichia coli sepsis | 0
    secondary to pneumonia | 0
    admitted to the intensive care unit | 0
    required ventilator respiratory support | 0
    systemic antibiotics | 0
    laboratory studies ruled out necrolytic acral erythema | 0
    imaging studies ruled out necrolytic acral erythema | 0
    laboratory studies ruled out pellagra | 0
    imaging studies ruled out pellagra | 0
    laboratory studies ruled out biotin deficiency | 0
    imaging studies ruled out biotin deficiency |' 0
    zinc levels low (28 μg/dL) | 0
    antitransglutaminase antibodies positive | 0
    antiendomysium antibodies positive | 0
    diagnosis of celiac disease | 0
    diagnosis of zinc deficiency | 0
    denied current alcohol abuse | 0
    history of excessive alcohol intake | 0
    chronic low zinc levels | 0
    deficiency dermatitis | 0
    distal duodenal biopsy | 0
    focal villi blunting | 0
    Brunner's gland hyperplasia | 0
    no significant intraepithelial lymphocytes | 0
    treated with gluten-free diet | 0
    treated with zinc sulfate 220-mg oral capsule twice daily | 0
    resolution of gastrointestinal symptoms | 168
    resolution of cutaneous symptoms | 168
    