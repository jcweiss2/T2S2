67 years old | 0
male | 0
admitted to the intensive care unit | 0
suspected sepsis | 0
alpha-hemolytic isolate from blood culture | 0
Gram stain revealed characteristic lanceolate diplococci | 0
capsule staining by India ink was positive for pneumococci | 0
optochin sensitivity test | 0
bile solubility test | 0
inulin fermentation test | 0
optochin-resistant | 0
bile soluble | 0
inulin fermentation positive | 0
identification by VITEK II | 0
identification by MALDI-TOF | 0
detection of lytA gene | 0
detection of ply gene | 0
synonymous single nucleotide polymorphism type of functional mutation in lytA gene | 0
treatment with ceftriaxone | 0
discharged | 24
complete recovery | 24
Gene sequencing | 0
lytA gene sequencing | 0
ply gene sequencing | 0
atp C, atpA and part of atp B from S. pneumoniae | -120
acquisition of atp C, atpA and part of atp B from S. pneumoniae | -120
open reading frame ant in 2 optochin sensitive viridians streptococci | -120
Southern blotting technique | -120
comparisons of the chromosomal framework of the atp operon regions | -120
nucleotide sequence of the atpC-atpA-atpB region | -120
recombinant origin of optochin-sensitive viridians streptococci | -120
point mutations in either a- or c-subunit of the H + ATPase | -120
optochin MICs 4- to 30-fold higher than susceptible isolates | -120
pneumolysin detection | -120
atypical presentation of pneumococci | -120
diminishing reliability of optochin sensitivity | -120
diminishing relevance of traditional optochin sensitivity testing | -120
optochin-resistant pneumococci | -120
bile insoluble S. pneumoniae isolates | -120
nontypeable, unencapsulated pneumococci | -120
optochin sensitivity testing | -120
sensitivity and specificity of optochin sensitivity testing | -120
patient consent | 0
financial support | 0
conflicts of interest | 0