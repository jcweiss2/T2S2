38 years old | 0
male | 0
admitted to the hospital | 0
complaining of long-term problems with food intake | 0
previous surgery for congenital pylorostenosis in childhood | -10000
native X-ray examination | -120
ultrasound examination | -120
CT scan | -120
suspicion of gastrostasis | -120
contrast-enhanced examination of the upper gastrointestinal tract | -120
barium sulphate as the contrast agent | -120
stenosis of the pylorus with gastrostasis | -120
repeated X-ray after 30 min | -90
stasis of all the contrast agent in the stomach | -90
suspected benign stenosis of the pylorus | -120
planned surgical intervention | -120
unplanned return to the surgeon’s office | 120
complaining of substantial and increasing pain in left epigastrium | 120
tender left epigastric region | 120
considerable pain on palpation | 120
X-ray examination | 120
evidence of the stasis of a large amount of contrast agent in the stomach | 120
inflammation parameters not elevated | 120
admitted to the surgery ward | 120
nasogastric tube inserted | 120
unsuccessful attempt to evacuate the contrast agent | 120
deterioration of the patient’s condition | 120
immediate laparotomy | 144
tumorous lesion on the pylorus | 144
dilated stomach and adhesions | 144
mobilizing the stomach and duodenum | 144
precipitated and sedimented barium sulphate scooped out | 144
BII partial stomach resection | 144
Roux-en-Y gastrojejunal anastomosis | 144
repeated lavage of the peritoneal cavity | 144
Tygon tube 27 drainage inserted | 144
intense antibiotics therapy initiated | 144
infusions and nutritional support | 144
worsening of the patient’s condition | 168
elevation of inflammation markers | 168
suspected leak of the anastomosis or contrast agent spillage with peritonitis | 168
CT scan | 168
no contrast agent spillage intraperitoneally and no anastomosis failure | 168
methylene blue administered through the nasogastric tube | 168
drained exudate observed for signs of methylene blue | 168
no hint of methylene blue | 168
drainage bags contained 200 mL of sanguinolent fluid | 168
another CT exam | 216
small amount of contrast agent identified in the paragastric intraperitoneal region | 216
previous CT exam reviewed | 216
same amount of contrast agent identified next to the stomach | 216
active leak not suspected | 216
laboratory results worsening | 216
increase in inflammation parameters | 216
sepsis suspected | 216
patient remained afebrile | 216
anastomosis dehiscence repeatedly unconfirmed on CT exams | 216
surgical revision not performed | 216
antibiotic therapy revised | 216
vasopressor support introduced | 216
improvement of the patient’s condition | 240
therapy with antibiotics and vasopressors continued | 240
amount of exudate drained significantly lower | 240
surgical wound dehiscent and phlegmonous | 240
local therapy applied | 240
stools being passed | 336
vasopressors discontinued | 336
inflammation parameters improved | 336
discharged | 336
histological exam of the resected tissue | 336
diagnosis of malignant stenosis of the pylorus | 336
resection margin positive for carcinoma | 336
repeated resection with the revision of the anastomosis | 504
surgical wound healed per secundam | 504
referred to the department of clinical oncology | 504
chemotherapy initiated | 504
last PET/CT exam | 1000
no metastatic lesions | 1000