65 years old | 0
    male | 0
    admitted to the hospital | 0
    melena | -24
    altered mental status | -24
    confusion | -24
    incoherent speech | -24
    progressive somnolence | -24
    profuse diarrhea | -24
    dark tarry stools | -24
    soiled clothing | -24
    no fevers | -24
    no chills | -24
    no abdominal pain | -24
    no nausea | -24
    no vomiting | -24
    chronic hepatitis C | 0
    polysubstance abuse | 0
    no recent travel | 0
    chronic alcoholism | -1680
    binge drinking | -1680
    blood pressure 125/100 mmHg | 0
    pulse 135 beats per minute | 0
    temperature 99.2ºF | 0
    O2 saturation 91% | 0
    respiratory rate 18 breaths per minute | 0
    dry mucous membranes | 0
    partially healed wound | 0
    surrounding erythema | 0
    no crepitus | 0
    no fluctuance | 0
    no jaundice | 0
    negative Murphy’s sign | 0
    lethargic | 0
    somnolent | 0
    Glasgow Coma Scale 8 | 0
    intubated | 0
    increased creatinine | 0
    decreased hemoglobin | 0
    cirrhosis | 0
    heterogeneous liver | 0
    nodular liver | 0
    portal hypertension | 0
    enlarged portal vein | 0
    gastric varices | 0
    cellulitis | 0
    no abscess | 0
    no gas formation | 0
    IV octreotide | 0
    packed red blood cells | 0
    platelets | 0
    broad-spectrum antibiotics | 0
    tachycardia | 0
    leukocytosis | 0
    SIRS | 0
    elevated lactate | 0
    hepatic encephalopathy | 0
    respiratory failure | 0
    bleeding varices | 0
    decompensated cirrhosis | 0
    admitted to ICU | 0
    upper endoscopy | 0
    non-bleeding esophageal varices | 0
    non-bleeding gastric varices | 0
    band ligation | 0
    no further melena | 0
    extubated | 72
    return to baseline mentation | 72
    dog bite | -504
    subjective fevers | -504
    subjective chills | -504
    blood culture positive | 0
    Pasteurella multocida | 0
    IV ceftriaxone | 0
    discharged | 360