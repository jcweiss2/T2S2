20 years old | 0
pregnant woman | 0
26 weeks gestation | 0
anti-epileptic therapy | -672
carbamazepine | -672
consumption of 4000 mg carbamazepine | -4
denied concomitant overdose | 0
gastric lavage | -4
transferred to hospital | -4
presentation | 0
glasgow coma score 3/15 | 0
pulse rate 138/min | 0
blood pressure 110/70 mmHg | 0
respiratory rate 25/min | 0
capillary blood glucose 109 mg/dl | 0
pupils dilated 6 mm bilaterally | 0
reacting to light | 0
deep tendon reflexes sluggish | 0
Babinski sign negative | 0
systemic examination unremarkable | 0
intubated | 0
multi-dose activated charcoal therapy | 0
shifted to ICU | 0
serum carbamazepine > 20 μg/ml | 0
hemoglobin 8 g/dl | 0
white count 15200/cumm | 0
renal function normal | 0
liver function test normal | 0
coagulation profile normal | 0
circulatory shock | 6
fluid resuscitation | 6
low dose vasopressors | 6
empiric antibiotic therapy | 6
discontinued antibiotics | 72
negative cultures | 72
low procalcitonin 0.34 | 72
absence of definite infection focus | 72
episodes of hypoglycemia | 72
managed with 50% dextrose bolus | 72
25% dextrose infusion | 72
hypoglycemia resolved | 144
other causes ruled out | 72
serum carbamazepine 17.3 μg/ml | 72
serum carbamazepine 2.97 μg/ml | 168
extubated | 168
vasoactive agents weaned | 168
serum carbamazepine normalized | 168
no further hypoglycemic episodes | 1344
