89 years old | 0
    male | 0
    atrial fibrillation | -4320
    valvular heart disease | -4320
    hypertension | -4320
    mitral bioprosthesis | -4320
    tricuspid valvuloplasty | -4320
    warfarin | -4320
    bisoprolol | -4320
    ramipril | -4320
    furosemide | -4320
    INR over 2 | -4320
    tested positive for SARS-CoV-2 | -240
    fever | -168
    cough | -168
    amoxicillin | -168
    spiramycin | -144
    azithromycin | -144
    admitted to emergency department | 0
    epistaxis | 0
    major bleeding | 0
    hypoxemia | 0
    pulse oxygen saturation 80% | 0
    systolic blood pressure 105 mmHg | 0
    diastolic blood pressure 59 mmHg | 0
    cardiac rate 104 per minute | 0
    INR > 10 | 0
    D-dimer 400 ng/mL | 0
    B-type natriuretic peptide 81 pg/mL | 0
    high-sensitivity troponin T 10 ng/L | 0
    ground-glass opacity | 0
    crazy paving | 0
    air space consolidation | 0
    dilatation of the colon | 0
    vitamin K administered | 0
    simple compression therapy | 0
    bleeding stopped | 0
    factor V 166 IU/dL | 0
    alanine aminotransferase 38 IU | 0
    aspartate aminotransferase 36 IU/L | 0
    fibrinogen 7.6 g/L | 0
    transferred to ICU | 0
    dexamethasone | 0
    cefotaxime | 0
    azithromycin continued | 0
    vitamin K administrations | 72
    INR fluctuations | 72
    enoxaparin | 168
    INR below 2 | 168
    hypoxemia worsened | 168
    D-dimer > 12000 ng/mL | 168
    acute proximal bilateral pulmonary embolism | 168
    NT-proBNP 2022 ng/L | 168
    high-sensitivity troponin T 48.9 ng/L | 168
    tinzaparin | 216
    discharged from ICU | 384
    oxygen therapy 2 L/min | 384
    clinical condition worsened | 432
    bacterial pneumonia | 432
    fever | 432
    increased biological inflammatory syndrome | 432
    new radiological infiltrates | 432
    broad-spectrum antibiotic therapy | 432
    septic shock | 504
    died | 504
    