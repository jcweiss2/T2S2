64 years old | 0
female | 0
right flank pain | -24
dysuria | -24
pollakuria | -24
diabetes | -672
hypertension | -672
hypothyroidism | -672
right renal pelvic stone | -24
PNL | 0
general anesthesia | 0
ureteral catheter placement | 0
nephrostomy tube placement | 0
respiratory distress | 0.75
hypotension | 0.75
hemorrhage | 0.75
hemoglobin 13 g/dl | -24
hemoglobin 11 g/dl | 0
hemoglobin 8.1 g/dl | 0.75
blood transfusion | 1
erythrocyte suspension transfusion | 1
fresh frozen plasma transfusion | 1
hemoglobin 10 g/dl | 2
AST elevation | 24
ALT elevation | 24
LDH elevation | 24
AST peak | 96
ALT peak | 96
LDH peak | 96
AST normalization | 192
ALT normalization | 192
LDH normalization | 192
discharge | 216
ischemic hepatitis diagnosis | 48
liver necrosis | 48
centrilobular hepatocytes damage | 48
hypoperfusion | 48
elevated serum aminotransferases | 48
elevated LDH | 48
normal serum bilirubin | 48
normal INR | 48
systemic hypotension | 0.75
hemorrhage after PNL | 0.75
insufficient hepatic perfusion | 48
routine serum biochemical parameters evaluation | 216