48 years old | 0
male | 0
admitted to the hospital | 0
nausea | -96
diffuse abdominal pain | -96
general weakness | -96
anorexia | -96
indigestion | -96
gastric ulcer perforation | -96
gastric cardia cancer | -96
peritoneal tumor seeding | -96
hypoactive bowel sounds | 0
direct tenderness in the epigastric area | 0
white blood cell counts 12.5 × 10^3/µL | 0
erythrocyte sedimentation rate 38 mm/h | 0
C-reactive protein 16.93 mg/dL | 0
free T4, T3, and T4 Levels exceeded the normal range | 0
thyroid stimulating hormone levels were below the normal range | 0
peritonitis | 0
gastric malignancy | 0
peritoneal carcinomatosis | 0
distal gastrectomy with Billroth II anastosis | 0
emergent surgery | 0
thyroid storm | 48
body temperature 41.3 °C | 48
tachycardia | 48
irritability | 48
abdominal pain | 48
Glasgow Coma Scale score of E3V1M5 | 48
severe pain | 48
propylthiouracil 800 mg | 48
intravenous glucocorticoids 40 mg | 48
oral acetaminophen 650 mg | 48
oral Lugol’s solution 1.5 mL | 48
bladder irrigation with cold saline | 48
hypothermic blanket | 72
propylthiouracil dose increased to 1200 mg/d | 72
PTU dose fixed at 200 mg, q6hd | 96
Lugol’s solution 0.5 mL, q8hd | 96
vital signs were stable | 192
clear mental status | 96
oral PTU dose decreased to 200 mg three times daily | 360
discharged | 696
asymptomatic status | 696
stable vital signs | 696