79 years old | 0
female | 0
admitted to the hospital | 0
high fever | -72
involuntary weight loss | -72
vomiting | -72
severe pain in the upper right abdomen | -72
diabetes | -672
hypertension | -672
atrial fibrillation | -672
cholestasis | -672
underweight | 0
BMI 17.8 kg/m2 | 0
fever | 0
nausea | 0
lack of appetite | 0
severe pain | 0
ciprofloxacin | 0
metronidazole | 0
intravenous rehydration therapy | 0
intravenous 0.5% glucose | 0
spasmolytic drugs | 0
gallbladder enlargement | 0
gallstones | 0
common bile duct expansion | 0
pancreas with finely inhomogeneous echostructure | 0
low concentrations of potassium | 0
low concentrations of phosphate | 0
low concentrations of magnesium | 0
respiratory failure | 72
cardiac failure | 72
enteral feeding | 72
confusion | 72
tachycardia | 72
respiratory insufficiency | 72
severe hypotension | 72
refeeding syndrome | 72
rapid fluid supplementation | 72
oxygen supplementation | 72
dopamine | 72
severe alterations of electrolytes | 72
severe alterations of vitamins | 72
hydric balance dysfunction | 72
parenteral feeding | 96
mild recovery | 96
oral feeding | 120
phosphorus supplementation | 120
potassium supplementation | 120
magnesium supplementation | 120
thiamine supplementation | 120
clinical improvement | 312
decrease in body temperature | 312
normalization of laboratory parameters | 312
low ejection fraction | 312
bilateral pleural effusion | 312
resumed eating | 336
hemodynamic status stabilized | 336
vasopressor therapy discontinued | 336
electrolyte imbalance disappeared | 336
discharged | 360