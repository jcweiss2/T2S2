38 years old | 0
man | 0
presented to the hospital | 0
abdominal pain | -3
nausea | -3
discharged from the hospital | -504
hospital course for COVID-19 pneumonia | -672
endotracheal intubation | -672
ventilatory support | -672
CT PE study | -672
no evidence of PE | -672
previous medical history significant for PE at age 16 | -168
PE provoked by trauma | -168
treated with 6 months of warfarin | -168
remained well until age 30 | -168
diagnosed with second PE | -168
chronic thromboembolic pulmonary hypertension | -168
thromboendarterectomy | -168
started on long-term warfarin therapy | -168
regular INR checks | -168
close follow-up visits | -168
hypercoagulable work-up after second PE negative | -168
reported with medication regimen | 0
INR levels consistently therapeutic | 0
blood pressure 129/86 mm Hg | 0
heart rate 99 bpm | 0
respiratory rate 16/min | 0
temperature 100.4 °F | 0
obesity | 0
moderate bilateral symmetrical lower extremity edema | 0
remained hemodynamically stable | 0
unremarkable basic metabolic panel | 0
negative high sensitivity troponins | 0
platelets within normal limit | 0
elevated white cell count 12.94×10^9/L | 0
INR therapeutic range | 0
PT elevated to 34.7 s | 0
PTT normal at 37.4 s | 0
CT abdomen | 0
no abnormalities in abdomen | 0
incidental finding of possible filling defect in dilated descending right pulmonary artery | 0
dedicated chest imaging with CTPE | 0
large filling defect within descending right main pulmonary artery | 0
filling defect not visualized during initial admission | 0
not evident on studies prior to COVID-19 infection | 0
echocardiogram | 0
dilated right atrium | 0
bowing of interatrial septum | 0
increased RA pressure 8 mm Hg | 0
severely dilated right ventricle | 0
severely reduced systolic function | 0
diastolic and systolic LV septal flattening | 0
dilated inferior vena cava | 0
lower extremity Doppler ultrasounds | 0
no deep vein thrombosis | 0
periumbilical abdominal pain | 0
nausea | 0
fever | 0
elevation in white cell count | 0
white cell count resolved by day 2 | 48
no diarrhea | 0
Clostridium difficile screen negative | 0
blood cultures negative | 0
CT abdomen and pelvis no infectious source | 0
stress ulcers considered | 0
no signs of gastrointestinal bleeding | 0
negative fecal occult blood test | 0
stable hemoglobin values | 0
acute pancreatitis ruled out | 0
normal serum amylase | 0
normal serum lipase | 0
normal appearance of pancreas on CT | 0
abdominal symptoms resolved | 0
fevers resolved | 0
leukocytosis resolved | 0
PE ruled in | 0
consideration of anticoagulation failure | 0
transiently on unfractionated intravenous heparin therapy | 0
decision to continue warfarin with higher INR target range | 0
advised to follow with hematology | 0
consideration of enoxaparin therapy after weight loss | 0
outcome decision to remain on warfarin | 0
close follow-up | 0
postdischarge attempts for follow-up | 0
no response to follow-up reminders | 0
recurrent pulmonary embolism | 0
COVID-19 disease | 0
therapeutic anticoagulation | 0
hypercoagulable state associated with COVID-19 | 0
challenges with treatment | 0
recurrent thrombosis despite therapeutic anticoagulation | 0
