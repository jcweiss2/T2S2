31 years old | 0
female | 0
pancreas-kidney transplant | -7872
diabetic nephropathy | -7872
End stage renal disease | -7872
chronic renal graft dysfunction | -1314
hemodialysis | -1314
PermCath | -1314
immunosuppressive therapy | -1314
mycophenolate | -1314
tacrolimus | -1314
prednisolone | -1314
type 1 diabetes | -7872
hypertension | -7872
bronchial asthma | -7872
glaucoma | -7872
depression | -7872
fever | -72
shortness of breath | -72
dry cough | -72
shivering | -72
high-grade fever | -72
admitted to hospital | 0
mild chest discomfort | 0
temperature 39.4 °C | 0
pulse 112 beats/min | 0
respiratory rate 24 breaths/min | 0
oxygen saturation 90% | 0
blood pressure 138/75 mmHg | 0
white blood cells 9.44 × 10^3/μL | 0
red blood cells 3.46 × 10^6/mcL | 0
hemoglobin 9.0 g/dL | 0
neutrophils 86% | 0
lymphocytes 8% | 0
absolute neutrophil count 7.17 × 10^3/mcL | 0
red cell distribution width 18.0 | 0
serum creatinine 541 μmol/L | 0
urea 11.66 mmol/L | 0
potassium 4.85 mmol/L | 0
sodium 139 mmol/L | 0
phosphorus 2.24 mmol/L | 0
eGFR 8.4 mL/min/1.73 m^2 | 0
total protein 51 g/L | 0
albumin 23.3 g/L | 0
C-reactive protein 78.0 mg/L | 0
procalcitonin 3.25 μg/L | 0
D-dimer 1.40 mg/L | 0
random blood sugar 7.5 mmol/L | 0
HbA1C 6.7% | 0
arterial blood gas pH 7.349 | 0
pCO2 40.9 mmHg | 0
pO2 115.4 mmHg | 0
HCO3 22.0 mmol/L | 0
chest CT widespread diffuse patchy areas | 0
ground glass veiling | 0
air space consolidations | 0
strandy reticulo-nodular infiltrates | 0
chest x-ray bilateral extensive multifocal pulmonary opacities | 0
line related sepsis | 0
immunosuppressive treatment curtailed | 0
tacrolimus 2 mg twice daily | 0
mycophenolate withheld | 0
prednisolone 20 mg/day | 0
empiric antibiotic therapy | 0
vancomycin 1 g every 48 h | 0
meropenem 500 mg every 24 h | 0
amikacin 400 mg every 48 h | 0
RT-PCR for COVID-19 | 0
blood culture | 0
pulmonology team consulted | 0
bronchoscopy refused | 0
chills | 168
shivering | 168
high-grade fever | 168
desaturating | 168
non-rebreather mask | 168
high-flow nasal cannula | 168
intensive care unit | 168
non-invasive continuous positive airway pressure | 168
hemodialysis | 168
repeat blood cultures | 168
sputum cultures | 168
TB workup | 168
oxygen requirements increased | 168
chest x-ray bilateral extensive multi-lobar air space filling | 168
ground glass opacities | 168
Pneumocystis pneumonia treatment | 192
trimethoprim/sulfamethoxazole | 192
vancomycin stopped | 192
meropenem stopped | 192
sputum analysis | 192
Pneumocystis jirovecii | 192
high-grade fever | 360
condition deteriorated | 360
pan-culture | 360
vancomycin | 360
meropenem | 360
yeast cells | 360
anidulafungin | 360
loading dose 200 mg | 360
maintenance dose 100 mg daily | 360
tachypneic | 360
respiratory rate 40/min | 360
severe respiratory distress | 360
chest X-ray | 360
extensive bilateral multifocal ground glass opacities | 360
obscured costophrenic angles | 360
severe hypoxemia | 360
intubated | 360
mechanical ventilation | 360
bradycardia | 360
asystole | 360
cardiopulmonary resuscitation | 360
advanced cardiac life support | 360
death | 360
blood culture | 432
Cryptococcus neoformans | 432