56 years old | 0
male | 0
admitted to the hospital | 0
dyspnea | -336
productive cough | -336
increasing dyspnea | -336
increasing productive cough | -336
blood pressure 127/93 mmHg | 0
heart rate 99 beats/min | 0
temperature 86.6°F | 0
respiratory rate 28/min | 0
97% saturation on 2L O2 | 0
anxious | 0
jugular venous distention | 0
bilateral rales | 0
wheezing | 0
regular cardiac rhythm | 0
no murmurs | 0
no S3 | 0
no S4 | 0
left lower extremity below the knee amputation | 0
right lower extremity with 1+ pitting edema | 0
furosemide 80 mg IV | 0
nebulized bronchodilator therapy | 0
methylprednisolone 125 mg IV | 0
respiratory status rapidly declined | 2
shock | 2
multisystem organ failure | 2
hypoxemic respiratory failure | 2
hypercapnic respiratory failure | 2
intubated | 2
vasopressor therapy | 2
nonischemic cardiomyopathy | -10000
left ventricular ejection fraction of 20%–25% | -10000
biventricular implantable cardioverter defibrillator | -10000
CarboMedics bi-leaflet mechanical aortic valve | -10000
paroxysmal atrial fibrillation | -10000
warfarin | -10000
intermittent noncompliance | -10000
labile INR values | -10000
chronic hypertension | -10000
hyperlipidemia | -10000
tobacco abuse | -10000
1.5 ppd use | -10000
chronic kidney disease stage IIIb | -10000
non-insulin-dependent diabetes mellitus | -10000
major depressive disorder | -10000
history of psychotic features | -10000
suicidal ideation | -10000
recurrent noncompliance | -10000
acute decompensated heart failure | 0
pulmonary thromboembolism | 0
decompensated chronic pulmonary disease | 0
cor pulmonale | 0
septic shock | 0
prosthetic valve dysfunction | 0
infectious endocarditis | 0
acute coronary syndrome | 0
transthoracic echocardiogram | 2
mechanical aortic valve stenosis | 2
peak velocity of 4.7 m/s | 2
acceleration time of 110 ms | 2
mean gradient of 52 mmHg | 2
Doppler velocity index of 0.25 | 2
mild aortic regurgitation | 2
Swan-Ganz placement | 4
intra-aortic balloon pump insertion | 4
fluoroscopy | 4
fixed nonmobile leaflet | 4
presumed thrombosis | 4
alteplase 10 mg IV bolus | 4
alteplase 90 mg IV infusion | 4
heparin infusion | 4
aPTT 1.5–2.0 times the control value | 4
serial transthoracic echocardiograms | 24
improvement of mechanical aortic valve function | 24
peak velocity of 3.6 m/s | 24
mean pressure gradient of 35 mmHg | 24
repeat fluoroscopic evaluation | 48
normal bi-leaflet motion | 48
successful thrombolysis | 48
restoration of function | 48
extubated | 72
discharged | 168
follow-up transthoracic echocardiogram | 2160
normal functioning mechanical aortic valve | 2160
peak velocity of 2.3 m/s | 2160
mean pressure gradient of 11 mmHg | 2160