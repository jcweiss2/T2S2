5 years old | 0
male | 0
admitted to the hospital | 0
fever | -48
neck pain | -48
odynophagia | -48
headache | -48
nasal congestion | -48
lethargy | -48
no cough | -48
no abdominal pain | -48
no vomiting | -48
no diarrhea | -48
no rash | -48
no sick contacts | -48
no recent travel | -48
COVID-19 infection | -336
unvaccinated against COVID-19 | -336
tachycardia | 0
fever | 0
full range of motion of the neck | 0
no respiratory distress | 0
no stridor | 0
shotty posterior cervical lymphadenopathy | 0
elevated inflammatory biomarkers | 0
lymphopenia | 0
mild hyponatremia | 0
rapid antigen testing for group A Streptococcus | 0
nasopharyngeal polymerase chain reaction (PCR) for SARS-CoV-2 | 0
influenza A and B | 0
respiratory syncytial virus | 0
blood cultures | 0
X-ray of the neck | 0
paravertebral soft tissue swelling | 0
computed tomography (CT) of the neck | 0
retropharyngeal phlegmonous changes | 0
possible early abscess | 0
bilateral reactive lymphadenopathy | 0
dexamethasone | 0
intravenous (IV) ampicillin–sulbactam | 0
maintenance IV fluids | 0
pediatric ear, nose, and throat (ENT) consultation | 0
persistent high-grade fevers | 24
tachycardia | 24
tachypnea | 24
worsening tachycardia | 72
worsening tachypnea | 72
borderline hypotension | 72
fluid resuscitation | 72
ongoing fevers | 72
softer voice | 72
facial edema | 72
increased pain with neck motion | 72
new prominent cardiac gallop | 72
1+ soft pulses | 72
mild hepatomegaly | 72
elevated CRP | 72
IV Vancomycin | 72
repeat CT neck | 72
retropharyngeal phlegmon | 72
persistent reactive cervical lymphadenopathy | 72
CT chest | 72
bilateral pleural effusions | 72
subsegmental atelectasis | 72
periportal edema | 72
mediastinal lymphadenopathy | 72
epinephrine infusion | 78
high-flow nasal cannula | 78
cardiac echocardiogram | 78
mild biventricular systolic dysfunction | 78
mild four-chamber dilated chambers | 78
positive SARS-CoV-2 serologies | 78
elevated troponin | 78
elevated brain natriuretic peptide (BNP) | 78
elevated D-dimer | 78
elevated ferritin | 78
elevated fibrinogen | 78
elevated international normalized ratio (INR) | 78
intravenous immune globulin (IVIG) | 78
methylprednisolone | 78
enoxaparin | 78
clinical status improvement | 126
laboratory findings improvement | 126
imaging findings improvement | 126
discharged | 192
prednisolone taper | 192
amoxicillin–clavulanate | 192
aspirin | 192
repeat cardiac echo | 336
normal cardiac function | 336
normal coronary arteries | 336