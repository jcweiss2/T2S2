60 years old | 0
male | 0
hypertension | -672
left ventricular dysfunction | -672
beta-blockers | -672
sartanic | -672
tiazidic diuretic | -672
chest pain | -4
alerted the emergency department | 0
morphine | 0
apirine | 0
dopamine infusion | 0
transferred to the nearest peripheral hospital | 0
angiographic study | 1
severe cardiogenic shock | 1
catecholamine | 1
IABP support | 1
angioplasty | 1
heparin bolus | 1
reopro | 1
bradi-asystolic cardiac arrest | 2.5
tracheal intubation | 2.5
transvenous pacing | 2.5
resuscitation manoeuvres | 2.5
cardiogenic shock | 2.5
high amines dosage | 2.5
IABP | 2.5
pacing | 2.5
mechanical ventilation | 2.5
anuria | 2.5
paO2 | 2.5
paCO2 | 2.5
pH | 2.5
lactates | 2.5
base excess | 2.5
echocardiography examination | 2.5
contractile reserve | 2.5
ECMO team | 3.5
percutaneous cannulation | 4.15
ECMO implantation | 4.15
perfusionist | 4.15
ECMO circuit | 4.15
blood flow | 4.15
gas flow | 4.15
FiO2 | 4.15
hemodynamic stabilization | 4.15
reduction of amines | 4.15
recovery of diuresis | 4.15
normalization of blood gas parameters | 4.15
reopro infusion | 4.15
transport to the cardiac surgery intensive care unit | 5.5
sedated | 5.5
muscle relaxant | 5.5
therapeutic hypothermia | 5.5
arterial catheter | 5.5
central venous catheter | 5.5
pulmonary artery catheter | 5.5
hemodynamic data | 5.5
dobutamine | 5.5
heparin infusion | 5.5
aspirin | 5.5
clopidogrel | 5.5
transe-sophageal echocardiography | 24
ejection fraction | 24
calcium-sensitizer | 72
weaning from ECMO | 72
reduction of blood flow | 72
Swan-Ganz catheter | 72
echocardiography | 72
cannulae removal | 96
hyperdynamic shock | 96
norepinephrine | 96
septic shock | 96
cultural examination | 96
empiric antibiotic therapy | 96
meropenem | 96
IABP removal | 120
nitrates | 120
echocardiography | 120
linezolid | 120
fever | 120
elevation of leukocytes | 120
inflammation indexes | 120
bronchial bleeding | 120
deterioration of blood gas parameters | 120
high PEEP | 120
heparin interruption | 120
clopidogrel interruption | 120
ecodoppler | 120
hypertensive crisis | 144
pulmonary oedema | 144
high pulmonary pressures | 144
mechanical ventilation | 144
PEEP | 144
FiO2 | 144
inhalatory nitric oxide | 144
negative water balance | 144
calcium-sensitizer | 144
diastolic dysfunction | 144
ACE-inhibitor | 144
beta-blockers | 144
extubation | 216
digoxin | 240
transfer to the hospital | 480
discharge | 480