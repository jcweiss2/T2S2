fever | -240
cough | -240
dyspnoea | -120
aggravated dyspnoea | -120
admission to hospital | 0
conscious of foetal movement | -196
foetal movement | -196
urine pregnancy test positive | -280
natural conception | -280
recurrent fever | -240
highest body temperature 39.2 ℃ | -240
decreased to normal after oral acetaminophen | -240
cough | -240
yellow viscous sputum | -240
chest distress | -240
shortness of breath | -240
no chills | -240
worsened symptoms | -120
dyspnoea | -120
admitted to hospital | 0
body temperature 36.4 ℃ | 0
blood pressure 117/87 mmHg | 0
heart rate 130 beats/min | 0
respiratory rate 20 times/min | 0
cyanosis of the lip | 0
thick breathing sounds in both lungs | 0
dry and wet rales in the right lower lung | 0
heart rate regular | 0
no noises heard in the auscultation area of each valve | 0
gestational and symmetric abdominal type | 0
height 166 cm | 0
pre-pregnancy weight 46.5 kg | 0
body mass index 16.87 | 0
weight gain 8.8 kg during pregnancy | 0
uterine height 34 cm | 0
abdominal circumference 89 cm | 0
contractions sporadic and weak | 0
head presentation | 0
foetal heart sounds 142 beats/min | 0
intrapelvic and extrapelvic measurements normal | 0
pH 7.472 | 0
partial pressure of carbon dioxide 34.0 mmHg | 0
partial pressure of oxygen 56 mmHg | 0
sulfur dioxide 88.6% | 0
C-reactive protein 186.33 mg/L | 0
erythrocyte sedimentation rate 69.00 mm/h | 0
procalcitonin 2.24 ng/mL | 0
White blood cell 18.29 × 10^9/L | 0
neutrophil % 90.10% | 0
lymphocyte 0.97 × 10^9/L | 0
Alkaline phosphatase 232 U/L | 0
total bilirubin 23.1 μmol/L | 0
albumin 33.9 g/L | 0
K+ 2.93 mmol/L | 0
sodium 129 mmol/L | 0
chloride 89 mmol/L | 0
cardiac markers normal | 0
D-dimer 3.50 mg/L | 0
chest computed tomography multiple plaques | 0
miliary foci | 0
nodular foci with partial consolidation and cavities | 0
obstetric ultrasound single viable foetus | 0
head presentation | 0
oligohydramnios | 0
cardiac ultrasound no significant abnormalities | 0
lower extremity vascular ultrasound no significant abnormalities | 0
caesarean section | 24
oxyhemoglobin saturation increased to 95%-98% | 24
high-flow nasal cannula oxygen therapy | 24
fraction of inspired oxygen 100% | 24
flow rate 50 L/min | 24
assisted ventilation by endotracheal intubation | 48
empirical antibiotic therapy | 48
meropenem | 48
vancomycin | 48
symptomatic treatment of fluid and ALB infusion | 48
irrigation solution collected and tested for metagenomic next-generation sequencing | 48
S. aureus combined with novel coronavirus infection | 48
no acid-fast bacilli in the sputum tuberculosis smear | 48
tubercle bacillus-polymerase chain reaction negative | 48
nontuberculosis mycobacterium-PCR negative | 48
galactomannan experiments normal | 48
vancomycin 1 g every 12 h | 72
meropenem 1 g every 8 h | 72
anticoagulant therapy | 72
treatments to relieve the cough and reduce the amount of sputum | 72
nasal tube oxygen with a flow rate of 3-4 L/min | 96
chest CT multiple areas of inflammation in both lungs | 96
mildly enlarged mediastinal lymph nodes | 96
small amount of bilateral pleural effusion | 96
CRP 38.54 mg/L | 96
WBC count 8.25 × 10^9/L | 96
PCT 0.129 ng/mL | 96
potassium 4.04 mmol/L | 96
D-dimer 2.44 mg/L | 96
TB-PCR negative | 96
chest CT inflammatory lesions | 216
pleural effusion absorbed | 216
antibiotics adjusted to sitafloxacin 50 mg twice daily | 216
discharged from hospital | 264
chest CT multiple lung inflammation absorbed | 720
chest CT multiple lung inflammation apparently absorbed | 744