49 years old|0
    male|0
    admitted to the hospital|0
    fever|-72
    chills|-72
    diarrhea|-72
    acute pancreatitis|-26280
    fatty liver|-26280
    liver cirrhosis|-432
    mild ascites|-432
    esophageal variceal ligation|-432
    acute variceal bleeding|-432
    alcohol consumption|0
    intermittently seditious|0
    confused|0
    disoriented|0
    yellowish skin|0
    shifting dullness positive|0
    moderate lower limb edema|0
    body temperature 38.7 °C|0
    heart rate 100 beats per minute|0
    blood pressure 100/54 mmHg|0
    WBC 6.0 × 10^9/L|0
    GR% 68.5%|0
    Hb 69 g/L|0
    TBIL 126.8 μmol/L|0
    DBIL 61.5 μmol/L|0
    ALT 37.39 U/L|0
    AST 54.7 U/L|0
    γ-GGT 72.05 U/L|0
    ALB 29 g/L|0
    BUN 9.77 mmol/L|0
    Cr 67.8 μmol/L|0
    PT 30.7 s|0
    INR 2.90|0
    procalcitonin 25.24 ng/mL|0
    PaO2 79 mmHg|0
    FiO2 29.0%|0
    pneumonia|0
    hydrothorax|0
    splenomegaly|0
    cholecystitis|0
    ascites|0
    right renal calculus|0
    ACLF grade 1|0
    Child-Pugh score 12|0
    MELD score 25.4|0
    ademetionine|0
    L#Ornithine#L#Aspartate|0
    montmorillonite powder|0
    bifidobacterium lactobacillus tripterygium|0
    ceftriaxone sodium|0
    fever persisted 38.5 °C|12
    blood pressure 59/23 mmHg|12
    heart rate 110 beats per minute|12
    oliguria 200 mL urine|12
    septic shock|12
    epidermal staphylococcus|12
    gram-positive bacteria|12
    WBC 9.9 × 10^9/L|12
    GR% 84.4%|12
    Hb 63 g/L|12
    TBIL 138.6 μmol/L|12
    DBIL 85.5 μmol/L|12
    AST 40.51 U/L|12
    γ-GGT 63.38 U/L|12
    BUN 15.76 mmol/L|12
    Cr 143.56 μmol/L|12
    PT 33.6 s|12
    INR 3.25|12
    AKI stage 2|12
    ACLF grade 2|12
    red blood cell transfusion|12
    dopamine|12
    meropenem|12
    terlipressin|12
    hematemesis 450 mL dark red blood|19
    esomeprazole|19
    somatostatin|19
    human albumin|19
    nutritional support|19
    blood pressure 86/57 mmHg|72
    heart rate 110 beats per minute|72
    body temperature 37 °C|72
    WBC 5.4 × 10^9/L|72
    GR% 78.4%|72
    Hb 94 g/L|72
    TBIL 155.9 μmol/L|72
    DBIL 90.4 μmol/L|72
    AST 32.52 U/L|72
    γ-GGT 52.3 U/L|72
    BUN 10.27 mmol/L|72
    Cr 42.04 μmol/L|72
    improved GR%|96
    improved C-reaction protein|96
    improved procalcitonin|96
    improved Cr|96
    improved urine volume|96
    no hematemesis|96
    no melena|96
    fecal occult blood test negative|312
    WBC 11.1 × 10^9/L|312
    GR% 65.5%|312
    Hb 84 g/L|312
    Cr 54.56 μmol/L|312
    C-reaction protein 16.5 mg/L|312
    procalcitonin 0.03 ng/mL|312
    no ACLF|312
    discharged|312
    mild distension of abdomen|2016
    mild lower limb edema|2016
    Hb 87 g/L|2016
    TBIL 77.4 μmol/L|2016
    DBIL 40.9 μmol/L|2016
    AST 54.77 U/L|2016
    ALT 28.05 U/L|2016
    γ-GGT 61.07 U/L|2016
    ALB 30.6 g/L|2016
    BUN 5.36 mmol/L|2016
    Cr 36.79 μmol/L|2016
    PT 19.7 s|2016
    INR 1.67|2016
    furosemide|2016
    spironolactone|2016

    