76 years old | 0
    female | 0
    hypertension | 0
    dyslipidaemia | 0
    intermittent palpitations | -336
    orthopnoea | -336
    New York Heart Association functional class III–IV shortness of breath | -336
    admitted to hospital for decompensated heart failure | 0
    uncontrolled atrial fibrillation | 0
    left bundle branch block | 0
    clinical evidence of decompensated heart failure | 0
    pulmonary oedema | 0
    bilateral pleural effusions | 0
    intravenous diuresis | 0
    furosemide 80 mg intravenous once | 0
    furosemide infusion 20 mg/h | 0
    metoprolol 5 mg intravenous once | 0
    oral metoprolol | 0
    intravenous digoxin load | 0
    increasingly diaphoretic | 24
    tachycardic | 24
    hypotensive 60/30 mmHg | 24
    high-sensitivity troponin 2040 ng/L | 24
    serum lactate 7.1 mmol/L | 24
    anuric acute kidney injury | 24
    serum creatinine 122 μmol/L | 24
    dual antiplatelet therapy | 0
    ASA 81 mg orally daily | 0
    clopidogrel 75 mg orally daily | 0
    fondaparinux 2.5 mg subcutaneously daily | 0
    vasopressors | 0
    significant biventricular systolic dysfunction | 0
    plethoric non-collapsible inferior vena cava | 0
    diastolic flattening of the interventricular septum | 0
    intubated for emergent cardiac catheterization | 24
    epinephrine | 24
    norepinephrine | 24
    vasopressin | 24
    left main coronary artery ectatic | 24
    left anterior descending ectatic | 24
    left circumflex arteries ectatic | 24
    right coronary artery emptying into pulmonary artery | 24
    transthoracic echocardiogram severe RV systolic dysfunction | 24
    right atrial dilatation | 24
    severe tricuspid regurgitation | 24
    positive cultures Streptococcus bovis | 24
    empiric antibiotics | 24
    Piperacillin/Tazobactam 4.5 g IV every 6 h | 24
    Vancomycin 1 g IV every 12 h | 24
    Doxycycline 100 mg orally twice daily | 24
    intermittent haemodialysis | 168
    transoesophageal echocardiogram dilated left main coronary artery | 168
    dilated right coronary artery draining into pulmonary artery | 168
    no vegetations | 168
    anomalous right coronary artery from the pulmonary artery diagnosis | 168
    reviewed at interdisciplinary heart team rounds | 168
    turned down for surgical intervention | 168
    bacteremic Streptococcus bovis | 192
    ceftriaxone | 192
    metronidazole | 192
    extubated | 216
    transferred to cardiology ward | 216
    dependent on intermittent haemodialysis | 216
    transferred to hospice care | 960
    deceased | 1800
    no flow-limiting stenoses | 24
    no murmurs | 0
    no rubs | 0
    no gallops | 0
    no prior electrocardiogram for comparison | 0
    no vegetations | 168
    no intra-cardiac left-to-right shunt | 24
    no pulmonary embolus | 24
    no fistula involving RVOT | 24
    no regional wall motion abnormalities | 24
    no gastrointestinal malignancy ruled out | 192
    no mechanical complication with RV infarction ruled out | 24
    no underlying cardiomyopathy ruled out | 24
    no pulmonary hypertension ruled out | 24
    no massive pulmonary embolism ruled out | 24
    no catecholaminergic state confirmed | 24
    no sepsis ruled out | 24
    no reversibility of disease | 192
    no surgical intervention | 168
    <|eot_id|>
    76 years old | 0
female | 0
hypertension | 0
dyslipidaemia | 0
intermittent palpitations | -336
orthopnoea | -336
New York Heart Association functional class III–IV shortness of breath | -336
admitted to hospital for decompensated heart failure | 0
uncontrolled atrial fibrillation | 0
left bundle branch block | 0
clinical evidence of decompensated heart failure | 0
pulmonary oedema |1 0
bilateral pleural effusions | 0
intravenous diuresis | 0
furosemide 80 mg intravenous once | 0
furosemide infusion 20 mg/h | 0
metoprolol 5 mg intravenous once | 0
oral metoprolol | 0
intravenous digoxin load | 0
increasingly diaphoretic | 24
tachycardic | 24
hypotensive 60/30 mmHg | 24
high-sensitivity troponin 2040 ng/L | 24
serum lactate 7.1 mmol/L | 24
anuric acute kidney injury | 24
serum creatinine 122 μmol/L | 24
dual antiplatelet therapy | 0
ASA 81 mg orally daily | 0
clopidogrel 75 mg orally daily | 0
fondaparinux 2.5 mg subcutaneously daily | 0
vasopressors | 0
significant biventricular systolic dysfunction | 0
plethoric non-collapsible inferior vena cava | 0
diastolic flattening of the interventricular septum | 0
intubated for emergent cardiac catheterization | 24
epinephrine | 24
norepinephrine | 24
vasopressin | 24
left main coronary artery ectatic | 24
left anterior descending ectatic | 24
left circumflex arteries ectatic | 24
right coronary artery emptying into pulmonary artery | 24
transthoracic echocardiogram severe RV systolic dysfunction | 24
right atrial dilatation | 24
severe tricuspid regurgitation | 24
positive cultures Streptococcus bovis | 24
empiric antibiotics | 24
Piperacillin/Tazobactam 4.5 g IV every 6 h | 24
Vancomycin 1 g IV every 12 h | 24
Doxycycline 100 mg orally twice daily | 24
intermittent haemodialysis | 168
transoesophageal echocardiogram dilated left main coronary artery | 168
dilated right coronary artery draining into pulmonary artery | 168
no vegetations | 168
anomalous right coronary artery from the pulmonary artery diagnosis | 168
reviewed at interdisciplinary heart team rounds | 168
turned down for surgical intervention | 168
bacteremic Streptococcus bovis | 192
ceftriaxone | 192
metronidazole | 192
extubated | 216
transferred to cardiology ward | 216
dependent on intermittent haemodialysis | 216
transferred to hospice care | 960
deceased | 1800
no flow-limiting stenoses | 24
no murmurs | 0
no rubs | 0
no gallops | 0
no prior electrocardiogram for comparison | 0
no vegetations | 168
no intra-cardiac left-to-right shunt | 24
no pulmonary embolus | 24
no fistula involving RVOT | 24
no regional wall motion abnormalities | 24
no gastrointestinal malignancy ruled out | 192
no mechanical complication with RV infarction ruled out | 24
no underlying cardiomyopathy ruled out | 24
no pulmonary hypertension ruled out | 24
no massive pulmonary embolism ruled out | 24
no catecholaminergic state confirmed | 24
no sepsis ruled out | 24
no reversibility of disease | 192
no surgical intervention | 168
