66 years old | 0
female | 0
admitted to the emergency department | 0
chills | -72
leukocytosis | -72
burning chest pain | -216
rigors | -24
febrile | 0
temperature of 102.2 | 0
essential hypertension | 0
dyslipidemia | 0
severe aortic stenosis | 0
atherosclerotic coronary artery disease | 0
coronary artery bypass grafting | -2628
surgical aortic valve replacement | -2628
bioprosthetic valve | -2628
infective endocarditis | 0
sepsis of unknown etiology | 0
intravenous antibiotics | 0
chest x-ray | 0
electrocardiogram | 0
urinalysis | 0
sputum cultures | 0
transthoracic echocardiogram | 0
large hyperechoic mass on the tricuspid valve | 0
tricuspid regurgitation | 0
elevated right ventricular systolic pressure | 0
hyperechoic mass on the lateral wall of the right atrium | 0
vegetations | 0
admitted to the cardiac unit | 0
mechanical thrombectomy | 24
remnant leads | 24
TEE imaging | 24
cardiac computed tomography | 24
CCT with 3D reconstruction | 24
atrial and ventricular epicardial wires | -2628
percutaneous lead removal | 48
cardiothoracic surgeon | 48
percutaneous extraction of the infected remnant lead | 48
right femoral vein accessed | 48
6 French sheath inserted | 48
EN Snare introduced | 48
CloverSnare introduced | 48
Amplatz Goose Neck Snare | 48
successful snaring and removal of the remnant lead | 48
absence of pericardial effusion | 48
peripherally inserted central catheter | 48
6 weeks of intravenous antibiotics | 48
follow-up by infectious disease specialist | 168
no recurrent bacteremia | 168
afebrile | 168
repeat transthoracic echocardiogram | 336
no vegetations in the tricuspid valve | 336
mild regurgitation | 336
discharged | 336