62 years old | 0
male | 0
hypertension | 0
smoking | 0
AICD implant | -9360
out of hospital ventricular fibrillation arrest | -9360
scheduled for AICD generator box change | 0
general anesthesia | 0
anesthetic pre assessment | 0
good ventricular function on echocardiogram | 0
break in the insulation of the AICD lead component | 0
generator box removed | 0
leads left in situ | 0
plan for laser extraction | 0
laser extraction of leads | 48
pericardial tamponade | 48
linear tear in the free wall of the right ventricle | 48
emergency surgery | 48
extubated | 48
central venous pressure | 48
intermittently hypoxemic | 72
PaO2 of 6.8–13.3 kPa | 72
high inspired oxygen via continuous positive airway pressure mask | 72
central venous pressure | 72
left basal collapse | 72
transthoracic echocardiogram | 72
computed tomography pulmonary angiography | 72
small right solitary pulmonary embolism | 72
small left pleural effusion | 72
atelectasis | 72
heparin infusion | 72
aneurysmal interatrial septum | 96
transesophageal echocardiography | 96
flail tricuspid valve | 96
severe eccentric TR | 96
large PFO with a bidirectional shunt | 96
dilatation of right atrial | 96
dilatation of right ventricular | 96
mild RV dysfunction | 96
preserved left ventricular function | 96
tricuspid valve replacement | 120
bovine pericardial patch closure of PFO | 120
good postoperative recovery | 144
discharged home | 144
follow-up | 1008
returned to normal activity | 1008
echocardiogram | 1008
well seated functioning tricuspid prosthesis | 1008
no residual shunt across the interatrial septum | 1008