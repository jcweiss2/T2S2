73 years old | 0
    female | 0
    arterial hypertension | 0
    calcium channel blocker | 0
    admitted to the emergency department | 0
    diffuse abdominal pain | 0
    abdominal pain more marked at the right hypochondrium | 0
    history of episodic hepatic colic | -168
    fever | -168
    hemodynamically unstable | 0
    blood pressure 80/50 mmHg | 0
    heart rate 135 bpm | 0
    cold extremities | 0
    prolonged reschooling time | 0
    respiratory rate 25 bpm | 0
    SpO2 92% on room air | 0
    G score 17 | 0
    temperature 39.2°C | 0
    BMI 32 kg/m² | 0
    oligo-anuric | 0
    tachycardia | 0
    normal pleuropulmonary auscultation | 0
    patient confused | 0
    GCS 14/15 | 0
    diffuse abdominal tenderness | 0
    defense in the right hypochondrium | 0
    positive Murphy sign | 0
    transferred to the intensive care unit | 0
    conditioning | 0
    vascular filling with 2L 0.9% saline solution | 0
    no hemodynamic response | 0
    no renal response | 0
    introduction of noradrenaline 0.4 μg/kg/min | 0
    central venous line | 0
    central venous pressure 1 mmHg | 0
    probabilistic bi8 antibiotic therapy with Ceftriaxon + Metronidazol | 0
    blood cultures performed | 0
    ECG regular sinus rhythm | 0
    heart rate 137 bpm | 0
    transthoracic echocardiography | 0
    no acute cor pulmonale | 0
    no disorders explaining shock | 0
    LVEF 50% | 0
    unremarkable chest X-ray | 0
    arterial blood gas showing uncompensated metabolic acidosis | 0
    hyperlactatemia 7.02 mmol/l | 0
    leukocytosis 15280/μl | 0
    platelet count 80000/μl | 0
    hemoglobin 8.2g/dl | 0
    CRP 336mg/l | 0
    PCT 45μg/l | 0
    ferritin 1500μg/l | 0
    TP 50% | 0
    elongated TCA | 0
    ASAT 73UI/l | 0
    ALAT 92UI/l | 0
    BT 27mg/l | 0
    BD 22mg/l | 0
    GGT 498 UI/l | 0
    PAL 425 UI/l | 0
    LDH 214UI/l | 0
    urea 4.5g/l | 0
    creatinine 100mg/l | 0
    potassium 7.2mEq/l | 0
    sodium 137mEq/l | 0
    corrected calcium 90mg/l | 0
    lipasemia 12 IU/l | 0
    ECBU sterile | 0
    acute cholangitis | 0
    abdominal ultrasound | 0
    distended gallbladder | 0
    thickened gallbladder wall 8mm | 0
    dilation of intrahepatic bile ducts | 0
    difficulty highlighting an obstacle | 0
    abdominal CT scan | 0
    diagnosis of Mirizzi syndrome | 0
    vitamin K 10mg IV | 0
    acute febrile angiocholitis | 0
    septic shock | 0
    acute renal failure | 0
    diagnosis of ictero-uremigenic angiocholitis | 0
    worsening hemodynamic state | 0
    increased norepinephrine doses | 0
    introduction of dobutamine | 0
    6-hour hemodialysis session | 0
    metabolic acidosis | 0
    threatening hyperkalemia | 0
    anuria | 0
    cardiorespiratory arrest during dialysis | 24
    unsuccessful resuscitation | 24
    death declared | 24
    