22 years old | 0
female | 0
dyspnea | -72
denied cough | -72
denied sputum | -72
denied chest pain | -72
denied other respiratory symptoms | -72
denied upper and lower extremity weakness | -72
denied blurred vision | -72
denied swallowing difficulty | -72
speech problem | -216
nasal speech | -216
treated by ENT surgeons | -216
treated by speech therapist | -216
no history of substance abuse | 0
no recent drug intake | 0
labored breathing | 0
respiratory rate of 40 breaths/minute | 0
confused | 0
SaO2 85% | 0
blood pressure 146/98 mm Hg | 0
pulse 104/minute | 0
regular | 0
body temperature 36.7°C | 0
pedal edema absent | 0
neck vein engorgement absent | 0
mild crackles at both lung fields | 0
arterial blood gas analysis | 0
pH 7.314 | 0
PaCO2 56.7 mm Hg | 0
PaO2 92.2 mmHg | 0
oxygen saturation 90% | 0
chest X-ray | 0
no definite infiltration | 0
lung volume reduced | 0
white blood cell count 6980 μL | 0
hemoglobin 12.5 g/dL | 0
platelet count 345 000 μL | 0
blood glucose 94 mg/dL | 0
BUN/Cr 12/0.8 mg/dL | 0
AST/ALT 24/25 units/L | 0
chest computed tomography scan | 0
no pulmonary thromboembolism | 0
ECG | 0
sinus tachycardia | 0
echocardiography | 0
normal systolic and diastolic heart function | 0
supplemental oxygen | 0
transferred to intensive care unit | 0
mechanically ventilated | 0
rapid sequence induction | 0
IV midazolam 3 mg | 0
succinylcholine 70 mg | 0
SaO2 improved to 100% | 0
unable to breathe without mechanical support | 24
assessment by ENT surgeon | 24
no upper airway obstruction | 24
considered other causes of respiratory failure | 24
Guillain–Barre syndrome | 24
myasthenia gravis | 24
physical and neurological examination | 24
cerebrospinal fluid analysis | 24
normal | 24
diagnosis of myasthenia gravis | 48
electromyography | 48
decremental response to repetitive nerve stimulation | 48
pharmacological Jolly test | 48
incremental responses of tidal volume of ventilation | 48
acetylcholine receptor antibody titer 12.4 nmol/L | 48
pyridostigmine bromide 720 mg/day | 48
prednisolone 30 mg/day | 48
intravenous gamma-globulin 400 mg/kg/day | 48
condition improved | 168
weaning from ventilator failed | 336
tracheostomy | 336
successfully weaned from ventilator | 720
discharged | 1440
advised to do thymectomy | 1440
developed respiratory distress | 2880
respiratory arrest | 2880
signs and symptoms of sepsis | 2880
successfully intubated | 2880
resuscitated | 2880
prednisolone stepped up | 2880
pyridostigmine stepped up | 2880
antibiotics | 2880
fluid | 2880
intravenous gamma-globulin 400 mg/kg/day | 2880
discharged | 3456
section of excised thymus | 3456
follicular hyperplasia | 3456
followed up | 3456
responded well with maintenance steroid | 3456
responded well with pyridostigmine | 3456