19 years old | 0
male | 0
admitted to the hospital | 0
severe pain in the nuchal area | -48
mild occipital headache | -48
mild sore throat | -72
headache started | -72
nuchal pain started | -72
fever up to 40 degrees Celsius | -24
chills | -24
nuchal rigidity | 0
opposition to passive anteflexion and rotation of the head | 0
mild redness and enlargement of tonsils | 0
limited straight leg raise maneuver | 0
afebrile | 0
normal blood pressure | 0
normal heart rate | 0
no edema | 0
no erythema | 0
no palpable mass of the neck | 0
leukocytosis (25,590 cells/mL) | 0
neutrophilia (23,180 cells/mL) | 0
elevated C-reactive protein (179.88 mg/L) | 0
elevated procalcitonin (17.38 ng/mL) | 0
CT head unremarkable | 0
chest radiogram without infiltrative or nodular changes | 0
no lateralization | 0
no limb paresis | 0
lumbar puncture performed | 0
borderline pleocytosis (10 mononuclear cells/μL) | 0
normal proteinorhachia (15.5 mg/dL) | 0
empiric antimicrobial therapy with ceftriaxone and vancomycin | 0
parenteral rehydration | 0
analgesic therapy | 0
headache disappeared | 24
pain in the nuchal area extended to left neck | 24
erythematous and tender left lateral neck skin | 24
generalized urticarial allergic exanthema | 24
antimicrobial therapy changed to piperacillin-tazobactam and clindamycin | 24
erythema and edema of left neck pronounced | 72
palpable mass in left neck | 72
CT neck revealed abscess | 72
thrombosis of left internal jugular vein | 72
CT scan revealed hypodense collection in spinal canal | 72
MRI cervical spine showed epidural effusion | 72
oropharyngeal swab culture positive for Klebsiella pneumoniae | 72
blood culture positive for Klebsiella pneumoniae | 72
diagnosed with tonsillopharyngitis | 72
cervical abscess | 72
epidural abscess | 72
treated with ceftriaxone and clindamycin | 72
CRP decline to 125 mg/L | 168
procalcitonin decline to 2.50 ng/L | 168
pain in neck area less severe | 168
local erythema fading | 168
transferred to Otorhinolaryngology | 168
surgical drainage of abscess | 168
pus culture positive for Klebsiella pneumoniae | 168
negative anaerobic culture | 168
postsurgical course unremarkable | 192
transferred back to intensive care | 192
afebrile | 192
minor pain near surgical wound | 192
no cervical pain | 192
no movement limitations | 192
CRP 26.00 mg/L | 192
clindamycin stopped | 192
continued piperacillin-tazobactam | 192
CT regression of cervical abscess | 504
partial recanalization of left internal jugular vein | 504
MRI regression of epidural effusion | 504
CRP 13.26 mg/L | 504
changed to moxifloxacin | 504
discharged | 504
asymptomatic after discharge | 672
CRP below 5 mg/L | 672
moxifloxacin discontinued | 672
