69 years old | 0
female | 0
presented to emergency room | 0
episodes of altered mental status | -24
hepatitis B-related liver cirrhosis/encephalopathy | -672
chronic kidney disease | -672
lactulose | 0
rifaximin | 0
hyperammonemia | 0
computed tomography scan of head | 0
no mass | 0
no hemorrhage | 0
no stroke | 0
admitted to the Intensive Care Unit | 0
intubated | 0
acute respiratory failure | 0
unresponsive | 0
magnetic resonance imaging (MRI) of the brain | 72
dark rim involving the globus pallidi bilaterally | 72
central high signal seen within the globus pallidi | 72
diffusion-weighted imaging (DWI) | 72
multiple areas of restricted diffusion | 72
lateral portion of the temporal lobes | 72
posterolateral portions of the parietal lobes | 72
medial portions of the frontal lobes | 72
thalami bilaterally | 72
centrally within the midbrain | 72
periaqueductal gray matter | 72
repeat MRI | 144
marked progression of diffuse cortical injury | 144
involving both cerebral hemispheres | 144
injury to the thalami and central structures | 144
partially pseudonormalized on DWI | 144
relative sparing of the perirolandic/motor-sensory cortex | 144
cerebellum | 144
mild, diffuse cerebral swelling | 144
sulcal effacement | 144
diffuse cortical injury | 144
without midline shift | 144
withdraw the life support | 216
terminally extubated | 216
died | 216
hyperammonemia | -24
hepatic failure | -672
liver cirrhosis | -672
encephalopathy | -672 
altered mental status | -24
acute hyperammonemic encephalopathy | 0
fatal condition | 0 
multiple medical complications | 216
unresponsiveness to medical management | 216
poor prognosis | 216