39 years old | 0
female | 0
admitted to the hospital | 0
carinal resection and reconstruction | 0
adenoid cystic carcinoma | -672
mild dyspnea | -672
chest computed tomography | -672
bronchoscopy | -672
obstructive pattern of the pulmonary function test | -672
forced expiratory volume in one second | -672
forced vital capacity | -672
ratio of 67% | -672
general anesthesia | -672
target-controlled infusion of propofol | -672
remifentanil | -672
rocuronium | -672
tracheal intubation | -672
35-Fr right-sided double-lumen tube | -672
right lateral position | -672
left bronchi and vasculature | -672
thoracoscopic surgery | -672
one-lung ventilation | -672
arterial oxygen tension | -672
inspired oxygen fraction | -672
left thoracoscopic surgery | -672
right-sided double-lumen tube | -672
single-lumen endotracheal tube | -672
bronchial blocker | -672
fiberoptic bronchoscope | -672
left lateral position | -672
right thoracotomy | -672
peak airway pressure | -672
tidal volume | -672
carinal resection | -672
sterile reinforced endotracheal tube | -672
airway pressure increased | -672
oxygen saturation by pulse oximetry | -672
SpO2 decreased | -672
two-lung ventilation | -672
SpO2 restored | -672
carina was removed | -672
anastomosis between the trachea and right main stem bronchus | -672
separated RMB | -672
anastomotic site | -672
no air leak | -672
left endobronchial tube | -672
non-dependent right lung | -672
ventilated by the transoral endotracheal tube | -672
low tidal volume | -672
airway pressure lower than 20 cmH2O | -672
SpO2 decreased | -672
tube was reinserted into the LMB | -672
both lungs were ventilated | -672
sufficient two-lung ventilation | -672
right OLV was reattempted | -672
SpO2 was gradually decreased | -672
left pulmonary artery was clamped | -672
SpO2 was maintained 100% | -672
left main pulmonary artery was ligated | -672
left endobronchial tube was removed | -672
right thoracotomy was closed | -672
patient was moved to the supine position | -672
tracheal extubation | -672
transferred to the intensive care unit | -672
discharged | 13