52 years old | 0
female | 0
scheduled for D10 neurofibroma excision | -7
pre-anaesthetic check-up | -7
no medical comorbidities | -7
no history of surgical or anaesthetic exposures | -7
baseline routine investigation | -7
random blood sugar 144 mg/dl | -7
pre-operative fasting period 7 h for solid food | -7
pre-operative fasting period 2 h for clear water | -2
laminectomy and tumour excision under general anaesthesia | 0
steroids not administered | 0
analgesia with intravenous fentanyl | 0
paracetamol administered | 3
reversal of neuromuscular blockade | 4
extubation of trachea | 4
shifted to Post-Anaesthesia Care Unit | 4
nausea | 4.5
abdominal pain | 4.5
agitation | 4.5
tachypnoea | 4.5
dry mouth, tongue and lips | 4.5
hypotension | 4.5
tachycardia | 4.5
afebrile | 4.5
blood sample for estimation of arterial blood gases and sugar | 4.5
blood glucose levels 464 mg/dl | 4.5
high anion gap metabolic acidosis | 4.5
pH 7.12 | 4.5
bicarbonate 8 mmol/L | 4.5
base deficit 18 | 4.5
anion gap 22 | 4.5
potassium 4.2 mmol/L | 4.5
sodium 132 mmol/L | 4.5
urinary sample tested using dipsticks | 5
presence of glucose and ketone bodies | 5
serum β-hydroxybutyrate elevated | 5
diagnosis of DKA | 5
fluid resuscitation with 0.9% normal saline | 5
insulin bolus administered | 5
electrolyte derangements corrected | 5
serum amylase level mildly elevated | 5
lipase within normal range | 5
resolution of ketoacidosis | 24
general condition of the patient improved | 24
subcutaneous insulin started | 24
cessation of IV insulin | 24
shifted to the ward | 72
glycosylated haemoglobin levels estimated | 72
HbA1c levels 7.2% | 72
blood and urine samples sent for culture | 72
culture results sterile | 72
blood glucose levels reasonably normal | 120
discharged | 168
advice to continue subcutaneous insulin therapy | 168
follow-up in the Endocrinology outpatient section | 168