78 years old | 0
male | 0
admitted to the hospital | 0
hydrocelectomy | -360
scrotal pain | -360
scrotal swelling | -360
temperature of 38 degrees C | 0
leukocytosis | 0
elevated CRP | 0
enlarged left testis | 0
swelling and fluids in the scrotal content | 0
enlarged epididymis | 0
initial diagnosis of orchidoepididymitis | 0
multiple abscesses | 0
surgical exploration of the scrotum | 0
left hemiscrotectomy | 0
placement of suprapubic catheter | 0
Actinomyces turicensis | 0
Streptococcus viridans | 0
Staphylococcus | 0
necrosis | 0
phlegmonous inflammation | 0
abscesses of the scrotum | 0
necrotizing fasciitis | 0
hyperbaric oxygen chamber | 24
parenteral administration of broad spectrum antibiotics | 24
Imipenem | 24
Cefotaxim | 24
Metronidazol | 24
intensive care unit | 24
resolution of critical condition | 48
referral to the department of plastic surgery | 48
Mesh-Grafting | 72
vacuum assisted closure | 72
skin auto transplantation | 72
recovered from the complication | 168