81 years old | 0
female | 0
admitted to the hospital | 0
fatigue | -72
lethargy | -72
fever | -72
chills | -72
phlegm | -72
wheezing | -72
coma | -24
oxygen saturation dropped | -24
admitted to the ICU | 0
progressive drop in blood pressure | 0
norepinephrine | 0
chronic obstructive pulmonary disease | -43800
bronchial asthma | -43800
chronic heart insufficiency | -43800
oral bisoprolol | -43800
body temperature 36 °C | 0
pulse 85 beats/min | 0
respiratory rate 18 breaths/min | 0
blood pressure 105/45 mmHg | 0
breath sounds decreased | 0
wet rales | 0
cardiac examination unremarkable | 0
abdominal examination unremarkable | 0
initial troponin level 0.05 ng/mL | 0
B-type natriuretic peptide 4164 pg/mL | 0
arterial blood gas analysis | 0
inflammatory indicators | 0
polymerase chain reaction-severe acute respiratory syndrome coronavirus 2 test negative | 0
blood cultures negative | 0
other blood tests normal | 0
fecal examinations normal | 0
coagulation function normal | 0
electrocardiogram findings | 0
echocardiography | 0
chest CT | 0
abdominal CT | 0
PCI | 24
diminished bowel sounds | 48
abdominal distension | 48
increased dose of norepinephrine | 48
abdominal wall swelling | 96
increased abdominal wall tension | 96
bowel sounds disappeared | 96
urgent abdominal CT scan | 96
extensive pneumatosis intestinalis | 96
extensive intestinal wall necrosis | 96
death | 120
AMI | 96
septic shock | 0
assisted ventilation | 0
vasoactive drugs | 0
anti-infection treatment | 0
PCI via left femoral artery approach | 24
no significant abnormalities in coronary arteries | 24
glycerin enema | 48
abdominal CT showed hepatic portal gas and intestinal necrosis | 96