67 years old | 0
    male | 0
    diabetes | 0
    hypertension | 0
    dyslipidemia | 0
    left foot pain | -48
    left foot swelling | -48
    left plantar ulcer | -48
    pus discharge | -48
    fever | -48
    generalized weakness | -48
    ill appearance | 0
    pale | 0
    febrile | 0
    temperature 38.7 | 0
    tachycardic | 0
    pulse 105 | 0
    left foot hotness | 0
    left foot redness | 0
    left foot tenderness | 0
    left plantar ulcer irregular shape | 0
    undermined edges | 0
    necrotic base | 0
    no abdominal distension | 0
    no abdominal tenderness | 0
    Foley catheter inserted | 0
    pus in urine | 0
    WBC 15.5 | 0
    HB 7.9 | 0
    CRP 41 | 0
    K 5.5 | 0
    Na 130 | 0
    random blood glucose 327 mg/dl | 0
    urine WBC | 0
    urine RBC | 0
    admitted | 0
    left plantar ulcer debridement | 0
    daily dressing | 0
    intravenous antibiotic | 0
    sudden onset severe abdominal pain | 72
    suprapubic pain | 72
    constant pain | 72
    fever | 72
    vomiting | 72
    abdominal distension | 72
    tense abdomen | 72
    tender abdomen | 72
    abdominal CT scan | 72
    pneumoperitoneum | 72
    abdomino-pelvic free fluid | 72
    hollow viscus perforation | 72
    diffuse mesentery haziness | 72
    small bowel dilatation | 72
    Foley catheter balloon in situ | 72
    partially distended urinary bladder | 72
    perforated viscus diagnosis | 72
    booked for surgery | 72
    exploratory laparotomy | 72
    intra-abdominal turbid fluid collection | 72
    pelvic pus pockets | 72
    right paracolic gutter pus | 72
    dilated congested bowel loops | 72
    no bowel perforation | 72
    mesentery edema | 72
    urinary bladder perforation 3x3 cm | 72
    inflamed bladder mucosa | 72
    pus from bladder | 72
    peritoneal lavage | 72
    biopsies taken | 72
    perforation edges refreshed | 72
    water-tight repair | 72
    suprapubic catheter inserted | 72
    Foley catheter inserted | 72
    histopathology nonspecific inflammation | 72
    no malignancy | 72
    post-operative recovery | 72
    SICU stay 3 days | 72
    transferred to surgical ward | 96
    oral fluids started | 96
    full diet commenced | 120
    intravenous antibiotics continued | 192
    discharged | 240
    spontaneous urinary bladder rupture | 72
    acute abdomen | 72
    septic shock | 72
    recurrent urinary tract infection | -48
    chronic infection | -48
    malignancy ruled out | 72
    diabetes complication | -48
    inflammation | 72
    infection | 72
    no enterocystoplasty | 72
    no bladder malignancy | 72
    no pelvic irradiation | 72
    neurologic bladder | 72
    obstructed labor | 72
    no alcoholism | 72
    no radiotherapy | 72
    no neurogenic bladder | 72
    no delayed postpartum complications | 72
    biochemical renal dysfunction | 72
    associated conditions ruled out | 72
    high index of suspicion | 72
    acute peritonitis | 72
    diagnostic laparoscopy | 72
    explorative laparotomy | 72
    biopsy for malignancy | 72
    conflict of interest | 240
    funding | 240
    consent | 240
    author contributions | 240
    <|eot_id|>
    