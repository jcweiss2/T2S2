31 years old | 0
female | 0
diagnosed with congenital bicuspid aortic valve | -133584
AV and ascending aortic root replacement | -43608
biventricular pacemaker inserted | -43608
presented with headaches | -168
presented with fevers | -168
presented with confusion | -168
aeromedical retrieval | -72
treated as meningoencephalitis | -72
blood cultures positive for methicillin-resistant Staphylococcus aureus | 0
transoesophageal echocardiogram confirming aortic prosthetic valve endocarditis | 0
cardiac case conference | 144
consensus for medical treatment | 144
craniotomy and drainage of brain abscess | 360
baseline PET-FDG consistent with PVE | 1008
imaging showing para-valvular abscess formation | 1080
imaging showing peri-aortic abscess formation | 1080
imaging showing bilateral pseudo0 aneurysms | 1080
aeromedical transfer to interstate cardiothoracic surgery facility | 1200
redo-bioprosthetic aortic valve replacement | 1344
aortic root replacement | 1344
PPM and leads explantation | 1344
PPM re-insertion | 1416
returned to NT hospital | 1776
discharged against medical advice | 2112
lost to follow-up | 2112
presented to remote community clinic | 2760
commenced high-dose oral dicloxacillin | 2760
commenced rifampicin | 2760
PET-FDG with no AVR uptake | 2976
CTCA showing pseudo-aneurysms | 2976
CTCA showing pseudo-aneurysms stable | 4656
transthoracic echocardiogram showing normal bioprosthetic valve function | 10008
diagnosed with bicuspid AV at age 15 | -133584
progression to severe stenosis | -43608
progression to regurgitation | -43608
development of 4.7 cm aneurysm of ascending aorta | -43608
bioprosthetic aortic valve replacement | -43608
replacement of ascending aorta with Dacron graft | -43608
dual-chamber pacemaker inserted | -43608
type 2 diabetes mellitus | 0
hypertension | 0
smoking | 0
suboptimal adherence to metformin | 0
suboptimal adherence to bisoprolol | 0
suboptimal adherence to aspirin | 0
hypotension | 0
pulse rate 80/min | 0
oxygen saturation 100% | 0
respiratory rate 22/min | 0
febrile at 40.1°C | 0
Glasgow Coma Scale 14 | 0
no peripheral stigmata of IE | 0
fluid resuscitation | 0
vasopressor support | 0
broad-spectrum antibiotics | 0
normocytic anaemia | 0
elevated CRP | 0
normal WCC | 0
neutrophilic pleocytosis | 0
multi-organ septic emboli | 0
cerebral septic emboli | 0
kidney septic emboli | 0
radial artery septic emboli | 0
intensive care unit admission | 0
septic shock management | 0
IV flucloxacillin | 0
hyperglycaemia treatment | 0
anaemia requiring transfusion | 0
diuresis for biventricular heart failure | 0
no evidence of bleeding | 0
chronic inflammation | 0
haemodilution | 0
sinus rhythm with ventricular pacing | 0
left bundle branch block | 0
mobile echodensity on AVR | 0
vegetation | 0
no aortic root abscess formation | 0
no para-valvular regurgitation | 0
no vegetations on PPM leads | 0
multiple cerebral infarcts | 144
meningeal enhancement | 144
non-surgical management recommendation | 144
evolving left frontal lobe cerebral abscess | 312
drainage of 30x40x20 mm abscess | 312
S. aureus culture | 312
unchanged TTE | 312
clinically stable | 312
rifampicin added | 312
interruptions to IV flucloxacillin | 0
interruptions to oral rifampicin | 0
FDG-PET performed | 984
new mild paravalvular aortic incompetence | 1080
abnormal Doppler flow external to aortic root | 1080
TOE demonstrating two pseudo-aneurysms | 1080
CTCA confirming abscess formation | 1080
CTCA confirming pseudo-aneurysms | 1080
repeat blood cultures negative | 1080
explantation of AV bioprosthesis | 1344
explantation of aortic graft | 1344
explantation of PPM | 1344
debridement | 1344
patch reconstruction of aortic root | 1344
AVR with Edwards LifeSciences Inspiris Resilia bioprosthesis | 1344
replacement of ascending aorta and hemi-arch | 1344
residual pseudo-aneurysm under left coronary sinus | 1344
PPM insertion | 1416
IV flucloxacillin post-AVR | 1344
rifampicin post-AVR | 1344
antibiotic duration shortened | 1344
high-dose oral dicloxacillin | 2760
high-dose rifampicin | 2760
no AVR uptake on PET-FDG | 2976
CTCA showing pseudo1 aneurysms | 2976
pseudo-aneurysms stable | 4656
normal bioprosthetic valve function | 10008
no follow-up attendance | 2112
inconsistent follow-up | 2112
last specialist review | 0
last TTE | 0
recent PPM interrogation | 0
CTCA overdue | 0
