67 years old | 0
    woman | 0
    backache | 0
    calculi in both kidneys | 0
    ureteral calculi | 0
    admitted | 0
    holmium laser lithotripsy | 0
    double J catheterization | 0
    purulent urine | 0
    severe fever | -30
    body temperature 39.5 °C | -30
    chill | -30
    low blood pressure | -30
    60/42 mmHg | -30
    empiric anti-infection drugs | -30
    imipenem | -30
    cilastatin sodium | -30
    fluid resuscitation | -30
    30 mL/kg | -30
    vasoactive agent | -30
    norepinephrine | -30
    hydrocortisone sodium succinate | -30
    symptoms progressively deteriorated | -48
    anuric | -48
    ARDS | -48
    invasive ventilatory support | -48
    endotracheal intubation | -48
    CRRT | -48
    transferred to ICU | 0
    sedated state | 0
    Richmond agitation-sedation scale -4 | 0
    blood pressure 80/62 mmHg | 0
    norepinephrine 1.5 μg/kg/min | 0
    epinephrine 1.0 μg/kg/min | 0
    heart rate 139 beats/min | 0
    transcutaneous oxygen saturation 80% | 0
    cold clammy extremities | 0
    loud bubbling sound in lung | 0
    oxygen partial pressure 50 mmHg | 0
    lactic acid 10.6 mmol/L | 0
    bicarbonate 10.8 mmol/L | 0
    central venous pressure 20 cmH20 | 0
    B lines in lung | 0
    diffuse dysfunction | 0
    severe damage in left ventricle | 0
    LVEF 20.3% | 0
    normal right ventricle function | 0
    sinus tachycardia | 0
    broad ST depression | 0
    troponin I 10.2 ng/mL | 0
    NT-BNP >35,000 pg/L | 0
    creatinine 356 μmol/L | 0
    anuria | 0
    multiple organ function failure | 0
    VA-ECMO initiated | 0
    ECMO catheter placement | 0
    arterial catheter placement | 0
    centrifugal pump Maquet Rotaflow RF 32 | 0
    3000 rpm | 0
    blood flow 3.5 L/min | 0
    arterial pressure 135 mmHg | 0
    venous pressure -29 mmHg | 0
    cyclic dynamics improved | 0.5
    norepinephrine stopped | 0.5
    epinephrine stopped | 0.5
    CRRT initiated | 0
    imipenem and cilastatin sodium | 0
    vancomycin | 0
    lactic acid declined | 2
    vasoactive drugs stopped | 10
    arterial lactate normal | 12
    extended-spectrum β-lactamase-positive E. coli | 48
    inflammatory indices diminished | 48
    vancomycin trough 15-20 μg/mL | 48
    LVEF 35% | 120
    necrotic skin in extremities | 120
    ECMO weaned | 144
    acute kidney injury grade 3 | 144
    CRRT discontinued | 144
    urinating | 144
    urine volume 1000 mL/day | 144
    vascular ultrasonography | 336
    computed tomography angiography | 336
    necrotic tissues amputated | 336
    tracheal intubation | 0
    spontaneous breathing | 120
    weaning failed | 120
    trachea opened | 240
    anti-infection regimen changed | 240
    cefoperazone sodium | 240
    sulbactam sodium | 240
    physical rehabilitation | 480
    ventilator weaned | 480
    tracheotomy tube sealed | 600
    discharged | 768
    intermittent hemodialysis | 768
    self-care at 6 months | 4320
    intermittent hemodialysis ongoing | 4320
    