57 years old | 0
male | 0
admitted to University Hospital | 0
paraparesis | -2160
sensory disturbances in both lower extremities | -2160
fall | -2160
diagnosed with CES | 0
L3 burst fracture | -2160
spinal canal compression | -2160
posterior lumbar interbody fusion | 0
neuropathic pain | 0
transferred to rehabilitation hospital | 0
fever | -168
general weakness | -168
leukocytosis | -168
Klebsiella pneumoniae isolated from blood and urine culture tests | -168
edema in bilateral renal parenchyma | -168
hyperechogenicity | -168
renal failure | -168
acute pyelonephritis | -168
sepsis | -168
meropenem administered intravenously | -168
vital signs stable | -120
laboratory findings returned to normal | -120
antibiotics stopped | -120
transferred to rehabilitation medicine department | 0
muscular weakness in both lower limbs | 0
tingling sensations | 0
allodynia | 0
hyperalgesia | 0
decreased sensations below the third lumbar segment | 0
sitting and standing up independently | 0
moderate assistance for balanced-level walking | 0
Modified Barthel Index 76 points | 0
deep tendon reflex decreased in both lower limbs | 0
anal sphincter tone decreased | 0
bulbocavernosus reflex decreased | 0
electrodiagnostic study | 0
somatosensory evoked potential | 0
needle electromyography | 0
bilateral lumbosacral polyradiculopathy | 0
sacral reflex arc lesion | 0
voided with an indwelling catheter | 0
self-voiding 100-200 mL | 0
residual urine volume 200-300 mL | 0
timed intermittent catheterization | 0
comprehensive rehabilitative managements | 0
drug therapy | 0
muscle strengthening exercises | 0
functional electrical stimulation | 0
gait training | 0
chills | 312
fever | 312
leukocytosis | 312
Klebsiella pneumoniae isolated from blood and urine culture tests | 312
recurrent acute pyelonephritis | 312
tazobactam administered intravenously | 312
meropenem administered intravenously | 312
pain and tenderness on the left flank | 315
mass palpated in left abdomen | 315
perirenal hemorrhage | 315
coil embolization | 315
conservative treatment for acute renal failure | 315
surgical hematoma removal | 318
voiding cystourethrography | 318
vesicoureteral reflux not observed | 318
urodynamic study | 318
detrusor areflexia | 318
oral medications | 318
intermittent self-catheterization | 318
transferred to rehabilitation hospital | 324