75 years old | 0
male | 0
admitted to the hospital | 0
resection of a ruptured abdominal aortic aneurysm | -20880
placement of an aortobifemoral bypass graft | -20880
Type 2 diabetes mellitus | 0
hypertension | 0
chronic thrombocytopenia | 0
chronic kidney injury | 0
postoperative renal failure | -20880
dialysis | -20880
rigors | -48
dysuria | -48
polyuria | -48
burning micturition | -48
fever | 0
weakness |-48
lethargy |0
denies cough | 0
denies chest pain | 0
denies palpitations | 0
denies nausea | 0
denies vomiting | 0
denies constipation | 0
blood pressure 70/35 mmHg | 0
blood pressure 90/48 mmHg | 0
temperature 101°F | 0
heart rate 90/min | 0
respiratory rate 20/min | 0
white blood cell count 18,000 | 0
lactic acid 4.1 | 0
20% bands | 0
platelet count 20,000 | 0
urinalysis white blood cells | 0
urinalysis red blood cells | 0
urinalysis moderate leukocyte esterase | 0
diffuse abdominal tenderness | 0
peri(peri-umbilical tenderness | 0
deep palpation without peritoneal signs | 0
diagnosis of severe sepsis | 0
secondary to urinary tract infection | 0
high anion gap metabolic acidosis | 0
secondary to lactic acidosis | 0
Eggerthella lenta septicemia | 0
Escherichia coli ESBL-positive urinary tract infection | 0
started on IV ertapenem | 0
abdominal CT with contrast | 24
induration with inflammatory changes around the graft | 24
stranding around the aorta near iliac components | 24
presence of an air bubble between components | 24
aortoenteric fistula | 24
recommended graft replacement surgery | 24
repair of the fistula | 24
refused surgery | 24
treated with IV antibiotics | 24
repeated negative blood cultures | 168
discharged home | 168
outpatient antibiotic treatment | 168
chronic antibiotic suppression | 168
