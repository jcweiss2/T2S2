46 years old | 0
male | 0
diagnosed with coccidioidomycosis | 0
presented to the emergency room | 0
shortness of breath | -2928
cough | -2928
pleuritic chest pain | -2928
malaise | -2928
diffuse joint pain | -2928
intermittent fevers | -2928
denied hemoptysis | 0
denied recent travel | 0
denied incarceration history | 0
denied homelessness | 0
worked as a farmer in Bakersfield for the past 3 years | 0
seen at an outside facility for fatigue | -672
seen at an outside facility for fevers | -672
seen at an outside facility for forearm lesions | -672
tested positive for Coccidioides antibody IgG | -672
tachycardic | 0
tachypneic | 0
afebrile | 0
normotensive | 0
hypoxic | 0
coarse bilateral breath sounds | 0
labored breathing | 0
palpable subcutaneous nodules in the forearms bilaterally | 0
no notable rashes | 0
no joint effusions | 0
no neurologic deficits | 0
transitioned to non-invasive mechanical ventilation | 0
admitted to the intensive care unit | 0
acute hypoxemic respiratory failure | 0
severe sepsis | 0
CT scan of the chest with IV contrast | 0
diffuse multifocal nodular consolidations | 0
ground glass opacities | 0
right upper lobe dense consolidations | 0
prominent mediastinal and hilar lymph nodes | 0
clear central airways | 0
no evidence of pulmonary embolism | 0
started on IV trimethoprim sulfamethoxazole | 0
started on IV cefepime | 0
started on oral fluconazole | 0
started on IV liposomal amphotericin B | 0
started on oral prednisone | 0
decompensated overnight | 0
required mechanical ventilation | 0
decompensated further into septic shock | 0
required norepinephrine | 0
blood cultures negative | 0
tuberculosis ruled out | 0
fungal studies negative for pneumocystis | 0
fungal studies negative for cryptococcus | 0
fungal studies negative for toxoplasmosis | 0
coccidiomycosis with titer levels of 1:64 in the blood | 0
coccidiomycosis with titer level of 1:1 in the cerebrospinal fluid | 0
infectious disease consulted | 0
antiretroviral therapy held | 0
declining mentation | 0
worsening respiratory status | 0
minimal response to proning | 0
intermittent severe metabolic acidosis | 0
renal failure | 0
improved with dialysis | 0
improved with bicarbonate drips | 0
CT scan of the head with IV contrast | 0
corpus callosum mass extending into the left lateral ventricle | 0
MRI of the brain showed hemorrhagic mass | 0
echocardiogram showed right ventricular mobile mass | 0
started on IV flucytosine | 0
switched to IV fluconazole | 0
placed on comfort care | 0
compassionately extubated | 0
expired | 0
