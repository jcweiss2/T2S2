72 years old | 0
woman | 0
urinary incontinence | 0
ground-level fall | -672
right frontal meningioma | -672
neurosurgery | -672
outpatient surgery scheduled | -672
dexamethasone 4 mg every 6 hours for 20 days | -672
outpatient surveillance | -672
second ground-level fall | -72
dyspnea | -72
nonproductive cough | -72
chest pain | -72
generalized weakness | -72
crackles in right lung base | 0
chest X-ray consolidation right lung base | 0
elevated white blood cell count | 0
elevated neutrophils | 0
thrombocytopenia | 0
normal renal function | 0
admitted for suspected community-acquired pneumonia | 0
admitted for meningioma management | 0
IV ceftriaxone | 0
IV azithromycin | 0
discontinued dexamethasone 3 days before admission | -72
restarted dexamethasone 4 mg IV every 6 hours | 0
tapered up to 6 mg IV every 6 hours | 168
chest pain continued | 168
productive cough | 168
hemoptysis | 168
repeat chest X-ray cavitary lesion | 168
CT scan cavitary mass right middle lobe 6x3.5 cm | 168
sputum samples for AFB stain and culture | 168
AFB stain negative | 168
AFB culture negative | 168
serum QuantiFERON gold test indeterminate | 168
repeat QuantiFERON gold test negative | 168
serum Aspergillus antigen enzyme immunoassay negative | 168
vancomycin | 168
piperacillin-tazobactam | 168
right-sided hydropneumothorax | 168
chest tube placement | 168
pneumothorax resolved | 168
pulmonary consult for diagnostic bronchoscopy | 168
bronchoscopy with bronchoalveolar lavage | 168
BAL culture grew Streptococcus viridans | 168
BAL culture grew Aspergillus fumigatus | 168
acute-angle hyphae septate consistent with A. fumigatus | 168
voriconazole 490 mg IV every 12 hours | 168
switched to isavuconazole 372 mg IV every 24 hours | 168
thrombocytopenia | 168
rash | 168
continued pleural leak | 168
persistent pneumothorax | 168
progressive pneumothorax | 168
prolonged ileus | 168
worsening renal function | 168
cardiothoracic surgery consult for lobectomy | 168
family declined surgical intervention | 168
Aspergillus cavitary lesion continued | 168
ongoing right pneumothorax | 168
bronchopulmonary fistula concern | 168
aspergilloma complications concern | 168
antifungal therapy continued | 168
supportive care continued | 168
severe septic shock | 168
multiorgan failure | 168
death | 168
