58 years old | 0
female | 0
admitted to the hospital | 0
hypertension | -6720
diabetes mellitus | -6720
Brugada syndrome | -6720
implantable cardioverter-defibrillator (ICD) implantation | -336
febrile illness | -72
syncopal episodes | 0
ventricular fibrillation (VF) | -72
nonsustained VF | -72
ICD shocks | -72
fever persisted | 0
antipyretics | 0
maximum temperature | 24
multiple episodes of VF | 0
rapid nasal swab testing | 0
SARS-CoV-2 positive | 0
isoproterenol infusion | 0
aggressive treatment of fever | 0
acetaminophen | 0
salsalate | 0
cooling blanket | 24
fever control | 48
hydroxychloroquine | 24
QTc prolongation | 48
discontinued hydroxychloroquine | 48
oxygenation | 0
respiratory status declined | 24
non-rebreather mask | 24
prone positioning | 24
chest radiograph | 0
multifocal airspace and interstitial opacities | 48
acute respiratory distress syndrome | 48
COVID-19-associated pneumonia | 48
isoproterenol discontinued | 72
atrial tachycardia | 72
broad-spectrum antibiotics | 120
remdesivir | 144
respiratory function declined | 144
intubation | 144
lymphopenia | 144
C-reactive protein increased | 144
D-dimer increased | 144
fibrinogen increased | 144
ferritin increased | 144
procalcitonin increased | 144
therapeutic anticoagulation | 144
low-molecular-weight heparin | 144
septic shock | 168
vasopressors | 168
atrial tachycardia | 168
no ventricular arrhythmias | 168
sedation holiday | 432
unarousable | 432
computed tomography imaging | 432
intracranial hemorrhage | 432
mass effect | 432
transition to comfort care | 432