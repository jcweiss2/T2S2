male | 0 | 0 | Factual
premature birth | -672 | -672 | Factual
emergency cesarean delivery | -672 | -672 | Factual
abruptio placenta | -672 | -672 | Factual
birth weight 1090g | -672 | -672 | Factual
Apgar 4 and 8 | -672 | -672 | Factual
respiratory distress | -672 | 0 | Factual
mild respiratory distress | -672 | 0 | Factual
respiration rate 65 breaths per min | -672 | 0 | Factual
chest retraction | -672 | 0 | Factual
CPAP machine | -672 | 0 | Factual
positive end expiratory pressures 6 | -672 | 0 | Factual
inspired oxygen 30% | -672 | 0 | Factual
cloudy eyes | 0 | 0 | Factual
ectropion | 0 | 0 | Factual
dry ichthyotic skin | 0 | 0 | Factual
typical male genitalia | 0 | 0 | Factual
bilateral undescended testicles | 0 | 0 | Factual
height 75th percentile | 0 | 0 | Factual
weight 25th percentile | 0 | 0 | Factual
head circumference 25th percentile | 0 | 0 | Factual
temperature 36.2°C | 0 | 0 | Factual
heart rate 167 beats per min | 0 | 0 | Factual
pulsations well felt | 0 | 0 | Factual
breath sounds equal | 0 | 0 | Factual
no organomegaly | 0 | 0 | Factual
normal blood count | 0 | 0 | Factual
normal electrolytes | 0 | 0 | Factual
normal liver function | 0 | 0 | Factual
respiratory distress syndrome | 0 | 0 | Factual
ground-glass opacity | 0 | 0 | Factual
minor respiratory acidosis | 0 | 0 | Factual
surfactant dosage | 0 | 0 | Factual
CPAP assistance | 0 | 0 | Factual
bowel movement at 12h | -12 | -12 | Factual
trophic feeding | -72 | 0 | Factual
breast milk | -72 | 0 | Factual
abdominal distension | 144 | 144 | Factual
tachycardia | 144 | 144 | Factual
tachypnea | 144 | 144 | Factual
thrombocytopenia | 144 | 144 | Factual
neutropenia | 144 | 144 | Factual
C-reactive protein 70 mg/L | 144 | 144 | Factual
meropenem | 144 | 168 | Factual
vancomycin | 144 | 168 | Factual
antibiotics discontinued | 216 | 216 | Factual
feeding restarted | 216 | 216 | Factual
high-flow oxygen treatment | 336 | 672 | Factual
relapses of unexplained apnea | 504 | 672 | Factual
CPAP | 504 | 672 | Factual
septic examination negative | 504 | 672 | Factual
brain MRI normal | 504 | 504 | Factual
nasogastric tube | 504 | 672 | Factual
conjugated hyperbilirubinemia | 504 | 672 | Factual
total bilirubin 69.8 umol/L | 504 | 504 | Factual
neonatal cholestasis workup | 504 | 672 | Factual
experts suspected hepatitis and TPN | 504 | 504 | Factual
genetic studies | 504 | 672 | Factual
X-ray of spine normal | 504 | 504 | Factual
echocardiogram normal | 504 | 504 | Factual
eye test normal | 504 | 504 | Factual
skull X-ray revealed craniosynostosis | 504 | 504 | Factual
hepatosplenomegaly not seen | 504 | 504 | Factual
biliary atresia not seen | 504 | 504 | Factual
albumin level decline | 504 | 672 | Factual
bilirubin, AST, and ALT levels rose | 504 | 672 | Factual
multiple albumin infusions | 504 | 672 | Factual
ursodeoxycholic acid 30 mg/kg/day | 504 | 672 | Factual
infectious etiology investigation | 504 | 672 | Factual
TSH, T3, T4, and cortisol normal | 504 | 504 | Factual
metabolic disorders negative | 504 | 504 | Factual
micropenis not detected | 504 | 504 | Factual
whole genomic sequence | 672 | 672 | Factual
NOTCH2 gene mutation | 1008 | 1008 | Factual
heterozygous variant c.1076c>T | 1008 | 1008 | Factual
pathogenic variant | 1008 | 1008 | Factual
severe cyanosis | 1008 | 1008 | Factual
apnea | 1008 | 1008 | Factual
bradycardia | 1008 | 1008 | Factual
cardio-respiratory resuscitation | 1008 | 1008 | Factual
intubation | 1008 | 1008 | Factual
mechanical breathing | 1008 | 1008 | Factual
epinephrine | 1008 | 1008 | Factual
septic shock | 1008 | 1008 | Factual
multiorgan failure | 1008 | 1008 | Factual
disseminated intravascular coagulation | 1008 | 1008 | Factual
acute renal damage | 1008 | 1008 | Factual
capillary leak syndrome | 1008 | 1008 | Factual
death | 2400 | 2400 | Factual
ALGS2 diagnosis | 2400 | 2400 | Factual
NOTCH2 mutation | 2400 | 2400 | Factual
craniosynostosis | 504 | 504 | Factual
ichthyosis | 0 | 0 | Factual
genetic counseling | 2400 | 2400 | Factual