26 years old | 0 | 0 
male | 0 | 0 
admitted to the hospital | 0 | 0 
new-onset headache | -24 | 0 
blurred vision | -24 | 0 
kidney transplant | -6048 | -6048 
end-stage kidney disease | -8736 | -6048 
immunosuppression | -24 | 0 
mycofenolate sodium | -24 | 0 
methylprednisolone | -24 | 0 
estimated glomerular filtration rate (eGFR) | 0 | 0 
proteinuria | 0 | 0 
chronic kidney transplant disease | 0 | 0 
status post vascular rejection | -6048 | -6048 
chronic calcineurin-inhibitor toxicity | -6048 | -6048 
contrast-enhancing intracerebral lesions | 0 | 0 
perifocal edema | 0 | 0 
methylprednisolone therapy stopped | 0 | 0 
dexamethasone administered | 0 | 24 
brain edema | 0 | 24 
transmitted to the university department of Nephrology | 24 | 24 
transmitted to the department of Neurosurgery | 24 | 48 
brain biopsy | 48 | 48 
diagnosis of cerebral PTLD | 48 | 48 
diffuse large B-cell lymphoma | 48 | 48 
positive for Ebstein-Barr virus | 48 | 48 
initial chemotherapy regime | 48 | 168 
high-dose cytarabin | 48 | 168 
Rituximab | 48 | 168 
complete remission of PTLD | 168 | 168 
impairment of the transplant function | 168 | 168 
cytomegalovirus (CMV) reactivated | 504 | 504 
pneumocystis jirovecii pneumonia | 504 | 504 
chemotherapy changed | 504 | 504 
Rituximab | 504 | 504 
antiviral and antibiotic therapy | 504 | 504 
mycofenolate sodium tapered | 504 | 504 
leukopenia | 504 | 504 
infections | 504 | 504 
generalized seizure | 720 | 720 
recurrence of PTLD | 720 | 720 
cerebral MRI scan | 720 | 720 
HDMTX | 720 | 720 
Leukovorine | 720 | 720 
Rituximab | 720 | 720 
vigorous hydration | 720 | 720 
alkalinization of the urine | 720 | 720 
high-flux hemodialysis (HFHD) | 744 | 912 
MTX-level measurements | 744 | 912 
dialysis sessions | 744 | 912 
nadir of leucocytes | 840 | 840 
granulocytes colony-stimulating factor | 840 | 840 
severe CMV- and E.coli pneumonia | 936 | 936 
sepsis | 936 | 936 
acute kidney transplant failure | 936 | 936 
transmission to an intensive care unit | 936 | 936 
invasive ventilation | 936 | 936 
sepsis managed | 936 | 1008 
mycofenolate sodium discontinued | 936 | 936 
antiviral and antibiotic therapy | 936 | 1008 
follow up cerebral MRI scan | 1092 | 1092 
small regredience of PTLD | 1092 | 1092 
cerebral radiation | 1092 | 1092 
no relevant response of the disease | 1092 | 1092 
dialysis parameters | 744 | 912 
MTX administration | 720 | 720 
Gambro machine AK 200 | 744 | 912 
high-flux dialyser (Polyflux 170H) | 744 | 912 
dialysate SelectBag One AX 450 G | 744 | 912 
unfractionated heparin | 744 | 912 
fluorescence polarization immunoassay | 744 | 912 
TDx analyser (Fa. Abbott) | 744 | 912 
MTX-level measurements | 744 | 912 
leucocytes measurements | 744 | 912 
estimated glomerular filtration rate (eGFR) measurements | 744 | 912 
hematological toxicities | 744 | 912 
infection developed | 936 | 936 
leucopenia | 840 | 840 
anemia | 840 | 840 
thrombocytes | 840 | 840 
CMV-colonization | -24 | 0 
CMV-activation | 504 | 504 
posttransplant immunosuppressive therapy | -24 | 0 
rituximab | 48 | 504 
impaired kidney function | 0 | 0 
high-flux hemodialysis (HFHD) | 744 | 912 
MTX clearance | 744 | 912 
MTX toxicity | 720 | 912 
MTX elimination | 744 | 912 
hemodialysis | 744 | 912 
hemodiafiltration | 744 | 912 
Charcoal hemoperfusion/hemofiltration | 744 | 912 
acute kidney failure | 936 | 936 
nephrotoxicity | 744 | 912 
granulocyte colony-stimulating factor | 840 | 840 
infection | 936 | 936 
sepsis | 936 | 936 
acute on chronic kidney failure | 936 | 936 
dialysis | 744 | 912 
MTX-level | 744 | 912 
leucocytes | 744 | 912 
eGFR | 744 | 912 
hematological toxicity | 744 | 912 
infection risk | 936 | 936 
CMV reactivation | 504 | 504 
pneumocystis jirovecii pneumonia | 504 | 504 
antiviral therapy | 504 | 504 
antibiotic therapy | 504 | 504 
mycofenolate sodium | 504 | 504 
Rituximab | 504 | 504 
high-dose cytarabin | 48 | 168 
cerebral radiation | 1092 | 1092 
PTLD | 48 | 1092 
diffuse large B-cell lymphoma | 48 | 48 
Ebstein-Barr virus | 48 | 48 
cerebral PTLD | 48 | 1092 
recurrence of PTLD | 720 | 720 
HDMTX therapy | 720 | 720 
MTX clearance | 744 | 912 
HFHD | 744 | 912 
MTX elimination | 744 | 912 
hemodialysis | 744 | 912 
hemodiafiltration | 744 | 912 
Charcoal hemoperfusion/hemofiltration | 744 | 912 
MTX toxicity | 720 | 912 
nephrotoxicity | 744 | 912 
hematological toxicity | 744 | 912 
infection risk | 936 | 936 
sepsis | 936 | 936 
acute on chronic kidney failure | 936 | 936 
dialysis | 744 | 912 
MTX-level | 744 | 912 
leucocytes | 744 | 912 
eGFR | 744 | 912 
hematological toxicity | 744 | 912 
infection | 936 | 936 
sepsis | 936 | 936 
acute kidney failure | 936 | 936 
cerebral radiation | 1092 | 1092 
PTLD | 48 | 1092 
diffuse large B-cell lymphoma | 48 | 48 
Ebstein-Barr virus | 48 | 48 
cerebral PTLD | 48 | 1092 
recurrence of PTLD | 720 | 720 
HDMTX therapy | 720 | 720 
MTX clearance | 744 | 912 
HFHD | 744 | 912 
MTX elimination | 744 | 912 
hemodialysis | 744 | 912 
hemodiafiltration | 744 | 912 
Charcoal hemoperfusion/hemofiltration | 744 | 912 
MTX toxicity | 720 | 912 
nephrotoxicity | 744 | 912 
hematological toxicity | 744 | 912 
infection risk | 936 | 936 
sepsis | 936 | 936 
acute on chronic kidney failure | 936 | 936 
dialysis | 744 | 912 
MTX-level | 744 | 912 
leucocytes | 744 | 912 
eGFR | 744 | 912 
hematological toxicity | 744 | 912 
infection | 936 | 936 
sepsis | 936 | 936 
acute kidney failure | 936 | 936 
cerebral radiation | 1092 | 1092 
PTLD | 48 | 1092 
diffuse large B-cell lymphoma | 48 | 48 
Ebstein-Barr virus | 48 | 48 
cerebral PTLD | 48 | 1092 
recurrence of PTLD | 720 | 720 
HDMTX therapy | 720 | 720 
MTX clearance | 744 | 912 
HFHD | 744 | 912 
MTX elimination | 744 | 912 
hemodialysis | 744 | 912 
hemodiafiltration | 744 | 912 
Charcoal hemoperfusion/hemofiltration | 744 | 912 
MTX toxicity | 720 | 912 
nephrotoxicity | 744 | 912 
hematological toxicity | 744 | 912 
infection risk | 936 | 936 
sepsis | 936 | 936 
acute on chronic kidney failure | 936 | 936 
dialysis | 744 | 912 
MTX-level | 744 | 912 
leucocytes | 744 | 912 
eGFR | 744 | 912 
hematological toxicity | 744 | 912 
infection | 936 | 936 
sepsis | 936 | 936 
acute kidney failure | 936 | 936 
cerebral radiation | 1092 | 1092 
PTLD | 48 | 1092 
diffuse large B-cell lymphoma | 48 | 48 
Ebstein-Barr virus | 48 | 48 
cerebral PTLD | 48 | 1092 
recurrence of PTLD | 720 | 720 
HDMTX therapy | 720 | 720 
MTX clearance | 744 | 912 
HFHD | 744 | 912 
MTX elimination | 744 | 912 
hemodialysis | 744 | 912 
hemodiafiltration | 744 | 912 
Charcoal hemoperfusion/hemofiltration | 744 | 912 
MTX toxicity | 720 | 912 
nephrotoxicity | 744 | 912 
hematological toxicity | 744 | 912 
infection risk | 936 | 936 
sepsis | 936 | 936 
acute on chronic kidney failure | 936 | 936 
dialysis | 744 | 912 
MTX-level | 744 | 912 
leucocytes | 744 | 912 
eGFR | 744 | 912 
hematological toxicity | 744 | 912 
infection | 936 | 936 
sepsis | 936 | 936 
acute kidney failure | 936 | 936 
cerebral radiation | 1092 | 1092 
PTLD | 48 | 1092 
diffuse large B-cell lymphoma | 48 | 48 
Ebstein-Barr virus | 48 | 48 
cerebral PTLD | 48 | 1092 
recurrence of PTLD | 720 | 720 
HDMTX therapy | 720 | 720 
MTX clearance | 744 | 912 
HFHD | 744 | 912 
MTX elimination | 744 | 912 
hemodialysis | 744 | 912 
hemodiafiltration | 744 | 912 
Charcoal hemoperfusion/hemofiltration | 744 | 912 
MTX toxicity | 720 | 912 
nephrotoxicity | 744 | 912 
hematological toxicity | 744 | 912 
infection risk | 936 | 936 
sepsis | 936 | 936 
acute on chronic kidney failure | 936 | 936 
dialysis | 744 | 912 
MTX-level | 744 | 912 
leucocytes | 744 | 912 
eGFR | 744 | 912 
hematological toxicity | 744 | 912 
infection | 936 | 936 
sepsis | 936 | 936 
acute kidney failure | 936 | 936 
cerebral radiation | 1092 | 1092 
PTLD | 48 | 1092 
diffuse large B-cell lymphoma | 48 | 48 
Ebstein-Barr virus | 48 | 48 
cerebral PTLD | 48 | 1092 
recurrence of PTLD | 720 | 720 
HDMTX therapy | 720 | 720 
MTX clearance | 744 | 912 
HFHD | 744 | 912 
MTX elimination | 744 | 912 
hemodialysis | 744 | 912 
hemodiafiltration | 744 | 912 
Charcoal hemoperfusion/hemofiltration | 744 | 912 
MTX toxicity | 720 | 912 
nephrotoxicity | 744 | 912 
hematological toxicity | 744 | 912 
infection risk | 936 | 936 
sepsis | 936 | 936 
acute on chronic kidney failure | 936 | 936 
dialysis | 744 | 912 
MTX-level | 744 | 912 
leucocytes | 744 | 912 
eGFR | 744 | 912 
hematological toxicity | 744 | 912 
infection | 936 | 936 
sepsis | 936 | 936 
acute kidney failure | 936 | 936 
cerebral radiation | 1092 | 1092 
PTLD | 48 | 1092 
diffuse large B-cell lymphoma | 48 | 48 
Ebstein-Barr virus | 48 | 48 
cerebral PTLD | 48 | 1092 
recurrence of PTLD | 720 | 720 
HDMTX therapy | 720 | 720 
MTX clearance | 744 | 912 
HFHD | 744 | 912 
MTX elimination | 744 | 912 
hemodialysis | 744 | 912 
hemodiafiltration | 744 | 912 
Charcoal hemoperfusion/hemofiltration | 744 | 912 
MTX toxicity | 720 | 912 
nephrotoxicity | 744 | 912 
hematological toxicity | 744 | 912 
infection risk | 936 | 936 
sepsis | 936 | 936 
acute on chronic kidney failure | 936 | 936 
dialysis | 744 | 912 
MTX-level | 744 | 912 
leucocytes | 744 | 912 
eGFR | 744 | 912 
hematological toxicity | 744 | 912 
infection | 936 | 936 
sepsis | 936 | 936 
acute kidney failure | 936 | 936 
cerebral radiation | 1092 | 1092 
PTLD | 48 | 1092 
diffuse large B-cell lymphoma | 48 | 48 
Ebstein-Barr virus | 48 | 48 
cerebral PTLD | 48 | 1092 
recurrence of PTLD | 720 | 720 
HDMTX therapy | 720 | 720 
MTX clearance | 744 | 912 
HFHD | 744 | 912 
MTX elimination | 744 | 912 
hemodialysis | 744 | 912 
hemodiafiltration | 744 | 912 
Charcoal hemoperfusion/hemofiltration | 744 | 912 
MTX toxicity | 720 | 912 
nephrotoxicity | 744 | 912 
hematological toxicity | 744 | 912 
infection risk | 936 | 936 
sepsis | 936 | 936 
acute on chronic kidney failure | 936 | 936 
dialysis | 744 | 912 
MTX-level | 744 | 912 
leucocytes | 744 | 912 
eGFR | 744 | 912 
hematological toxicity | 744 | 912 
infection | 936 | 936 
sepsis | 936 | 936 
acute kidney failure | 936 | 936 
cerebral radiation | 1092 | 1092 
PTLD | 48 | 1092 
diffuse large B-cell lymphoma | 48 | 48 
Ebstein-Barr virus | 48 | 48 
cerebral PTLD | 48 | 1092 
recurrence of PTLD | 720 | 720 
HDMTX therapy | 720 | 720 
MTX clearance | 744 | 912 
HFHD | 744 | 912 
MTX elimination | 744 | 912 
hemodialysis | 744 | 912 
hemodiafiltration | 744 | 912 
Charcoal hemoperfusion/hemofiltration | 744 | 912 
MTX toxicity | 720 | 912 
nephrotoxicity | 744 | 912 
hematological toxicity | 744 | 912 
infection risk | 936 | 936 
sepsis | 936 | 936 
acute on chronic kidney failure | 936 | 936 
dialysis | 744 | 912 
MTX-level | 744 | 912 
leucocytes | 744 | 912 
eGFR | 744 | 912 
hematological toxicity | 744 | 912 
infection | 936 | 936 
sepsis | 936 | 936 
acute kidney failure | 936 | 936 
cerebral radiation | 1092 | 1092 
PTLD | 48 | 1092 
diffuse large B-cell lymphoma | 48 | 48 
Ebstein-Barr virus | 48 | 48 
cerebral PTLD | 48 | 1092 
recurrence of PTLD | 720 | 720 
HDMTX therapy | 720 | 720 
MTX clearance | 744 | 912 
HFHD | 744 | 912 
MTX elimination | 744 | 912 
hemodialysis | 744 | 912 
hemodiafiltration | 744 | 912 
Charcoal hemoperfusion/hemofiltration | 744 | 912 
MTX toxicity | 720 | 912 
nephrotoxicity | 744 | 912 
hematological toxicity | 744 | 912 
infection risk | 936 | 936 
sepsis | 936 | 936 
acute on chronic kidney failure | 936 | 936 
dialysis | 744 | 912 
MTX-level | 744 | 912 
leucocytes | 744 | 912 
eGFR | 744 | 912 
hematological toxicity | 744 | 912 
infection | 936 | 936 
sepsis | 936 | 936 
acute kidney failure | 936 | 936 
cerebral radiation | 1092 | 1092 
PTLD | 48 | 1092 
diffuse large B-cell lymphoma | 48 | 48 
Ebstein-Barr virus | 48 | 48 
cerebral PTLD | 48 | 1092 
recurrence of PTLD | 720 | 720 
HDMTX therapy | 720 | 720 
MTX clearance | 744 | 912 
HFHD | 744 | 912 
MTX elimination | 744 | 912 
hemodialysis | 744 | 912 
hemodiafiltration | 744 | 912 
Charcoal hemoperfusion/hemofiltration | 744 | 912 
MTX toxicity | 720 | 912 
nephrotoxicity | 744 | 912 
hematological toxicity | 744 | 912 
infection risk | 936 | 936 
sepsis | 936 | 936 
acute on chronic kidney failure | 936 | 936 
dialysis | 744 | 912 
MTX-level | 744 | 912 
leucocytes | 744 | 912 
eGFR | 744 | 912 
hematological toxicity | 744 | 912 
infection | 936 | 936 
sepsis | 936 | 936 
acute kidney failure | 936 | 936 
cerebral radiation | 1092 | 1092 
PTLD | 48 | 1092 
diffuse large B-cell lymphoma | 48 | 48 
Ebstein-Barr virus | 48 | 48 
cerebral PTLD | 48 | 1092 
recurrence of PTLD | 720 | 720 
HDMTX therapy | 720 | 720 
MTX clearance | 744 | 912 
HFHD | 744 | 912 
MTX elimination | 744 | 912 
hemodialysis | 744 | 912 
hemodiafiltration | 744 | 912 
Charcoal hemoperfusion/hemofiltration | 744 | 912 
MTX toxicity | 720 | 912 
nephrotoxicity | 744 | 912 
hematological toxicity | 744 | 912 
infection risk | 936 | 936 
sepsis | 936 | 936 
acute on chronic kidney failure | 936 | 936 
dialysis | 744 | 912 
MTX-level | 744 | 912 
leucocytes | 744 | 912 
eGFR | 744 | 912 
hematological toxicity | 744 | 912 
infection | 936 | 936 
sepsis | 936 | 936 
acute kidney failure | 936 | 936 
cerebral radiation | 1092 | 1092 
PTLD | 48 | 1092 
diffuse large B-cell lymphoma | 48 | 48 
Ebstein-Barr virus | 48 | 48 
cerebral PTLD | 48 | 1092 
recurrence of PTLD | 720 | 720 
HDMTX therapy | 720 | 720 
MTX clearance | 744 | 912 
HFHD | 744 | 912 
MTX elimination | 744 | 912 
hemodialysis | 744 | 912 
hemodiafiltration | 744 | 912 
Charcoal hemoperfusion/hemofiltration | 744 | 912 
MTX toxicity | 720 | 912 
nephrotoxicity | 744 | 912 
hematological toxicity | 744 | 912 
infection risk | 936 | 936 
sepsis | 936 | 936 
acute on chronic kidney failure | 936 | 936 
dialysis | 744 | 912 
MTX-level | 744 | 912 
leucocytes | 744 | 912 
eGFR | 744 | 912 
hematological toxicity | 744 | 912 
infection | 936 | 936 
sepsis | 936 | 936 
acute kidney failure | 936 | 936 
cerebral radiation | 1092 | 1092 
PTLD | 48 | 1092 
diffuse large B-cell lymphoma | 48 | 48 
Ebstein-Barr virus | 48 | 48 
cerebral PTLD | 48 | 1092 
recurrence of PTLD | 720 | 720 
HDMTX therapy | 720 | 720 
MTX clearance | 744 | 912 
HFHD | 744 | 912 
MTX elimination | 744 | 912 
hemodialysis | 744 | 912 
hemodiafiltration | 744 | 912 
Charcoal hemoperfusion/hemofiltration | 744 | 912 
MTX toxicity | 720 | 912 
nephrotoxicity | 744 | 912 
hematological toxicity | 744 | 912 
infection risk | 936 | 936 
sepsis | 936 | 936 
acute on chronic kidney failure | 936 | 936 
dialysis | 744 | 912 
MTX-level | 744 | 912 
leucocytes | 744 | 912 
eGFR | 744 | 912 
hematological toxicity | 744 | 912 
infection | 936 | 936 
sepsis | 936 | 936 
acute kidney failure | 936 | 936 
cerebral radiation | 1092 | 1092 
PTLD | 48 | 1092 
diffuse large B-cell lymphoma | 48 | 48 
Ebstein-Barr virus | 48 | 48 
cerebral PTLD | 48 | 1092 
recurrence of PTLD | 720 | 720 
HDMTX therapy | 720 | 720 
MTX clearance | 744 | 912 
HFHD | 744 | 912 
MTX elimination | 744 | 912 
hemodialysis | 744 | 912 
hemodiafiltration | 744 | 912 
Charcoal hemoperfusion/hemofiltration | 744 | 912 
MTX toxicity | 720 | 912 
nephrotoxicity | 744 | 912 
hematological toxicity | 744 | 912 
infection risk | 936 | 936 
sepsis | 936 | 936 
acute on chronic kidney failure | 936 | 936 
dialysis | 744 | 912 
MTX-level | 744 | 912 
leucocytes | 744 | 912 
eGFR | 744 | 912 
hematological toxicity | 744 | 912 
infection | 936 | 936 
sepsis | 936 | 936 
acute kidney failure | 936 | 936 
cerebral radiation | 1092 | 1092 
PTLD | 48 | 1092 
diffuse large B-cell lymphoma | 48 | 48 
Ebstein-Barr virus | 48 | 48 
cerebral PTLD | 48 | 1092 
recurrence of PTLD | 720 | 720 
HDMTX therapy | 720 | 720 
MTX clearance | 744 | 912 
HFHD | 744 | 912 
MTX elimination | 744 | 912 
hemodialysis | 744 | 912 
hemodiafiltration | 744 | 912 
Charcoal hemoperfusion/hemofiltration | 744 | 912 
MTX toxicity | 720 | 912 
nephrotoxicity | 744 | 912 
hematological toxicity | 744 | 912 
infection risk | 936 | 936 
sepsis | 936 | 936 
acute on chronic kidney failure | 936 | 936 
dialysis | 744 | 912 
MTX-level | 744 | 912 
leucocytes | 744 | 912 
eGFR | 744 | 912 
hematological toxicity | 744 | 912 
infection | 936 | 936 
sepsis | 936 | 936 
acute kidney failure | 936 | 936 
cerebral radiation | 1092 | 1092 
PTLD | 48 | 1092 
diffuse large B-cell lymphoma | 48 | 48 
Ebstein-Barr virus | 48 | 48 
cerebral PTLD | 48 | 1092 
recurrence of PTLD | 720 | 720 
HDMTX therapy | 720 | 720 
MTX clearance | 744 | 912 
HFHD | 744 | 912 
MTX elimination | 744 | 912 
hemodialysis | 744 | 912 
hemodiafiltration | 744 | 912 
Charcoal hemoperfusion/hemofiltration | 744 | 912 
MTX toxicity | 720 | 912 
nephrotoxicity | 744 | 912 
hematological toxicity | 744 | 912 
infection risk | 936 | 936 
sepsis | 936 | 936 
acute on chronic kidney failure | 936 | 936 
dialysis | 744 | 912 
MTX-level | 744 | 912 
leucocytes | 744 | 912 
eGFR | 744 | 912 
hematological toxicity | 744 | 912 
infection | 936 | 936 
sepsis | 936 | 936 
acute kidney failure | 936 | 936 
cerebral radiation | 1092 | 1092 
PTLD | 48 | 1092 
diffuse large B-cell lymphoma | 48 | 48 
Ebstein-Barr virus | 48 | 48 
cerebral PTLD | 48 | 1092 
recurrence of PTLD | 720 | 720 
HDMTX therapy | 720 | 720 
MTX clearance | 744 | 912 
HFHD | 744 | 912 
MTX elimination | 744 | 912 
hemodialysis | 744 | 912 
hemodiafiltration | 744 | 912 
Charcoal hemoperfusion/hemofiltration | 744 | 912 
MTX toxicity | 720 | 912 
nephrotoxicity | 744 | 912 
hematological toxicity | 744 | 912 
infection risk | 936 | 936 
sepsis | 936 | 936 
acute on chronic kidney failure | 936 | 936 
dialysis | 744 | 912 
MTX-level | 744 | 912 
leucocytes | 744 | 912 
eGFR | 744 | 912 
hematological toxicity | 744 | 912 
infection | 936 | 936 
sepsis | 936 | 936 
acute kidney failure | 936 | 936 
cerebral radiation | 1092 | 1092 
PTLD | 48 | 1092 
diffuse large B-cell lymphoma | 48 | 48 
Ebstein-Barr virus | 48 | 48 
cerebral PTLD | 48 | 1092 
recurrence of PTLD | 720 | 720 
HDMTX therapy | 720 | 720 
MTX clearance | 744 | 912 
HFHD | 744 | 912 
MTX elimination | 744 | 912 
hemodialysis | 744 | 912 
hemodiafiltration | 744 | 912 
Charcoal hemoperfusion/hemofiltration | 744 | 912 
MTX toxicity | 720 | 912 
nephrotoxicity | 744 | 912 
hematological toxicity | 744 | 912 
infection risk | 936 | 936 
sepsis | 936 | 936 
acute on chronic kidney failure | 936 | 936 
dialysis | 744 | 912 
MTX-level | 744 | 912 
leucocytes | 744 | 912 
eGFR | 744 | 912 
hematological toxicity | 744 | 912 
infection | 936 | 936 
sepsis | 936 | 936 
acute kidney failure | 936 | 936 
cerebral radiation | 1092 | 1092 
PTLD | 48 | 1092 
diffuse large B-cell lymphoma | 48 | 48 
Ebstein-Barr virus | 48 | 48 
cerebral PTLD | 48 | 1092 
recurrence of PTLD | 720 | 720 
HDMTX therapy | 720 | 720 
MTX clearance | 744 | 912 
HFHD | 744 | 912 
MTX elimination | 744 | 912 
hemodialysis | 744 | 912 
hemodiafiltration | 744 | 912 
Charcoal hemoperfusion/hemofiltration | 744 | 912 
MTX toxicity | 720 | 912 
nephrotoxicity | 744 | 912 
hematological toxicity | 744 | 912 
infection risk | 936 | 936 
sepsis | 936 | 936 
acute on chronic kidney failure | 936 | 936 
dialysis | 744 | 912 
MTX-level | 744 | 912 
leucocytes | 744 | 912 
eGFR | 744 | 912 
hematological toxicity | 744 | 912 
infection | 936 | 936 
sepsis | 936 | 936 
acute kidney failure | 936 | 936 
cerebral radiation | 1092 | 1092 
PTLD | 48 | 1092 
diffuse large B-cell lymphoma | 48 | 48 
Ebstein-Barr virus | 48 | 48 
cerebral PTLD | 48 | 1092 
recurrence of PTLD | 720 | 720 
HDMTX therapy | 720 | 720 
MTX clearance | 744 | 912 
HFHD | 744 | 912 
MTX elimination | 744 | 912 
hemodialysis | 744 | 912 
hemodiafiltration | 744 | 912 
Charcoal hemoperfusion/hemofiltration | 744 | 912 
MTX toxicity | 720 | 912 
nephrotoxicity | 744 | 912 
hematological toxicity | 744 | 912 
infection risk | 936 | 936 
sepsis | 936 | 936 
acute on chronic kidney failure | 936 | 936 
dialysis | 744 | 912 
MTX-level | 744 | 912 
leucocytes | 744 | 912 
eGFR | 744 | 912 
hematological toxicity | 744 | 912 
infection | 936 | 936 
sepsis | 936 | 936 
acute kidney failure | 936 | 936 
cerebral radiation | 1092 | 1092 
PTLD | 48 | 1092 
diffuse large B-cell lymphoma | 48 | 48 
Ebstein-Barr virus | 48 | 48 
cerebral PTLD | 48 | 1092 
recurrence of PTLD | 720 | 720 
HDMTX therapy | 720 | 720 
MTX clearance | 744 | 912 
HFHD | 744 | 912 
MTX elimination | 744 | 912 
hemodialysis | 744 | 912 
hemodiafiltration | 744 | 912 
Charcoal hemoperfusion/hemofiltration | 744 | 912 
MTX toxicity | 720 | 912 
nephrotoxicity | 744 | 912 
hematological toxicity | 744 | 912 
infection risk | 936 | 936 
sepsis | 936 | 936 
acute on chronic kidney failure | 936 | 936 
dialysis | 744 | 912 
MTX-level | 744 | 912 
leucocytes | 744 | 912 
eGFR | 744 | 912 
hematological toxicity | 744 | 912 
infection | 936 | 936 
sepsis | 936 | 936 
acute kidney failure | 936 | 936 
cerebral radiation | 1092 | 1092 
PTLD | 48 | 1092 
diffuse large B-cell lymphoma | 48 | 48 
Ebstein-Barr virus | 48 | 48 
cerebral PTLD | 48 | 1092 
recurrence of PTLD | 720 | 720 
HDMTX therapy | 720 | 720 
MTX clearance | 744 | 912 
HFHD | 744 | 912 
MTX elimination | 744 | 912 
hemodialysis | 744 | 912 
hemodiafiltration | 744 | 912 
Charcoal hemoperfusion/hemofiltration | 744