49 years old | 0
male | 0
admitted to the hospital | 0
spider bite | -120
backed up into a spider web | -120
mild elevation in AST | -72
mild elevation in ALT | -72
elevation in total bilirubin | -72
elevation in white blood cell count | -72
elevation in hemoglobin | -72
elevation in platelet count | -72
orange urine | -72
no blood in urine | -72
prescription for doxycycline | -72
did not get doxycycline | -72
worsening rash | -48
fever | -48
body aches | -48
discoloration of urine | -48
febrile | -48
elevated heart rate | -48
elevated blood pressure | -48
elevated respirations | -48
elevated oxygen saturation | -48
normal creatinine | -48
elevated total bilirubin | -48
elevated AST | -48
elevated ALT | -48
elevated creatinine kinase | -48
elevated white blood cell count | -48
elevated hemoglobin | -48
elevated platelet count | -48
elevated lactic acid | -48
sepsis criteria met | -48
recommended admission | -48
refused admission | -48
pain around the bite | -24
extension to chest | -24
fevers | -24
body aches | -24
shortness of breath | -24
nausea | -24
vomiting | -24
black colored urine | -24
admitted to the hospital | 0
intravenous vancomycin | 0
intravenous piperacillin/tazobactam | 0
admitted to intensive care unit | 0
nephrology consultation | 0
acute renal failure | 0
hemolysis | 0
elevated bicarbonate level | 0
elevated BUN | 0
elevated creatinine | 0
elevated total bilirubin | 0
elevated AST | 0
elevated ALT | 0
elevated creatinine kinase | 0
elevated lactate dehydrogenase | 0
elevated haptoglobin | 0
elevated white blood cell count | 0
elevated hemoglobin | 0
elevated platelet count | 0
elevated reticulocyte count | 0
direct Coombs test positive for C3 | 0
direct Coombs test negative for IgG | 0
peripheral smear showed normocytic anemia | 0
peripheral smear showed spherocytes | 0
peripheral smear showed nucleated red blood cells | 0
peripheral smear showed leukocytosis | 0
peripheral smear showed left shifted neutrophil series | 0
peripheral smear showed eosinophilia | 0
transfused two units packed red blood cells | 0
hematology consultation | 0
supportive care recommended | 0
transfusions recommended | 0
plasmapheresis recommended | 24
initiation of plasmapheresis | 48
one-to-one exchange with albumin | 48
transfused one unit packed red blood cells | 48
improvement in laboratory evaluation | 72
continuation of plasmapheresis | 72
broadened antibiotics | 72
repeat ultrasound | 72
no evidence of fluid collection or abscess | 72
second treatment of plasmapheresis | 96
improvement in laboratory evaluation | 120
no additional blood transfusions needed | 120
no additional plasmapheresis recommended | 120
started folic acid | 120
underwent three sessions of hemodialysis | 120
stopped hemodialysis | 120
supportive management recommended | 120
discharged | 168
close follow-up recommended | 168
outpatient labs recommended | 168