31 years old | 0
male | 0
motor vehicle accident | -12000
severe head injury | -12000
cervical spine fracture | -12000
intubated | -12000
spine fixed with plate and screw | -12000
discharged from hospitalization | -12000
paraplegic | -12000
recurrent chest infections | -12000
treated conservatively with antibiotics | -12000
referred to cardiothoracic unit | -24
chest x-ray showed widened mediastinum | -24
initial laboratory investigations | -24
Hemoglobin 11.3 g/dL | -24
hematocrit 35% | -24
Mean corpuscular volume 67.7 fL | -24
mean corpuscular hemoglobin 21.8 pg | -24
albumin 2.7 g/L | -24
creatinine 0.5 μmol/L | -24
Na 135 mmol/L | -24
erythrocyte sedimentation rate 93 mm/h | -24
further radiological assessment | -24
computed tomography of the neck, cervical spine, and chest | -24
superior mediastinal collection | -24
chronic esophageal perforation | -24
swallowing test | -24
upper gastroesophageal endoscopy | -24
upper esophageal perforation | -24
erosion of the cervical spine plate and screw into the esophagus | -24
surgical approach | -24
neck exploration | -24
plate removed | -24
perforation repaired | -24
limited thoracotomy | -24
extensive pleural adhesions | -24
feeding jejunostomy tube created | -24
surgical site infection | 168
exploration and drainage | 168
antimicrobial therapy | 168
lengthy post-operative course | 168
repeated episodes of sepsis | 168
admissions to intensive care unit | 168
bronchoscopies | 168
exchanging the tracheostomy | 168
acute surgical abdomen | 168
exploration and drainage of multiple intra-abdominal abscess collections | 168
persistent status epilepticus | 168
cardiac arrest | 720
XDR-P. aeruginosa strain isolated | 1296
elevated resistance to antimicrobial agents | 1296
ceftolozane-tazobactam | 1296
ceftazidime-avibactam | 1296
whole genome sequencing | 1296
genomic islands | 1296
mobile genetic elements | 1296
resistance determinants | 1296
virulence genes | 1296
phageomics | 1296
blaOXA-10 | 1296
blaOXA-50 | 1296
blaVEB-9 | 1296
blaPAO | 1296
PDC-11 | 1296
Metallo-β-lactamases | 1296
aminoglycoside resistant determinants | 1296
fluoroquinolone-related resistance genes | 1296
phenicol resistance gene | 1296
tetracycline resistance genes | 1296
efflux pump proteins | 1296
MexCD-OprJ | 1296
CorC | 1296
MacA | 1296
KefA | 1296
MexX | 1296
MexA | 1296
MexE | 1296
virulence factor identification | 1296
VFDB | 1296
VFanalyser | 1296
type secretion system proteins | 1296
T1SS | 1296
T2SS | 1296
T3SS | 1296
T4SS | 1296
T5SS | 1296
T6SS | 1296
T7SS | 1296
bacteriophages | 1296
PHAST | 1296
CRISPR | 1296
CRISPR-Cas systems | 1296
genomic islands | 1296
Island Viewer | 1296
mobile genetic elements | 1296
integrons | 1296
conjugative transposons | 1296
resistance genes | 1296
virulence factors | 1296
secretion systems | 1296
biofilm-specific antibiotic resistance | 1296
T6SS-deficient P. aeruginosa mutants | 1296
prophages | 1296
phage therapy | 1296
P. aeruginosa blood steam infections | 1296
whole genome sequencing | 1296
AMR surveillance systems | 1296
resistant foci | 1296
genomic basis of resistance | 1296
virulence | 1296
clone dissemination | 1296
mobile genetic elements | 1296
AMR vehicles | 1296
pandrug-resistant | 1296
colistin BMD | 1296
CLSI | 1296
VITEK 2 | 1296
novel cephalosporins | 1296
cefiderocol | 1296
carbapenem-beta-lactamase | 1296
imipenem-cilastatin-relebactam | 1296
mechanism of potential resistance | 1296
cross-resistance | 1296
existing drugs | 1296
clinical use | 1296
intense preventive measures | 1296
healthcare facilities | 1296
debilitated patients | 1296
infections | 1296
virulent | 1296
drug-resistant strains | 1296