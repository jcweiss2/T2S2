73 years old | 0
    man | 0
    hypertension | 0
    diabetes mellitus | 0
    percutaneous coronary intervention | -17520
    aspirin 100 mg daily | -17520
    COVID-19 | -672
    SARS-CoV-2 positive RT-PCR | -672
    admitted to Pohang Medical Center | -672
    fever 37.7℃ | -672
    cough | -672
    chest radiography hazy streaky density both lungs | -672
    hydroxychloroquine treatment | -672
    pneumonia | -672
    hypotension | -672
    melena | -672
    transferred to Samsung Medical Center | -672
    vital signs stabilized | -672
    observation without additional treatment | -672
    expelled large quantity of melena | 0
    hypotension | 0
    tachycardia | 0
    SpO2 80% | 0
    hemoglobin 6.3 mg/dl | 0
    blood transfusion | 0
    endotracheal intubation | 0
    arterial catheter insertion | 0
    central venous catheter insertion | 0
    esophagogastroduodenoscopy | 0
    duodenal ulcer without active bleeding | 0
    risk of re-bleeding | 0
    computed tomography not possible | 0
    embolization not possible | 0
    transferred to our hospital | 24
    COVID-19 patient care environment prepared | 24
    endoscopic hemoclipping | 24
    embolization | 24
    surgery considered | 24
    abdominal pain | 24
    chest X-ray subphrenic free air | 24
    pneumoperitoneum | 24
    suspected duodenal ulcer perforation | 24
    emergency surgery planned | 24
    fever 37.8℃ | 24
    preoperative vital signs stable | 24
    ECG normal sinus rhythm | 24
    chest radiography peripheral lung consolidation | 24
    aggravated pneumonia | 24
    hemoglobin 11.1 mg/dl | 24
    C-reactive protein 103 mg/L | 24
    arterial blood gas analysis | 24
    mechanical ventilation | 24
    remifentanil infusion | 24
    intravenous antibiotics | 24
    SARS-CoV-2 positive RT-PCR | 24
    severe pneumonia | 24
    persistent SARS-CoV-2 detection | 24
    nosocomial transmission risk | 24
    PPE worn | 24
    negative-pressure operating room | 24
    PAPR hood | 24
    N95 masks | 24
    protective suits | 24
    double gloves | 24
    boots | 24
    shoe covers | 24
    aprons | 24
    face shields | 24
    sedated patient transferred to operating room | 24
    portable ventilator with HEPA filter | 24
    anesthesiologist and nurse standby | 24
    patient transferred to operating room | 24
    stretcher disinfected | 24
    invasive monitoring commenced | 24
    endotracheal tube clamped | 24
    anesthesia machine connected | 24
    end-tidal carbon dioxide monitoring | 24
    general anesthesia induced | 24
    propofol 0.5 mg/kg | 24
    rocuronium 0.6 mg/kg | 24
    esophageal temperature probe placed | 24
    temperature monitoring | 24
    sevoflurane 2.0% | 24
    remifentanil infusion | 24
    rocuronium infusion 0.15 mg/kg/h | 24
    lung-protective mechanical ventilation | 24
    operating room pressure maintained | 24
    items delivered via anteroom | 24
    arterial blood gas sample sent | 24
    operation duration 120 min | 24
    perforated ulcer found | 24
    pyloric exclusion | 24
    primary closure | 24
    gastrojejunostomy | 24
    midazolam 0.07 mg/kg | 24
    rocuronium 0.3 mg/kg | 24
    sedation during transfer | 24
    closed in-line tracheal suction | 24
    ventilator switched to manual mode | 24
    adjustable pressure-limiting valve opened | 24
    tracheal tube clamped | 24
    stretcher cart placed in anteroom | 24
    monitoring continued | 24
    oxygen supplied via Ambu bag | 24
    patient transferred to ICU | 24
    disposable equipment discarded | 24
    reusable equipment disinfected | 24
    patient monitored in ICU | 24
    antibiotics administered | 24
    hydroxychloroquine administered | 24
    no surgical complications | 24
    pneumonia treatment continued | 168
    C-reactive protein elevated | 168
    fever 37.3-38.8℃ | 168
    SARS-CoV-2 positive RT-PCR | 168
    chest radiography increased pneumonic infiltration | 168
    pleural effusion | 168
    vital signs stable | 168
    fever 39.5℃ | 216
    hypotension | 216
    fluid administration | 216
    norepinephrine administration | 216
    septic shock diagnosed | 216
    patient expired | 240