79 years old | 0
male | 0
German descent | 0
admitted to the hospital | 0
abdominal pain | -1
collapsed | -1
pale | -1
hypotensive | -1
bradycardic | -1
slow atrial fibrillation | -1
ruptured infrarenal abdominal aortic aneurysm | -1
open repair of the aneurysm | 0
significant blood loss | 0
cell saver returning 5.5 L of blood | 0
received 6 units of packed cells | 0
received 4 units of fresh-frozen plasma | 0
received 6 units of cryoprecipitate | 0
received 1 pooled bag of platelets | 0
received 4 L of crystalloids | 0
intubated | 0
requiring a high dose of vasopressors | 0
hypertension | -672
benign prostatic hypertrophy | -672
atorvastatin | -672
amlodipine | -672
dutasteride-tamsulosin | -672
allergy to penicillin | -672
rash | -672
unstable postoperatively | 0
acute kidney injury | 24
mild abdominal hypertension | 24
sedation | 24
paralysis | 24
enteral feeding not tolerated | 24
total parenteral nutrition | 24
extubated | 240
re-intubated | 240
respiratory failure | 240
sepsis | 240
fever | 240
leukocytosis | 240
vasopressors | 240
meropenem commenced | 240
vancomycin commenced | 240
Serratia marcescens isolated | 240
hemodynamic improvement | 288
renal function improvement | 288
ventilator-dependent | 288
encephalopathic | 288
tracheostomy | 336
hyperbilirubinemia | 336
mildly deranged liver transaminase levels | 336
biochemical markers of cholestasis | 336
bile duct obstruction | 336
cholelithiasis not found | 336
dilation of the biliary ducts not found | 336
bilirubin increased to 200 µmol/L | 336
endoscopic retrograde cholangiopancreatography | 336
transcutaneous hepatic cholangiography | 336
widely patent right and left hepatic and common biliary ducts | 336
smooth tapering toward the ampulla | 336
cystic duct patent | 336
stent inserted in the common bile duct | 336
8.5-French external biliary drain inserted | 336
no improvement after cholangiography and insertion of the external biliary drain | 336
bilirubin level continued to rise | 336
biliary drain producing up to 600 mL of bile | 336
direct bilirubin level reached 300 µmol/L | 432
conjugated bilirubin level of 169 µmol/L | 432
no evidence of an intra-abdominal collection | 432
no bleeding | 432
no new pathology | 432
stent and bile ducts remained widely patent | 432
meropenem changed to ciprofloxacin | 432
decrease in bilirubin level | 456
meropenem restarted | 504
increase in serum bilirubin level | 504
meropenem discontinued | 552
ciprofloxacin and metronidazole commenced | 552
dramatic decrease in bilirubin level | 552
bilirubin level normalized | 720
biliary drain plugged and removed | 720
prolonged ICU stay | 720
ventilator-dependent | 720
decannulated | 2160
discharged from ICU | 2160
discharged from hospital | 2160