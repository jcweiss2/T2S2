69 years old | 0
male | 0
admitted to the hospital | 0
local recurrence of a prostate carcinoma metastatic to bone | -4320
endoscopic prostatectomy | -4320
adjuvant radiotherapy | -4320
chemotherapy with docetaxel | 0
deterioration of general condition | 0
tumor induced anemia | 0
Hgb 7.2 g/dL | 0
serum prostate specific antigen levels > 200 ng/mL | 0
upper stomach pain | 168
diarrhea | 168
cholecystitis | 168
increased CRP: 280 mg/L | 168
increased procalcitonin: 6.52 ng/mL | 168
open cholecystectomy | 168
calculated anti-infective therapy with metronidazole | 168
calculated anti-infective therapy with ceftriaxone | 168
blood cultures obtained | 168
purulent gangrenous gallbladder | 168
ileostomy performed | 168
multiple adhesions | 168
necrotizing/gangrenous cholecystitis | 168
ulcero-phlegmonous cholecystitis | 168
fibrinous pericholecystitis | 168
cholecystolithiasis | 168
intraoperative culture taken | 168
transferred to intensive care unit | 168
extubated | 168
vasopressor therapy ended | 168
postoperative course uneventful | 336
transferred to ward | 336
discharged | 336
blood cultures taken | 168
F. plautii detected in anaerobic blood culture | 216
gram positive rod | 216
identified via MALDI-TOF | 216
cultured on Columbia agar | 216
slow growth | 288
Maldi-TOF repeated with score > 2.0 | 288
16S rRNA sequencing confirmed F. plautii | 288
grey glassy colonies formed | 288
resistance testing results | 336
penicillin MIC 0.5 mg/L | 336
ampicillin MIC 0.5 mg/L | 336
cefuroxime MIC 4.0 mg/L | 336
ceftriaxone MIC 0.75 mg/L | 336
piperacillin/tazobactam MIC 0.19 mg/L | 336
meropenem MIC 0.023 mg/L | 336
imipenem MIC 0.064 mg/L | 336
ertapenem MIC 0.023 mg/L | 336
gentamicin MIC 4.0 mg/L | 336
cotrimoxazole MIC ≥32 mg/L | 336
ciprofloxacin MIC ≥32 mg/L | 336
levofloxacin MIC 2.0 mg/L | 336
moxifloxacin MIC 0.5 mg/L | 336
vancomycin MIC 2.0 mg/L | 336
teicoplanin MIC 0.25 mg/L | 336
daptomycin MIC 8.0 mg/L | 336
linezolid MIC 3.0 mg/L | 336
metronidazole MIC 0.25 mg/L | 336
clindamycin MIC 0.38 mg/L | 336
tetracyclin MIC 0.094 mg/L | 336
tigecyclin MIC 0.0160 mg/L | 336
chloramphenicol MIC 0.125 mg/L | 336
rifampicin MIC 3.0 mg/L | 336
intraabdominal cultures showed no growth | 168
additional blood cultures remained sterile | 168
immunosuppression due to prostate cancer | 0
immunosuppression due to docetaxel treatment | 0
acute gangrenous cholecystitis | 168
F. plautii bloodstream infection | 216
