72 years old | 0
male | 0
high-grade fever | -96
influenza B virus infection | -96
wife diagnosed with influenza B virus infection | -168
daughters diagnosed with influenza B virus infection | -168
rapid test positive for influenza B antigens | -96
oseltamivir administered | -96
persistent fever | -48
dyspnea at rest | -48
admitted to hospital | 0
temperature 38.7°C | 0
blood pressure 117/80 mmHg | 0
heart rate 76 beats/min | 0
oxygen saturation level 88% | 0
fine crackles in lung fields | 0
white blood cell count 7400/mm3 | 0
C-reactive protein 18.1 mg/dL | 0
aspartate transaminase 91 IU/L | 0
L-lactate dehydrogenase 362 IU/L | 0
creatine kinase 793 IU/L | 0
Krebs von den Lungen-6 1772 U/mL | 0
hypoxemia | 0
PaO2 = 72 Torr | 0
nasal oxygen inhalation | 0
ground-glass opacity in lung fields | 0
chest computed tomography showed diffuse ground-glass opacity | 0
Gram staining negative | 0
Ziehl-Neelsen staining negative | 0
periodic acid-Schiff stain negative | 0
sputum culture negative | 0
blood cultures negative | 0
high-flow nasal oxygen support | 0
intravenous peramivir | 0
antibiotics administered | 0
piperacillin/tazobactam | 0
levofloxacin | 0
reticular shadow on chest CT worsened | 72
PaO2/FiO2 ratio deteriorated | 72
diagnosed with severe ARDS | 72
mechanical ventilation proposed | 72
high levels of positive end-expiratory pressure proposed | 72
patient refused intubation | 72
polymyxin B-immobilized fiber column hemoperfusion | 72
intravenous methylprednisolone | 144
noninvasive positive pressure ventilation support | 144
immunosuppressant therapy | 144
intravenous cyclophosphamide | 144
patient's condition worsened | 129*24
died | 129*24
autopsy performed | 129*24
diffuse alveolar damage | 129*24
prominent hyaline membranes | 129*24
no specific abnormality in other organs | 129*24