33 years old | 0
female | 0
admitted to the hospital | 0
recurrent episodes of headache | -4320
myalgia | -4320
occasional episodes of nausea | -4320
vomiting | -4320
hypotension | -4320
leucocytosis | -4320
treated with broad-spectrum antibiotics | -4320
anasarca | -720
no hematuria | -720
no reduction in urine output | -720
afebrile | 0
blood pressure 110/70 mmHg | 0
no postural hypotension | 0
nephrotic range proteinuria | 0
microscopic hematuria | 0
hypoalbuminemia | 0
hypercholesterolemia | 0
hypertriglyceridemia | 0
serum creatinine 1.08 mg/dl | 0
leucocytosis | 0
started on diuretics | 0
intravenous albumin | 0
blood culture | 0
no pathogen growth | 0
renal biopsy | 0
mesangial matrix increase | 0
hypercellularity | 0
immunofluorescence negative | 0
idiopathic unsampled focal and segmental glomerulosclerosis | 0
started on prednisolone | 0
discharged | 0
myalgia | 120
giddiness | 120
weakness | 120
no fever | 120
tachycardia | 120
tachypnea | 120
hypotension | 120
leucocytosis | 120
neutrophilic predominance | 120
elevated serum procalcitonin | 120
started on meropenem | 120
leukocyte count increased | 144
imaging chest and abdomen | 144
no focus of sepsis | 144
managed in ICU | 144
inotropic support | 144
clinical improvement | 192
reduction of inotropic requirement | 192
normalization of leukocyte count | 288
blood culture grew non-O1, non-O139 V. cholerae | 288
stool culture | 288
no pathogen growth | 288
sea-water exposure | -2688
completed meropenem | 432
repeat blood culture sterile | 432
discharged | 432
continue prednisolone | 432
