65 years old | 0 | 0 
female | 0 | 0 
admitted to the hospital | 0 | 0 
recurrent fever | -744 | 0 
nausea | -168 | 0 
vomiting | -168 | 0 
neutrophil count 6.96×10^9/L ↑ | 0 | 0 
monocyte count 0.86×10^9/L ↑ | 0 | 0 
lymphocyte percentage 14.9% ↓ | 0 | 0 
red blood cell count 3.17×10^12/L ↓ | 0 | 0 
hemoglobin content 87 g/L ↓ | 0 | 0 
hematocrit 0.28 L/L ↓ | 0 | 0 
average red blood cell hemoglobin concentration 312 g/L ↓ | 0 | 0 
platelet count 363×10^9/L ↑ | 0 | 0 
platelet distribution width 8.3 fl ↓ | 0 | 0 
C-reactive protein (CRP) 52.01 mg/L ↑ | 0 | 0 
diagnosed with secondary infectious thrombocytopenia | 0 | 0 
diagnosed with gram-negative bacilli septicemia (Klebsiella pneumoniae) | 0 | 0 
diagnosed with liver abscess | 0 | 0 
diagnosed with bilateral lung inflammation | 0 | 0 
diagnosed with type 2 diabetes | 0 | 0 
diagnosed with hypertension grade 3 (extremely high risk) | 0 | 0 
treated with vancomycin | 0 | 168 
treated with caspofungin | 0 | 168 
treated with dexamethasone | 0 | 168 
treated with posaconazole oral suspension | 0 | 168 
liver abscess puncture and drainage treatment | 0 | 168 
inflammatory indexes decreased | 168 | 168 
light perception disappeared in the left eye | 168 | 168 
eyelid redness and pain | 168 | 168 
purulent secretion | 168 | 168 
repeated fever | 168 | 168 
left-sided headache | 168 | 168 
diagnosed with endogenous endophthalmitis (left) | 168 | 168 
diagnosed with orbital cellulitis (left) | 168 | 168 
diagnosed with rubeosis iridis (left) | 168 | 168 
diagnosed with exudative retinal detachment (left) | 168 | 168 
diagnosed with diabetic retinopathy (right) | 168 | 168 
intravitreal injection with vancomycin | 168 | 336 
intravitreal injection with ceftazidime | 168 | 336 
symptoms relieved | 336 | 336 
systemic infection under control | 336 | 336 
left eyeball enucleation | 336 | 336 
fever again after the operation | 336 | 336 
treated with moxifloxacin | 336 | 504 
treated with sulperazon | 336 | 504 
temperature elevated again | 504 | 504 
CT examination | 504 | 504 
inflammation of both lungs | 504 | 504 
pericardial effusion | 504 | 504 
bilateral pleural thickening and effusion | 504 | 504 
atelectasis in right inferior lobe | 504 | 504 
liver cyst | 504 | 504 
liver abscess | 504 | 504 
right renal cyst | 504 | 504 
myoma of the uterus | 504 | 504 
history of hypertension | -8760 | 0 
highest blood pressure of 180/100 mmHg | -8760 | 0 
oral valsartan | -8760 | 0 
blood pressure controlled at 140/80 mmHg | -8760 | 0 
no special history of other systematic diseases | 0 | 0 
no history of surgery | 0 | 0 
no history of blood transfusion | 0 | 0 
no history of drug allergy | 0 | 0 
diagnosed with sepsis | 0 | 0 
diagnosed with secondary thrombocytopenia | 0 | 0 
diagnosed with liver abscess | 0 | 0 
diagnosed with gram-negative bacilli sepsis (Klebsiella pneumoniae) | 0 | 0 
diagnosed with infection of lumbar vertebrae | 0 | 0 
diagnosed with mesenteric panniculitis | 0 | 0 
diagnosed with pelvic effusion | 0 | 0 
diagnosed with pericardial effusion | 0 | 0 
diagnosed with suppurative endophthalmitis (left) | 0 | 0 
diagnosed with orbital cellulitis (left) | 0 | 0 
diagnosed with retinal detachment (left) | 0 | 0 
diagnosed with choroidal detachment (left) | 0 | 0 
diagnosed with type 2 diabetes retinopathy (right) | 0 | 0 
diagnosed with cortical senile cataract (right, immature stage) | 0 | 0 
diagnosed with type 2 diabetes | 0 | 0 
diagnosed with type 2 diabetes nephropathy stage I | 0 | 0 
diagnosed with type 2 diabetic peripheral neuropathy | 0 | 0 
diagnosed with hypertension grade 3 (extremely high risk) | 0 | 0 
diagnosed with hepatic cyst | 0 | 0 
diagnosed with renal cyst | 0 | 0 
diagnosed with hypoproteinemia | 0 | 0 
diagnosed with coronary atherosclerotic heart disease | 0 | 0 
diagnosed with lacunar cerebral infarction | 0 | 0 
diagnosed with moderate anemia | 0 | 0 
diagnosed with risk of malnutrition | 0 | 0 
convulsion with unconsciousness | 504 | 504 
transferred to the respiratory intensive care unit | 504 | 504 
CT examination | 504 | 504 
lacunar infarction | 504 | 504 
encephalomalacia | 504 | 504 
bilateral pleural effusion | 504 | 504 
lower lobe of the right lung insufficiently inflated | 504 | 504 
coma | 504 | 504 
unresponsive | 504 | 504 
slight neck resistance | 504 | 504 
weak light response of the eye | 504 | 504 
uncooperative physical examination of limb muscle strength | 504 | 504 
low muscle tension | 504 | 504 
suspicious left Babinski sign (+) | 504 | 504 
right Babinski sign (−) | 504 | 504 
diagnosed with intracranial infection | 504 | 504 
lumbar puncture | 504 | 504 
cerebrospinal fluid (CSF) sent for biochemistry analysis and microbial metagenomic next-generation sequencing (mNGS) | 504 | 504 
biochemistry analysis | 504 | 504 
glucose <1.1 mmol/L ↓ | 504 | 504 
chlorine 108 mmol/L ↓ | 504 | 504 
CSF protein >3,000 mg/L ↑ | 504 | 504 
microbial mNGS results | 504 | 504 
high sequence of Klebsiella pneumoniae with drug-resistant gene SHV-type beta-lactamases (blaSHV) | 504 | 504 
treated with 2 g meropenem q8h prolonged for 3 hours | 504 | 744 
body temperature improved | 744 | 744 
blood routine improved | 744 | 744 
CRP improved | 744 | 744 
CT examination | 744 | 744 
pulmonary edema and pleural effusion dissipated and absorbed | 744 | 744 
CSF analyses | 744 | 744 
chlorine 119 mmol/L ↓ | 744 | 744 
micro amount of proteins 1,107 mg/L ↑ | 744 | 744 
microalbumin 816.3 mg/L ↑ | 744 | 744 
immunoglobulin G 308.5 mg/L ↑ | 744 | 744 
α2-macroglobulin 18.5 mg/L ↑ | 744 | 744 
β2-microglobulin 2.67 mg/L ↑ | 744 | 744 
discharged from the hospital | 744 | 744 
close follow-up | 744 | 744