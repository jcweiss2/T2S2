55 years old | 0
female | 0
admitted to the emergency department | 0
abdominal pain | -240
diabetes mellitus | -21600
coronary bypass operation | -87600
left infrapatellar amputation | -35040
chronic renal failure | -17520
hemodialysis treatment | -8760
no history of abdominal trauma | 0
white blood cell: 15,100/mm³ | 0
hemoglobin: 8.5 g/dL | 0
C-reactive protein: 40 mg/dL | 0
urea: 37.9 mg/dL |&lt;no_output&gt;
