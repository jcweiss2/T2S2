56 years old | 0
female | 0
Hispanic | 0
admitted to the clinic | 0
blurred vision | 0
floaters in both eyes | 0
septic shock | -744
bilateral pneumonia | -744
leptospirosis | -744
hospitalized | -744
elevated bilirubin | -744
elevated liver enzymes | -744
anemia | -744
severe thrombocytopenia | -744
platelet count of 37,000 | -744
treated with blood transfusions | -744
treated with intravenous ceftriaxone | -744
retinal hemorrhages | -744
visual loss | -744
visual acuity 20/200 OD | 0
visual acuity 20/30 OS | 0
intraocular pressure 14 OU | 0
anterior segment quiet | 0
2+ nuclear sclerosis | 0
sub-internal limiting membrane hemorrhage | 0
dot hemorrhages in the superior retina | 0
posterior vitreous detachment | 0
optical coherence tomography | 0
fluorescein angiography | 0
no improvement in visual acuity | 168
minimal hemorrhage resolution | 168
pars-plana vitrectomy | 672
internal limiting membrane removal | 672
blood aspiration | 672
best corrected visual acuity 20/60 OD | 744
dot hemorrhages resolved | 744
follow-up 8 months post vitrectomy | 2304
best corrected visual acuity 20/60 OD | 2304