30 years old | 0
Caucasian | 0
female | 0
gravida 2 | 0
para 1 | 0
admitted to the hospital | 0
preterm labor | 0
onset of preterm labor | 0
no significant past medical history | 0
postpartum depression | -672
denies recent international travel | 0
last travel 2 months prior to delivery | -336
denies any illnesses in the 3 months prior to delivery | 0
no sick contacts in the last month prior to delivery | 0
no known positive COVID-19 contacts | 0
denies any recent fever | 0
denies respiratory symptoms | 0
denies fatigue | 0
denies myalgia | 0
denies anosmia | 0
denies cough | 0
received adequate prenatal care | 0
no maternal or fetal concerns during pregnancy | 0
prenatal tests unremarkable | 0
group B Streptococcus status unknown | 0
SARS-CoV-2 testing not done | 0
precipitous vaginal delivery | 0
spontaneous rupture of membranes | 0
no respiratory symptoms before delivery | 0
no respiratory symptoms during delivery | 0
no respiratory symptoms after delivery | 0
no concerns for chorioamnionitis | 0
placental pathology assessment not done | 0
newborn vigorous at birth | 0
1-minute Apgar score 8 | 0
5-minute Apgar score 9 | 0
skin-to-skin care with mother | 0
mild respiratory distress | 0
grunting | 0
taken to radiant warmer | 0
transferred to newborn nursery | 0
noninvasive respiratory support | 0
Vapotherm at 4 liters per minute | 0
capillary blood gas unremarkable | 0
chest X-ray with hazy lung fields | 0
no clear infiltrates or effusions | 0
complete blood count with differential normal | 0
transferred to level III NICU | 5
worsening hypercarbia | 5
respiratory support escalated | 5
continuous positive airway pressure | 5
noninvasive positive pressure ventilation | 5
21% FiO2 | 5
SARS-CoV-2 testing by RT-PCR | 24
nasal pharyngeal swab | 24
test result positive | 48
repeat testing for SARS-CoV-2 | 96
repeat test result positive | 144
parents afebrile and asymptomatic | 0
parents allowed at bedside | 0
breastfeeding not done | 0
expressed breast milk | 0
parental visitation restricted | 48
parents tested for SARS-CoV-2 | 48
parents tested negative | 48
parents tested negative again | 120
respiratory support weaned off | 24
treated with empiric antibiotics | 24
ampicillin and gentamicin | 24
antibiotics discontinued | 72
feedings provided via gavage support | 24
discharged home | 216
indirect hyperbilirubinemia | 24
phototherapy | 24
newborn screen for congenital adrenal hyperplasia | 24
congenital adrenal hyperplasia ruled out | 216
NICU transport team notified | 48
no known COVID-19 cases among caretakers | 48
NICU transport team members tested for SARS-CoV-2 antibodies | 168
NICU transport team members tested negative | 168