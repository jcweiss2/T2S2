Here is the table of events and timestamps:

15 years old | 0
female | 0
acute myelogenous leukemia (AML) | 0
received standard induction treatment | 0
pancytopenia | -168
developed tachycardia | -168
developed hypotension | -168
developed lactic acidosis | -168
admitted to the pediatric intensive care unit | -168
transthoracic echocardiography | -168
severely impaired left ventricular ejection fraction | -168
sinus tachycardia with incomplete right bundle branch block | -168
N-terminal prohormone of brain natriuretic peptide (NT-proBNP) | -168
high-sensitive troponin T | -168
fluid therapy | -168
noradrenaline | -168
dobutamine | -168
milrinone | -168
deep sedation | -168
mechanical ventilation | -168
lactate acidosis worsened | -168
hypotonic | -168
heart rate of 160/min | -168
va-ECMO was initiated | -168
cannulation of the left femoral artery and vein | -168
13 Fr/15 cm arterial and 21 Fr/55 cm venous HLS Cannula | -168
Seldinger technique under sonographic guidance | -168
9 Fr sheath | -168
left superficial femoral artery | -168
Cardiohelp System with a 7.0 HLS Set Advanced Bioline Coating | -168
blood flow of 3.3 l/min at 3800 rpm | -168
extracorporeal blood flow (ECBF) | -168
mean arterial pressure (MAP) | -168
noradrenaline (80 µg/min) | -168
vasopressin (2 units/h) | -168
levosimendan (0.5 mg/h) | -168
hydrocortisone (200 mg/d) | -168
Continuous venovenous hemodiafiltration (CVVHDF) | -168
anti-infective therapy | -168
dose-adjustment of meropenem | -168
ciprofloxacin | -168
metronidazole | -168
cotrimoxazole | -168
liposomal amphotericin B | -168
acyclovir | -168
linezolid was replaced by vancomycin | -168
Procalcitonin (PCT) | -168
C-reactive protein (CRP) | -168
MAP declined to 40 torr | -24
increasing doses of vasopressors | -24
LVEF further decreased below 10% | -24
levosimendan infusion was stopped | -24
acute ischemic injury of the non-cannulated leg | -24
right femoral artery was dissected | -24
insufficient blood inflow due to low cardiac output | -24
lactate levels rose to 25 mmol/l | -24
Dacron conduit was sewed on the right femoral artery | -24
second arterial cannula (13 Fr/15 cm) | -24
Y-connector | -24
ECBF could be enhanced to 4–5 l/min | -24
MAP could be maintained at 40–50 torr | -24
venous drainage pressures could be reduced | -24
sufficient preload within the right atrium and vena cava | -24
echocardiography | -24
inspiratory oxygen fraction of the respirator was increased | -24
arterial oxygen partial pressure in blood drawn from the right radial artery was normal | -24
PCT levels rose to 42.5 ng/ml | -24
Hickman catheter was explanted | -24
broad-complex tachycardia | -24
esmolol and metoprolol | -24
left ventricular function further decreased | -24
aortic valve ceased to open | -24
pulmonary edema | -24
intracardiac clot formation | -24
second venous cannula (21 Fr/55 cm) | -24
percutaneous atrioseptostomy | -24
left atrium | -24
ECBF now reached 5–6 l/min | -24
lactate levels peaked at 29 mmol/l | -24
MAP rose from a nadir of 30 torr | -24
cerebral oximetry by near infrared spectroscopy | -24
sufficient regional oxygen saturation | -24
therapeutic anticoagulation | -24
unfractionated heparin | -24
target partial thrombin time of 60–80 s | -24
PCT peaked with 80.4 ng/ml | -24
CRP peaked with 7.23 mg/dl | -24
leukocytes remained low | -24
high-sensitive troponin T increased | -24
creatine kinase MB increased | -24
all microbial specimens collected remained negative | -24
viral myocarditis was excluded | -24
myocardial biopsy | -24
cardiac systolic function gradually recovered | -24
ECMO cannulas in the left femoral vessels were removed | -72
ECMO was completely removed | -72
LVEF had recovered to approximately 30% | -72
mean arterial pressures of 60–70 torr | -72
CVVHDF could be stopped | -72
renal function was normal | -72
leucocyte count recovered to 1000/µl | -72
normal values were reached spontaneously | -72
respirator weaning was reached | -72
successful allogenic stem cell transplantation | -72
allogenic stem cell transplantation | -72
severe critical illness | -72
polyneuropathy | -72
LVEF recovered to approximately 40% | -72