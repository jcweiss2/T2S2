25 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
autoimmune hepatitis | -672 | 0 | Factual
acetaminophen | -672 | 0 | Factual
ibuprofen | -672 | 0 | Factual
azathioprine | -672 | -168 | Factual
prednisone | -672 | -168 | Factual
unprotected sexual intercourse | -336 | -336 | Factual
influenza vaccination | -672 | -672 | Factual
COVID-19 vaccination | -672 | -672 | Factual
admitted to the hospital | 0 | 0 | Factual
bilateral lower extremity pain | -72 | 0 | Factual
edema | -72 | 0 | Factual
ascites | -72 | 0 | Factual
fever | -72 | 0 | Factual
chills | -72 | 0 | Factual
nausea | -72 | 0 | Factual
dizziness | -72 | 0 | Factual
heavy menorrhagia | -72 | 0 | Factual
hemodynamically unstable | 0 | 0 | Factual
blood pressure 67/39 mmHg | 0 | 0 | Factual
heart rate 129 beats per minute | 0 | 0 | Factual
respirations 33 per minute | 0 | 0 | Factual
temperature 35.1 degrees Celsius | 0 | 0 | Factual
jaundice | 0 | 0 | Factual
scleral icterus | 0 | 0 | Factual
abdominal ascites with fluid wave | 0 | 0 | Factual
anasarca | 0 | 0 | Factual
erythematous vaginal vault | 0 | 0 | Factual
minimal discharge | 0 | 0 | Factual
no vesicles | 0 | 0 | Factual
no lesions | 0 | 0 | Factual
no retained foreign objects | 0 | 0 | Factual
fine reticular violaceous patches | 0 | 16 | Factual
lactic acidosis | 0 | 0 | Factual
lactic acid 13.1 mmol/L | 0 | 0 | Factual
creatinine 1.49 mg/dL | 0 | 0 | Factual
aspartate transaminase 56 units/L | 0 | 0 | Factual
alanine transaminase 62 units/L | 0 | 0 | Factual
total bilirubin 3.7 mg/dL | 0 | 0 | Factual
direct bilirubin 3.19 mg/dL | 0 | 0 | Factual
alkaline phosphatase 213 units/L | 0 | 0 | Factual
total protein 5.3 g/dL | 0 | 0 | Factual
albumin 1.4 g/dL | 0 | 0 | Factual
hemoglobin 5.2 g/dL | 0 | 0 | Factual
leukocytes 1.3 k/uL | 0 | 0 | Factual
platelets 90 k/uL | 0 | 0 | Factual
prothrombin time 37.9 s | 0 | 0 | Factual
international normalized ratio 3.9 | 0 | 0 | Factual
beta-human chorionic gonadotropin test negative | 0 | 0 | Factual
occasional schistocytes | 0 | 0 | Factual
peritoneal fluid analysis | 0 | 0 | Factual
leukocyte count 9821 | 0 | 0 | Factual
neutrophilic predominance | 0 | 0 | Factual
CT angiography | 0 | 0 | Factual
cirrhosis with portal hypertension | 0 | 0 | Factual
large volume abdominal ascites | 0 | 0 | Factual
splenomegaly | 0 | 0 | Factual
generalized edematous wall thickening of the colon and rectum | 0 | 0 | Factual
intubation | 0 | 0 | Factual
intravenous fluids | 0 | 48 | Factual
blood products | 0 | 48 | Factual
vasopressors | 0 | 48 | Factual
broad-spectrum antibiotic therapy | 0 | 48 | Factual
vancomycin | 0 | 48 | Factual
piperacillin-tazobactam | 0 | 48 | Factual
doxycycline | 0 | 48 | Factual
clindamycin | 0 | 48 | Factual
intravenous immunoglobulin | 0 | 0 | Factual
large violaceous non-blanching ecchymoses | 16 | 16 | Factual
flaccid bullae | 16 | 16 | Factual
dusky and violaceous skin | 36 | 36 | Factual
bullae | 36 | 36 | Factual
lactate dehydrogenase 298 units/L | 16 | 16 | Factual
fibrinogen 187 mg/dL | 16 | 16 | Factual
D-dimer > 20 mcg/mL | 16 | 16 | Factual
urinalysis without signs of infection | 16 | 16 | Factual
salicylate level negative | 16 | 16 | Factual
acetaminophen level negative | 16 | 16 | Factual
Chlamydia trachomatis and Neisseria gonorrhea nucleic acid amplification tests negative | 16 | 16 | Factual
urine toxicology screen negative | 16 | 16 | Factual
peritoneal fluid culture negative | 16 | 16 | Factual
blood culture positive for Streptococcus pneumoniae | 16 | 16 | Factual
progressive hypoxia | 16 | 48 | Factual
shock | 16 | 48 | Factual
death | 48 | 48 | Factual
autopsy | 48 | 48 | Factual
cirrhotic liver | 48 | 48 | Factual
diffuse alveolar damage | 48 | 48 | Factual
serous fluid in the abdominal compartment | 48 | 48 | Factual