101 years old|0
    male|0
    admitted with pulmonary oedema|0
    mechanical ventilation|0
    weaning from mechanical ventilation unsuccessful|0
    tracheostomy performed|0
    gram-negative bacteraemia|0
    sepsis|0
    haemodynamic instability|0
    oliguric|168
    acidemic|168
    creatinine rise from 177 micromole/L to 335 micromole/L|168
    abdominal aortic aneurysm|0
    ischaemic heart disease|0
    tricuspid regurgitation|0
    pulmonary hypertension|0
    congestive heart failure|0
    pacemaker insertion|0
    chronic kidney disease|0
    diabetes|0
    cardiorenal syndrome|0
    preserved intellectual capacity|0
    active rabbi and teacher|0
    extremely frail|0
    unable to speak due to tracheostomy tube|0
    respiratory instability precluding speech valve use|0
    decreased level of consciousness|168
    uraemic encephalopathy|168
    haemodialysis initiated|168
    cuffed tunneled catheter placed in right internal jugular vein|168
    dialysis initiated ∼1 month before 102nd birthday|168
    56 haemodialysis treatments over ∼4 months|168
    death|672
    worsening heart failure|672
    recurrent sepsis|672
    pulmonary oedema|0
    chronic kidney disease|0
    acute kidney injury|0
    gram-negative bacteraemia|0
    sepsis|0
    haemodynamic instability|0
    oliguric|168
    acidemic|168
    creatinine rise|168
    preserved intellectual capacity|0
    active rabbi and teacher|0
    extremely frail|0
    unable to speak|0
    respiratory instability|0
    decreased consciousness|168
    uraemic encephalopathy|168
    haemodialysis initiated|168
    catheter placement|168
    dialysis initiation|168
    haemodialysis treatments|168
    death|672
    worsening heart failure|672
    recurrent sepsis|672<|eot_id|>
    
    101 years old|0
    male|0
    admitted with pulmonary oedema|0
    mechanical ventilation|0
    weaning from mechanical ventilation unsuccessful|0
    tracheostomy performed|0
    gram-negative bacteraemia|0
    sepsis|0
    haemodynamic instability|0
    oliguric|168
    acidemic|168
    creatinine rise from 177 micromole/L to 335 micromole/L|168
    abdominal aortic aneurysm|0
    ischaemic heart disease|0
    tricuspid regurgitation|0
    pulmonary hypertension|0
    congestive heart failure|0
    pacemaker insertion|0
    chronic kidney disease|0
    diabetes|0
    cardiorenal syndrome|0
    preserved intellectual capacity|0
    active rabbi and teacher|0
    extremely frail|0
    unable to speak due to tracheostomy tube|0
    respiratory instability precluding speech valve use|0
    decreased level of consciousness|168
    uraemic encephalopathy|168
    haemodialysis initiated|168
    cuffed tunneled catheter placed in right internal jugular vein|168
    dialysis initiated ∼1 month before 102nd birthday|168
    56 haemodialysis treatments over ∼4 months|168
    death|672
    worsening heart failure|672
    recurrent sepsis|672
    pulmonary oedema|0
    chronic kidney disease|0
    acute kidney injury|0
    gram-negative bacteraemia|0
    sepsis|0
    haemodynamic instability|0
    oliguric|168
    acidemic|168
    creatinine rise|168
    preserved intellectual capacity|0
    active rabbi and teacher|0
    extremely frail|0
    unable to speak|0
    respiratory instability|0
    decreased consciousness|168
    uraemic encephalopathy|168
    haemodialysis initiated|168
    catheter placement|168
    dialysis initiation|168
    haemodialysis treatments|168
    death|672
    worsening heart failure|672
    recurrent sepsis|672