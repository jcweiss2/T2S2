57 years old | 0
male | 0
lepromatous leprosy | -336
treatment with rifampicin/clofazimine/dapsone | -336
admitted to the hospital | 0
abdominal distension | 0
constipation | 0
vomiting | 0
10-kg weight loss | 0
peripheral lymphadenopathy | 0
distended abdomen | 0
positive shifting dullness | 0
mural thickening of the terminal ileum | 0
enlarged mesenteric lymph nodes | 0
mesenteric fat stranding | 0
intra-abdominal free fluid | 0
abdominal granulomatous infection | 0
neoplastic process | 0
abdominal paracentesis | 24
atypically large lymphocytes | 24
high-grade lymphoma | 24
flow cytometry | 24
abnormal CD4/CD8 double-negative T-cell population | 24
cervical lymph node biopsy | 48
high-grade peripheral T-cell lymphoma | 48
bone marrow examination | 48
no involvement of T-cell NHL | 48
stage IV lymphoma | 48
dexamethasone | 48
tumor-lysis syndrome precautions | 48
severe sepsis | 72
transfer to the medical intensive care unit | 72
antibiotics | 72
antifungals | 72
ICU care | 168
recovered | 168
transferred to the national cancer center | 168
EPOCH chemotherapy protocol | 168
CNS prophylaxis | 168
intrathecal methotrexate | 168
complete metabolic remission | 336
positron emission tomography/computed tomography | 336
febrile neutropenia episodes | 336
recurrent bacteremia | 336
generalized weakness | 336
no sensory changes | 336
no clear fatigability | 336
decreased power in all proximal and distal muscles | 336
critical illness myopathy-neuropathy | 336
toxic neuropathy | 336
paraneoplastic syndrome | 336
electromyogram/nerve conduction study | 336
normal distal latencies | 336
normal compound muscle action potential | 336
normal conduction velocities | 336
normal F waves | 336
normal sensory nerve studies | 336
needle electromyogram | 336
normal insertional activity | 336
no spontaneous activity | 336
normal motor unit action potential | 336
poor recruitment effects | 336
repetitive nerve stimulation | 336
significant incremental response | 336
presynaptic neuromuscular junction disorder | 336
Lambert-Eaton myasthenic syndrome | 336
intravenous immunoglobulins | 336
significant improvement of motor function | 360
ambulate | 360
consolidation by autologous bone marrow transplant | 360
recurrent bacteremia | 360
sepsis | 360
multiorgan failure | 360
re-admitted to the medical ICU | 360
passed away | 432