52 years old | 0
male | 0
Caucasian | 0
admitted to the hospital | 0
jaundice | -96
darkening of urine color | -96
fatigue | -96
dyspnea | -96
tachycardia | 0
heart rate up to 150 beats per minute | 0
normal blood pressure | 0
respiratory rate of 50 breaths per minute | 0
oxygen saturation as low as 80% | 0
15 L of O2 support from a non-rebreather mask | 0
admitted to the medical intensive care unit (ICU) | 0
computed tomography (CT) of the chest | -96
tested for COVID-19 with a polymerase chain reaction (PCR) | -96
PCR test came back negative | 0
chest CT was consistent with COVID-19 pneumonia | 0
toxoplasma serology | 0
rubella serology | 0
HSV serology | 0
EBV serology | 0
CMV serology | 0
HIV serology | 0
hantavirus serology | 0
Leptospira serology | 0
ANA | 0
ANCA | 0
anti-dsDNA | 0
haptoglobin | 0
IGG | 0
IGM | 0
IGA | 0
IGE | 0
direct coombs | 0
indirect coombs | 0
complements C3 | 0
complements C4 | 0
peripheral blood smear demonstrated no schistocytes | 0
abdominal ultrasonography revealed a mild hepatomegaly | 0
high-flow nasal cannula | 0
empirical treatment with meropenem | 0
empirical treatment with doxycycline | 0
femoral central venous catheter was inserted | 0
plasmapheresis was initiated | 0
60 units of fresh frozen plasma was used during five sessions of plasmapheresis | 0
total bilirubin level had dropped down to 19.6 mg/dL | 24
Leptospira test using real-time PCR came back positive | 96
medical treatment was continued with both meropenem and doxycycline | 96
patient showed significant clinical improvement | 96
weaned off of oxygen | 192
laboratory values and chest X-ray greatly improved | 192
transferred to the infectious diseases ward | 192
discharged from the hospital | 192
uneventful recovery | 192
no further complications | 192
catastrophic floods in the west of the Black Sea region of Turkey | -336
patient’s initial symptoms | -96
incubation period of leptospirosis | -168
plasmapheresis played a vital role in the patient’s rapid recovery | 192