60 years old | 0
hypertensive | 0
diabetic | 0
Asian | 0
male | 0
admitted | 0
recent onset fever (38.6 °C) | 0
persistent productive cough | 0
chest pain |, 0
myalgias | 0
fatigue | 0
respiratory distress | 0
past history of TB | 0
unprotected contact with cousin | -672
cousin recently recovered from COVID-19 | -672
decreased breath sounds at lung bases | 0
saturation of peripheral oxygen (SpO2) 72% | 0
no respiratory distress | 0
portable chest X-ray bilateral interstitial infiltrates | 0
electrocardiogram normal | 0
cardiac enzymes normal | 0
coagulation profile normal | 0
echocardiography normal | 0
lymphocytopenia (0.59 × 10⁹/L) | 0
increased C-reactive protein (243.3 mg/liter) | 0
increased lactate dehydrogenase (944 units/liter) | 0
increased ferritin (876 ng/ml) | 0
admission chest CT diffuse bilateral ground-glass opacities | 0
nasopharyngeal swabs confirmed COVID-19 | 0
admitted to isolation chamber | 0
full diagnostic work-up | 0
higher level of respiratory support via HFNC | 0
awake prone positioning (16–20 hours daily) | 0
ROX maintained over 6 for 48 hours | 0
empiric therapy with lopinavir/ritonavir | 0
empiric therapy with ribavirin | 0
dexamethasone | 0
prophylactic anticoagulation | 0
NAAT on sputum specimens revealed Mycobacterium tuberculosis | 0
started on isoniazid | 0
started on pyridoxal phosphate | 0
started on rifampicin | 0
started on pyrazinamide | 0
started on ethambutol | 0
no side effects | 0
ratio of partial arterial pressure of oxygen to fractional inspired concentration of oxygen >250 | 168
HFNC discontinued | 288
awake prone positioning discontinued | 288
oxygen therapy (2–4 L) administered | 288
oxygen supportive care discontinued | 384
RT-PCR test negative | 480
microbiology negative | 480
discharged to home isolation | 648
followed-up by outreach team | 648
increased inflammation biomarkers | 0
lymphocytopenia | 0
extensive lung parenchymal disease | 0
poor prognosis | 0
drug-susceptible TB | 0
standard first-line regimen | 0
combination of anti-TB therapy and antiviral treatment | 0
risk for side-effects | 0
no side-effects recorded | 0
uneventful recovery | 648
application of HFNC effective | 0
application of awake prone positioning effective | 0
increased C-reactive protein | 0
increased lactate dehydrogenase | 0
increased ferritin | 0
lymphocytopenia upon admission | 0
laboratory abnormalities | 0
correlation with TB uncertain | 0
