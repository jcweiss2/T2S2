34 years old | 0
male | 0
admitted to the hospital | 0
alcohol dependence | 0
1-day history of left-sided, cramping abdominal pain | -24
abdominal pain radiating to the back | -24
denied prior episodes | -24
denied any inciting incidents | -24
denied known history of diabetes mellitus | -24
denied medication use | -24
denied pancreatitis | -24
denied family history of genetic dyslipidemias | -24
not obese (BMI 24.4) | 0
no acute distress | 0
tachycardia (112/min) | 0
moderate tenderness to palpation in the right upper quadrant | 0
moderate tenderness to palpation in the left upper quadrant | 0
moderate tenderness to palpation in the left lower quadrant | 0
leukocytes 12 k/µL | 0
neutrophils 81.8% | 0
potassium 3.2 mEq/L | 0
random glucose 136 mg/dL | 0
calcium 6.8 mg/dL | 0
alanine aminotransferase 73 U/L | 0
aspartate aminotransferase 80 U/L | 0
alkaline phosphatase 135 IU/L | 0
TGs 9708 mg/dL | 0
low-density lipoprotein 373 mg/dL | 0
lipase 245 U/L | 0
computed tomography revealing acute interstitial pancreatitis | 0
peripancreatic fluid surrounding the pancreatic tail | 0
fatty infiltration of the terminal ileum submucosa | 0
concern for inflammatory bowel disease | 0
admitted to the medical ICU | 0
nil per os | 0
insulin drip | 0
dextrose 10% in water drip | 0
high-volume intravenous fluids | 0
electrolyte replenishment | 0
analgesia | 0
serum TG level 4025 mg/dL | 0
plasmapheresis initiated | 0
fresh frozen plasma replacement (1250 cm3) | 0
5% albumin replacement (1250 cm3) | 0
TG level 603 mg/dL after one cycle | 0
continued insulin drip | 0
continued treatments | 0
TG level 304 mg/dL after 1 day | 24
transferred to the medical floors | 24
HTGP diagnosed | 0
initial conservative management | 0
aggressive intravenous hydration | 0
bowel rest | 0
insulin therapy | 0
heparin therapy | 0
plasmapheresis with albumin replacement | 0
reduced TG levels by 58.5% over 2 days | 48
further reduction of TGs by 85% after plasmapheresis | 48
ICU stay of 2 days | 48
hospital stay duration | 48
rapid alleviation of symptoms | 48
reduction of lab abnormalities | 48
discharge in stable condition | 48
written informed consent obtained | 0
