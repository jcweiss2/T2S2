45 years old | 0
male | 0
admitted to the hospital | 0
shortness of breath | 0
confusion | 0
severe asthenia | 0
arterial blood pressure 75/50 mmHg | 0
heart rate 120 beats per minute | 0
peripheral oxygen saturation 85% | 0
diffuse bilateral reduction in vesicular breath sounds | 0
tachypnoea | 0
axillary temperature 37.8°C | 0
sinus tachycardia | 0
diffuse repolarization abnormalities | 0
low peripheral voltages | 0
mild leukocytosis | 0
thrombocytopenia | 0
high sensitive troponin T increased | 0
NT-proBNP increased | 0
C-reactive protein increased | 0
fever | -72
mild dyspnoea | -72
fatigue | -72
nasopharyngeal swab for SARS-CoV-2 negative | -24
computed tomography of the thorax showed mild ground-glass opacities | -24
cardio-septic shock | 0
pyretic | 0
hypoxic | 0
severe biventricular impairment | 0
metabolic acidosis | 0
non-invasive mechanical ventilation | 0
inotropic support with noradrenaline | 0
inotropic support with adrenaline | 0
empiric antibiotic therapy | 0
intra-aortic balloon pump | 4
worsening hypotension | 4
persistent metabolic acidosis | 4
bronchoscopy | 24
bronchoalveolar lavage tested positive for SARS-CoV-2 | 24
clinical stabilization | 120
IABP removed | 120
complete weaning from inotropic support | 120
transferred to the Cardiology department | 144
cardiac magnetic resonance imaging | 144
severe biventricular dysfunction | 144
augmented T1 mapping | 144
signs of acute myocarditis | 144
myocardial biopsy | 168
mild lymphohistiocytic infiltrate | 168
diffuse platelet clots | 168
Parvovirus B-19 DNA detected | 168
SARS-CoV-2 RNA not detected | 168
levosimendan administered | 168
Anakinra started | 168
echocardiography showed significant improvement | 168
discharged | 216
optimal medical therapy for heart failure | 216
IL-1 inhibitor | 216
follow-up | 744
good clinical conditions | 744
mild effort dyspnoea | 744
stable improvement of biventricular function | 744
normalization of T1 mapping | 744
follow-up | 1296
good clinical conditions | 1296
no more dyspnoea | 1296
complete recovery of biventricular function | 1296