54 years old | 0
male | 0
alcoholic cirrhosis | 0
diabetes mellitus | 0
admitted to the hospital | 0
altered sensorium | -48
fever | -48
no prior history of headache | 0
no prior history of vomiting | 0
no prior history of seizures | 0
no prior history of decreasing urine output | 0
febrile | 0
disoriented | 0
pulse rate was 100/min | 0
blood pressure was 150/70 mmHg | 0
mild icterus | 0
pedal edema | 0
no evidence of focal neurological deficit | 0
no signs of meningism | 0
no features of papilledema or retinitis | 0
bilateral pupils were equal and reacting to light | 0
free fluid | 0
no organomegaly | 0
Hb 9.6 gm/dL | 0
total leukocyte count (TLC) 16 800/ mm3 | 0
normal eosinophil counts | 0
platelet count 1.1lac/mm3 | 0
normal coagulation profile | 0
INR of 1.3 | 0
serum bilirubin was 3.0 mg/dL | 0
AST/ALT of 87/96 IU/L | 0
arterial ammonia was 239 μg/dL | 0
IgM anti-HEV positive | 0
HBsAg negative | 0
anti-HCV negative | 0
IgM anti-HAV negative | 0
HIV negative | 0
high ascites | 0
high serum-ascites albumin gradient | 0
normal cell counts | 0
chronic liver disease | 0
coarse echotexture | 0
normal bilateral kidneys | 0
1+ proteinuria | 0
full field leucocytes | 0
8-10 RBC/high-power field | 0
urine culture positive for enterococcus faecalis | 0
sensitive to linezolid | 0
hepatic encephalopathy | 0
uro-sepsis | 0
lactulose | 0
supportive care for liver failure | 0
linezolid 600 mg twice a day | 0
pruritus | 72
erythematous macular rash | 72
eosinophilia | 72
absolute eosinophil count of 2125 cells/mm3 | 72
elevated serum IgE levels | 72
2+ proteinuria | 72
15-20 leukocytes | 72
WBC casts | 72
RBC cast | 72
no evidence of eosinophils | 72
renal functions deranged | 72
serum creatinine rising to 5.2 mg/dL | 72
decreasing urine output | 72
dialytic support | 72
DRESS syndrome | 72
linezolid stopped | 72
rash subsided | 120
fever subsided | 120
renal functions remained deranged | 120
recovered from hepatic encephalopathy | 120
liver functions improved | 120
ANA negative | 120
ANCA negative | 120
normal complement levels | 120
renal biopsy | 168
normal glomeruli | 168
interstitium showed edema | 168
moderate inflammatory infiltrate | 168
mononuclear cells | 168
few eosinophil | 168
proximal tubular dilatation | 168
patchy necrosis | 168
birefringent oxalate crystals | 168
foreign body giant cell reaction | 168
no granuloma formation | 168
no immune complex deposition | 168
acute tubulointerstitial nephritis | 168
patchy tubular necrosis | 168
prednisolone | 168
renal functions improved | 240
serum creatinine level decreasing to 1.4 mg/dL | 240
estimated creatinine clearance of 56 mL/min | 240
follow-up | 720