6 years old | 0
female | 0
admitted to the emergency department | 0
severe headache | -48
nausea | -48
vomiting | -48
mumps infection | -240
spontaneous resolution of mumps infection | -240
altered consciousness level | 0
mildly confused | 0
Glasgow Coma Scale = E4 V4 M6 | 0
trunk and gait ataxia | 0
bilateral dysmetria on finger-nose tests | 0
body temperature 37.5 °C | 0
normal heart rate | 0
normal breath rate | 0
dysautonomic troubles | 2
heart rate decreased to 55 beats/min | 2
arterial pressure dropped to 80/50 mmHg | 2
transferred to the Pediatric Intensive Care Unit | 2
brain computed tomography scan | 2
cerebellar ill-defined hypodense lesion | 2
mass effect on the fourth ventricle | 2
dilation of the upper ventricular system | 2
multimodal magnetic resonance imaging | 4
cerebellar high-intensity areas on T2-weighted and FLAIR images | 4
diffuse edema | 4
mass effect on the fourth ventricle and brainstem | 4
tonsillar herniation | 4
supratentorial hydrocephalus | 4
Gadolinium-enhanced T1-weighted sequence | 4
leptomeningeal enhancement along the cerebellar folia | 4
mildly reduced level of N acetyl aspartate (NAA)/Creatine | 4
normal Choline/Creatine ratios | 4
doublet of lactate-lipid peak | 4
hemoglobin concentration of 12.7 g/dL | 4
white blood cell count of 14280/mm3 | 4
platelet count | 4
erythrocyte sedimentation rate showed moderate increase | 4
C-reactive protein level above 2 mg/L | 4
serological test for mumps virus positive with IgM and IgG | 4
post-infectious acute hemicerebellitis diagnosed | 4
treated with mannitol and corticosteroid | 4
IV methylprednisolone 30 mg/kg per day | 4
oral prednisone 1 mg/kg per day | 4
tapered within 1 mo | 672
favorable evolution | 24
partial resolution of signal alterations in the cerebellar hemispheres | 432
complete resolution confirmed by brain MRI | 720
discharged | 24