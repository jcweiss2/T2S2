60 years old | 0
female | 0
admitted to the hospital | 0
back pain | -96
leg weakness | -96
loss of consciousness | 0
head injury | 0
preceding symptoms | 0
sharp back pain | -96
lower back pain | -96
falls | -96
sore throat | -96
earache | -96
chills | -96
mildly productive cough | -96
atrioventricular node dysfunction | -672
dual-chamber pacemaker placement | -672
hypercoagulable state | -672
pulmonary emboli | -672
type two diabetes mellitus | -672
hypertension | -672
ill appearance | 0
no acute distress | 0
blood pressure 102/51 mm Hg | 0
heart rate 72 beats per minute | 0
temperature 97.2 degrees Fahrenheit | 0
breathing 16 breaths per minute | 0
oxygen saturation 100% | 0
systolic murmur | 0
moderate right lumbar paraspinal tenderness | 0
poor dentition | 0
multiple dental caries | 0
lactic acid 2.9 mmol/L | 0
procalcitonin > 100 | 0
platelet count 57 | 0
creatinine 1.44 | 0
Gram-positive cocci in chains | 0
abscess in right psoas muscle | 0
mobile echodensity attached to the tricuspid valve | 0
mobile echodensity on the pacemaker lead | 0
infective endocarditis | 0
vancomycin | 0
cefepime | 0
cardiology consultation | 0
infectious diseases consultation | 0
Streptococcus agalactiae | 0
ceftriaxone | 0
pacemaker extraction | 24
temporary pacing wire placement | 24
hypotensive | 24
vasopressors | 24
Gram-negative, anaerobic rods | 24
meropenem | 24
Prevotella bivia | 24
ertapenem | 48
new pacemaker device placement | 168
clearance of P. bivia bacteremia | 168
right psoas muscle abscess evaluation | 168
discharged home | 336
home health | 336
6-week course of intravenous ertapenem | 336
follow-up | 504
no complications | 504
no adverse events | 504