76 years old | 0
female | 0
end-stage kidney disease | 0
lambda light chain multiple myeloma | 0
multiple myeloma diagnosis | -25920
fatigue | -25920
bone pain | -25920
weight loss (22 kg) | -25920
hemodialysis replacement | -25920
international staging system III | 0
durie salmon stage IIIB | 0
systemic arterial hypertension | 0
glucose intolerance | 0
fragile (myeloma frailty score: 3) | 0
hypercalcemia | 0
anemia | 0
renal impairment | 0
lytic lesions | 0
bortezomib | 0
dexamethasone | 0
admitted to emergency service | -216
confusion | -216
hip pain | -216
respiratory distress | -192
COVID-19 diagnosis (RT-PCR) | -192
plasmacytoma in left hip | -192
clinical support | 0
transfusion support | 0
pain control support | 0
ceftriaxone | 0
vancomycin | 0
discharged | 168
RT-PCR test | 384
RT-PCR SARS-COV-2 detected | 384
partial recovery of symptoms | 384
sporadic delirium | 384
radiotherapy referral | 432
radiotherapy 3000cGy | 432
daratumumab monotherapy | 432
daratumumab infusion delayed | 564
chills | 564
tremors | 564
hemodialysis | 564
recovered symptoms | 588
negative blood culture | 588
daratumumab infused | 588
dyspnea | 588
emergency room visit | 600
acute respiratory failure | 600
hypoxemia | 600
COVID-19 positive (RT-PCR) | 600
COVID-19 reinfection | 600
negative SARS-COV-2 IgG | 600
negative SARS-COV-2 IgM | 600
close family members infected | 600
shilley catheter-related bloodstream infection | 600
pseudomonas aeruginosa | 600
extended spectrum beta-lactamase | 600
meropenem | 600
vancomycin | 600
dexamethasone | 600
catheter exchanged | 600
clinical stability | 600
worse chest CT | 600
febrile event | 672
antibiotics escalated (polymixicin, linezolid) | 672
RT-PCR SARS-COV-2 undetectable | 720
hemodynamic instability | 768
refractory septic shock | 768
klebsiella pneumonia | 768
carbapenemase | 768
intensive care | 768
mechanical ventilation | 768
high-dose vasoactive drugs | 768
death | 816
