66 years old| 0
male| 0
presented to the hospital with a 1-month history of dyspnoea on exertion| -720
dyspnoea on exertion| -720
orthopnoea| -720
paroxysmal nocturnal dyspnoea| -720
4 kg unintentional weight loss| -720
blood pressure of 103/81 mmHg| 0
heart rate 90 b.p.m.| 0
respiratory rate 20 b.p.m.| 0
oxygen saturation of 98% on room air| 0
jugular venous pressure elevated at +4 cm| 0
bilateral peripheral oedema to the knees| 0
pansystolic murmur at the apex| 0
third heart sound| 0
bilateral crackles at the lung bases| 0
elevated N-terminal pro-brain natriuretic peptide| 0
normal troponin I| 0
sinus rhythm| 0
left axis deviation| 0
inferior Q-waves| 0
no ST changes| 0
dilated left and right ventricles| 0
LV internal diameter end diastole 64 mm| 0
LV internal diameter end systole 61 mm| 0
LV ejection fraction (LVEF) 17%| 0
moderate mitral regurgitation| 0
moderate tricuspid regurgitation| 0
pulmonary artery systolic pressure 34 mmHg| 0
estimated mean right atrial pressure 10–15 mmHg| 0
inferior vena cava (IVC) diameter 17 mm which collapses less than 50% on inspiration| 0
masses in both apices| 0
two further masses in the right atrium suspicious for type B thrombi| 0
intracardiac masses had high signal intensity on T1- and T2-weighted sequences| 0
low-signal on first pass imaging following gadolinium administration| 0
LV end-diastolic volume 385 mL| 0
RV end-diastolic volume 305 mL| 0
calculated LVEF 19%| 0
RV ejection fraction (RVEF) 20%| 0
small bilateral pleural effusions| 0
IVC diameter 29 mm| 0
delayed enhancement sequences showed near full thickness scars in the lateral and inferior walls| 0
occlusion of the left circumflex artery| 0
occlusion of the right coronary artery| 0
severe stenosis of the mid-left anterior descending artery| 0
suspected right heart thrombi| 0
elevated liver enzymes| 0
aspartate aminotransferase 106 U/L| 0
alanine aminotransferase 406 U/L| 0
gamma-glutamyl transferase 64 U/L| 0
hyperbilirubinemia 60 μmol/L| 0
prolonged prothrombin time 24 s| 0
prothrombin ratio 2.0| 0
activated partial thromboplastin time 43 s| 0
started on warfarin| 0
bridging enoxaparin| 0
lisinopril 10 mg daily| 0
frusemide 40 mg daily| 0
carvedilol 12.5 mg twice daily| 0
discharged | 432
repeat cardiac MRI showed complete resolution of intracardiac masses| 432
LVEF 22%| 432
RVEF 46%| 432
out of hospital cardiac arrest| 648
admitted to intensive care unit| 648
percutaneous coronary intervention to left anterior descending artery| 768
implantable cardioverter defibrillator inserted| 792
patient discharged home| 1032
