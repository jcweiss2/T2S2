24 years old | 0
female | 0
admitted to the hospital | 0
fever | 0
constitutional symptoms | 0
preterm labor | 0
leukocytosis | 0
elevated C-reactive protein | 0
vaginal hyperthermia | 0
warm amniotic fluid | 0
treatment for chorioamnionitis | 0
delivered vaginally | 0
preterm infant | 0
mild respiratory distress | 0
treatment with ampicillin and gentamycin | 0
normal laboratory examinations | 0
negative blood cultures | 0
completed 7 days of antibiotics | 168
discharged | 168
fever | 0
abdominal pain | 0
foul smelling lochia | 0
acute abdomen | 0
antimicrobial therapy | 0
computed tomographic scan of the abdomen | 0
peritonitis | 0
exploratory laparotomy | 192
hysterectomy | 192
left salpingectomy | 192
appendectomy | 192
febrile | 192
worsening respiratory distress | 192
bilateral alveolar infiltrates | 192
pleural effusion | 192
broad spectrum antibiotics | 192
transferred to the intensive care unit | 408
ventilator support | 408
histopathology | 408
chronic granulomatous inflammation | 408
necrotic changes | 408
acid-fast bacilli positive | 408
miliary TB | 408
treatment with a four-drug regimen for TB | 408
isoniazid | 408
rifampin | 408
pyrazinamide | 408
ethambutol | 408
bronchoalveolar lavage | 408
Mycobacterium tuberculosis isolated | 408
newborn infant readmitted | 456
good condition | 456
no fever | 456
no respiratory distress | 456
no hepatosplenomegaly | 456
adequate weight gain | 456
normal chest X-ray | 456
normal laboratory tests | 456
normal tuberculin test | 456
negative gastric aspirates | 456
apnea | 480
desaturations | 480
leukocytosis | 480
neutrophil predominance | 480
platelets | 480
CRP | 480
bilateral alveolar infiltrates | 480
antibiotics | 480
suspected nosocomial pneumonia | 480
cultures | 480
negative CSF | 480
normal CSF indices | 480
gastric aspirates | 480
AFB positive | 480
treatment for TB | 480
isoniazid | 480
rifampin | 480
pyrazinamide | 480
amikacin | 480
lumbar puncture | 480
normal CSF indexes | 480
negative AFB stain | 480
positive PCR for M. tuberculosis | 480
M. tuberculosis isolated | 480
magnetic resonance imaging of the brain | 480
normal | 480
susceptibility to isoniazid | 480
susceptibility to rifampin | 480
susceptibility to ethambutol | 480
susceptibility to streptomycin | 480
steady improvement | 504
resolution of fever | 504
resolution of oxygen requirements | 504
follow-up chest X-ray | 720
significant improvement | 720
follow-up gastric aspirates | 720
negative for AFB | 720
no mycobacteria isolated | 720
discharged home | 720
completed 12 months of anti-TB therapy | 8760
mild hepatotoxicity | 8760
clinical resolution of disease | 8760