62 years old | 0
male | 0
gastroesophageal reflux disease | 0
benign prostatic hyperplasia | 0
elevated prostate-specific antigen | 0
transrectal ultrasound–guided prostate biopsy | 0
septic shock | 0
admitted to the intensive care unit | 0
urosepsis | 0
extended spectrum beta lactamase Escherichia coli | 0
pyelonephritis | 0
continuous high-dose vasopressors | 0
phenylephrine | 0
vasopressin | 0
norepinephrine | 0
hypoxemic respiratory failure | 12
shock liver | 12
acute renal failure | 12
acalculous cholecystitis | 12
bilateral upper and lower extremities underwent distal pressor-induced ischemia | 12
gangrene | 12
topical nitroglycerin | 108
hyperbaric oxygen therapy | 288
bilateral amputations of all fingers | 216
tissue demarcation at the level of the metatarsal heads | 216
loss of all plantar skin on the left foot | 216
weight-bearing skin on the right foot | 216
partial loss of both calcanei | 216
multiple debridement | 216
intravenous antibiotics | 216
wound bed preparation | 216
bilayered bovine collagen | 216
porcine xenografts | 216
bilateral transmetatarsal amputations | 432
removal of both necrotic calcanei and soft tissues | 432
INTEGRATM Bilayer Matrix Wound Dressing | 432
skin grafts to the dorsum of his TMAs | 432
free flap planning | 1092
angiography | 1092
sensate anterolateral thigh flap to his left foot | 1092
end-to-side anastomosis to the inframalleolar posterior tibial artery | 1092
end-to-end venous anastomosis to the saphenous vein and deep vena comitantes | 1092
neurotization via the lateral femoral cutaneous nerve to the posterior tibial nerve | 1092
Integra | 1092
split-thickness skin graft from the left thigh | 1105
neurotized ALT flap to the right foot | 1105
end-to-side anastomosis to the inframalleolar posterior tibial artery | 1105
2-vein anastomosis and coaptation of the lateral circumflex femoral nerve to the posterior tibial nerve | 1105
non–weight-bearing for 6 weeks | 1105
ankle foot orthoses and custom braces | 1105
intensive physical therapy | 1105
protective sensation of bilateral heels | 1105
walking 2 months after free tissue transfer | 1512
retained sensation of both free flaps | 2184
functionally ambulatory with an ExoSymTM prosthesis | 2184