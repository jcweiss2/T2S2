48 years old | 0
male | 0
chronic renal failure | -96
ischemic stroke | -96
insulin-dependent diabetes | -96
fever | -96
malaise | -96
oliguria | -96
haematuria | -96
nausea | -96
vomiting | -96
febrile (38°C) | 0
normal blood pressure (110/80 mmHg) | 0
depressible abdomen | 0
painful prostate | 0
leukocytosis (12,900) | 0
renal failure (creatinine 399 μmol/l) | 0
high C-reactive protein (137 mg/l) | 0
urea (30 mg/l) | 0
hyperglycemia | 0
acidosis | 0
positive acetonuria | 0
male urinary tract infection suspected | 0
diabetic ketoacidosis suspected | 0
abdominopelvic CT scan | 0
emphysematous lesions in prostate | 0
emphysematous lesions in seminal vesicles | 0
normal kidneys | 0
no dilatation of excretory cavities | 0
cytobacteriological examination of urine | 0
blood culture | 0
empirical intravenous antibiotics (cefotaxime and ciprofloxacine) | 0
antibiotics changed to imipenem and ciprofloxacin | 24
Enterobacter cloacae isolated | 24
suprapubic catheterization | 24
apyretic | 72
aggravation of inflammatory syndrome | 72
white blood cells increased to 20,000 | 72
CRP increased to 200 mg/l | 72
severe metabolic acidosis | 72
emergency hemodialysis | 72
abdominopelvic control scan | 72
prostatic hydroaeric collections | 72
trans-rectal aspiration | 72
purulent liquid (50 ml) | 72
bacteriological examination same germ | 72
generalized convulsive seizures | 96
apyretic | 96
regression of inflammatory syndrome | 96
white blood cells 16,000 | 96
CRP 123 mg/l | 96
correct metabolic balance | 96
chronic renal failure | 96
head CT scan normal | 96
seizures attributed to antibiotics | 96
antibiotics changed to piperacillin and flagyl | 96
antibiotic adaptation | 168
worsening state of consciousness | 336
septic shock | 336
transfer to intensive care | 336
orotracheal intubation | 336
norepinephrine in high dose | 336
death | 336
multi-organ failure | 336
