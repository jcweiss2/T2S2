72 years old | 0
female | 0
admitted to the hospital | 0
general weakness | -336
poor oral intake | -336
bilateral knee joint pain | -672
osteoarthritis | -672
intra-articular steroid injections | -672
triamcinolone acetonide | -672
weight gain | -336
mild systemic edema | -336
cushing's syndrome | -336
fever | 0
acute ill appearance | 0
sleepy | 0
multiple ulcers | 0
whitish patches | 0
mild crackle sound | 0
hemoglobin level of 15.3 g/dL | 0
white blood cell count of 13×10^3/mL | 0
platelet count of 349×10^3/µL | 0
mild hyperglycemia | 0
random blood glucose level of 174 mg/dL | 0
Hb A1C level of 7.7% | 0
fasting plasma C-peptide level of 6.1 ng/mL | 0
serum albumin level of 2.4 g/dL | 0
C-reactive protein level of 13.37 mg/dL | 0
human immunodeficiency virus test negative | 0
sick euthyroid state | 0
basal cortisol level of 0.55 µg/dL | 0
30 minute cortisol level of 6.3µg/dL | 0
90 minute cortisol level of 5.5µg/dL | 0
adrenal insufficiency | 0
multiple cavitary nodules in both lungs | 0
mass and cavitary nodules with mild homogenous enhancement | 0
percutaneous needle biopsy | 72
aggregate of fungal hypae | 72
invasive aspergillosis | 120
amphotericin B | 120
unconscious | 144
brain magnetic resonance imaging | 144
cerebrospinal fluid tapping | 144
numerous thin peripheral enhancing cystic nodules | 144
brain involvement | 144
voriconazole | 192
ventilator care | 192
respiratory failure | 336
septic shock | 336
death | 336