60 years old | 0
female | 0
presented to the emergency department | 0
back pain | -96
leg weakness | -96
fall | -96
denied loss of consciousness | 0
denied head injury | 0
denied preceding symptoms | 0
persistent sharp back pain | 0
back pain radiating across lower back | 0
multiple similar falls | -96
weakness | -96
legs giving out | -96
recent sore throat | -96
recent earache | -96
recent chills | -96
recent mildly productive cough | -96
atrioventricular node dysfunction | 0
dual-chamber pacemaker placement | 0
hypercoagulable state | 0
prior pulmonary emboli | 0
type two diabetes mellitus | 0
hypertension | 0
ill appearance | 0
no acute distress | 0
blood pressure 102/51 mm Hg | 0
heart rate 72 beats per minute | 0
temperature 97.2 degrees Fahrenheit | 0
breathing 16 breaths per minute | 0
oxygen saturation 100% on room air |$|0
2/6 systolic murmur | 0
lower left sternal border | 0
moderate right lumbar paraspinal tenderness | 0
reproducible with hip flexion | 0
poor dentition | 0
multiple dental caries | 0
lactic acid 2.9 mmol/L | 0
procalcitonin >100 ng/mL | 0
platelet count 57 K/uL | 0
creatinine 1.44 mg/dL | 0
blood cultures growth of Gram-positive cocci in chains | 0
CT scan of lumbar spine with contrast | 0
small abscess in right psoas muscle | 0
transthoracic echocardiogram | 0
transesophageal echocardiogram | 0
mobile echodensity attached to tricuspid valve | 0
mobile echodensity on pacemaker lead in right ventricle | 0
confirmed infective endocarditis | 0
prescribed empiric antimicrobials | 0
vancomycin | 0
cefepime | 0
initial blood cultures grew Streptococcus agalactiae | 0
antibiotics de-escalated to ceftriaxone | 0
pacemaker extraction | 24
temporary pacing wire placement | 24
hypotensive | 24
transfer to cardiovascular intensive care unit | 24
hemodynamic support with vasopressors | 24
cultures of cardiac device | 24
repeat blood cultures | 24
growth of Gram-negative anaerobic rods | 24
antibiotics broadened to meropenem | 24
Gram-negative rods identified as Prevotella bivia | 24
P. bivia CIED related endocarditis | 24
Streptococcus agalactiae bacteremia | 24
antimicrobial therapy changed to ertapenem | 24
placement of new pacemaker device | 24
clearance of P. bivia bacteremia | 24
right psoas muscle abscess evaluated | 24
deemed too small for percutaneous drainage | 24
discharged home with home health | 240
completed 6-week course of intravenous ertapenem | 240
followed up regularly without complications | 240
