female | 0
infant | 0
born via vaginal delivery | 0
33 0/7 weeks gestation | 0
mother with hypertension | -672
mother with preeclampsia | -672
mother with poorly controlled type 2 diabetes mellitus | -672
mother with previous postpartum deep vein thrombosis | -672
mother with small pulmonary embolism | -672
birth weight 1744 g | 0
Apgar scores 9 and 9 | 0
transferred to neonatal intensive care unit | 0
severe persistent hypoglycemia | 48
umbilical venous catheter placed | 48
glucose infusion rate 21 mg/kg/min | 48
systolic murmur | 120
echocardiogram showed small patent ductus arteriosus | 120
UVC tip at foramen ovale | 120
removal of UVC | 120
fever | 168
tachypnea | 168
grunting | 168
thrombocytopenia | 168
platelets 81 000 bil/L | 168
blood culture collected | 168
cerebrospinal fluid studies collected | 168
started on gentamicin | 168
started on vancomycin | 168
started on acyclovir | 168
peripherally inserted central catheter attempted | 168
peripherally inserted central catheter failed | 168
bilious emesis | 192
abdominal ultrasound negative | 192
upper gastrointestinal studies negative | 192
cranial ultrasound showed bilateral grade 1 intraventricular hemorrhages | 192
Broviac catheter inserted | 192
blood culture grew methicillin-sensitive Staphylococcus aureus | 192
cerebrospinal fluid yielded no growth | 192
acyclovir discontinued | 192
cefotaxime added | 192
repeat echocardiogram showed 5 × 5 mm mass in atrial septum | 240
mass in contact with tip of central line | 240
Broviac pulled back under echo guidance | 240
anticoagulation withheld | 240
repeat echocardiogram showed questionable increase in size of mass | 264
gradual decrease in size of mass | 264
mass no longer seen on DOL 23 | 552
repeated cranial ultrasounds stable | 264
debridement of 1-cm nodules on scalp and leg | 408
nafcillin started | 408
gentamicin continued | 408
Broviac removed | 1008
echocardiograms 1 month after discharge stable | 1248
no other sites of infection | 1248