29 years old | 0
male | 0
penetrating stab wound to the anterior left second intercostal space | -1
right tibia-fibula fracture with intra-medullary nailing | -6048
haemodynamically unstable | -1
grade 3 haemorrhagic shock | -1
resuscitation | -1
left-sided intercostal drain inserted | -1
large haemothorax | -1
heart rate 100 | 0
respiratory rate 14 | 0
saturating at 95% on room air | 0
blood pressure 101/64 | 0
no angina | 0
no features of cardiac failure | 0
central cyanosis | 0
bruits | 0
murmurs | 0
no ST or other rhythm abnormalities | 0
chronic septic hardware of the right lower limb | -1
microbiological workup of the local septic limb deferred | 0
preliminary diagnosis of local septic hardware | 0
screening for methicillin-resistant Staphylococcus aureus | 0
antibiotic prophylaxis with broad-spectrum coverage | 0
Focused Assessment with Sonography for Trauma scan | 1
1 cm pericardial effusion | 1
contrasted computed tomographical scan of the chest | 2
cardiac TTE | 2
right ventricular outflow tract injury | 2
associated suspected thrombus | 2
small aortic root injury | 2
small pseudo-aneurysm | 2
intimal flap | 2
injury tract extended to the medial superior vena cava | 2
high index of suspicion for an SVC injury | 2
transthoracic cardiac ECHO | 3
no valvulopathies | 3
clear flow reversal or shunting | 3
regional wall motion abnormalities | 3
tamponade | 3
features of infective endocarditis | 3
preserved left ventricular ejection fraction | 3
large dense lesion | 3
beat to beat movement | 3
highly suggestive of a clot | 3
normal renal and liver function | 4
normocytic normochromic anaemia | 4
haemoglobin = 10.9 | 4
no coagulation abnormalities | 4
intubated under general anaesthesia | 5
single lumen endotracheal tube | 5
femoral cardiopulmonary bypass initiated | 6
median sternotomy performed | 7
no active bleeding | 7
aorta clamped | 8
heart arrested with cold blood cardioplegia | 8
cardioplegia given every 20 min | 8
large clot found | 9
defect in the medial wall of the RVOT | 9
clot removed | 10
RVOT repaired with continuous 3/0 prolene sutures | 11
aorta opened via a transverse ‘J’ incision | 12
0.5 cm laceration in the aortic wall | 12
repaired primarily | 13
plane between the main pulmonary artery and ascending aorta dissected | 14
right coronary artery not injured | 14
contralateral side of the ascending aorta had a defect | 14
small point injury to the base of the SVC | 14
defects primarily repaired | 15
patient weaned off of cardiopulmonary bypass | 16
closure of the femoral cannulation site | 17
sternum closed | 18
patient remained intubated | 19
transported to intensive care unit | 20
complete recovery | 120
no residual thrombus or intracardiac shunt | 120
no cardiac, respiratory, or neurological sequelae | 720