59 years old | 0
male | 0
non-obstructive hypertrophic cardiomyopathy | 0
cardiac insufficiency | 0
inotropic therapy | 0
intra-aortic balloon | 0
prioritized for cardiac transplantation | 0
blood cultures collected 24 h before transplantation | -24
blood cultures collected 48 h before transplantation | -48
negative blood cultures | -24
negative blood cultures | -48
bicaval–bipulmonary heart transplantation | 0
mechanical ventilation | 0
vasoactive drugs | 0
intra-aortic balloon | 0
immunosuppressive regimen | 0
mycophenolate mofetil | 0
cyclosporine | 0
prednisone | 0
blood culture from the donor positive for Gram-negative bacilli | 72
piperacillin–tazobactam | 72
blood cultures and surveillance cultures collected | 72
final identification turned out ColR KPC-Kp | 120
blood cultures from the recipient positive for ColR KPC-Kp | 168
surveillance cultures negative | 168
afebrile | 168
hemodynamically stable | 168
leukocyte count 26,000 cells/mm3 | 168
C-reactive protein levels 6.5 mg/dL | 168
double-carbapenems | 168
meropenem | 168
ertapenem | 168
amikacin | 168
pericarditis | 216
drainage of 1000 mL of exudate | 216
pericardial fluid cultures positive for ColR KPC-Kp | 216
surgical approach to clean the pericardium | 216
repeated surgery | 224
sternum bone fragment collected | 224
sternum bone fragment positive for ColR KPC-Kp | 224
worsening respiratory signs | 888
chest computed tomography exhibiting consolidation with lung fluid levels | 888
pulmonary cavitation due to necrosis | 888
histopathology of lung fragments | 888
pulmonary abscess with liquefactive necrosis and necrotizing arteritis | 888
septic shock | 888
antibiotic coverage extended to linezolid and fluconazole | 888
multiple organ failure | 1200
death | 1200
donor 17 years old | -72
donor male | -72
donor died from traumatic brain injury | -72
donor hospitalized in the intensive care unit for seven days | -72
piperacillin/tazobactam | -72
vancomycin | -72
blood cultures and surveillance cultures negative | -72
culture collected from the splenic artery | -72
culture positive for ColR KPC-Kp | -72
recipients of other organs did not present any infectious complications | 0
recipients of other organs did not receive specific antimicrobial treatment | 0
liver not used for transplantation | 0