68 years old | 0
male | 0
admitted to the emergency room | 0
progressive bullous and erosive skin lesions | 0
painful oral ulcer | -168
bilateral enlarged supraclavicular lymph nodes | -168
metastatic squamous cell carcinoma | -168
diabetes | -7200
diabetic nephropathy | -2880
blood pressure 93/64 mmHg | 0
heart rate 91/min | 0
respiration rate 20/min | 0
flaccid blisters | 0
exfoliated skin | 0
crusted erosions | 0
anemia | 0
thrombocytopenia | 0
white blood count 5,170/mm3 | 0
hemoglobin 7.7 mg/dL | 0
platelets 426,000/mm3 | 0
azotemia | 0
blood urea nitrogen 52.3 mg/dL | 0
creatinine 2.98 mg/dL | 0
multiple cervical and mediastinal lymph node enlargement | 0
increased fluorodeoxyglucose uptake | 0
deep ulcerative mass | 0
moderately differentiated squamous cell carcinoma | 0
suprabasal acantholysis | 0
bullous cleft formation | 0
C3 deposits in the basal layer of mucosa | 0
PNP associated with esophageal cancer | 0
palliative combination chemotherapy | 0
fluorouracil | 0
carboplatin | 0
intravenous methylprednisolone | 0
neutropenic fever | 144
broad spectrum antibiotics | 144
overwhelming sepsis | 216
death | 216