62 years old | 0
    male | 0
    chronic obstructive pulmonary disease | 0
    tobacco abuse | 0
    hypertension | 0
    former alcoholism | 0
    admitted to the hospital | 0
    abdominal pain | -96
    bloating | -96
    elevated liver function tests | 0
    elevated total bilirubin | 0
    elevated alkaline phosphatase | 0
    elevated AST | 0
    elevated ALT | 0
    acetaminophen use | -96
    bilateral leg swelling | -96
    denied dyspnea | 0
    denied chest pain | 0
    denied urinary retention | 0
    denied urinary frequency | 0
    denied headache | 0
    denied fever | 0
    denied night sweats | 0
    leukocytosis | 0
    normocytic anemia | 0
    elevated lipase | 0
    elevated lactate | 0
    elevated CRP | 0
    normal troponin | 0
    normal PTT | 0
    normal PT | 0
    normal INR | 0
    clear urinalysis | 0
    chest x-ray mass | 0
    CT abdomen findings | 0
    hepatomegaly | 0
    adrenal enlargement | 0
    lymphadenopathy | 0
    bilateral lower extremity duplex scan | 0
    right upper quadrant ultrasound | 0
    liver biopsy | 24
    CT chest | 24
    MRI brain | 24
    left upper lobe tumor | 24
    palliative radiation | 24
    small cell lung cancer diagnosis | 24
    port placement | 24
    chemotherapy started | 24
    carboplatin | 24
    etoposide | 24
    furosemide started | 24
    acute kidney injury | 72
    furosemide stopped | 72
    gentle hydration started | 72
    worsening leukocytosis | 72
    post-obstructive pneumonia | 72
    lethargy | 72
    hypotension | 72
    hypoxic respiratory failure | 72
    transfer to ICU | 72
    chest x-ray congestion | 72
    septic shock | 72
    tachycardia | 72
    low systolic blood pressure | 72
    Levophed started | 72
    colloid administration | 72
    antibiotic switch | 72
    levofloxacin | 72
    meropenem | 72
    renal failure worsened | 96
    intubation | 96
    norepinephrine use | 96
    vasopressin started | 96
    bronchoscopy | 96
    Enterobacter aerogenes culture | 96
    negative blood cultures | 96
    sinus tachycardia | 96
    supraventricular tachycardia | 96
    vasopressor requirement increase | 96
    troponin elevation | 96
    fever | 96
    ECG showing Brugada syndrome | 96
    heparin started | 96
    antiplatelet therapy | 96
    echocardiogram findings | 96
    defervescence | 120
    ECG resolution of Brugada wave | 120
    extubation | 120
    dialysis started | 120
    lethargy increased | 120
    comfort care elected | 120
    patient deceased | 120
    