62 years old| 0
female | 0
aortobifemoral bypass | -2640
abdominal aortic aneurysm | -2640
coronary artery stenting | -240
unstable angina | -240
presentation to emergency department | 0
fatigue | -24
myalgia | -24
left flank pain | -24
left flank pain irradiating to left thigh | -24
acute pain | -96
severe pain | -96
partial pain relief | -72
temporary pain relief | -72
no fever | 0
no urinary symptoms | 0
soft abdomen | 0
severe leukocytosis (27,000 cells/mm3) | 0
elevated CRP (300 mg/L) | 0
altered liver function test | 0
positive urinalysis | 0
leukocyturia | 0
microscopic hematuria | 0
bacteriuria | 0
CT-urography | 0
large left retroperitoneal hematoAurinoma | 0
6 mm left proximal ureteral stone | 0
ureteral rupture | 0
urinary extravasation | 0
renal pelvis blood clots | 0
calyceal blood clots | 0
medical treatment | 0
supportive treatment | 0
intravenous hydration | 0
antibiotics | 0
analgesics | 0
urgent endoscopic drainage | 0
JJ stent insertion | 0
Foley urinary catheter | 0
urine culture showing multi-sensitive Escherichia Coli | 0
discharged home | 240
Foley catheter kept for 10 days | 240
ciprofloxacin | 240
follow-up meeting in 3 weeks | 240
scanographic control scheduled | 240
return to emergency department | 408
septic shock | 408
intensive care unit admission | 408
imaging showed previous findings | 408
JJ stent in place | 408
CT-guided left 8F nephrostomy insertion | 408
10F left percutaneous drain insertion | 408
retroperitoneal collection drainage | 408
fungal infection (Candida Kefyr) | 408
treated fungal infection | 408
recovered from infectious process | 408
percutaneous catheter draining urine | 408
persistent ureteral fistula | 408
quadruple drainage | 408
Foley catheter | 408
JJ stent | 408
nephrostomy tube | 408
percutaneous drain | 408
complicated renal colic episode | -1440
laparoscopic nephrectomy | 1440
subtotal ureterectomy | 1440
necrotic ureter | 1440
inflamed ureter | 1440
stone extraction | 1440
aortobifemoral bypass effect on ureteral fragility | 0
ureteral rupture mechanism | 0
stone migration | 0
impaction | 0
ureteral wall injury | 0
erosion | 0
weakening | 0
intrarenal pressure elevation | 0
intraureteric pressure elevation | 0
ureteral dilatation | 0
genitofemoral nerve irritation | 0
persistent ureteral extravasation | 408
failure of conservative management | 1440
ureteral necrosis | 1440
bacterial infection | 408
severe inflammatory process | 408
delay in presentation | 408
delay in urinary drainage | 408
fibrotic retroperitoneum | 408
adherent retroperitoneum | 408
friable ureteral tissue | 408
urinoma | 408
sepsis | 408
kidney loss | 1440
