58 years old|0
female|0
presented to the emergency department|0
unresponsive|-24
sudden onset headache|-24
urinary tract infection|-72
unspecified oral treatment|-72
discharged (from ED)|-72
mid-stream urine sample positive for E. coli|-72
samples from previous years positive for E. coli|0
Glasgow Coma Score 6/15|0
right-sided weakness|0
facial droop|0
afebrile|0
no neck stiffness|0
myoclonic jerks in both arms|0
anxiety|0
sertraline treatment|0
smoked thirty cigarettes per day|0
alcohol intake seven units per day|0
no recent history of travel|0
no recent history of trauma|0
no recent history of surgery|0
intubated in the ED|0
transferred to the Intensive Care Unit|0
working diagnosis of stroke|0
possible CNS infection|0
ceftriaxone 2 grams 12-hourly|0
aciclovir 640 milligrams 12-hourly|0
white cell count 9.8 10^9/L|0
neutrophils 8.8 10^9/L|0
lymphocytes 0.2 10^9/L|0
platelets 62 10^9/L|0
C-reactive protein 643 mg/L|0
creatinine 232 μmol/L|0
urea 19.7 mmol/L|0
CT brain showing left-sided MCA infarct|0
MRI brain showing right internal capsule infarct|0
debris in the ventricles|0
blood cultures positive for E. coli|0
lumbar puncture performed|0
CSF turbid|0
CSF white cell count 15,680 10^6/L|0
CSF polymorphs 95%|0
CSF lymphocytes 5%|0
CSF red blood cells 220 10^6/L|0
CSF protein 4.26 g/L|0
CSF glucose 0.4 mmol/L|0
serum glucose 7.0 mmol/L|0
CSF gram-negative organisms|0
E. coli culture|0
unenhanced CT brain confirming right internal capsule infarct|168
repeat lumbar puncture on day 11|264
CSF clear and colorless|264
CSF white cell count 14 10^6/L|264
CSF polymorphs 30%|264
CSF lymphocytes 70%|264
CSF red blood cells 1 10^6/L|264
CSF protein 0.55 g/L|264
CSF glucose 4.1 mmol/L|264
serum glucose 6.8 mmol/L|264
no bacterial growth in CSF|264
prolonged ICU stay|0
mechanical ventilation for 27 days|648
reliable neurological examination after sedation hold|648
left-sided hemiparesis|648
ceftriaxone continued until day 25|600
ceftriaxone dose reduced to 2 grams daily|600
aciclovir stopped|0
Strongyloides serology negative|0
HIV serology negative|0
Hepatitis B serology negative|0
Hepatitis C serology negative|0
renal tract ultrasound showing no hydronephrosis|0
renal tract ultrasound showing no collection|0
transthoracic echocardiogram normal|0
MRI brain with contrast on day 27|648
persistent ventriculitis|648
subacute infarct in right internal capsule|648
trapped occipital horn of right lateral ventricle|648
tracheostomy performed|648
marked global weakness|648
successfully decannulated|648
stepped-down to Stroke ward|696
intensive physiotherapy|696
neuro-rehabilitation|696
MRI brain on day 41|984
mild reduction of ring-enhancing lesion|984
persistent ventricular debris|984
discharged to rehabilitation facility|1392
eight weeks of intravenous antibiotics|1392
follow-up imaging at four months|1392
significant regression of findings|1392
no evidence of hydronephrosis|0
no evidence of collection|0
