67 years old | 0 | 0 
male | 0 | 0 
admitted to the hospital | 0 | 0 
left leg swelling | -168 | 0 
cactus plant injury | -168 | -168 
Primary Sclerosing Cholangitis | 0 | 0 
mild Ulcerative Colitis | 0 | 0 
deranged liver function tests | 0 | 0 
progressive left leg swelling | -48 | 0 
worsening of erythema | -48 | 0 
pain | -48 | 0 
felt generally unwell | -48 | 0 
paramedic assistance | -24 | -24 
presentation to ED | 0 | 0 
Blood Pressure (BP): 71/41mmHg | 0 | 0 
Mean Arterial Pressure (MAP): 48mmHg | 0 | 0 
Respiratory Rate: 36 breaths per minute | 0 | 0 
Heart Rate (HR): 125 beats per minute | 0 | 0 
sinus tachycardia | 0 | 0 
Temperature: 39°C | 0 | 0 
Oxygen Saturation: 86% with 0.21 FiO2 | 0 | 0 
admitted to the intensive care unit (ICU) | 0 | 0 
pH 7.15 | 0 | 0 
PO2 84 | 0 | 0 
HCO3 15 | 0 | 0 
Lactate 7.6 | 0 | 0 
Sodium (Na) 134 | 0 | 0 
Urea 7.6 | 0 | 0 
Creatinine (sCr) 173 | 0 | 0 
eGFR 27 | 0 | 0 
White Cell Count (WCC) 13.8 | 0 | 0 
C-reactive protein (CRP) 22 | 0 | 0 
Hemoglobin (Hb) 114 | 0 | 0 
Platelet (Plt) 81 | 0 | 0 
Liver Function Test (LFT)- Total Bilirubin (Bili) 99 | 0 | 0 
Alanine transaminase (ALT) 61 | 0 | 0 
Aspartate aminotransferase (AST) 83 | 0 | 0 
Alkaline Phosphatase (ALP) 96 | 0 | 0 
Triple vasopressor support initiated | 0 | 0 
Noradrenaline 20mcg/min | 0 | 24 
Adrenaline 20mcg/min | 0 | 24 
Vasopressin 0.04units/min | 0 | 24 
Piperacillin-Tazobactam IV 4.5g | 0 | 0 
Meropenem IV 2g | 0 | 168 
Lincomycin IV 600mg | 0 | 168 
Vancomycin IV 2g | 0 | 168 
Emergency left lower limb fasciotomy | 0 | 0 
debridement | 0 | 0 
below knee amputation | 0 | 0 
LRINEC Score of 5 | 0 | 0 
extensive left foot and below knee tissue necrosis | 0 | 0 
dishwasher fluid | 0 | 0 
liquefied fat | 0 | 0 
unviable skin and muscle | 0 | 0 
Histopathology | 0 | 0 
post operatively | 24 | 24 
oliguria | 24 | 168 
blood gas showed severe acidosis | 24 | 24 
left internal jugular vascath insertion | 24 | 24 
continuous renal replacement therapy (CRRT) | 24 | 168 
Ventilation sedation | 24 | 168 
Propofol 170mg/hr | 24 | 168 
Fentanyl 40mcg/hr | 24 | 168 
CRRT (Day 1) | 24 | 24 
heparin circuit | 24 | 24 
Renal dose | 24 | 24 
Triple vasopressor support continued | 24 | 168 
Noradrenaline 23mcg/min | 24 | 168 
Adrenaline 18mcg/min | 24 | 168 
Vasopressin 0.04units/min | 24 | 168 
Antibiotics (MLV) | 24 | 168 
Meropenem IV 2g TDS | 24 | 168 
Lincomycin IV 600mg TDS | 24 | 168 
Vancomycin IV 2g BD | 24 | 168 
Intravenous Immunoglobin G (IVIgG) therapy 100g | 24 | 24 
taken back to theatre | 48 | 48 
source control | 48 | 48 
viability of the left stump | 48 | 48 
no evidence of necrotic tissue | 48 | 48 
Rapid Atrial Fibrillation (RAF) | 48 | 168 
HR 110bpm | 48 | 48 
oliguric | 48 | 168 
pH 7.40 | 48 | 48 
Lactate 3.9 | 48 | 48 
Sodium (Na) 131 | 48 | 48 
sCr 116 | 48 | 48 
WCC 26 | 48 | 48 
CRP 105 | 48 | 48 
Procalcitonin (PCT) 21.18 μg/L | 48 | 48 
Hb 83 | 48 | 48 
Plt 63 | 48 | 48 
INR 3.1 | 48 | 48 
Fibrinogen 2.4 | 48 | 48 
Echocardiography | 48 | 48 
Moderate segmental left ventricular dysfunction | 48 | 48 
Ejection Fraction 40-45% | 48 | 48 
Dilated atria bilaterally | 48 | 48 
Raised Right Atrial Pressure | 48 | 48 
Amiodarone loading dose 300mg | 48 | 48 
maintenance dose 900mg | 48 | 168 
Antibiotics remained unchanged (MLV) | 48 | 168 
CRRT (Day 2) | 48 | 48 
AN69 anti-inflammatory heparin laden adsorbing filter | 48 | 48 
Oxiris Filter | 48 | 48 
Citrate based anticoagulation circuit | 48 | 168 
Sepsis Induced Coagulopathy (ISTH -SIC criteria) | 72 | 72 
bedside surgical debridement | 72 | 72 
pH 7.31 | 72 | 72 
Lactate 2.4 | 72 | 72 
Sodium (Na) 135 | 72 | 72 
sCr 79 | 72 | 72 
WCC 27 | 72 | 72 
CRP 127 | 72 | 72 
Hb 78 | 72 | 72 
Plt 50 | 72 | 72 
INR 2.0 | 72 | 72 
Histopathology consistent with NF | 72 | 72 
Wound culture for microscopy culture and sensitivity (MCS) | 72 | 72 
medium growth of GBSPn | 72 | 72 
Tissue culture (intraoperatively) | 72 | 72 
medium growth of GBSPn | 72 | 72 
Vasopressor support - weaning | 72 | 168 
Noradrenaline 20mcg/min | 72 | 168 
Adrenaline weaned off | 72 | 72 
Vasopressin 2.4units/min | 72 | 168 
Antibiotics remained unchanged (MLV) | 72 | 168 
CRRT (Day 3) | 72 | 72 
oliguric | 96 | 168 
Furosemide IV 250mg | 96 | 96 
renal response | 96 | 96 
Citrate based CRRT | 96 | 168 
new onset purpura | 96 | 96 
multiple weeping skin tears | 96 | 96 
RAF HR 130 | 96 | 168 
pH 7.36 | 96 | 96 
Lactate 1.5 | 96 | 96 
Sodium (Na) 130 | 96 | 96 
sCr 116 | 96 | 96 
WCC 33 | 96 | 96 
CRP 103 | 96 | 96 
PCT 15.37 | 96 | 96 
Hb 91 | 96 | 96 
Plt 53 | 96 | 96 
INR 1.7 | 96 | 96 
LFT - Bili 131 | 96 | 96 
AST 127 | 96 | 96 
ALP 121 | 96 | 96 
Double inotropic support | 96 | 168 
Noradrenaline 20mcg/min | 96 | 168 
Vasopressin 2.4units/min | 96 | 168 
Antibiotics remained unchanged (MLV) | 96 | 168 
CRRT (Day 4) | 96 | 96 
Amiodarone infusion | 96 | 168 
fulminant hepatic failure | 120 | 120 
encephalopathy | 120 | 120 
refractory oliguria | 120 | 168 
pH 7.39 | 120 | 120 
Lactate 1.2 | 120 | 120 
Sodium (Na) 134 | 120 | 120 
sCr 124 | 120 | 120 
WCC 39.5 | 120 | 120 
CRP 74 | 120 | 120 
Hb 116 | 120 | 120 
Plt 49 | 120 | 120 
INR 1.5 | 120 | 120 
LFT- Bili 139 | 120 | 120 
AST 69 | 120 | 120 
ALT 97 | 120 | 120 
ALP 140 | 120 | 120 
Dual inotropic support | 120 | 168 
Noradrenaline 20mcg/min | 120 | 168 
Vasopressin weaned off | 120 | 120 
Antibiotics remained unchanged (MLV) | 120 | 168 
CRRT (Day 5) | 120 | 120 
severely deconditioned | 144 | 144 
ICU acquired weakness | 144 | 144 
unarousable | 144 | 144 
no response to noxious stimuli | 144 | 144 
intubated and ventilated | 144 | 168 
Pressure Support Ventilation | 144 | 168 
refractory oliguria | 144 | 168 
PH 7.44 | 144 | 144 
Lactate 1.1 | 144 | 144 
WCC 43.5 | 144 | 144 
CRP 109 | 144 | 144 
Hb 90 | 144 | 144 
Plt 57 | 144 | 144 
INR 1.5 | 144 | 144 
LFT - Bili 150 | 144 | 144 
AST 95 | 144 | 144 
ALP 154 | 144 | 144 
Sedation weaned off | 144 | 144 
off vasopressor | 144 | 144 
Noradrenaline weaned off | 144 | 144 
Antibiotic de-escalation | 144 | 168 
Lincomycin and Vancomycin ceased | 144 | 144 
Meropenem IV 2g TDS continued | 144 | 168 
CRRT (Day 6) | 144 | 144 
Hyper-Ammonium Therapy initiated | 144 | 168 
Rifaximin NGT 550mg BD | 144 | 168 
Lactulose NGT 20ml TDS | 144 | 168 
2 units of PRBCs transfusion | 144 | 144 
jaundice | 168 | 168 
Hypoactive delirium | 168 | 168 
deeply sedated | 168 | 168 
RASS -5 | 168 | 168 
new onset lateralizing signs | 168 | 168 
CT Brain | 168 | 168 
No acute intracranial pathology | 168 | 168 
Ultrasound abdomen | 168 | 168 
Acute Calculous Cholecystitis | 168 | 168 
pH 7.44 | 168 | 168 
Lactate 1.1 | 168 | 168 
WCC 44.3 | 168 | 168 
CRP 109 | 168 | 168 
Hb 129 | 168 | 168 
Plt 66 | 168 | 168 
INR 1.3 | 168 | 168 
LFT - Bili 235 | 168 | 168 
AST 75 | 168 | 168 
ALP 175 | 168 | 168 
Conjugated Bilirubin 142 | 168 | 168 
Meropenem IV 2g TDS | 168 | 168 
CRRT (Day 7) | 168 | 168 
Heparin circuit | 168 | 168 
Anuria | 192 | 192 
Hypotensive BP 71/33 | 192 | 192 
MAP 51mmHg | 192 | 192 
Febrile 39°C | 192 | 192 
RAF HR 160 | 192 | 192 
Significant deterioration | 192 | 192 
palliative care pathway | 192 | 192 
deceased | 192 | 192 
Family was involved | 192 | 192 
consent for critical care supportive therapy was withdrawn | 192 | 192 
not deemed to be a coroner's case | 192 | 192 
Troponin 616 | 192 | 192 
Ammonia 158 | 192 | 192 
LFT - Bili 352 | 192 | 192 
AST 100 | 192 | 192 
ALP 299 | 192 | 192 
CRRT (Day 8) | 192 | 192 
Renal recovery assessment | 192 | 192 
Furosemide IV 250mg | 192 | 192 
Acetazolamide IV 500mg | 192 | 192 
Vasopressor support | 192 | 192 
Noradrenaline 2.5mcg/min | 192 | 192 
Antibiotic regimen | 192 | 192 
Lincomycin IV 600mg TDS | 192 | 192 
Meropenem IV 2g TDS | 192 | 192 
Digoxin IV 500mcg | 192 | 192 
Metoprolol IV 15mg | 192 | 192