65 years old | 0
male | 0
diabetic | 0
transhiatal oesophagectomy | 0
gastric resection | 0
adenocarcinoma of the gastro-oesophageal junction | 0
progressive breathlessness | 240
severe breathlessness | 264
reduced air entry on the left hemithorax | 264
diaphragmatic hernia | 264
emergency thoracolaparotomy | 264
severe respiratory distress | 264
inability to lie down | 264
nasal flaring | 264
active accessory muscles | 264
sweating | 264
dilated neck veins | 264
respiratory rate 40/min | 264
thready pulse | 264
pulse rate 180/min | 264
blood pressure 90/60 mmHg | 264
oxygen saturation 85-90% | 264
supplemental oxygen 6 l/min | 264
preoxygenated | 264
induced in sitting position | 264
fluid resuscitation | 264
rapid sequence induction technique | 264
haemodynamic instability | 264
noradrenaline infusion | 264
airway pressures 42 cm of water | 264
reduction of herniated colon | 264
improvement in haemodynamic parameters | 264
resolution of high airway pressures | 264
noradrenaline infusion weaned off | 264
ventilatory support | 264
severe mixed acidosis | 264
weaned off and extubated | 288
septic shock | 288
anastomotic leak | 288 
death | 288