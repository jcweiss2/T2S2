45 years old | 0
    male | 0
    low backache | -17520
    weakness of both lower limbs | -17520
    urinary retention | -48
    constipation | -48
    full power in upper limbs | 0
    Grade 3 power in lower limbs | 0
    thickened ligamentum flavum | 0
    cord oedema | 0
    distended abdomen | 0
    soft abdomen | 0
    no ascites | 0
    no organomegaly | 0
    bowel sounds present | 0
    urinary bladder catheterized | 0
    laminectomy | 0
    decompression of the spine | 0
    invasive blood pressure monitoring | 0
    arterial blood gas (ABG) monitoring | 0
    propofol | 0
    fentanyl citrate | 0
    rocuronium bromide | 0
    tracheal intubation | 0
    mechanical prophylaxis for deep vein thrombosis | 0
    warm air blanket | 0
    sevoflurane | 0
    propofol infusion | 0
    vecuronium bromide | 0
    surgery duration 5 hours | 0
    intermittent fentanyl | 0
    intravenous saline | 0
    colloid (tetra starch) | 0
    noradrenaline | 0
    blood loss 250 ml | 0
    urine output 250 ml | 0
    metabolic acidosis (2 hours post-induction) | 120
    severe canal stenosis | 0
    methylprednisolone bolus | 0
    methylprednisolone infusion | 0
    inadequate motor power | 0
    inadequate respiratory effort | 0
    metabolic acidosis (post-surgery) | 300
    blood sugar 246 mg% | 0
    urine ketone negative | 0
    insulin infusion | 0
    elective ventilation | 0
    central venous line inserted | 0
    central venous pressure 1-2 cm H2O | 0
    fluid therapy resolved acidosis | 24
    fluid therapy resolved oliguria | 24
    extubated | 24
    high normal kidney function test values | 24
    normal serum sodium | 24
    normal serum potassium | 24
    normal thyroid status | 24
    upper limb power almost normal | 24
    lower limbs power 1/5 | 24
    continuation of methylprednisolone | 24
    tense abdominal distension | 30
    respiratory distress | 30
    respiratory alkalosis | 30
    reintubation | 30
    ventilation | 30
    normal chest X-ray | 30
    normal echocardiogram | 30
    inconclusive abdominal ultrasound | 30
    computerized tomography of abdomen | 30
    colonic gaseous distension | 30
    no free fluid in abdomen | 30
    Ryle's tube inserted | 30
    neostigmine started | 30
    deranged kidney function test (POD 2) | 48
    high-grade fever (POD 2) | 48
    cultures sent | 48
    antibiotics upgraded | 48
    sepsis | 48
    hypocalcaemia (serum calcium 4.1 mg%) | 48
    hypoalbuminemia (2 g%) | 48
    normal serum amylase | 48
    normal serum lipase | 48
    factitious hypocalcaemia ruled out | 48
    hyperphosphatemia | 48
    low parathormones | 48
    normal magnesium levels | 48
    IV albumin started | 48
    IV calcium started | 48
    oral calcitriol started | 48
    renal functions resolving (POD 3) | 72
    acidosis resolving (POD 3) | 72
    neostigmine trial | 72
    prokinetics | 72
    laxatives | 72
    persistent abdominal symptoms | 72
    no faecal impaction | 72
    decompressive sigmoidoscopy | 72
    total parenteral nutrition (TPN) started | 72
    GI symptoms decreasing | 96
    procalcitonin decreasing | 96
    total leucocyte count decreasing | 96
    serum calcium 7.7 mg% | 96
    extubated (POD 9) | 216
    reintubation (18 hours later) | 234
    severe tachypnoea | 234
    decreased consciousness | 234
    pulmonary embolism ruled out | 234
    no fresh MRI spine changes | 234
    cerebrospinal fluid analysis normal | 234
    tracheostomised (POD 13) | 312
    steady improvement | 336
    ventilator weaned | 336
    full consciousness | 336
    good power in all limbs | 336
    normal calcium levels | 336
    normal albumin levels | 336
    no GI symptoms | 336
    decannulated | 336
    discharged | 336
    