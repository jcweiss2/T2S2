47 years old | 0
female | 0
cirrhosis | -8760
intestinal failure associated liver disease | -8760
short bowel syndrome | -8760
small intestinal bacterial overgrowth | -8760
gastrointestinal dysmotility | -8760
multivisceral transplantation | 0
liver biopsy | -8760
advanced cirrhosis | -8760
methylprednisolone | 0
alemtuzumab | 0
prednisolone | 0
tacrolimus | 0
cyclosporine | 40
meropenem | 0
vancomycin | 0
liposomal amphotericin B | 0
co-trimoxazole | 0
acyclovir | 0
Candida glabrata | -72
increased dose of liposomal amphotericin B | -72
cutaneous drug reaction | -96
voriconazole | -96
pyrexia | -96
intermittent bacteremia | -96
enterococci | -96
Elizabethkingia meningoseptica | -96
Staphylococcus haemolyticus | -96
Escherichia coli | -96
no fungemia | -96
micafungin | -96
low serum voriconazole levels | -96
diffuse maculopapular rash | -79
graft-versus-host disease | -79
peripheral blood chimerism analysis | -79
bone marrow failure | -90
frequent red cell and platelet transfusions | -90
bone marrow examination | -90
immunosuppression increased | -90
high-dose methylprednisolone | -90
basiliximab | -90
alemtuzumab | -90
immunosuppression withdrawn | -120
haplo-identical bone marrow transplant | -168
granulocyte infusion | -168
dysarthria | -168
unilateral isolated upper motor neurone facial nerve palsy | -168
cranial computed tomography scan | -168
acute frontal infarct | -168
extensive and catastrophic infarcts | -24
treatment withdrawn | -24
death | 0
post mortem examination | 0
invasive mucormycosis | 0
lung involvement | 0
brain involvement | 0
heart involvement | 0
liver involvement | 0
left ventricular fungal thrombus | 0