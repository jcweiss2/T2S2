preterm | -216 
male | 0 
born | -216 
gestation 29 + 3 weeks | -216 
spontaneous vaginal delivery | -216 
uncomplicated pregnancy | -216 
healthy 33-year-old G2P1 mother | -216 
birth weight 1650 g | -216 
90th percentile | -216 
ventilatory support | -216 
surfactant | -216 
infant respiratory distress syndrome | -216 
umbilical artery catheter | -216 
monitoring blood pressure | -216 
no umbilical venous catheter | -216 
transferred to local hospital | -192 
readmitted | -168 
suspected septicaemia | -168 
cardiac arrhythmias | -168 
alternating tachycardia | -168 
bradycardia | -168 
mean blood pressure 33 mm Hg | -168 
weak peripheral pulses | -168 
prolonged capillary refill | -168 
mild respiratory distress | -168 
grunting | -168 
oxygen saturation 90% | -168 
no heart murmur | -168 
lungs clear | -168 
abdomen soft | -168 
no hepatosplenomegaly | -168 
circulatory support | -168 
intravenous fluids | -168 
antibiotics | -168 
suspected septicaemia | -168 
blood cultures negative | -168 
rectal culture positive | -168 
sputum culture positive | -168 
Coxsackie B III virus | -168 
chest X-ray no significant abnormalities | -168 
electrocardiogram | -168 
ST-depression | -168 
ST elevation | -168 
increased cardiac enzymes | -168 
myocardial damage | -168 
echocardiography | -168 
left-ventricular dysfunction | -168 
severely hypokinetic posterolateral wall | -168 
hyperkinetic septum | -168 
pericardial effusion | -168 
abnormal coronary anatomy excluded | -168 
no sources for thromboemboli | -168 
clotting studies normal | -168 
respiratory distress increased | -156 
mechanical ventilation | -156 
inotropics | -156 
diuretic therapy | -156 
milrinone | -156 
captopril | -156 
necrotizing enterocolitis | -156 
antibiotics | -156 
parental nutrition | -156 
discharged | 0 
nasogastric tube feeding | 0 
medication for chronic heart failure | 0 
diuretics | 0 
beta blocker | 0 
ACE inhibitor | 0 
echocardiographic follow-up | 0 
persisting pattern of decreased left-ventricular function | 0 
increased right ventricle pressure | 0 
no compensatory hypertrophy | 0 
global impairment of ventricular function | 0 
post–myocarditis cardiomyopathy | 0 
progressive left-ventricle dilatation | 120 
suprasystemic pressure in right ventricle | 120 
heart transplantation evaluation | 120 
heart function deteriorated | 216 
died | 216 
progressive heart failure | 216 
medication-resistant | 216 
autopsy | 216 
increased heart weight | 216 
intracardiac anatomy normal | 216 
coronary arteries normal | 216 
focal intima hyperplasia | 216 
global subendocardial fibroelastosis | 216 
scar tissue | 216 
loss of myocytes | 216 
hypertrophy of residual myocytes | 216 
thickened right ventricle | 216 
dilated pulmonary trunk | 216 
alveolar and septal hemorrhage | 216 
hemosiderophages | 216 
venous congestion | 216 
no pulmonary arterial hypertension | 216