81 years old | 0
male | 0
ischemic stroke | 0
hypertension | 0
stage 3 nephropathy | 0
multiple myeloma type IgA lambda | 0
symptomatic anemia | -17520
monoclonal gammaglobulinemia | -17520
melphalan | -17520
prednisone | -17520
bortezomib | -17520
paraproteinemia decrease | -17520
anemia recovery | -17520
lenalidomide | -12960
dexamethasone | -12960
poorly tolerated | -12960
clinically stable condition | 0
low paraproteinemia | 0
mild anemia | 0
hemoglobin 6.8 mmol/L | 0
admitted to Department of Internal Medicine | 0
dyspnea | 0
general discomfort | 0
muscle weakness | 0
poor performance status (WHO 3–4) | 0
tachypnea | 0
normal body temperature | 0
normal blood pressure | 0
no pneumonia | 0
no cardiac decompensation | 0
respiratory compensated metabolic acidosis | 0
anion gap increased | 0
arterial lactate level elevated | 0
lactic acidosis | 0
normal vital parameters | 0
normal ECG | 0
contrast enhancement of major vessels | 0
no pulmonary embolism | 0
normal liver function | 0
stable kidney function | 0
eGFR 41 mL/min | 0
elevated PSA level | 0
no toxic cause | 0
enlarged prostate | 0
hydronephrosis right kidney | 0
liver nodules | 0
enlarged mediastinal lymph nodes | 0
enlarged paratracheal lymph nodes | 0
sclerotic bone metastases | 0
metastatic prostate cancer | 0
cyproterone acetate | 0
prednisone | 0
thiamine | 0
no chemotherapy | 0
clinically deteriorated | 24
lactate levels increased | 24
pH levels lowered | 24
unconscious | 24
admitted to ICU | 24
NaHCO3 | 24
cardiac arrest | 72
DNR | 72
locally advanced prostate cancer | 72
metastatic prostate cancer | 72
encasement right ureter | 72
metastases thoracic spine | 72
metastases lumbar spine | 72
metastases liver | 72
metastases lungs | 72
metastases peritoneum | 72
bilateral tumor thrombi | 72
no multiple myeloma activity | 72
no cardiac ischemia | 72
TP53 mutation | 72
PIK3CA mutation | 72
no PTEN mutations | 72
no IDH1 mutations | 72
