33 years old | 0
female | 0
left leg pain | 0
admitted to the hospital | 0
cardiac arrest | 0
attempted suicide by hanging | 0
incarcerated | 0
advanced cardiovascular life support initiated | 0
emergent left leg IO needle placement | 0
intubated | 0
admitted to the neurologic intensive care unit | 0
postextubation | 48
hospital day 2 | 48
complained of left leg pain | 48
severe tenderness at the left shin IO site | 48
decreased strength on ankle dorsal and plantar flexion | 48
mild dorsal foot swelling | 48
conventional radiograph (CR) of the left leg obtained | 48
small, shallow, linear cortical defect in the proximal diaphysis of the lateral tibial cortex | 48
no associated fracture line | 48
moderate localized soft tissue swelling of the left knee and lower leg | 48
hospital day 4 | 96
increased swelling of the left leg | 96
erythema of the left leg | 96
differential considerations: deep venous thrombosis (DVT) | 96
differential considerations: infection | 96
differential considerations: sequela of possible blunt soft tissue trauma | 96
elevated D-dimer | 96
pulmonary CT angiography (CTA) negative for pulmonary embolism (PE) | 96
ultrasound for DVT negative | 96
CT delayed venous phase extended from the pelvis through bilateral lower extremities | 96
small, shallow, linear cortical defect in the anterolateral tibia | 96
no penetration into the medullary cavity | 96
asymmetric soft tissue swelling of the left tibialis anterior muscle | 96
left lower extremity magnetic resonance imaging (MR) ordered | 96
small, partial-thickness cortical defect along the anterior lateral aspect of the proximal tibia | 96
marked distention of the anterior muscle compartment | 96
less conspicuous distention of the deep posterior and proximal aspect of the lateral compartments | 96
anterior compartment: abnormally increased T1 and T2 signal | 96
early subacute intramuscular hemorrhage | 96
normal marrow signal of the tibia and fibula | 96
patient elected to prematurely terminate the MR exam | 96
contrast portion of the study not performed | 96
surgical consultation for potential fasciotomy obtained | 96
clinical signs and symptoms of compartment syndrome deemed equivocal | 96
watchful waiting approach adopted | 96
intracompartmental pressure measurements not obtained | 96
pain and swelling gradually decreased | 120
discharged from the hospital | 120
