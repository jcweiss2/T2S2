18 years old | 0
male | 0
hypertension | 0
insulin-dependent diabetes | 0
diabetic retinopathy | 0
weight loss | -336
iron deficiency anemia | -336
colon ascendens tumor | -336
liver metastases | -336
right hemicolectomy | -336
adenocarcinoma | -336
activated BRAF mutation | -336
mismatch repair-deficient (MMR-D)/microsatellite-instable (MSI) tumor | -336
pembrolizumab | 0
cold | -7
leukocytosis | -7
C-reactive protein | -7
fever | -22
coughing | -22
AST | -22
ALT | -22
ICI-induced hepatitis grade 2 | -22
prednisolone | -22
dyspnea | -29
myocardial infarction | -29
septal hypokinesia | -29
somnolence | -30
dysarthria | -30
hoarseness | -30
pain in neck and right leg | -30
difficulty raising right leg | -30
CK | -30
myoglobin | -30
MG | -30
albumin in cerebrospinal fluid | -30
pain in neck and shoulders | -34
severe dysarthria and dysphagia | -34
absent reflexes | -34
intubated | -35
methylprednisolone | -35
intravenous immunoglobulins | -35
infliximab | -37
carbon dioxide retention | -39
sinus bradycardia | -39
death | -39
autopsy | -39
significant stenosis of the right coronary artery | -39
fibrosis or signs of recent myocardial infarction | -39
tongue softened | -39
metastasis in the right liver lobe | -39
pronounced inflammatory infiltration of lymphocytes | -39
fibrosis | -39
myocardial infarction | -39
inflammatory infiltrate | -39
HCC | -39
fibrosis stage 2–3 | -39
respiratory insufficiency | -39