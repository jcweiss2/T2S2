66 years old | 0
male | 0
dual-chamber pacemaker | -10512
sick sinus syndrome | -10512
paroxysmal atrial fibrillation | -10512
severe lumbar back pain | 0
mental status changes | 0
hypotension | 0
acute renal failure | 0
hypoxemic respiratory failure | 0
emergent intubation | 0
severe sepsis | 0
hemodynamic support | 0
vasopressin | 0
norepinephrine | 0
blood cultures | 0
methicillin-sensitive Staphylococcus aureus | 0
vancomycin | 0
nafcillin | 0
transthoracic echocardiogram | 0
left ventricular ejection fraction | 0
patent foramen ovale | 0
Doppler of the intra-atrial septum | 0
computed tomography scan | 0
osteomyelitis | 0
magnetic resonance imaging | 0
septic emboli | 0
transesophageal echocardiogram | 0
vegetation | 0
right atrium | 0
pacemaker lead | 0
tricuspid valve | 0
right ventricle | 0
cardiothoracic surgery | 0
surgical intervention | 0
laser lead extraction | 0
Indigo Penumbra system | 0
intracardiac echocardiography | 0
aspiration | 0
vegetation removal | 0
RA lead extraction | 0
RV lead extraction | 0
pocket inspection | 0
suture | 0
hemostasis | 0
procedure time | 0
blood loss | 0
pathology | 0
gram-positive cocci | 0
culture-positive | 0
methicillin-sensitive Staphylococcus aureus | 0
condition improved | 48
condition worsened | 72
tissue necrosis | 72
lactic acidosis | 72
renal failure | 72
withdraw care | 72
extubation | 72
death | 72