87 years old | 0
    male | 0
    presented to the emergency department | 0
    generalized weakness | 0
    diabetic ketoacidosis | 0
    uncontrolled diabetes mellitus | 0
    chronic renal failure | 0
    left below knee amputation | 0
    penetrating keratoplasty procedure in the right eye | -240
    afebrile | 0
    confused | 0
    generally weak | 0
    incoherent | 0
    complete ophthalmoplegia | 0
    no marked signs of inflammation | 0
    non-reactive pupils | 0
    no view of the posterior fundus | 0
    reduction in right visual acuity | 0
    ophthalmic B scan revealed infiltration of the right globe | 0
    computed tomography scan of the orbit and brain | 0
    cavernous sinus thrombosis | 0
    orbital cellulitis | 0
    intravenous meropenem | 0
    vancomycin | 0
    heparin | 0
    level of consciousness deteriorated | 24
    seizures | 24
    orbital involvement of the infection worsened | 24
    CT brain venography | 24
    poor enhancement of the right cavernous sinus | 24
    lumbar puncture sample negative for microorganisms | 24
    provisional diagnosis of mucormycosis | 24
    presence of micronasal abscesses | 24
    right alar blackish discoloration | 24
    intravenous amphotericin B | 24
    caspofungin | 24
    rapid progression to the orbit | 48
    gangrenous area on the tip of the nose | 48
    suspicion of mucormycosis confirmed | 48
    surgical debridement | 48
    right orbital exenteration | 48
    widespread deep excision of the necrotic area | 48
    peri-operative intravenous antibiotics | 48
    antifungals | 48
    transferred to the intensive care unit | 48
    Glasgow Coma Score of three post-operatively | 48
    clinically septic | 72
    clear extension of necrotic tissue | 72
    right ear involved | 72
    left eye involved | 72
    family refused further surgical intervention | 72
    blood cultures negative | 72
    microscopic examination of tissue samples | 72
    invasive broad fungal hyphae yeast cells | 72
    acute and chronic inflammatory cells | 72
    necrotic tissue | 72
    suppurative microabscesses | 72
    confirmed clinical suspicion | 72
    extensive tissue debridement | 72
    antifungal therapy | 72
    rapid fungal invasion of the tissues | 72
    died | 96
    