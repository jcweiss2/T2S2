57 years old | 0
male | 0
recent dental work | -672
altered mental status | 0
urinary incontinence | 0
generalized weakness | 0
malaise | -336
fever | -336
emesis | -336
diarrhea | -336
computed tomography of the head | 0
intracranial hemorrhage | 0
dissection flap within the aortic arch | 0
transfer to Stanford Hospital | 0
CT angiography of the chest, abdomen, and pelvis | 0
Stanford Type A aortic dissection | 0
temperature 39.1°C | 0
heart rate 106 beats/min | 0
blood pressure 67/32 mm Hg | 0
SaO2 97% | 0
alert and oriented | 0
slow to respond | 0
right upper and lower extremity weakness | 0
increased WBC count | 0
thrombocytopenia | 0
anemia | 0
elevated BUN | 0
elevated creatinine | 0
elevated D-dimer | 0
coagulopathy | 0
disseminated intravascular coagulation | 0
sepsis | 0
vancomycin | 0
piperacillin-tazobactam | 0
blood cultures sent | 0
Gram stain showed Gram-positive cocci | 0
infective endocarditis | 0
neurocritical care consultation | 0
neurosurgery consultation | 0
bedside transthoracic echocardiography | 0
mobile mass in the left ventricular outflow tract | 0
subarachnoid hemorrhage | 0
no midline shift | 0
no elevated intracranial pressure | 0
international normalized ratio (INR) normalization | 0
platelet transfusion | 0
fresh frozen plasma transfusion | 0
packed red blood cells transfusion | 0
cryoprecipitate transfusion | 0
activated prothrombin complex concentrate | 0
cardiopulmonary bypass | 0
surgical repair of Type A aortic dissection | 0
aortic valve replacement | 0
bioprosthetic aortic valve | 0
composite-valve-graft | 0
hemi-arch replacement | 0
dissection flap extending into the aneurysmal root | 0
purulent thrombus within the false lumen | 0
vegetation on the aortic valve | 0
Streptococcus equi (S. equi) | 0
bacteremia | 0
endocarditis | 0
penicillin | 0
intravenous penicillin | 0
postoperative day (POD) 1 | 24
spontaneous movement of all extremities | 24
stable SAH | 24
extubation | 48
transfer to the ward | 192
mentation improvement | 720
dysarthria improvement | 720
mild word-finding difficulty | 720
mobility improvement | 720
platelet normalization | 720
discharge to rehabilitation facility | 720
peripherally inserted central catheter placement | 720
penicillin G | 720
readmission for pleuritic chest pain | 2880
contrast extravasation within a perigraft fluid collection | 2880
redo sternotomy | 2880
replacement of aortic and mitral valves | 2880
dehiscence of the aorto-mitral curtain | 2880
recurrent endocarditis | 2880
lifelong amoxicillin-clavulanate | 3000
follow-up appointment | 4032