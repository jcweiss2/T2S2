50 years old | 0
male | 0
presented with L5 nerve root radiculopathy | 0
nonsteroidal anti-inflammatory drugs | 0
physiotherapy | 0
epidural administration of 80 mg of methylprednisolone | 0
severe pain in both lower limbs | 0
pruritus | 0
severe cramps | 0
profuse sweating | 0
progressive weakness of both lower limbs | 0
complete flaccid paraplegia below T11 level | 0
absent reflexes below T11 | 0
blood pressure 210/110 mmHg | 0
heart rate 124 beats per minute | 0
shifted to medicine emergency | 0
labetalol given | 0
refractory blood pressure | 0
continued sweating | 0
continued agitation | 0
electrocardiography showing hyperkalemia | 0
tachycardia | 0
absent P-wave | 0
tall T-wave | 0
accidental use of 15% KCl instead of NS | 0
shifted to Intensive Care Unit | 0
supportive measures | 0
calcium gluconate | 0
raised potassium levels (7 mg/dL) | 0
potassium chelating agent (Ksylate) | 0
blood pressure normal | 120
heart rate normal | 120
return of sensory modalities | 360
spasticity | 360
exaggeration of deep tendon reflexes | 360
extensor plantar reflex | 360
neurologically normal | 480
discharged from Intensive Care Unit | 576
