22 years old | 0
White | 0
G2P1001 | 0
admitted to the hospital | 0
cerebrovascular accident tenderness | 0
malaise | 0
polysubstance abuse | -8760
MSSA bacteremia | -8760
hepatitis C virus | -8760
endocarditis | -8760
IV antibiotics | -8760
COVID-19 pneumonia | 0
pyelonephritis | 0
MSSA bacteremia | 0
thrombocytopenia | 0
respiratory failure | 0
intubated | 0
transesophageal echocardiogram | 0
severe TV regurgitation | 0
large TV vegetations | 0
flail TV leaflets | 0
severe valve malcoaptation | 0
betamethasone | 0
fetal lung maturation | 0
transferred to a tertiary care hospital | 0
cardiothoracic surgery team recommended medical management | 0
IV antibiotics | 0
valve surgery after delivery | 0
extubated | 0
transferred to the MFM unit | 48
Subutex initiation | 48
continuation of IV antibiotics | 48
ID team recommended continuation of IV cefazolin | 48
tachypneic | 168
tachycardic | 168
increasing oxygen supplementation | 168
computed tomography angiogram | 168
septic emboli | 168
pericardial effusion | 168
multidisciplinary discussion | 168
AngioVac procedure recommended | 168
counseled on the risks of the AngioVac procedure | 168
informed consent | 168
preprocedure echocardiogram | 216
ejection fraction of 60% | 216
moderate TV regurgitation | 216
mobile vegetation on the TV | 216
AngioVac procedure performed | 216
general anesthesia | 216
continuous fetal monitoring | 216
obstetrician present | 216
NICU on standby | 216
Foley catheter | 216
external fetal heart monitor | 216
access obtained to both the femoral veins and the right internal jugular vein | 216
intracardiac echocardiogram | 216
vegetations on both the posterior and anterior leaflets of the TV | 216
eustachian valve | 216
AngioVac cannula introduced | 216
venous bypass circuit activated | 216
multiple passes made | 216
vegetations debulked | 216
vegetations grew S aureus | 216
postoperative echocardiogram | 216
ejection fraction of 57% | 216
mobile vegetations on the TV | 216
flail TV | 216
severe TV regurgitation | 216
clinical status improved | 216
blood cultures negative | 504
nonreassuring fetal heart tracing | 504
cesarean delivery | 504
live-born male infant | 504
Apgar scores of 9 and 9 | 504
placental pathology | 504
perivillous fibrin deposition | 504
calcification | 504
neonate admitted to the NICU | 504
respiratory distress syndrome | 504
prematurity | 504
neonate discharged on day 35 of life | 1008
preeclampsia with severe features | 504
magnesium | 504
long-acting nifedipine | 504
postpartum course complicated | 504
repeat echocardiogram | 672
severe TV regurgitation | 672
TV vegetations | 672
flail leaflet | 672
Chiari network | 672
dilated right atrium | 672
normal ventricular function | 672
patent foramen ovale | 672
blood cultures showed no growth | 672
TV replacement with a porcine valve | 672
primary closure of the patent foramen ovale | 672
antibiotics course completed | 1008
discharged on postpartum day 24 | 1008