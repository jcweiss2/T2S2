25 years old | 0
    female | 0
    nausea | -120
    vomiting | -120
    dizziness | -120
    abdominal pain | -120
    altered sensorium | -120
    weighing 55 kg | 0
    ingestion of two bottles (refills) of mosquito repellent | -120
    each refill containing 45 ml (396 mg) transfluthrin | -120
    conscious | 0
    semi constricted pupils | 0
    sluggishly reactive pupils | 0
    crepitations in lungs | 0
    respiratory rate 28/min | 0
    blood pressure 110/70 mmHg | 0
    gastric lavage | 0
    continuous gastric aspiration | 0
    oral syrup charcoal 10 ml | 0
    Ryles tube closed | 0
    aspiration through Ryles tube continued | 0
    atropine 0.6 mg | 0
    pantoprazole 40 mg | 0
    ondansetron 4 mg | 0
    tonic-clonic convulsions | 60
    phenytoin 700 mg bolus | 60
    diazepam 10 mg | 60
    hydrocortisone 100 mg | 60
    frusemide 20 mg | 60
    oxygen enrichment | 60
    uncontrolled convulsions | 60
    shifted to intensive care unit | 60
    midazolam 5 mg | 60
    propofol 100 mg | 60
    endotracheal intubation | 60
    cuff inflated | 60
    oxygen enrichment 4–6 L/min | 60
    midazolam 4 mg/h infusion | 60
    propofol 200 mg/h infusion | 60
    SpO2 100% | 60
    blood pressure 94/62 mmHg | 60
    pulse rate 74/min | 60
    ABG normal | 60
    IV mannitol (20%)100 ml twice a day | 60
    IV phenobarbitone (SOS) | 60
    seizure free for few hours | 60
    seizures restarted | 60
    blood pressure 80/40 mmHg | 60
    respiratory rate 35/min | 60
    pulse rate 190/min | 60
    SpO2 95% | 60
    serum potassium 2.98 mmol/L | 60
    serum calcium 2.5 mmol/L | 60
    serum sodium 129 mmol/L | 60
    dopamine 10 μg/kg/min | 60
    potassium chloride 1.5 g | 60
    hypertonic saline | 60
    uncontrolled seizures | 60
    elective ventilation planned | 60
    vecuronium 4 mg bolus | 60
    vecuronium 4 mg/h infusion | 60
    controlled mechanical ventilation | 60
    blood pressure decreased | 60
    dopamine dose increased | 60
    propofol infusion stopped | 60
    ABG normal | 60
    computed tomography scan normal | 60
    chest X-ray normal | 60
    input/output charting | 60
    central venous pressure 5-8 cm H2O | 60
    ventilator for 48 hours | 60
    weaning started | 108
    vecuronium infusion stopped | 108
    midazolam infusion stopped | 108
    SIMV mode | 108
    airway pressure support 15 cm H2O | 108
    PEEP 4 cm H2O | 108
    pulse rate 102/min | 108
    blood pressure 132/82 mmHg | 108
    SpO2 96% | 108
    total leucocyte count 7200/mm³ | 24
    leucocyte count 22,000/mm³ | 48
    leucocyte count 32,000/mm³ | 72
    leucocyte count 13,000/mm³ | 96
    neutrophilia | 24
    antibiotics continued | 24
    leucocyte count 4000/mm³ | 144
    dopamine infusion tapered | 108
    dopamine stopped | 114
    spontaneous respiration 16 breaths/min | 114
    neostigmine 2.5 mg | 114
    glycopyrrolate 0.4 mg | 114
    spontaneous breathing | 114
    adequate tidal excursion | 114
    followed verbal commands | 114
    extubated | 114
    oxygen mask 4–5 L/min | 114
    respiratory rate 25/min | 114
    blood pressure 108/72 mmHg | 114
    pulse rate 119/min | 114
    pupils reactive to light | 114
    nebulised with mistabron 3 mg | 114
    referred to psychiatrist | 114
    shifted to ward | 96
    discharged | 168
    