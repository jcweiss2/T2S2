45 years old | 0
    male | 0
    admitted to the hospital | 0
    hepatic echinococcosis | -105216
    right abdominal distension pain | -105216
    pulmonary echinococcosis | -87600
    surgery | -87600
    pulmonary hypertension | 0
    filling defects of the pulmonary artery | 0
    peripheral blood cells normal | 0
    bilirubin normal | 0
    prescribed enoxaparin | 0
    prescribed torsemide | 0
    prescribed spironolactone | 0
    prescribed albendazole | 48
    prescribed praziquantel | 192
    increased bilirubin | 168
    severe myelosuppression | 432
    WBC 1.35 | 432
    NEUT 0.73 | 432
    Hgb 97 | 432
    febrile | 432
    diarrhea | 432
    stomachache | 432
    severe hair loss | 432
    WBC 0.46 | 456
    NEUT 0.13 | 456
    Hgb 88 | 456
    stopped albendazole | 456
    stopped praziquantel | 456
    treated with parenteral nutrition | 456
    treated with omeprazole | 456
    treated with glutathione | 456
    treated with meropenem | 456
    treated with granulocyte colony-stimulating factor | 456
    gastrointestinal tract reaction recovered gradually | 528
    WBC 0.86 | 528
    NEUT 0.25 | 528
    PLT 78 | 528
    Hgb 92 | 528
    very high risk for severe infection | 528
    blood count began to increase slowly | 672
    discharged | 672
    