27 years old | 0
female | 0
Mayer Rokitansky Syndrome | -0
Mullerian agenesis | -0
sigmoid neovaginoplasty | -6480
lower abdominal pain | 0
bilateral pelvic pain | 0
denied routinely irrigating or dilating her neovagina | 0
penetrative sexual intercourse | 0
CT imaging of the abdomen | 0
tubular, heterogenous, fluid-filled structure | 0
blind ending | 0
abdominal pain acutely worsened | 24
diaphoresis | 24
significant distress due to pain | 24
leukocytosis | 24
absolute neutrophils | 24
increasing inflammatory process | 24
empiric intravenous piperacillin-tazobactam | 24
transferred emergently to our children’s hospital | 24
hypotensive | 24
tachycardic | 24
afebrile | 24
tachypneic | 24
oxygen saturation | 24
IV fluid boluses | 24
antimicrobials were empirically changed | 24
exploratory laparotomy | 24
cystoscopy | 24
vaginoscopy | 24
normal bladder | 24
urethra | 24
obliterated introitus | 24
diffuse intra-abdominal spillage | 24
mucus | 24
perforated sigmoid neovagina | 24
purulent fluid | 24
intrabdominal drains | 24
intubated | 24
mechanical ventilation | 24
septic shock | 24
vasopressor agents | 24
antimicrobials were transitioned | 24
preliminary peritoneal culture | 24
gram-negative rods | 24
blood cultures | 24
peritoneal cultures | 24
Bacterioides thetaioaomicron | 24
Bacteroides caccae | 24
Actinomyces species | 24
weaned off vasopressors | 192
extubated | 192
transferred to the general floor | 288
Infectious Diseases team | 288
antimicrobial management | 288
susceptibilities | 288
discharged home | 360
abdominal wound vacuum | 360
IV piperacillin-tazobactam | 360
generalized malaise | 432
diffuse abdominal pain | 432
readmitted | 432
sepsis | 432
white blood count | 432
absolute neutrophil count | 432
d-dimer | 432
lactate | 432
CT of the chest | 432
abdomen | 432
pelvis | 432
bilateral pleural effusions | 432
loculated left pleural effusion | 432
multiple new abdominal abscesses | 432
transcutaneous drainage catheter | 432
open anterior midline wound | 432
wound vacuum | 432
hypoxemia | 432
transferred to the intensive care unit | 432
IV piperacillin-tazobactam | 432
placement of a right perihepatic drain | 432
aspiration of purulence | 432
unsuccessful drainage | 432
peri-splenic collection | 432
interventional radiology | 432
drained fluid | 432
right perinephric abscess | 432
perisplenic abscess | 432
Broad-spectrum PCR | 432
improved clinically | 768
antimicrobials were narrowed | 768
IV ampicillin-sulbactam | 768
discharge | 768
Broad spectrum PCR | 768
Gleimia europaea | 768
Alistipes onderdonkil | 768
Varibaculum timonense | 768
Jonquetella anthropi | 768
followed up | 1056
adult infectious diseases clinic | 1056
continued on ampicillin-sulbactam | 1056
plans to reimage | 1056
clinically improved | 1056
repeat CT abdomen | 1056
decreased in the size | 1056
right and left sub-phrenic abscesses | 1056
transitioned from IV ampicillin-sulbactam | 1056
oral amoxicillin-clavulanate | 1056