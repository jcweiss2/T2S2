35 years old | 0
gravida 3 | 0
para 1–0-1–1 | 0
admitted to the hospital | 0
diagnosis of early midtrimester oligohydramnios | -98
routine anatomical survey ultrasound examination | -98
18 weeks of gestation | -98
preterm prelabor rupture of membranes | -98
pooling of amniotic fluid in posterior vaginal fornix | -98
arborization ferring testing | -98
nitrazine testing | -98
evaluation for preterm prelabor rupture of membranes | -98
intra-amniotic dye infusion testing | -98
declined intra-amniotic dye infusion testing | -98
ultrasound at 20 6/7 weeks of gestation | -56
single live fetus | -56
amniotic fluid index of 2.8 cm | -56
membrane separation | -56
possible membrane rupture distal to the cervical opening | -56
high amniotic leak | -56
fetal kidneys and bladder seen on ultrasound | -56
normal fetal kidneys and bladder | -56
history of gestational diabetes | 0
history of loop electrical excision procedure | 0
herpes simplex type 2 | 0
maternal obesity | 0
prepregnancy body mass index 34 kg/m2 | 0
episode of domestic violence | 0
early genetic screening with cell free fetal DNA | -56
appropriate fetal fraction | -56
sex chromosomes XY | -56
low risk for trisomy 13, 18, and 21 | -56
second trimester maternal serum α-fetoprotein | -56
2.16 MoM | -56
prenatal counseling with neonatology and maternal-fetal medicine | -28
wishes for full neonatal resuscitation at 22 weeks | -28
understanding of the prognosis | -28
amnioinfusion and intra-amniotic dye instillation testing | -14
counseling | -14
amnioinfusion | -14
intra-amniotic dye installation | -14
22-gauge-needle inserted into the intra-amniotic cavity | -14
15 mL of clear yellow fluid removed | -14
genetic and infection testing | -14
40 mL of warmed 0.9% sodium chloride solution containing 1,000 mg/L oxacillin infused | -14
5 mL of indigo carmine added | -14
intra-amniotic dye instillation test | -14
400 mL of warmed 0.9% sodium chloride solution containing 1,000 mg/L oxacillin infused | -14
ambulated for 30 minutes | -14
tampon testing confirmed rupture of fetal membranes | -14
admitted to the hospital for latency antibiotics and serial intra-amniotic infusions | 0
acyclovir prophylaxis started | 0
no active herpes lesions seen | 0
7-day-course of latency antibiotics consisting of ampicillin and azithromycin | 0
completed 7-day-course of latency antibiotics | 7
betamethasone administered at 23 weeks of gestation | 7
second amnioinfusion | 14
800 mL of warmed 0.9% sodium chloride solution containing 1,000 mg/L oxacillin infused | 14
normal maximum vertical pocket | 14
plan for serial intra-amniotic infusions until 26 weeks of gestation | 14
denied continued leakage of fluid | 21
MVP was normal | 21
amnion resealed | 21
decision to cease further intra-amniotic infusions | 21
amniotic fluid testing returned with no evidence of intra-amniotic infection | 21
genetic testing with karyotype and microarray confirmed no genetic abnormalities in the fetus | 21
gestational hypertension without clinical or laboratory evidence for preeclampsia | 28
expectantly managed in the hospital | 28
fetal status remained reassuring | 28
appropriate fetal growth on serial ultrasounds | 28
MVP remained normal for the duration of her pregnancy | 28
second course of betamethasone | 49
external cephalic version performed at 34 weeks | 49
breech presentation | 49
induction of labor at 34 2/7 weeks | 56
penicillin in labor for group B streptococcus prophylaxis | 56
delivered a vigorous male infant | 56
birth weight of 2,160 g | 56
Apgar's scores of 9 at 1 and 5 minutes of life | 56
placenta weighed 390 g | 56
evidence of moderate acute inflammation at the chorion | 56
no evidence of inflammation elsewhere on the amnion or umbilical cord | 56
newborn's initial white blood cell count was 11.7 × 1,000 μL | 56
ampicillin and gentamycin for 48 hours | 56
negative blood cultures | 58
newborn stayed in the hospital for 9 days | 65
no immediate complications | 65