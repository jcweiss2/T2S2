diagnosed with papillary thyroid carcinoma | -9720
treated by resection and radiotherapy | -9720
developed a stenosis of the esophagus | -8760
repeated aspiration led to several episodes of respiratory insufficiency due to pneumonia and purulent pleurisy | -8760
treated by pleurectomy | -8760
developed a restrictive ventilation pattern and a recurrent nerve palsy | -8760
treated by percutaneous endoscopic gastrostomy and tracheostoma | -8760
put on home ventilation | -8760
mobility decreased | -8760
developed secondary depression | -8760
stopped talking | -8760
mandible was nearly fixed | -8760
could not open her mouth over a maximum of 20 degrees | -8760
left axis vertebralis was stented | -4380
developed stenosis of the internal axis carotis on both sides | -4380
diagnosed with arterial hypertension and secondary lactase deficiency | -4380
esophageal stenosis was dilated | -120
referred to the University of Erlangen due to a decreasing general condition | 0
fistula between the esophagus and tracheal membrane had occurred | 0
examined by several chiefs and consultants | 0
deemed too unstable for open surgery | 0
inability to open the mouth and the recurrent nerve palsy | 0
referred to our hospital on the surgical intensive care unit | 15
suffering from pneumonia by 4-multiresistente gramnegative Pseudomonas aeruginosa in the right lung | 15
put on veno-venous extracorporeal membrane oxygenation (vv-ECMO) | 15
thoracic computed tomography confirmed a big fistula of the tracheal membrane | 16
decision to try endobronchial stenting was made | 16
procedure was performed | 17
vv-ECMO began to be partly ineffective due to rising septical issues | 17
high volume input of physiological saline was needed | 17
oral approach would only allow a small flexible bronchoscope | 17
approach for the upper part of the trachea had to be performed through the percutaneous tracheostoma in a retrograde manner | 17
trying different Dumon and one-hybrid self expandable metalic y-stent | 17
plan was to changeover to a more floppy Freitag stent (FS) | 17
successful retrograde stenting was performed in four steps | 17
Step I: manually compressed “y” of the FS was successfully pushed downward on the main carina | 17
Step II: frontal surface of the stent was cut with at least 1 cm opening in the longitudinal axis | 17
Step III: jagwire was introduced through the mouth into the trachea | 17
Step IV: regular tracheal cannula was introduced for ventilation | 17
lungs were not aerated at that point of time | 17
spontaneous breathing work increased and the vv-ECMO support was reduced | 120
lungs became re-aerated again | 120
patient woke up again and could communicate with her family by writing and her eyes | 120
infections continued to be very severe | 120
spontaneous work of breathing never exceeded a tidal ventilation of 170 mL per breath | 120
reduction of intravenous saline injection was limited | 120
patient along with her family decided actively to reduce the vv-ECMO support | 360
patient died on 18 November 2016 due to pulmonary infection | 420