68 years old | 0
female | 0
admitted to the hospital | 0
diagnosed with AML | -30
FLT3-itd positive | -30
normal karyotype | -30
full blood count | -30
pancytopenia | -30
blast count of 30% | -30
DA-chemotherapy | -20
refractory to DA-chemotherapy | -20
FLAG-IDA | -18
complete remission | -16
2nd course of FLAG-IDA | -14
HLA-mismatched allogeneic transplant | 0
Fludarabine/Busulphan/Alemtuzumab | 0
Enterobacter and E.coli bacteremias | 0
treated with meropenem | 0
neutrophil engraftment | 18
platelet engraftment | 20
discharged | 26
febrile episode | 26
mild skin graft versus host disease | 42
topical steroids | 42
clostridium difficile diarrhea | 60
oral vancomycin | 60
3-month bone marrow aspirate | 90
100% donor chimerism | 90
99% donor chimerism in CD3+ T cells | 90
ciclosporin tapered | 120
ongoing diarrhea | 120
flexible sigmoidoscopy | 150
inflammation | 150
no gut GVHD | 150
ciclosporin stopped | 210
mild chronic skin GVHD | 365
vaccination program | 365
relapse | 540
reduction in neutrophil count | 540
viral screen | 540
bone marrow arranged | 540
relapsed disease | 540
20% blasts detected | 540
mixed chimerism | 540
48% donor in whole sample | 540
92% donor in CD3+ T cells | 540
azacitadine | 540
donor lymphocyte infusion | 560
access to AC220 and Crenolanib | 560
compassionate access declined | 560
1st cycle of azacitadine | 560
2nd cycle of azacitadine | 570
1st DLI | 580
red cell and platelet transfusion | 580
cycles 3 and 4 azacitadine | 600
2nd DLI | 620
3rd DLI | 660
gastrointestinal symptoms | 720
azacitadine dose reduced | 720
9th cycle of azacitadine | 730
gram-negative sepsis | 740
E.coli | 740
intensive care admission | 740
inotropic support | 740
recovered | 750
bone marrow aspirate | 780
complete morphological remission | 780
FLT3-itd negativity | 780
no further treatment | 780
monthly monitoring | 780
100% donor chimerism | 960
100% donor chimerism in CD3+ T cells | 960
100% donor chimerism | 1200
100% donor chimerism in CD3+ T cells | 1200