25 years old | 0
female | 0
transferred to the Emergency Department | 0
head-on motor vehicle collision | -72
located in the center rear passenger seat | -72
single transverse band seat belt | -72
hemodynamically stable | 0
patent airway | 0
Glasgow Coma Scale of 15 | 0
Focused Abdominal Sonography for Trauma (FAST) scan | 0
small amount of perisplenic and pelvic fluid | 0
no solid organ injury | 0
no pneumoperitoneum | 0
computerized tomography | 0
lower left rib fractures (7th–11th) | 0
compression fractures with anterior wedging of L1 and L2 | 0
transverse process fracture of the same vertebra levels | 0
managed conservatively | 0
admitted to the Intensive Care Unit (ICU) | 0
acutely hemodynamically unstable | 72
physical examination findings concerning for an acute abdomen | 72
repeat FAST scan | 72
increase in free intraperitoneal fluid | 72
septic shock | 72
taken back to the operative theater | 72
retroperitoneal hematoma in bilateral Zone II | 72
steatonecrosis plaques throughout the peritoneal cavity | 72
incomplete jejunal laceration 40 cm from the Treitz angle | 72
complete section of the pancreas at the body-tail level | 72
peripancreatic hematoma | 72
necrohemorrhagic pancreatitis | 72
distal pancreatectomy | 72
splenectomy | 72
jejunal enterorraphy | 72
open abdomen | 72
catastrophic abdomen | 72
numerous complex enterocutaneous fistulas | 72
open abdomen management | 72
~40 interventions performed | 72
negative pressure systems not available | 72
aspiration probes | 72
placement of Goretex™ mesh | 72
linitud films | 72
progressed favorably | 72
multiple established enterocutaneous fistulas | 72
short-gut syndrome | 72
discharged with home parenteral nutrition | 2880
3 months in the ICU | 2880
4 months of admission in the ward | 2880
strategy of abdominal reconstruction | 8760
elective surgery | 8760
re-establish the intestinal transit | 8760
study to identify the different fistulous openings | 8760
reconstruction of the abdominal wall | 8760
Plastic Surgery Service support | 8760
en bloc excision of the midlaparotomy scar | 8760
subtotal colectomy up to the descending-sigmoid junction | 8760
resection of the intestinal ileostomy | 8760
excision of three segments of the small intestine | 8760
reconstruction of the intestinal transit | 8760
four anastomoses | 8760
three mechanical latero-lateral entero4-enteric anastomosis | 8760
mechanical lateral-lateral ileosigmoid anastomosis | 8760
repair of the abdominal wall | 8760
permacol mesh plasty | 8760
wide skin flap | 8760
discharged on Day 16 | 8760
follow-up control for 12 years | 105120
no incidents to date | 105120
