68 years old | 0
woman | 0
admitted to the hospital | 0
laparoscopic tension-free hernioplasty | 0
incisional hernia | 0
repair of sigmoid perforation | -672
platelet count 224.1×109/L | -672
postoperative day 4 | -96
low platelet count 70.8×109/L | -96
test tubes containing EDTA | -96
erythrocyte counts obtained on automated analyzer | -96
disease progressed | -96
sudden development of shortness of breath | -96
chest tightness | -96
dizziness | -96
abdominal distension | -96
nausea | -96
laboratory investigation | -96
low platelet count 36.9×109/L | -96
low white blood cell count 3.32×109/L | -96
culture from purulent secretion | -96
growth of Escherichia coli | -96
serum endotoxin 54.51 pg/mL | -96
sepsis | -96
abdominal computed tomography scan | -96
extensive gas-fluid levels in intestinal tract | -96
intestinal wall swelling | -96
acute intestinal obstruction | -96
exploratory laparotomy | -96
intra-abdominal infections | -96
arterial blood gas analyses | -96
PaO2 51 mmHg | -96
PaCO2 45 mmHg | -96
respiratory failure | -96
transferred to intensive care unit | 144
postoperative day 6 | 144
fresh-frozen plasma | 144
platelet transfusions | 144
teicoplanin | 144
ornidazole | 144
imipenem | 144
cilastatin sodium | 144
failure to respond to platelet transfusions | 144
postoperative day 10 | 240
blood collected with EDTA | 240
blood collected with sodium citrate | 240
platelet count 7.20×109/L (EDTA) | 240
platelet count 136.00×109/L (sodium citrate) | 240
platelet clumps identified by microscopic examination | 240
pseudothrombocytopenia | 240
resolution of infection | 240
EDTA-PTCP disappeared | 240
