56 years old | 0
female | 0
admitted to the hospital | 0
high-grade fever | -48
shortness of breath | -48
hypotensive | 0
tachycardic | 0
tachypneic | 0
mottled cold extremities | 0
multilobar pneumonia | 0
intubated | 0
transferred to the medical Intensive care unit | 0
IV norepinephrine | 0
IV vasopressin | 0
IV dopamine | 0
haemodynamic support | 0
blood cultures | 0
IV vancomycin | 0
IV ceftriaxone | 0
IV azithromycin | 0
prothrombin time prolonged | 0
partial thromboplastin time prolonged | 0
fibrin degradation products elevated | 0
disseminated intravascular coagulopathy | 0
urine Streptococcus pneumonia antigen positive | 0
blood cultures grew Streptococcus pneumoniae | 0
diffuse petechial rash | 24
non-blanching purpuric ecchymotic skin lesions | 24
flaccid bullae | 48
extensive skin sloughing | 72
skin biopsy | 72
non-inflammatory vascular occlusion | 72
skin necrosis | 72
purpura fulminans | 72
broad-spectrum antibiotics | 0
heparin drip | 0
blood products | 0
hyperbaric oxygen therapy | 72
anuric renal failure | 120
haemodialysis | 120
bedside incisional fasciotomy | 120
no muscle necrosis | 120
no compartment syndrome | 120
transferred to the burns unit | 168
comfort measures only | 240
dismal prognosis | 240
no meaningful recovery | 240