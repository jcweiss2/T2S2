34 years old | 0
male | 0
admitted to the hospital | 0
hematemesis | -96
dyspnea | -96
hemoptysis | -96
fever | -96
tachycardia | 0
blood pressure 100/58 mmHg | 0
tachypnea | 0
diaphoresis | 0
Glasgow scale 15 | 0
pulse oximetry 70% | 0
rales in the left base | 0
hemorrhagic pangastritis | 0
moderate duodenitis | 0
sparse mucosal bleeding | 0
diffuse and bilateral reticulo-nodular pattern | 0
HIV serology positive | 0
viral load >500,000 copies | 0
CD4 count 58 cells/mm3 | 0
increased WBC count | 0
leukocytes 20.4 × 103/mm3 | 0
myelocytes 1% | 0
metamyelocytes 3% | 0
rods 34% | 0
eosinophils 0% | 0
basophils 0% | 0
lymphocytes 2% | 0
monocytes 7% | 0
platelets 283 × 103/mm3 | 0
AST 79 U/L | 0
ALT 84 U/L | 0
LDH 405 U/L | 0
amylase 106 U/L | 0
albumin 3.1 g/dL | 0
lactate 7.4 mg/dL | 0
CRP 140 mg/L | 0
empirical antimicrobial therapy | 0
trimethoprim-sulfamethoxazole | 0
ceftriaxone | 0
clarithromycin | 0
prednisone | 0
petechiae | 72
bronchoscopy | 72
refractory shock | 76
fever 41.9 °C | 76
cardiac arrest | 76
death | 76
autopsy | 76
mild meningeal inflammatory infiltrate | 76
filariform larva of Strongyloides stercoralis | 76
intra-alveolar hemorrhage | 76
diffuse alveolar damage | 76
hyaline membrane | 76
healing process | 76
fragments of Strongyloides stercoralis larvae | 76
eggs of Schistosoma mansoni | 76
ischemic areas of the centrilobular zone III | 76
microvesicular steatosis | 76
infective larvae of S. stercoralis | 76
eggs of S. mansoni | 76
granuloma | 76
hemorrhagic gastritis | 76
adult females of S. stercoralis | 76
hemorrhagic enteritis | 76
mucosal necrosis | 76
larvae of S. stercoralis | 76
eggs of S. mansoni | 76
calcified eggs of S. mansoni | 76
adult worms of S. mansoni | 76
generalized visceral congestion | 76
reactive bone marrow | 76