62 years old | 0
male | 0
COPD Gold II | 0
Hashimoto's disease | 0
admitted to the hospital | 0
shortness of breath | -240
coughing | -240
fever | -240
myalgia | -240
tested positive for SARS-CoV-2 | -168
treatment with remdesivir | 0
treatment with dexamethasone | 0
treatment with high-dose prophylactic low molecular weight heparin | 0
severe hypoxia | 0
high-flow nasal cannula support | 0
increased events of paroxysmal hypoxia | 192
chest pain | 192
stable macrocirculation | 192
mono-organ failure | 192
SOFA score of 2 | 192
electrocardiogram showed no abnormalities | 192
cardiac markers showed no abnormalities | 192
echocardiography showed no abnormalities | 192
increased D-dimer | 192
CTPA showed large vessel thrombosis | 192
thrombosis of pulmonary arteries | 192
thrombosis of thoracic aorta | 192
renal infarction | 192
spleen infarction | 192
sublingual microcirculation measurements | 192
hyperdynamic circulation | 192
increased total vessel density | 192
increased functional capillary density | 192
increased proportion of perfused vessels | 192
increased red blood cell velocity | 192
treatment with continuous high molecular weight heparin infusion | 198
respiratory status deteriorated | 216
mechanical ventilation | 216
Staphylococcus Aureus pneumosepsis | 504
progressive multi-organ failure | 504
death | 504