46 years old | 0
female | 0
admitted to the emergency ward | 0
severe trauma | 0
collapse of a brick kiln | 0
burns (II°, 18% TBSA) | 0
multiple lacerations (scalp, right canthus, right eyelid) | 0
acute traumatic craniocerebral injury | 0
superficial skin contusion (right zygomatic, left frontal) | 0
multiple fractures (right sacral promontory, bilateral superior pubic ramus, right inferior pubic ramus, right 1–5th rib) | 0
debridement | 0
analgesics | 0
anti-infection (levofloxacin 0.4 QD + cefazolin 1.0 Q12H, I.V.) | 0
hemostasis | 0
tetanus prevention | 0
wound exposure | 0
rehydration | 0
blood pressure drop to 85/50mmHg | 24
HGB 104g/L | 24
hemorrhagic shock | 24
transferred to ICU | 24
enhanced dilatation | 24
anti-infection (ceftazidime 1.0 Q8H + levofloxacin 0.4 QD, I.V.) | 24
analgesia | 24
nutritional support | 24
single room isolation | 24
appropriate braking | 24
wound disinfection | 24
external application of burn cream | 24
exposure treatments | 24
intermittent moderate fever (38.2°C) | 24
wound exudation | 24
blood culture (aerobic and anaerobic) | 168
WBC 3.75×109/L | 168
CRP 145 mg/L | 168
PCT 0.81 ng/mL | 168
first blood culture positive for Pandoraea species | 264
in vitro susceptibility testing | 264
body temperature 38.9°C | 288
second blood culture | 288
WBC 4.21×109/L | 288
CRP 93.7 mg/L | 288
PCT 0.74 ng/mL | 288
CT scan (chest and abdomen) | 288
anti-infection changed to imipenem 1.0 Q8H + tigecycline 50 mg Q12H I.V. | 312
second blood culture positive for Pandoraea species | 384
wound secretion culture | 432
Staphylococcus epidermidis | 432
Candida parapsilosis | 432
16S rRNA sequencing confirmed Pandoraea sputorum | 432
MALDI-TOF MS confirmed Pandoraea sputorum | 432
no bacteria in blood on days 17 and 23 | 408, 552
normal body temperature | 336
CRP 6.0mg/L | 336
PCT 0.11ng/mL | 336
scanty wound exudation | 336
shifted to Burn and Plastic Surgery | 336
discharged | 1440
wounds healed | 1440
fractures healed | 1440
