60 years old | 0
female | 0
elective percutaneous nephrolithotomy | 0
pre-diabetes | -672
chronic obstructive pulmonary disease | -672
morbid obesity | -672
obstructive sleep apnea | -672
heart failure with preserved ejection fraction | -672
febrile | 24
tachycardic | 24
leukocytosis | 24
vancomycin | 24
piperacillin/tazobactam | 24
meropenem | 24
respiratory distress | 24
hypoxemia | 24
non-invasive positive pressure ventilation | 24
endotracheal intubation | 48
lung protective ventilation | 48
bilateral pulmonary ground glass opacities | 48
infectious process | 48
acute respiratory distress syndrome | 48
pulmonary edema | 48
pulmonary embolism | 48
normal ejection fraction | 48
ventricular size | 48
paralysis | 48
ventilator desynchrony | 48
refractory hypoxemia | 48
bronchoalveolar lavage | 120
nasopharyngeal swab | 120
rhinovirus pneumonia | 120
antibiotics discontinued | 120
no antivirals | 120
high airway pressures | 120
peak inspiratory pressure | 120
positive end-expiratory pressure | 120
FiO2 | 120
PaO2 to FiO2 ratio | 120
moderate to severe ARDS | 120
LPV strategy | 120
APRV | 144
mechanical ventilation settings adjusted | 144
PHigh | 144
PLow | 144
expiratory duration adjusted | 144
TLow | 144
peak expiratory flow rate | 144
weaned to extubation | 216
diuresis | 216
discharged home | 312