65 years old | 0
    male | 0
    admitted to the hospital | 0
    non-ischaemic cardiomyopathy | 0
    left ventricular ejection fraction 20% | 0
    guideline-directed medical therapy | 0
    bisoprolol 5 mg PO o.d. | 0
    candesartan 4 mg PO o.d. | 0
    primary prevention implantable cardioverter-defibrillator | 0
    New York Heart Association class II | -120
    paroxysmal atrial fibrillation | 0
    treated with apixaban | 0
    previous cerebrovascular accident | 0
    hypertension | 0
    dyslipidaemia | 0
    depression | 0
    presented with persistent epigastric abdominal pain | 0
    presented with fatigue | 0
    blood pressure 112/81 mmHg | 0
    heart rate 70 b.p.m. | 0
    respiratory rate 18 breaths per minute | 0
    jugular venous pressure 5–6 cm | 0
    peripheral oedema 1+ | 0
    lactate 5.6 mmol/L | 0
    creatinine 125 µmol/L | 0
    eGFR 60 mL/min/1.73 m2 | 0
    alanine transaminase 174 IU/L | 0
    transthoracic echocardiography | 0
    left ventricular function 11% | 0
    mild right ventricular dysfunction | 0
    intravenous furosemide infusion | 0
    home medications held | 0
    bisoprolol held | 0
    candesartan held | 0
    acute kidney injury | 192
    creatinine 176 µmol/L | 192
    eGFR 41 mL/min/1.73 m2 | 192
    alanine transaminase 350 IU/L | 192
    aspartate transaminase 913 IU/L | 192
    international normalized ratio 4.4 | 192
    lactate normalized to 1.7 mmol/L | 192
    heart rate 86 b.p.m. | 192
    blood pressure 103/66 mmHg | 192
    started bisoprolol 2.5 mg PO o.d. | 192
    started sacubitril/valsartan 24/26 mg PO b.i.d. | 192
    developed progressive shock | 216
    creatinine 476 µmol/L | 216
    eGFR 12 mL/min/1.73 m2 | 216
    hypotension | 216
    norepinephrine 0.28 µg/kg/min | 216
    dobutamine 18.7 µg/kg/min | 216
    transferred to tertiary academic centre | 240
    right heart catheterization | 240
    pulmonary capillary wedge pressure 24 mmHg | 240
    cardiac index 5.7 L/min/m2 | 240
    systemic vascular resistance 297 dyne/s/cm5 | 240
    diagnosed vasoplegic shock secondary to sacubitril/valsartan | 240
    sepsis ruled out | 240
    adrenal insufficiency ruled out | 240
    fulminant liver failure ruled out | 240
    neurogenic cause ruled out | 240
    vasoplegic shock resolved | 336
    creatinine normalized to 95 µmol/L | 336
    eGFR 84 mL/min/1.73 m2 | 336
    norepinephrine weaned off | 336
    right heart catheterization shows resolving vasodilatory shock | 360
    predominant cardiogenic shock | 360
    dobutamine continued | 360
    intravenous furosemide infusion started | 360
    dobutamine weaned off | 408
    hydralazine uptitration | 408
    spironolactone uptitration | 408
    bisoprolol initiated | 624
    ramipril initiated | 768
    discharged | 816
    net 25 kg weight loss | 816
    creatinine 148 µmol/L | 816
    eGFR 53 mL/min/1.73 m2 | 816
    sacubitril/valsartan discontinued | 816
    hyperkalaemia | 816
    New York Heart Association class II | 20160
