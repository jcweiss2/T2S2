80 years old | 0
    woman | 0
    non-smoker | 0
    hypertension | 0
    acute dyspnea | 0
    fecal incontinence | -1320
    left hemiplegia | -1320
    dextroversion | -1320
    dysarthria | -1320
    vomiting | -1320
    impaired consciousness | -1320
    right thalamus bleeding | 0
    right putamen bleeding | 0
    systolic blood pressure 91 mmHg | 0
    respiratory rate 24/min | 0
    SpO2 86% | 0
    poor oral hygiene | 0
    diminished breath sounds left side | 0
    coarse crackles right lung | 0
    decreased breath sounds front chest | 0
    respiratory deterioration | 0
    SpO2 not maintained at 90% | 0
    endotracheal intubation | 0
    mechanical ventilation | 0
    bilateral infiltration | 0
    admission to ICU | 0
    decreased leukocyte count (1900/μL) | 0
    elevated CRP 3.6 mg/dL | 0
    PaO2 64 mmHg | 0
    normal hepatorenal function | 0
    extensive infiltration chest radiography | 0
    cerebral edema | 0
    consolidations chest CT | 0
    ground-glass opacities chest CT | 0
    A-DROP score | 0
    negative coronavirus test | 0
    chemical pneumonitis | 0
    Mendelson's syndrome | 0
    sputum culture Streptococcus agalactiae | 0
    sputum culture Klebsiella oxytoca | 0
    aspiration bacterial pneumonia | 0
    leukocytopenia | 0
    low serum CRP | 0
    respiratory viral pneumonia considered | 0
    WBC elevation | 0
    CRP elevation | 0
    ventilator management started | 0
    meropenem | 0
    levofloxacin | 0
    P/F ratio 128.75 | 0
    prednisolone started | 0
    no fever | 0
    temperature never exceeded 37°C | 0
    improvement infiltration shadows | 288
    P/F ratio improved ≥250 | 288
    extubated | 288
    transferred to neurosurgery | 528
    transferred to rehabilitation | 528
    successful extubation | 288
    steroid use | 0
    antibiotic use | 0
    ARDS management | 0
    radiographic resolution | 288
    clinical recovery | 288
    Streptococcus agalactiae infection | 0
    Klebsiella oxytoca infection | 0
    cerebral hemorrhage | 0
    bilateral lung injury | 0
    invasive mechanical ventilation | 0
    lung-protection strategies | 0
    Sivelestat sodium hydrate | 0
    Berlin definition ARDS | 0
    spontaneous respiration permitted | 0
    low tidal volume strategy | 0
    permissive hypercapnia | 0
    intracranial hypertension considered | 0
    moderate severity pneumonia | 0
    prednisolone 1 mg/kg/day | 0
    stable vital signs | 288
    clinical stability achieved | 288
    comprehensive treatment | 0
    corticosteroids effectiveness | 0
    antibiotics effectiveness | 0
    bacterial pneumonia treatment | 0
    chemical lung injury | 0
    combined bacterial and chemical injury | 0
    consent for publication obtained | 0
    Ethics Committee approval | 0
    Declaration of Helsinki compliance | 0
