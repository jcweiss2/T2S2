73 years old | 0
male | 0
admitted to the hospital | 0
symptoms began | -120
meteorism | -120
diarrhea | -120
vomiting | -120
fever | -120
low blood pressure | -120
history of ischemic stroke | 0
history of untreated type II diabetes | 0
enlarged abdomen | 0
abdomen slightly painful with palpation in the right iliac fossa | 0
abdominal radiography | 0
paraumbilical hydroaerial levels | 0
white blood cell count abnormal | 0
hemoglobin abnormal | 0
glucose abnormal | 0
creatinine abnormal | 0
urea abnormal | 0
creatinine phosphokinase abnormal | 0
potassium abnormal | 0
sodium abnormal | 0
chloride abnormal | 0
bicarbonate abnormal | 0
PCT measured | 0
PCT value >32 µg/L | 0
CRP measured | 0
CRP value 1228.5 nmol/L | 0
septic shock suspected | 0
empirical intravenous antibiotic therapy started | 0
emergency surgery performed | 0
exploratory laparotomy | 0
agglutinated intestinal loops found | 0
false membranes found | 0
purulent-appearing fluid found | 0
acute gangrenous appendicitis with perforation found | 0
suppurative omentitis found | 0
jejunum and ileum overdistended | 0
occlusive appearance | 0
appendectomy performed | 0
segmental omentectomy performed | 0
lavage and drainage of peritoneal cavity performed | 0
neglected peritonitis diagnosed | 0
intraoperative diagnosis confirmed | 0
histopathological examination performed | 0
acute fibrinopurulent peritonitis confirmed | 0
bacterial culture and sensitivity performed | 0
Escherichia coli found | 0
antibiotic resistance found | 0
antibiotic sensitivity found | 0
postoperative care started | 0
acute pancreatitis developed | 24
paroxysmal atrial fibrillation developed | 24
low blood pressure | 24
complex drug treatment started | 24
antibiotics administered | 24
anticoagulants administered | 24
analgesics administered | 24
corticosteroids administered | 24
vasopressors administered | 24
fluid volume replacement performed | 24
electrolyte and acid-base rebalancing performed | 24
patient's condition improved | 120
patient discharged | 456
follow-up at 3 months | 2160
patient in good general health | 2160
resumption of activities of daily living | 2160