45 years old|0
    woman|0
    malaise|-72
    upper respiratory tract infection|-72
    use of over-the-counter remedy containing ibuprofen and pseudoephedrine|-72
    temperature 38.5°C|0
    hypotension|0
    heart rate 250 bpm|0
    vagal maneuvers|0
    escalating doses of intravenous adenosine|0
    narrow QRS complex tachycardia|0
    crystalloid administration|0
    IV diltiazem|0
    sedation|0
    unsuccessful electrical cardioversion|0
    IV esmolol|0
    digoxin|0
    magnesium sulfate|0
    loading dose of 150 mg amiodarone|0
    increasing oxygen requirements|0
    pulmonary edema|0
    IV furosemide|0
    transfer to tertiary hospital cardiac intensive care unit|0
    second loading dose of IV amiodarone|0
    additional unsuccessful attempts at electrical cardioversion|0
    IV lidocaine|0
    procainamide|0
    transient reductions in heart rate|0
    worsening respiratory status|0
    general anesthetic|0
    intubation|0
    cooling to target temperature of 35.5°C|0
    esmolol infusion|0
    lidocaine infusion|0
    procainamide infusion|0
    heart rate slowed to 130 bpm|0
    AV dissociation|0
    heart rate gradually increased over next 12 hours|12
    infusion of vasopressin|12
    mean arterial pressure 50 mm Hg|12
    discontinuation of antiarrhythmic infusions|0
    multipolar catheters placed in coronary sinus|0
    His bundle region|0
    right ventricular apex|0
    tachycardia cycle length 504 ms|0
    reinitiation spontaneous|0
    premature ventricular contractions from RV catheter|0
    atrial beats timed to septal refractoriness|0
    sinus P waves advancing immediate His potential|0
    ventricular overdrive pacing from RV apical catheter|0
    VHHV response|0
    electroanatomic mapping|0
    earliest local potentials in mid-septal region|0
    catheter pressure terminating tachycardia|0
    radiofrequency ablation|0
    termination of tachycardia after 26 seconds|0
    slower junctional beats|0
    insurance lesions|0
    transient AH prolongation|0
    temporary atrial pacing wire|0
    sinus node suppression|0
    Streptococcus pneumoniae sputum culture|0
    IV antibiotics|0
    discharge|216
    no recurrence of tachycardia|216
    9 months of follow-up|6480
    previous medical contacts with unstable tachycardia|N/A
    prolonged admission to intensive care unit|N/A
    supraventricular tachycardia|N/A
    supportive medical treatment|N/A
    administration of beta blockade|N/A
    <|eot_id|>
    