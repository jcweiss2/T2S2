history of untreated hypertension | -168
history of morbid obesity | -168
history of chronic back pain | -168
history of IVDU | -168
back pain | -336
diffuse abdominal pain | -336
lower extremity weakness | -336
anorexia | -336
fever | -336
chills | -336
shortness of breath | -336
dizziness | -336
constipation | -336
use of acetaminophen | -336
use of gabapentin | -336
use of hydrocodone | -336
use of methamphetamines | -336
use of marijuana | -336
admission | 0
blood pressure of 79/53 mmHg | 0
heart rate of 149 bpm | 0
lactic acid of 4.2 mg dl-1 | 0
white blood cell count 37 500 u l-1 | 0
erythrocyte sedimentation rate 75 mm h-1 | 0
urine toxicology positive for cannabis | 0
urine toxicology positive for amphetamines | 0
midline tenderness of the lumbar spine | 0
3/5 strength in bilateral lower extremities | 0
bilateral shoulder warmth | 0
bilateral shoulder erythema | 0
bilateral shoulder tenderness | 0
limited range of motion | 0
multiple needle puncture sites on the antecubital fossas | 0
puncture wounds on the right foot | 0
collection of blood cultures | 0
start of vancomycin | 0
start of metronidazole | 0
start of aztreonam | 0
start of IV fluids | 0
growth of MRSA in blood cultures | 24
sensitivity of MRSA to vancomycin | 24
sensitivity of MRSA to rifampin | 24
sensitivity of MRSA to levofloxacin | 24
sensitivity of MRSA to clindamycin | 24
sensitivity of MRSA to daptomycin | 24
sensitivity of MRSA to linezolid | 24
bilateral shoulder plain radiographs | 24
arthrocentesis of the AC joints | 48
WBC of 93 137 u l-1 in one shoulder | 48
WBC of 32 043 u l-1 in the other shoulder | 48
growth of MRSA in aspirates | 48
emergent surgical debridement of the shoulders | 72
intubation | 72
MRI of the lumbar spine | 96
L3-L5 osteomyelitis | 96
facet septic arthritis | 96
dorsal paraspinous myositis | 96
L2-L5 epidural abscess | 96
bilateral psoas myositis | 96
bilateral psoas abscesses | 96
MRI of the bilateral shoulders | 120
septic arthritis of the AC joints | 120
right distal trapezius abscess | 120
left supraclavicular abscess | 120
MRI of the brain | 120
no acute intracranial processes | 120
TTE | 120
no valvular vegetations | 120
repeat surgical debridement of the shoulders | 144
evaluation by neurosurgery | 144
leukocytosis | 144
peak WBC of 52 100 u l-1 | 168
trough levels of vancomycin | 168
repeat blood cultures positive for MRSA | 168
escalation of antibiotics to daptomycin | 240
escalation of antibiotics to ceftaroline | 240
clearance of bacteraemia | 336
addition of rifampin | 336
surgical drainage of the epidural abscess | 432
intraoperative wound cultures positive for MRSA | 432
intraoperative wound cultures positive for Proteus mirabilis | 432
removal of all drains | 504
discharge | 504
prescription of oral levofloxacin | 504
prescription of oral rifampin | 504
loss to follow-up | 672