87 years old | 0
male | 0
admitted to the hospital | 0
epigastric discomfort | -24
burning sensation | -24
radiating to chest | -24
radiating to left upper quadrant | -24
nausea | -24
watery, nonbloody emesis | 0
hiccupping | 0
denied chest pain | 0
denied fever | 0
denied diarrhea | 0
denied constipation | 0
denied sneezing | 0
denied coughing | 0
denied Valsalva maneuvers | 0
coronary artery disease | 0
angina | 0
valvular heart disease | 0
hypertension | 0
hyperlipidemia | 0
gout | 0
gastro-esophageal reflux disease | 0
recent hospital admission for constipation | -168
furosemide | 0
atenolol | 0
doxazosin | 0
nifedipine | 0
simvastatin | 0
nitroglycerin | 0
omeprazole | 0
oxybutynin | 0
denied smoking | 0
denied alcohol usage | 0
hypertension | 0
afebrile | 0
abdominal distention | 0
sluggish bowel sounds | 0
soft abdomen | 0
nontender abdomen | 0
negative cardiac enzymes | 0
no acute electrocardiogram changes | 0
normal serum lactate | 0
normal creatinine | 0
contrast-enhanced CT | 0
diffuse dilation of small bowel | 0
diffuse dilation of stomach | 0
diffuse dilation of mid-to-distal esophagus | 0
esophageal pneumatosis | 0
no pneumomediastinum | 0
no pneumoperitoneum | 0
upper gastrointestinal and small bowel ileus | 0
nondiagnostic esophagram | 2
nasogastric tube placement | 2
decompression | 2
drained 1700 ccs of nonbloody fluid | 2
bowel rest | 2
intravenous fluids | 2
close observation | 2
esophagram through NG tube | 4
negative for perforation | 4
additional nasogastric tube decompression | 4
repeat CT examination | 11
resolution of esophageal pneumatosis | 11
interval improvement of upper gastrointestinal ileus | 11
septic | 48
broad-spectrum antibiotics | 48
tracheal aspirates grew Klebsiella pneumoniae | 48
acute kidney injury | 48
antibiotic regimen adjustment | 48
resolution of acute kidney injury | 120
discharged home | 288
tolerating regular oral diet | 288