54 years old | 0
male | 0
Caucasian | 0
admitted to the emergency department | 0
progressive pain | -168
swelling of the right lower extremity | -168
permanent redness | -168
petechial haemorrhage | -168
hit his leg | -168
septic shock | 0
tachycardia | 0
dyspnoea | 0
arterial hypotension | 0
transfer to the ICU | 0.5
blood pressure 81/42 mmHg | 0
heart rate 128 bpm | 0
temperature 39.2°C | 0
respiratory rate 38 breaths per minute | 0
SpO2 96% | 0
paO2 114 mmHg | 0
moderately impaired left ventricular ejection fraction | 0
white blood cell count 20.23 × 10^9/L | 0
C-reactive protein 3362 nmol/L | 0
procalcitonin 43.5 µg/L | 0
lactate 8.8 mmol/L | 0
platelet count 160 × 10^9/L | 0
total bilirubin 42.75 µmol/L | 0
aspartate aminotransferase 950 nmol/s*L | 0
alanine aminotransferase 850 nmol/s*L | 0
blood glucose level 20.8 mmol/L | 0
undiagnosed and untreated diabetes mellitus | 0
necrotising fasciitis | 0
severe sepsis | 0
multiple organ failure | 0
liver failure | 0
renal failure | 0
elevated renal values | 0
absent urine output | 0
acute renal failure | 0
myoglobin level 125 nmol/L | 0
continuous veno-venous haemodialysis | 0
intubation | 2
acidosis | 2
paO2 179 mmHg | 2
Horowitz Index 256 mmHg | 2
mild acute respiratory distress syndrome | 2
wound debridement | 6
excision of the fascia | 6
microbiological biopsy sampling | 6
haemodynamic situation deteriorated | 24
catecholamine therapy | 24
whole-body computed tomography scan | 24
subcutaneous fluid retention | 24
perifascial air | 24
indication for immediate transfemoral amputation | 24
amputation | 24
stump revision | 96
wound closure | 216
pathologic findings | 216
necrotising florid inflammation | 216
antibiotic therapy | 0
piperacillin/tazobactam | 0
clindamycin | 0
Streptococcus pyogenes | 48
penicillin G | 48
immunoglobulin therapy | 48
Pentaglobin | 48
weaning from mechanical ventilation | 168
extubation | 168
inflammatory parameters decreased | 168
transfer to the normal ward | 384
prosthesis for the right thigh | 384
discharge to rehabilitation | 624
discharge home | 720