32 years old | 0
Hispanic | 0
female | 0
presented to the Emergency Department | 0
fever | -72
chills | -72
generalized weakness | -72
malaise | -72
body aches | -72
symptoms progressed in severity | -72
reported to the Emergency Department on two separate occasions | 0
initial presentation | -96
physical exam revealed fever | -96
maximum temperature of 103.3 °F | -96
tachycardia | -96
heart rate of 120 beats per minute | -96
blood pressure of 128/82 mmHg | -96
respiratory rate of 18 breaths per minute | -96
oxygen saturation of 99% on room air | -96
physical exam unremarkable | -96
patient denied chest pain | -96
denied cough | -96
denied shortness of breath | -96
denied abdominal pain | -96
resided in a rural community in coastal South Texas | 0
had dogs and cats at home | 0
no recent exposure to communicable diseases | 0
no recent travel outside of the country | 0
no tobacco use | 0
no alcohol use | 0
no illicit drug use | 0
complete blood count showed white blood cells 4300 cells/mm³ | -96
neutrophils 85% | -96
lymphocytes 11.4% | -96
monocytes 3% | -96
hemoglobin 12.4 g/dL | -96
hematocrit 37.2% | -96
platelets 230,000 per cubic mm | -96
aspartate aminotransferase 38 U/L | -96
alanine aminotransferase 28 U/L | -96
alkaline phosphatase 62 U/L | -96
rapid influenza A and B test normal | -96
urinalysis normal | -96
lactic acid normal | -96
thyroid-stimulating hormone normal | -96
chest radiograph indicated mild peribronchial cuffing consistent with bronchitis | -96
received one liter of 0.9% normal saline intravenously | -96
received one oral dose of ibuprofen 800 mg | -96
diagnosed with viral bronchitis | -96
discharged home | -96
patient deteriorated clinically | -72
returned to the Emergency Department four days later | 0
fever | 0
body aches | 0
temperature of 101.2 °F | 0
tachycardia with heart rate of 125 beats per minute | 0
respiratory rate of 17 breaths per minute | 0
blood pressure of 118/56 mmHg | 0
oxygen saturation of 99% at room air | 0
physical examination remarkable for diminished breath sounds to bilateral lung fields | 0
tachycardia | 0
dry mucous membranes | 0
decreased skin turgor | 0
laboratory data showed white blood cells 3600 cell/mm³ | 0
neutrophils 82.8% | 0
lymphocytes 11% | 0
monocytes 5% | 0
hemoglobin 11.6 g/dL | 0
hematocrit 33.2% | 0
platelets 64,000 per cubic mm | 0
aspartate aminotransferase 226 U/L | 0
alanine aminotransferase 138 U/L | 0
alkaline phosphatase 182 U/L | 0
D-dimer >5000 ng/mL | 0
lactic acid 2.4 mmol/L | 0
normal fibrinogen | 0
chest radiograph identified bilateral alveolar infiltrates | 0
computed tomographic angiogram of the chest negative for pulmonary embolism | 0
confirmed bilateral lower lobe consolidation | 0
admitted to the medical-surgical floor | 0
diagnosis of sepsis secondary to community-acquired pneumonia | 0
sepsis protocol initiated | 0
meropenem | 0
voriconazole | 0
blood cultures obtained | 0
urine cultures obtained | 0
resuscitation with 3 liters of intravenous 0.9% normal saline fluid | 0
remained tachypneic | 0
remained tachycardic | 0
condition deteriorated | 6
became hypotensive | 6
blood pressure of 87/53 mmHg | 6
heart rate of 137 beats per minute | 6
respiratory rate of 36 breaths per minute | 6
transferred to the Intensive Care Unit | 6
requiring two more liters of intravenous fluid of 0.9% normal saline | 6
initial impression was atypical pneumonia | 6
serology panel for suspected zoonoses collected | 6
developed a dry cough | 24
progressed to acute hypoxemic respiratory failure | 24
heart rate of 144 beats per minute | 24
respiratory rate of 33 breaths per minute | 24
oxygen saturation of 82% | 24
echocardiogram revealed mild right heart chamber dilatation | 24
normal left ventricular systolic function | 24
ejection fraction of 65% | 24
arterial blood gases showed PaO2/FiO2 of 102 | 24
consistent with moderately severe ARDS | 24
managed with non-invasive positive pressure ventilation | 24
voriconazole discontinued | 24
meropenem continued | 24
doxycycline continued | 24
awaiting final serology panel and culture results | 24
all bacterial cultures yielded negative results | 24
developed a nontender pink maculopapular rash to the bilateral lower extremities | 96
no associated lymphadenopathy | 96
zoonoses serology panel confirmed acute infection of murine typhus | 168
Typhus Fever group IgM titer of 1:128 | 168
murine typhus IgG titer of 1:258 | 168
meropenem discontinued | 168
antimicrobials deescalated to doxycycline monotherapy | 168
weaning process from non-invasive positive pressure ventilation | 168
weaning to high flow oxygen nasal cannula | 168
weaning to low flow oxygen nasal cannula at 2 liters per minute | 168
discharged home | 192
no oxygen supplementation | 192
treatment completed with minocycline for 11 additional days | 192
nationwide shortage of doxycycline | 192
generalized weakness at discharge | 192
no other complaints | 192
