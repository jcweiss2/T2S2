67 years old | 0
male | 0
admitted to the hospital | 0
malaise | -96
anorexia | -96
dry cough | -96
dyspnea | -96
severe respiratory distress | 0
oxygen saturation of 79% | 0
bilateral interstitial infiltrates | 0
right lower lobe consolidation | 0
shock | 0
elevated lactic acid of 7.8 mmol/L | 0
endotracheal intubation | 0
mechanical ventilation | 0
fluid resuscitation | 0
antibiotics | 0
vasopressor support | 0
septic shock secondary to presumed community-acquired pneumonia | 0
hepatocellular carcinoma | -720
rectal adenocarcinoma | -720
non-small-cell lung cancer | -720
surgical resections | -720
chemoradiation therapy | -720
remission | -720
chronic obstructive lung disease | -720
chronic kidney disease (stage 3) | -720
diabetes mellitus | -720
SARS-CoV-2 infection | 0
positive real-time polymerase chain result for SARS-CoV-2 | 0
preserved left ventricular ejection fraction | 0
severely dilated right ventricle | 0
reduced RV function | 0
flattening of the interventricular septum | 0
severe tricuspid regurgitation | 0
estimated systolic pulmonary artery pressure of 56 mm Hg | 0
normal RV function | -35040
elevated D-dimer >4.0 mg/L | 0
high-sensitivity troponin at baseline of 275 ng/L | 0
subsequent 6-hour high-sensitivity troponin of 255 ng/L | 6
normal sinus rhythm | 0
no significant ST-T-wave changes | 0
therapeutic anticoagulation | 0
elevated d-dimer level | 0
acute deep vein thrombosis in the left posterior tibial vein | 0
subsegmental right upper lobe pulmonary embolism | 0
neuromuscular blockade | 0
prone-position ventilation | 0
respiratory failure from ARDS due to COVID-19 | 0
tidal volumes between 5 and 7 ml/kg of ideal body weight | 0
positive end-expiratory pressure between 10 and 14 cm H2O | 0
plateau pressure between 26 and 32 cm H2O | 0
vasopressor support with norepinephrine | 0
vasopressor support with vasopressin | 0
acute kidney injury | 0
continuous renal replacement therapy | 0
shock liver | 0
gastrointestinal hemorrhage | 0
Escherichia coli pneumonia | 0
bacteremia | 0
poor prognosis | 0
comfort measures | 0
withdrawal of life-support interventions | 0
passed away after 22 days in the ICU | 528
