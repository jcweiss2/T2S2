78 years old | 0
male | 0
admitted to the hospital | 0
pacemaker implantation | -6120
advanced atrioventricular block | -6120
transient loss of pacing capture | -120
septic cholangitis | -120
cardiologist assessment | -120
pacemaker interrogation | -120
pulse generator upgrade | -60
Medtronic Advisa | -60
DDD mode | -60
dual chamber pacing and sensing | -60
dual response to sensing | -60
lower rate limit of 70 beats/min | -60
gastrectomy | -unknown
gastroduodenal ulcer | -unknown
type 2 diabetes mellitus | -unknown
glargine | 0
vildagliptin | 0
moderate distress | 0
blood pressure of 176/73 mm Hg | 0
abdominal tenderness | 0
right upper quadrant tenderness | 0
electrocardiogram | 0
dual-chamber atrial and ventricular pacing | 0
capture at 70 beats/min | 0
hematocrit of 32.5% | 0
anesthesia induction | 0
remifentanil | 0
propofol | 0
rocuronium | 0
sevoflurane | 0
pacemaker interrogation | 0
DOO mode | 0
asynchronous atrial and ventricular pacing | 0
70 beats/min | 0
adhesiolysis | 0
small bowel obstruction | 0
cholecystectomy | 0
ultrasound-guided rectus sheath block | 0
40-mL 0.25% levobupivacaine | 0
pacemaker reinterrogation | 0
pacemaker reprogramming | 0
DDD mode | 0
ventricular pacing threshold of 1.25 V | 0
emergence from anesthesia | 0
extubation | 0.5
asystole | 0.5
cardiopulmonary resuscitation | 0.5
ventricular pacing output increase | 0.5
stable hemodynamics | 0.5
ventricular pacing threshold of 3.0 V | 0.5
arterial blood gas analysis | 1
pH 7.29 | 1
Pco2 46 mm Hg | 1
Po2 112 mm Hg | 1
HCO3 22.5 mmol/L | 1
sodium 142 mmol/L | 1
potassium 4.4 mmol/L | 1
tranthoracic echocardiography | 1
good left ventricular systolic function | 1
no regional wall motion abnormalities | 1
ICU admission | 0
ventricular pacing threshold of 1.75 V | 8
discharge | 288
ventricular pacing threshold of 0.75 V | 288
ventricular pacing output of 2.5 V | 288