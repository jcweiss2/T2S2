23 years old | 0
    female | 0
    admitted for induction of labour | 0
    cervical ripening balloon catheter inserted | -12
    cervical ripening balloon catheter removed | 0
    artificial rupture of membranes | 0
    clear liquor observed | 0
    intravenous oxytocin infusion commenced | 0
    epidural anaesthesia requested | 0
    indwelling catheter inserted | 0
    full dilatation reported | 6
    passive descent of fetal head allowed | 6
    active pushing commenced | 7
    pathological cardiotocograph | 7
    late decelerations | 7
    prolonged decelerations | 7
    instrumental delivery decision | 7
    indwelling catheter balloon deflated | 7
    rosé-coloured haematuria noted | 7
    no significant vaginal bleeding | 7
    low cavity vacuum delivery | 8
    right mediolateral episiotomy | 8
    baby delivered occiput-anterior | 8
    McRoberts manoeuvre required | 8
    healthy male neonate delivered | 8
    Apgar scores 9 at 1 minute postpartum | 8
    Apgar scores 10 at 5 minutes postpartum | 8
    postpartum haemorrhage secondary to atony | 8
    local haemorrhage at episiotomy site | 8
    syntocinon infusion administered | 8
    ergometrine administered | 8
    episiotomy laceration suture repair | 8
    estimated blood loss 600 mL | 8
    indwelling catheter reinserted | 8
    clear urine noted | 8
    epidural catheter removed | 8
    well overnight | 8
    no concerns of pain | 8
    no haemodynamic instability | 8
    indwelling catheter removed on day 1 postpartum | 24
    one normal micturition | 26
    acute right-flank pain developed | 27
    right-flank pain radiating to right iliac fossa | 27
    constant severe pain | 27
    opioid analgesia required | 27
    rebound tenderness at right iliac fossa | 27
    rebound tenderness at right renal angle | 27
    indwelling catheter re-inserted | 27
    1000 mL clear urine drained | 27
    no improvement in pain after bladder decompression | 27
    febrile 38.4 °C | 27
    tachycardic | 27
    hypotensive | 27
    haemoglobin level 86 | 27
    white cell count 6 | 27
    venous lactate 1.9 | 27
    creatinine 58 | 27
    CRP 87 | 27
    uterine rupture considered | 27
    puerperal sepsis considered | 27
    renal calculi considered | 27
    appendicitis considered | 27
    IV crystalloid administered | 27
    ceftriaxone administered | 27
    metronidazole administered | 27
    gentamicin administered | 27
    urine output >100 mL/h | 27
    remained hypotensive | 27
    remained tachycardic | 27
    CT abdomen and pelvis with contrast performed | 27
    free fluid in right retroperitoneal space | 27
    free fluid involving inferior perinephric space | 27
    free fluid extending into lateral pelvic side wall | 27
    no signs of uterine rupture | 27
    simple fluid suspected | 27
    fluid suspected to be urine | 27
    haemoglobin stable at 86 | 27
    haematocrit 0.265 | 27
    CRP 76 | 27
    creatinine 50 | 27
    urine microscopy presence of organisms | 27
    sepsis from urinary tract source considered | 27
    transudative fluid considered | 27
    lower urinary tract injury considered unlikely | 27
    haemodynamically unstable | 27
    transferred to intensive care | 28
    IV metaraminol commenced | 28
    packed red blood cells administered | 28
    urology team consulted | 28
    CT IV pyelogram recommended | 28
    CT IV pyelogram performed | 28
    contrast extravasation at right mid ureter | 28
    no hydronephrosis bilaterally | 28
    no collection amenable to drainage | 28
    ureteric injury unexpected | 28
    maintaining urine output >100 mL/h | 28
    urine clear | 28
    emergency cystoscopy performed | 51
    posterior bladder wall ecchymosis noted | 51
    normal mucosa | 51
    normal ureteral orifice | 51
    guide wire could not be passed | 51
    right rigid ureteroscopy performed | 51
    grade III incomplete proximal ureteric rupture | 51
    ureteric stent placed | 51
    postoperative monitoring in ICU | 51
    persistent fevers | 51
    antibiotics upgraded to piperacillin/tazobactam | 51
    urine microscopy positive for E. coli | 51
    stepped down to ward-based care | 51
    remained well | 51
    discharged home 10 days after delivery | 360
    follow-up cystoscopy planned | 360
    retrograde pyelogram planned | 360
    stent removal or exchange planned | 360
    intra-operative pyelogram demonstrated no contrast leak | 1008
    stent removed | 1008
    no complications | 1008
    