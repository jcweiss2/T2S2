57 years old | 0
post-menopausal female | 0
admitted to the hospital | 0
bleeding per vaginum | -48
diabetes mellitus Type 2 | 0
dyslipidaemia | 0
hypothyroidism | 0
hysteroscopic myomectomy | 0
general anaesthesia | 0
morphine | 0
glycopyrrolate | 0
ondansetron | 0
propofol | 0
succinylcholine | 0
endotracheal intubation | 0
nitrous oxide | 0
isoflurane | 0
vecuronium | 0
normal saline solution | 0
electrocardiography | 0
non-invasive blood pressure | 0
end tidal carbon dioxide | 0
pulse oximetry | 0
temperature | 0
hysteroscopic examination | 0
submucous fibroid | 0
resection of fibroid | 0
1.5% glycine | 0
Karl Storz hysteroscope | 0
intrauterine pressure | 0
SpO2 fell | 45
airway pressure rose | 45
breath sounds diminished | 45
NIBP 90/70 mmHg | 45
pulse rate 100/min | 45
pink frothy secretions | 45
crackles | 45
acute pulmonary oedema | 45
lasix | 45
morphine | 45
nasogastric tube | 45
bladder catheterized | 45
urine output 100 mL | 45
12 lead ECG | 45
arterial blood gas | 45
pO2: 165.3 mmHg | 45
pCO2: 50.5 mmHg | 45
pH: 7.17 | 45
K+: 5.3 mmol/L | 45
Na+: 100 mmol/L | 45
HCO3-: 17.8 mmol/L | 45
BE: –8.2 mmol/L | 45
O2 Sat: 98.6% | 45
portable chest radiograph | 45
perihilar interstitial infiltrates | 45
pulmonary vasculature | 45
glycine deficit | 45
fluid overload | 45
hyponatraemia | 45
metabolic acidosis | 45
pulmonary oedema | 45
right internal jugular vein cannulated | 45
left radial artery cannulated | 45
haemodynamic monitoring | 45
ABG analysis | 45
central venous pressure | 45
elective mechanical ventilation | 45
IV morphine sedation | 45
soda bicarbonate | 45
3% sodium chloride | 45
inotropes | 45
urgent echocardiogram | 45
serial ABG | 45
Na+ levels | 45
3% NaCl stopped | 45
profuse bleeding per vaginum | 12
endometrial tamponade | 12
Foley's catheter | 12
Disseminated intravascular coagulation | 12
oozing from other sites | 12
nasogastric tube | 12
coffee ground aspirate | 12
coagulation profile | 12
Haemoglobin 5 gm% | 12
platelet count 90,000/mm3 | 12
prothrombin time 22 s | 12
partial thromboplastin time 68 s | 12
International Normalized Ratio 1.94 | 12
d-dimer positive | 12
hypocalcaemia | 12
fresh blood | 12
blood products | 12
fresh frozen plasma | 12
cryoprecipitate | 12
IV calcium | 12
coagulation profile improved | 48
inotropic support tapered off | 48
SIMV mode ventilation | 48
pressure support | 48
FiO2 reduction | 48
continuous positive airway pressure trial | 48
extubation | 48
tachypnoeic | 72
respiratory rate 36/min | 72
bilateral wheeze | 72
SpO2 85% | 72
chest X-ray | 72
opacities in left lower zone | 72
pneumonitis | 72
fibreoptic bronchoscopy | 72
long tubular casts | 72
left bronchial tree | 72
asthalin nebulization | 72
chest physiotherapy | 72
BIPAP support | 72
broad-spectrum antibiotics | 72
Pseudomonas aeruginosa | 72
cramps in both legs | 120
bilateral foot drop | 120
nerve conduction studies | 120
common peroneal nerve palsy | 120
physiotherapy | 120
discharged to home | 336