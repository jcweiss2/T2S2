69 years old | 0
    male | 0
    scheduled for repeated arthroscopic lavage of the right knee | 0
    unimproved septic arthritis | -336
    previous arthroscopic lavage procedure | -336
    peripheral arterial occlusive disease in the lower extremities | -336
    no evidence of deep vein thrombosis | -336
    hypertension | 0
    type 2 diabetes | 0
    new onset atrial fibrillation with rapid ventricular response | -336
    transthoracic echocardiography showing left atrial enlargement, normal left ventricular function, ejection fraction 61.3%, no intracardiac thrombus | -336
    flecainide | -336
    aspirin | -336
    preoperative electrocardiogram showing normal sinus rhythm | 0
    intramuscular injection of glycopyrrolate 0.2 mg | 0
    anesthesia induced with propofol | 0
    anesthesia induced with rocuronium | 0
    airway secured with cuffed 7.5 mm endotracheal tube | 0
    monitoring electrocardiogram | 0
    monitoring pulse oxygen saturation | 0
    monitoring capnogram | 0
    monitoring esophageal temperature |=
    monitoring invasive arterial pressure | 0
    anesthesia maintained with sevoflurane | 0
    anesthesia maintained with 50% nitrous oxide in oxygen | 0
    arterial blood gas analysis 10 minutes after induction | 0
    arterial blood gas analysis showing pH 7.38 | 0
    arterial blood gas analysis showing PaCO2 45.1 mmHg | 0
    arterial blood gas analysis showing PaO2 85.7 mmHg | 0
    arterial blood gas analysis showing HCO3- 26.0 mEq/L | 0
    arterial blood gas analysis showing SaO2 95.5% | 0
    end tidal CO2 24 mmHg | 0
    tidal volume increased to 750 ml from 650 ml | 0
    arterial blood gas analysis 20 minutes after changing ventilator setting | 20
    arterial blood gas analysis showing pH 7.31 | 20
    arterial blood gas analysis showing PaCO2 47.0 mmHg | 20
    arterial blood gas analysis showing PaO2 75.1 mmHg | 20
    arterial blood gas analysis showing HCO3) 23.6 mEq/L | 20
    arterial blood gas analysis showing SaO2 92.8% | 20
    phenylephrine 100 µg injected intravenously at 30 minutes after induction | 30
    blood pressure dropped to 90/60 mmHg | 30
    heart rate increased to 100 beats per minute | 30
    arterial blood pressure dropped to 65/45 mmHg at 40 minutes after induction | 40
    heart rate 48 beats per minute at 40 minutes after induction | 40
    epinephrine 30 µg administered intravenously | 40
    additional 50 µg epinephrine administered intravenously | 40
    atropine sulfate 0.5 mg administered intravenously | 40
    vital signs deteriorated | 40
    pulsatile activity disappeared in arterial line | 40
    cardiopulmonary resuscitation (CPR) started | 40
    surgery completed | 40
    nitrous oxide turned off | 40
    sevoflurane turned off | 40
    epinephrine 1 mg administered intravenously | 40
    atropine sulfate 0.5 mg administered intravenously | 40
    vital signs not improved despite intermittent epinephrine administration | 40
    arterial blood gas analysis during CPR | 40
    arterial blood gas analysis showing pH 7.37 | 40
    arterial blood gas analysis showing PaCO2 27.8 mmHg | 40
    arterial blood gas analysis showing PaO2 63.9 mmHg | 40
    arterial blood gas analysis showing HCO3- 15.8 mEq/L | 40
    arterial blood gas analysis showing SaO2 90.8% | 40
    FiO2 1.0 during CPR | 40
    external cardiac massage stopped 8 minutes after starting CPR | 48
    arterial blood gas analysis after stopping external cardiac massage | 48
    arterial blood gas analysis showing pH 6.96 | 48
    arterial blood gas analysis showing PaCO2 63.9 mmHg | 48
    arterial blood gas analysis showing PaO2 221.4 mmHg | 48
    arterial blood gas analysis showing HCO3- 13.9 mEq/L | 48
    arterial blood gas analysis showing SaO2 98.5% | 48
    vital signs fluctuating severely | 48
    CPR intermittently continued | 48
    administration of epinephrine during CPR | 48
    administration of sodium bicarbonate during CPR | 48
    emergency transthoracic echocardiogram performed 10 minutes after CPR initiation | 50
    echocardiogram showing massive thrombus in right atrium | 50
    echocardiogram showing dilated hypokinetic right ventricle | 50
    echocardiogram showing D-shaped left ventricle | 50
    preliminary diagnosis of massive pulmonary embolism | 50
    decision to proceed with fibrinolysis during CPR | 50
    alteplase 20 mg administered intravenously 37 minutes after CPR initiation | 77
    alteplase 100 mg continuously infused over 90 minutes | 77
    echocardiogram after r-tPA injection showing improved D-shaped left ventricle | 77
    echocardiogram after r-tPA injection showing remaining thrombi in right atrium | 77
    hemodynamic performance stabilized | 77
    no sign of bleeding at operation site | 77
    external cardiac massage stopped 26 minutes after r-tPA injection | 103
    patient transferred to intensive care unit intubated | 103
    blood pressure 110/60 mmHg upon transfer | 103
    heart rate 100 beats per minute upon transfer | 103
    mechanical ventilation upon transfer | 103
    heparin administered 12 hours after r-tPA injection | 192
    PT INR 1.65 | 192
    aPTT 50-70 seconds | 192
    patient's consciousness became alert 18 hours after r-tPA | 180
    endotracheal tube extubated | 180
    thrombi completely disappeared on echocardiogram 3 days after surgery | 288
    dilated hypokinetic right ventricle returned to normal | 288
    heparin infusion stopped 5 days after surgery | 360
    patient recovered completely without hemorrhagic episodes | 360
    transferred from intensive care unit to medical ward | 360

    69 years old | 0  
    male | 0  
    scheduled for repeated arthroscopic lavage of the right knee | 0  
    unimproved septic arthritis | -336  
    previous arthroscopic lavage procedure | -336  
    peripheral arterial occlusive disease in the lower extremities | -336  
    no evidence of deep vein thrombosis | -336  
    hypertension | 0  
    type 2 diabetes | 0  
    new onset atrial fibrillation with rapid ventricular response | -336  
    transthoracic echocardiography showing left atrial enlargement, normal left ventricular function, ejection fraction 61.3%, no intracardiac thrombus | -336  
    flecainide | -336  
    aspirin | -336  
    preoperative electrocardiogram showing normal sinus rhythm | 0  
    intramuscular injection of glycopyrrolate 0.2 mg | 0  
    anesthesia induced with propofol | 0  
    anesthesia induced with rocuronium | 0  
    airway secured with cuffed 7.5 mm endotracheal tube | 0  
    monitoring electrocardiogram | 0  
    monitoring pulse oxygen saturation | 0  
    monitoring capnogram | 0  
    monitoring esophageal temperature | 0  
    monitoring invasive arterial pressure | 0  
    anesthesia maintained with sevoflurane | 0  
    anesthesia maintained with 50% nitrous oxide in oxygen | 0  
    arterial blood gas analysis 10 minutes after induction | 0  
    arterial blood gas analysis showing pH 7.38 | 0  
    arterial blood gas analysis showing PaCO2 45.1 mmHg | 0  
    arterial blood gas analysis showing PaO2 85.7 mmHg | 0  
    arterial blood gas analysis showing HCO3- 26.0 mEq/L | 0  
    arterial blood gas analysis showing SaO2 95.5% | 0  
    end tidal CO2 24 mmHg | 0  
    tidal volume increased to 750 ml from 650 ml | 0  
    arterial blood gas analysis 20 minutes after changing ventilator setting | 20  
    arterial blood gas analysis showing pH 7.31 | 20  
    arterial blood gas analysis showing PaCO2 47.0 mmHg | 20  
    arterial blood gas analysis showing PaO2 75.1 mmHg | 20  
    arterial blood gas analysis showing HCO3- 23.6 mEq/L | 20  
    arterial blood gas analysis showing SaO2 92.8% | 20  
    phenylephrine 100 µg injected intravenously at 30 minutes after induction | 30  
    blood pressure dropped to 90/60 mmHg | 30  
    heart rate increased to 100 beats per minute | 30  
    arterial blood pressure dropped to 65/45 mmHg at 40 minutes after induction | 40  
    heart rate 48 beats per minute at 40 minutes after induction | 40  
    epinephrine 30 µg administered intravenously | 40  
    additional 50 µg epinephrine administered intravenously | 40  
    atropine sulfate 0.5 mg administered intravenously | 40  
    vital signs deteriorated | 40  
    pulsatile activity disappeared in arterial line | 40  
    cardiopulmonary resuscitation (CPR) started | 40  
    surgery completed | 40  
    nitrous oxide turned off | 40  
    sevoflurane turned off | 40  
    epinephrine 1 mg administered intravenously | 40  
    atropine sulfate 0.5 mg administered intravenously | 40  
    vital signs not improved despite intermittent epinephrine administration | 40  
    arterial blood gas analysis during CPR | 40  
    arterial blood gas analysis showing pH 7.37 | 40  
    arterial blood gas analysis showing PaCO2 27.8 mmHg | 40  
    arterial blood gas analysis showing PaO2 63.9 mmHg | 40  
    arterial blood gas analysis showing HCO3- 15.8 mEq/L | 40  
    arterial blood gas analysis showing SaO2 90.8% | 40  
    FiO2 1.0 during CPR | 40  
    external cardiac massage stopped 8 minutes after starting CPR | 48  
    arterial blood gas analysis after stopping external cardiac massage | 48  
    arterial blood gas analysis showing pH 6.96 | 48  
    arterial blood gas analysis showing PaCO2 63.9 mmHg | 48  
    arterial blood gas analysis showing PaO2 221.4 mmHg | 48  
    arterial blood gas analysis showing HCO3- 13.9 mEq/L | 48  
    arterial blood gas analysis showing SaO2 98.5% | 48  
    vital signs fluctuating severely | 48  
    CPR intermittently continued | 48  
    administration of epinephrine during CPR | 48  
    administration of sodium bicarbonate during CPR | 48  
    emergency transthoracic echocardiogram performed 10 minutes after CPR initiation | 50  
    echocardiogram showing massive thrombus in right atrium | 50  
    echocardiogram showing dilated hypokinetic right ventricle | 50  
    echocardiogram showing D-shaped left ventricle | 50  
    preliminary diagnosis of massive pulmonary embolism | 50  
    decision to proceed with fibrinolysis during CPR | 50  
    alteplase 20 mg administered intravenously 37 minutes after CPR initiation | 77  
    alteplase 100 mg continuously infused over 90 minutes | 77  
    echocardiogram after r-tPA injection showing improved D-shaped left ventricle | 77  
    echocardiogram after r-tPA injection showing remaining thrombi in right atrium | 77  
    hemodynamic performance stabilized | 77  
    no sign of bleeding at operation site | 77  
    external cardiac massage stopped 26 minutes after r-tPA injection | 103  
    patient transferred to intensive care unit intubated | 103  
    blood pressure 110/60 mmHg upon transfer | 103  
    heart rate 100 beats per minute upon transfer | 103  
    mechanical ventilation upon transfer | 103  
    heparin administered 12 hours after r-tPA injection | 192  
    PT INR 1.65 | 192  
    aPTT 50-70 seconds | 192  
    patient's consciousness became alert 18 hours after r-tPA | 180  
    endotracheal tube extubated | 180  
    thrombi completely disappeared on echocardiogram 3 days after surgery | 288  
    dilated hypokinetic right ventricle returned to normal | 288  
    heparin infusion stopped 5 days after surgery | 360  
    patient recovered completely without hemorrhagic episodes | 360  
    transferred from intensive care unit to medical ward | 360  
    