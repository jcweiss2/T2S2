40 years old | 0
male | 0
diabetic for 4 years | 0
COVID-19 | -2928
hospitalized for 6 days | -2928
ventilator support | -2928
unilateral swelling (post-COVID) left side of the face | -216
loosening of teeth | -216
diagnosed with mucormycosis | -216
surgical debridement | -216
amphotericin B drug therapy | -216
oroantral communication | 0
oronasal communication | 0
mastication difficulties | 0
nasal regurgitations | 0
absence of the left orbit | 0
total maxilla absence | 0
concave profile | 0
obliterated nasolabial fold | 0
drooped corners of mouth | 0
insufficient upper lip support | 0
porcelain-fused ceramic full-veneer crown on right molar | 0
slightly supraerupted malaligned anterior teeth | 0
normal tongue movement | 0
normal temporomandibular joint movement | 0
left total maxillectomy | 0
right subtotal maxillectomy | 0
left orbital decompression | 0
resection of left zygomatic arch | 0
resection of left zygomatic rim | 0
implant-supported removable prosthesis | 0
general anesthesia | 0
custom-made subperiosteal zygomatic implants | 0
healing after 15 days | 360
impression-making process | 360
open-tray impression copings | 360
polyvinyl siloxane impression material | 360
inter arch records | 360
titanium metal bar | 360
obturator fabrication | 360
heat-cured acrylic resin | 360
metal mesh reinforcement | 360
bilateral balanced occlusion | 360
semianatomic teeth | 360
prosthesis insertion | 360
lacking seal on left posterior tooth region | 360
soft relining material | 360
follow-up visits after 15 days | 360
follow-up visits after 30 days | 720
follow-up visits after 45 days | 1080
follow-up visits after 60 days | 1440
follow-up visits after 90 days | 2160
occlusal refinements | 360
speech quality evaluation | 360
peripheral seal evaluation | 360
patient satisfied with prosthesis | 2160
