73 years old | 0
male | 0
medical history of multiple thromboses | -2160
deep vein thrombosis | -2160
deep vein thrombosis | -24
pulmonary embolism | -2160
pulmonary embolism | -108
admitted to cardiology department | 0
acute thoracic pain | 0
electrocardiogram evidenced inferior Q waves with ST elevation | 0
echography revealed antero-inferior akinesia | 0
coronary catheterization showed a thrombosis in the right coronary artery | 0
balloon angioplasty | 0
antiplatelet therapy with acetylsalicylic acid and clopidogrel | 0
fluidione | 0
fever | 0
inflammatory syndrome | 0
fatigue | 0
signs of anemia | 0
hemoglobin level was 90 g/L | 0
reticulocytes were 52 × 10^9/L | 0
white blood cells 6.6 × 10^9/L | 0
platelet count was 52 × 10^9/L | 0
C-reactive protein level was 147 mg/L | 0
serum haptoglobin was decreased | 0
lactate dehydrogenase level was markedly elevated | 0
direct antiglobulin test was negative | 0
computerized tomography scan showed a thrombosis of the hepatic vein | 0
flow cytometry test disclosed a big-sized PNH clone | 0
diagnosis of classical PNH | 0
eculizumab treatment started | 24
prophylaxis including vaccination against meningococcal and pneumococcal infection | 24
penicillin V therapy | 24
recovery | 48
fever resolved | 48
abdominal pain resolved | 48
inflammatory syndrome resolved | 48
severe thrombocytopenia occurred | 216
new BM examination showed a normocellular BM with dysplasia | 216
diagnosis of refractory anemia with excess blast-2 | 216
vitamin K antagonists stopped | 216
antiplatelet treatment maintained | 216
platelet and red blood cell transfusions | 216
hypomethylating treatment with 5-azacytidine added | 216
septic shock due to the infection of his implantable chamber by Aeromonas veronii | 312
multiorgan failure | 312
death | 312