51 years old | 0
male | 0
end-stage renal disease | -6720
polycystic kidney disease | -6720
renal transplant | -3456
renal transplant | -2880
sepsis | 0
E coli bacteremia | 0
acute renal failure | 0
hemodialysis | 0
intubation | 0
pressors | 0
broad-spectrum antibiotics | 0
stabilized | 0
weaned off pressor support | 144
extubated | 144
poor urine output | 144
dialysis | 144
transplant ultrasound | 144
abdominal X-ray | 144
new renal parenchymal gas | 144
emphysematous pyelonephritis | 144
percutaneous drain | 168
increasing pressor support | 168
re-intubated | 168
nephrectomy | 192
infected kidney | 192
soft and boggy | 192
infarcted | 192
liquefaction necrosis | 192
endarteritis | 192
chronic transplant arteriopathy | 192
arterial thrombi | 192
cortical infarctions | 192
thrombotic microangiopathy | 192
micro abscess formation | 192
extubated | 216
pressor support discontinued | 216
progressive ischemia | 216
peripheral artery disease | 216
bilateral amputation | 240
transmetatarsal amputation | 240
bilateral knee amputation | 720
worsening sepsis | 720
lower limb extremity tissue necrosis | 720
cardiopulmonary arrest | 720 
death | 720