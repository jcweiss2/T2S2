55 years old | 0
male | 0
diagnosed with Hodgkin lymphoma | -43800
received chemotherapy | -1464
autologous peripheral blood stem cell transplantation | -1440
fever | -168
marked dyspnea | -168
hospitalized | 0
increased serum lactate dehydrogenase | 0
increased C-reactive protein | 0
marked hypoxemia | 0
ground-glass opacities in bilateral lower lung fields | 0
consolidation with GGO in bilateral lung fields | 0
negative urinary pneumococcal antigen test | 0
negative Legionella antigen test | 0
no significant bacteria in sputum culture | 0
no significant bacteria in blood culture | 0
drug-induced lung injury diagnosis | 0
methylprednisolone pulse therapy | 0
CRP decrease | 72
lung involvement improvement | 72
CRP elevation | 240
progressive bilateral diffuse extensive infiltrates | 240
tazobactam/piperacillin use | 240
micafungin use | 240
respiratory failure worsening | 336
death | 336
Corynebacterium spp. detected in tracheal sputum culture | 336
diffuse alveolar damage | 336
extensive fibrosis | 336
no evidence of bacterial pneumonia | 336
neutrophilic infiltration in tracheal epithelium | 336
mucosal hemorrhage | 336
ARDS diagnosis | 336
VAT diagnosis | 336
septic ARDS due to VAT conclusion | 336
