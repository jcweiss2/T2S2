33 years old | 0
    female | 0
    generalized anxiety disorder | 0
    right ankle pain | -48
    edema | -48
    fall | -72
    edema increased | -24
    edema migrated proximally to involve right leg | -24
    pain exacerbated by elevation | -24
    pain exacerbated by range of motion of ankle | -24
    pain exacerbated by weight-bearing | -24
    paresthesia throughout entire foot | -24
    denied fever | -24
    denied chills | -24
    denied shortness of breath | -24
    denied systemic symptoms | -24
    X-rays obtained | -24
    no evidence of acute osseous pathology | -24
    no soft-tissue gas | -24
    edema | 0
    erythema | 0
    tenderness to palpation | 0
    ecchymosis over lateral malleolus | 0
    compartments firm but compressible | 0
    mild pain with passive stretch | 0
    triphasic dorsalis pedis pulses | 0
    triphasic posterior tibial artery pulses | 0
    sensation intact but diminished | 0
    motor function intact | 0
    referred to emergency department | 0
    venous duplex ultrasound | 0
    no deep venous thrombosis | 0
    admitted to emergency room observation unit | 0
    serial compartment checks | 0
    improvement in emergency room | 0
    became hypotensive | 12
    became tachycardic | 12
    emergent trip to operating room | 12
    dual incision fasciotomy | 12
    dishwater fluid encountered | 12
    weakened fascia | 12
    tissue biopsy sent to pathology | 12
    fasciotomy sites copiously irrigated | 12
    wound VAC placed | 12
    transferred to SICU | 12
    requiring norepinephrine pressors | 12
    blood cultures positive for Gram-positive cocci | 18
    vancomycin started | 18
    clindamycin started | 18
    penicillin started | 18
    continued to deteriorate | 18
    hemodynamically unstable | 18
    requiring vasopressin | 18
    reevaluation 5 h post-operative | 23
    necrotic right foot | 23
    biopsy results revealed acute inflammation | 23
    biopsy results revealed necrosis | 23
    taken to operative room | 23
    necrosis of fascia | 23
    necrosis of subcutaneous fat | 23
    necrosis of muscle | 23
    guillotine amputation through tibia | 23
    incision over medial thigh | 23
    ascending infection | 23
    necrotic muscle | 23
    necrotic fat | 23
    necrotic fascia | 23
    guillotine amputation through mid-thigh | 23
    stabilized | 23
    managed on ceftriaxone | 23
    repeat irrigation and debridement | 24
    finalized above-knee amputation | 72
    ambulating with prosthesis | 5760
    