70 years old | 0
male | 0
admitted to ICU | 0
acute respiratory distress | 0
fever | 0
cerebrovascular accident | -2160
hemorrhagic stroke | -2160
anticoagulation therapy | -2160
acute pulmonary embolism | -2160
implantation of vena cava filter | -2160
hospital-acquired pneumonia | 0
severe sepsis | 0
hemodynamic collapse | 0
hypotension | 0
cold sweating | 0
hypoxia | 0
transthoracic echocardiography | 0
massive tricuspid insufficiency | 0
papillary muscle rupture | 0
suspected endocardial vegetation | 0
transesophageal echocardiography | 0
pericardial effusion | 0
cava filter migration into cardiac cavity | 0
open heart surgery | 12
tricuspid valve insufficiency | 12
metallic fragments between leaflets | 12
800 ml of blood in the pericardium | 12
migration of cava filter fragments | 12
tricuspid valve and vena cava filter fragments removed | 12
prosthetic tricuspid valve implanted | 12
recovered successfully | 24
discharged | 168