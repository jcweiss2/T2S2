52 years old | 0
male | 0
visit emergency department | 0
diffuse vesicular skin rash | 0
headache | 0
sore throat | 0
nausea | 0
contact with varicella zoster patients | -96
immunosuppressants | -6720
methotrexate | -6720
azathioprine | -6720
prednisolone | -6720
cutaneous leukocytoclastic vasculitis | -6720
denied prior history of chicken pox | 0
Vesicle Tzank smear | 0
Multinucleated giant cells | 0
herpes virus infection | 0
white blood cell count 4100/uL | 0
hemoglobin 14.8 gm/dL | 0
platelets 13,4000/uL | 0
serum creatinine 0.62 mg/dL | 0
Aspartate transaminase (AST) 782 U/L | 0
Alanine transaminase (ALT) 603 U/L | 0
total bilirubin 0.4 mg/dL | 0
prothrombin time 12.6 s | 0
C reactive protein 1.45 mg/L | 0
varicella zoster complicated with hepatitis | 0
oral famciclovir 500 mg | 0
discontinued immunosuppressive drugs | 0
discharged home | 48
outpatient clinics follow up | 48
visit emergency department again | 48
general malaise | 48
nausea | 48
acute ill looking | 48
alert | 48
temperature 36.2 °C | 48
blood pressure 54/46 mmHg | 48
pulse rate 102 beats/minute | 48
respiratory rate 20 cycles/min | 48
white blood cell 12700/uL | 48
hemoglobin 15.4 g/dL | 48
platelets 61000/uL | 48
prothrombin time 35.7 s | 48
actived partial thrombin time 44.5 s | 48
fibrinogen <50 mg/dL | 48
AST 8989 U/L | 48
ALT 6048 U/L | 48
total bilirubine 2.0 mg/dL | 48
indirect total bilirubin 1.5 mg/dL | 48
serum creatinine 2.99 mg/dL | 48
Blood arterial gas analysis | 48
PH 7.31 | 48
CO2 23 mmHg | 48
O2 83 mmHg | 48
HCO3 15.1 mm/L | 48
nasal cannula oxgen flow 5 L/min | 48
serum tests for possible causes of acute hepatitis | 48
Hepatitis B surface antigen (HbsAg) | 48
antibodies against hepatitis C (anti-HCV) | 48
anti-hepatitis A immunoglobulin M (IgM) antibody | 48
Epstein-Barr virus (EBV) viral capsid antigen IgM | 48
immunoglobulin G (IgG) | 48
serum Cytomegalovirus (CMV) IgM | 48
CMV IgG | 48
CMV pp65 antigen test | 48
serum Herpes simplex virus IgM | 48
serum HSV DNA PCR | 48
PCR test for VZV | 48
Vesicular base and serum viral isolation | 48
VZV | 48
serum VZV IgM | 48
serum VZV IgG | 48
admitted to an intensive care unit | 48
septic shock | 48
multiple organ failure | 48
disseminated intravascular coagulopathy | 48
aggressive fluid resuscitation | 48
broad-spectrum empirical antibiotics | 48
glycopeptide | 48
carbapenem | 48
blood transfusion | 48
intravenous acyclovir | 48
intubated | 50
comatose consciousness | 50
dyspnea | 50
profound shock | 50
lactate acidosis | 50
multiple organ failure | 50
expired | 72