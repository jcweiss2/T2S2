37 years old | 0
    male | 0
    healthcare worker | 0
    close contact with COVID-19 patient | -144 to -120
    high-grade fever | -168 to -144
    myalgia | -168 to -144
    dry cough | -168 to -144
    tested positive for COVID-19 | -168
    self-isolate at home | -168
    worsening shortness of breath | -144 to -120
    admitted to the hospital | 0
    bibasal crackles | 0
    gallop rhythm | 0
    resting tachycardia | 0
    no pedal oedema | 0
    lymphopaenia | 0
    raised CRP (74 mg/L) | 0
    lactate dehydrogenase (303 U/L) | 0
    BNP (247 pg/mL) | 0
    deranged liver function tests | 0
    normal haemoglobin | 0
    normal WBC count | 0
    normal electrolytes | 0
    normal renal function | 0
    negative cardiac troponins | 0
    sinus tachycardia on ECG | 0
    minimal bibasal infiltrates on chest X-ray | 0
    echocardiography (LVEF 10-15%) | 0
    dilated left ventricle | 0
    LV internal diameter end diastole (7.1 cm) | 0
    LV internal diameter end systole (6.3 cm) | 0
    high-grade temperature spikes (39°C-40°C) | 0
    CRP <100 mg/L | 0
    prescribed ceftriaxone | 0
    negative blood cultures | 0
    negative urine cultures | 0
    CRP increasing | 72
    no improvement in fever spikes | 72
    switched to piperacillin/tazobactam | 72
    vancomycin added | 72
    renal functions deteriorating | 72
    vancomycin levels normal | 72
    creatinine clearance worsening | 96
    GFR <10 mL/min/1.73 m² | 96
    creatinine (657 μmol/L) | 96
    oliguric | 96
    intermittent haemodialysis | 96
    renal biopsy planned | 96
    acute tubular injury | 96
    granular casts | 96
    localised inflammation | 96
    vancomycin discontinued | 96
    low-dose beta blocker | 0
    ACE inhibitor started | 0
    ACE inhibitor held | 72
    serial ECGs | 0
    serial TTEs | 0
    intravenous antibiotics | 0
    intermittent RRT (haemodialysis) | 96
    intensive care admission | 96
    symptom improvement | 336
    ejection fraction improved (25-30%) | 336
    renal function improving | 336
    no longer oliguric | 336
    dialysis discontinued | 336
    discharged | 336
    follow-up cardiac MRI (EF 46%) | 2064
    renal function normal | 4032
    advised to self-isolate | 336
    heart failure clinic follow-up | 720
    renal clinic follow-up | 1080
    negative cardiac troponins (days 0, 5, 21) | 0, 120, 504
    sinus tachycardia on ECGs (days 0, 5, 21) | 0, 120, 504
    premature ventricular contractions | 504
    no ischaemia | 504
    gradual EF improvement | 336
    cardiac MRI ordered | 504
    moderate LV impairment | 504
    no myocardial fibrosis | 504
    pre-COVID-19 cardiomyopathy considered | 504
    CRP creeping up | 72
    ceftriaxone changed | 72
    vancomycin discontinued (after 3 days) | 96
    vancomycin levels monitored | 96
    renal biopsy results | 96
    acute tubular necrosis/tubular injury | 96
    no glomerular change | 96
    AKI related to vancomycin exposure | 96
    intermittent haemodialysis for 8 days | 96
    volume input-output monitoring | 96
    symptom free at discharge | 336
    ejection fraction 25-30% at discharge | 336
    creatinine clearance recovery | 336
    advised follow-up in clinics | 720, 1080
    cardiac MRI at follow-up (EF 46%) | 2064
    renal function normal at follow-up | 4032