25 years old | 0
female | 0
returned from Ghana | -48
no prophylactics taken | -48
febrile | -48
diarrhea | -48
hypotension | -48
blood smear positive for malaria | -48
suspected Plasmodium falciparum | -48
normal hemoglobin | -48
high lactate dehydrogenase | -48
discharged with doxycycline | -48
returned to emergency department | -120
worsening symptoms | -120
inability to tolerate oral medications | -120
chills | -120
nausea and vomiting | -120
dizziness | -120
generalized malaise | -120
admitted to intensive care unit | -120
diagnosed with septic malaria | -120
diagnosed with influenza | -120
acute kidney injury | -120
elevated creatine | -120
elevated BUN | -120
elevated lactate | -120
received intravenous artesunate | 0
thrombocytopenic | 24
anemic | 24
received blood transfusions | 24
hemolytic anemia | 72
elevated reticulocyte count | 72
elevated LDH | 72
low haptoglobin | 72
discharged from hospital | 168
followed up with weekly labs | 168
elevated reticulocyte count | 336
elevated hemoglobin | 336
low haptoglobin | 336
low lactate dehydrogenase | 336
recovered from hemolytic anemia | 672