32 years old | 0
primigravida | 0
spontaneous dichorionic twin pregnancy | 0
admitted to emergency department | 0
preterm rupture of membranes of the first fetus | 0
20 weeks of gestation | 0
no relevant personal medical history | 0
blood type O Rh-positive | 0
ultrasound revealed two viable twins | 0
normal growth for gestational age | 0
oligohydramnios of the first fetus | 0
normal cervical length | 0
subserous uterine fibroid with 10 cm | 0
spontaneous onset of labor | -6
female baby weighing 340 g was vaginally delivered | -6
fetal death occurred within 1 h | -5
histopathological examination of the aborted fetus | -5
multi-organic congestion | -5
uterine contractions ceased | 0
cervix was reconstituted | 0
no signs of chorioamnionitis | 0
amniotic membrane of the second twin remained intact | 0
ultrasonography showed a healthy remaining fetus | 0
informed consent was obtained from parents | 0
umbilical cord of the first fetus was ligated high up in the cervix | 0
placenta was left inside the uterus | 0
cervical cultures were taken | 0
mother's perineum and vagina were disinfected with chlorhexidine | 0
patient remained in the hospital | 0
treated with bed rest | 0
low-molecular-weight heparin | 0
broad-spectrum antibiotics | 0
Ampicillin | 0
Gentamycin | 0
Amoxicillin | 11
no signs of infection | 0
serial ultrasonography revealed normal fetal growth | 0
wellbeing of the second twin | 0
digital vaginal examinations were avoided | 0
antenatal corticosteroids | -72
Betamethasone | -72
urgent cesarean section | 32*24
breech presentation | 32*24
onset of spontaneous labor | 32*24
685 g female neonate was delivered | 32*24
Apgar scores of 1/8/9 | 32*24
neonate received full resuscitation | 32*24
immediate life-support intervention | 32*24
admitted to the Neonatal Intensive Care Unit | 32*24
extreme prematurity | 32*24
extreme low birth weight | 32*24
Hyaline membrane disease | 32*24
patent ductus arteriosus | 32*24
satisfactory evolution | 90
spontaneous respiration | 90
mother developed postpartum sepsis | 32*24
endometritis | 32*24
admitted in the Intensive Care Unit | 32*24
remained for 4 days | 32*24+4
discharged | 32*24+12
child exhibited normal cognitive and neurological development | 15*30*24
low weight | 15*30*24
deficient physical development for age | 15*30*24
patent ductus arteriosus | 15*30*24