49 years old | 0
    male | 0
    presented to emergency department | 0
    worsening fever | -168
    cough | -168
    shortness of breath | -168
    febrile | 0
    temperature of 100.9°F | 0
    tachycardic | 0
    heart rate of 94 | 0
    hypoxic | 0
    SpO2 of 70% | 0
    chest X-ray revealed patchy opacities | 0
    placed on nasal cannula oxygen | 0
    SpO2 improved to 92%-95% | 0
    white blood cell count of 11.3 × 10^9/L | 0
    lactate dehydrogenase of 3,147 units/L | 0
    C-reactive protein of 265.9 mg/L | 0
    ferritin of 1,760 ng/mL | 0
    D-dimer of 124,802 ng/mL | 0
    admitted for acute hypoxic respiratory failure | 0
    suspected COVID-19 virus infection | 0
    SARS-CoV-2 RNA test positive | 0
    initial treatment with ceftriaxone | 0
    azithromycin | 0
    enoxaparin | 0
    dexamethasone | 0
    remdesivir | 0
    convalescent plasma therapy refused | 0
    inflammatory markers increased | 24
    started on tocilizumab | 24
    became acutely dyspneic | 336
    required nonrebreather mask | 336
    chest X-ray noted large right pneumothorax | 336
    mediastinal shift | 336
    CT-guided chest tube placement | 336
    8.5-French pigtail catheter inserted | 336
    repeat chest X-ray showed persistent right pneumothorax | 336
    second 22-French chest tube placed | 336
    chest X-ray showed mildly improved right pneumothorax | 336
    transferred to intensive care unit | 336
    antibiotic therapy broadened | 336
    immunosuppressive therapy continued | 336
    chest tube advanced to 36-French | 336
    CT chest noted large air-filled bullous process | 336
    suspicious for bronchopulmonary fistula | 336
    intubated | 336
    recommended right middle invasive thoracotomy | 336
    bronchopleural fistula repair | 336
    pleurodesis | 336
    large bronchopleural fistula documented | 336
    necrotic empyema | 336
    affected area repaired | 336
    resected | 336
    intraoperative specimens sent for pathological evaluation | 336
    initial cultures concerning for fungal process | 336
    started on amphotericin B | 336
    worsening respiratory failure | 504
    septic shock | 504
    marked bradycardia | 504
    asystole | 504
    microbiological analysis positive for Rhizopus species | 672
    <|eot_id|>
    