67 years old | 0
male | 0
admitted to the hospital | 0
malaise | -96
anorexia | -96
dry cough | -96
dyspnea | -96
severe respiratory distress | 0
oxygen saturation of 79% | 0
bilateral interstitial infiltrates | 0
right lower lobe consolidation | 0
shock | 0
elevated lactic acid | 0
endotracheal intubation | 0
mechanical ventilation | 0
fluid resuscitation | 0
antibiotics | 0
vasopressor support | 0
septic shock | 0
hepatocellular carcinoma | -672
rectal adenocarcinoma | -672
non-small-cell lung cancer | -672
surgical resections | -672
chemoradiation therapy | -672
remission | -720
chronic obstructive lung disease | 0
chronic kidney disease | 0
diabetes mellitus | 0
SARS-CoV-2 infection | 0
nasopharyngeal swab specimen | 0
real-time polymerase chain reaction | 0
positive result | 0
echocardiography | 0
preserved left ventricular ejection fraction | 0
severely dilated right ventricle | 0
reduced RV function | 0
flattening of the interventricular septum | 0
severe tricuspid regurgitation | 0
estimated systolic pulmonary artery pressure | 0
elevated D-dimer | 0
high-sensitivity troponin | 0
electrocardiogram | 0
normal sinus rhythm | 0
therapeutic anticoagulation | 0
venous thromboembolism | 0
venous duplex studies | 0
acute deep vein thrombosis | 0
computed tomographic angiography | 0
subsegmental right upper lobe pulmonary embolism | 0
neuromuscular blockade | 0
prone-position ventilation | 0
ARDS | 0
mechanical ventilatory support | 0
vasopressor support | 0
norepinephrine | 0
vasopressin | 0
acute kidney injury | 24
continuous renal replacement therapy | 24
shock liver | 24
gastrointestinal hemorrhage | 24
Escherichia coli pneumonia | 24
bacteremia | 24
comfort measures | 528
withdrawal of life-support interventions | 528
death | 528
acute RV dysfunction | 0
increased RV afterload | 0
acute cor pulmonale | 0
RV dilation | 0
septal dyskinesis | 0
RV dysfunction | 0
thrombolytic use | 0
extracorporeal support | 0
echocardiography | 0
point-of-care ultrasound | 0
transthoracic echocardiography | 0
POCUS examinations | 0
personal protective equipment | 0
disinfecting protocols | 0