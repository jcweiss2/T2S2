55 years old | 0
    man | 0
    alcohol use | 0
    necrotizing biliary pancreatitis | 0
    hospitalized 2 times over 3 months | -2160
    acute portal vein thrombus | -2160
    anticoagulation with therapeutic enoxaparin | -2160
    large multiloculated peripancreatic fluid collections | -2160
    WON | -2160
    EUS-guided cystogastrostomy procedures | -2160
    lumen-apposing metal stent placed | -2160
    double-pigtail catheter placed | -2160
    color Doppler imaging confirmed absence of interposed blood vessels | -2160
    underwent 2 endoscopic necrosectomies | -2040
    removal of initial lumen-apposing metal stent | -2040
    removal of pigtail catheter | -2040
    placement of 2 double-pigtail catheters | -2040
    subsequent necrosectomy | -1680
    replacement of double-pigtail catheters | -1680
    computed tomography imaging showed persistent WON | -1680
    worsening abdominal pain | 0
    fevers | 0
    admitted for sepsis from necrotizing pancreatitis | 0
    white blood cell count 29.6 | 0
    hemoglobin 8.7 g/dL | 0
    international normalized ratio 1.3 | 0
    became hypotensive | 120
    tachycardic | 120
    lactic acidosis | 120
    worsening anemia (hemoglobin 5.3 g/dL) | 120
    international normalized ratio 1.9 | 120
    activated partial thromboplastin time 26 | 120
    escalation to intensive care unit | 120
    retroperitoneal hematoma | 120
    intraperitoneal hemorrhage | 120
    enoxaparin discontinued | 120
    massive transfusion protocol | 120
    administration of protamine sulfate | 120
    temporary improvement in blood pressure | 120
    anemia continued to worsen | 120
    computed tomography angiography | 168
    small serpiginous area of internal arterial enhancement | 168
    active arterial bleeding into hematoma | 168
    angiogram identified L2 and L3 distal lumbar artery focal pseudoaneurysms | 168
    extravasation | 168
    coil embolization performed | 168
    additional angiographic evaluation | 168
    selective catheterization | 168
    imaging of celiac axis | 168
    imaging of right upper quadrant | 168
    imaging of superior mesenteric artery | 168
    imaging of right internal iliac artery | 168
    no focal pseudoaneurysm | 168
    no evidence of vasculitis | 168
    no active extravasation | 168
    blood pressure stabilized | 168
    transferred to tertiary care center | 168
    critical condition | 168
    continued blood transfusion requirements | 168
    exploratory laparotomy | 168
    evacuation of retroperitoneal hematomas | 168
    evacuation of intraperitoneal hematomas | 168
    large clots | 168
    active arterial bleeding | 168
    controlled with electrical cautery | 168
    subsequent surgeries for re-exploration | 168
    cholecystectomy | 168
    transfers to intensive care unit | 168
    hospital course complicated by nonobstructive ileus | 168
    pleural effusion | 168
    thoracentesis | 168
    bacteremia | 168
    hydronephrosis | 168
    4-week hospital stay | 672
    esophagogastroduodenoscopy performed | 672
    dilation of posterior cystogastrostomy | 672
    necrosectomy performed | 672
    2 double-pigtail stents left in place | 672
    no further complications | 672