73 years old | 0
male | 0
admitted to the hospital | 0
smoking 20 cigarettes a day | 0
occasional alcoholism to drunkenness | 0
recently diagnosed diabetes mellitus | 0
hypertension | 0
allergy to paracetamol | 0
no family history of hypertension | 0
no family history of diabetes mellitus | 0
no known genetic history | 0
no previous surgeries | 0
moderate to severe respiratory distress | -168
fever | -168
general malaise | -168
rapid test positive for SARS CoV-2 (IgM +, IgG +) | -168
management with oxygen | -168
management with steroids | -168
no anticoagulation | -168
severe abdominal pain | -48
nausea | -48
fecal emesis | -48
fever of 39.5 °C | -48
peritoneal irritation | -48
distention of intestinal loops | -48
inter-loop edema | -48
intestinal pneumatosis | -48
hemoglobin 15 g/dl | 0
leukocytes 17 thousand/cm3 | 0
platelets 120 thousand/cm3 | 0
procalciton of 26 ng/ml | 0
D-dimer>5000 ng/ml | 0
laparotomy | 0
resect 3-meter segment of small intestine (terminal jejunum and proximal ileon) | 0
end to end anastomosis | 0
purulent collection drained in the pelvis | 0
placement of drains | 0
management with antibiotics | 24
analgesic | 24
enoxaparin (60 mg/0.6 ml) every 24 h | 24
mechanical ventilation | 24
atrial fibrillation | 168
treated with amiodarone | 168
slight leakage of intestinal fluid | 240
intestinal fistula | 240
conservative treatment | 240
parenteral nutrition | 240
closing fistula at 3 weeks | 504
pathology report on ischemia and necrosis of the intestinal mucosa | 120
significant deterioration in lung function | 720
multi-organ failure | 720
dying 30 days after the procedure | 720
