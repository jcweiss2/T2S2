64 years old | 0
female | 0
admitted to the clinic | 0
cardiac evaluation | 0
increasing dyspnoea | -72
oedema of the lower limbs | -72
elevated NT-proBNP | 0
right axis deviation | 0
signs of right atrial enlargement | 0
history of carcinoid tumour | -10080
carcinoid tumour of the terminal ileum | -10080
hepatic metastasis | -10080
lymphatic metastasis | -10080
osseous metastasis | -10080
partial ileum resection | -10080
treated with somatostatin analogue | -10080
partial remission | -10080
computed tomography | 0
severe pulmonary stenosis | 0
torrential tricuspid regurgitation | 0
thickening and retraction of leaflets of the valves | 0
surgical valve replacement | 24
surgery | 24
postoperative course | 48
cardiac complications | 72
carcinoid crises | 72
pneumogenic sepsis | 72
broad-spectrum targeted anti-infective therapy | 72
intensive care measures | 72
therapy-refractory multi-organ failure | 120
death | 120