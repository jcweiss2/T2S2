41 years old | 0
male | 0
admitted to the hospital | 0
loss of olfactory sense | -504
loss of gustatory sense | -504
RT-PCR test for SARS-CoV-2 positive | -504
isolated at home | -504
returned to work | -462
annual medical checkup | -168
normal chest X-ray findings | -168
normal biochemical panel | -168
painful swelling of the left cervical lymph nodes | -144
high fever | -144
admitted to a local hospital | -144
computed tomography (CT) revealed an enlargement of the left cervical lymph nodes | -144
intravenous ceftriaxone | -144
oral prednisolone | -144
fever persisted | -144
painful cervical lymphadenopathy persisted | -144
fatigue | -120
poor appetite | -120
diarrhea | -120
dyspneic | -48
drowsy | -48
arterial oxygen saturation (SpO2) less than 90% | -48
hypotension | -48
oxygen supplementation | -48
noradrenaline | -48
contrast-enhanced CT revealed airspace consolidation | -48
enlargement of the right cervical and supraclavicular lymph nodes | -48
transferred to our hospital | 0
high fever | 0
hypotension | 0
enlarged right cervical lymph nodes | 0
bilateral conjunctivitis | 0
severe anasarca | 0
white blood cell count of 13.6×10^3 /mm^3 | 0
hemoglobin level of 11.9 g/dL | 0
platelet count of 28×10^3/mm^3 | 0
C-reactive protein (CRP) level of 34.62 mg/dL | 0
albumin level of 1.9 g/dL | 0
total bilirubin level of 4.8 mg/dL | 0
direct bilirubin level of 4.0 mg/dL | 0
aspartate aminotransferase level of 29 U/L | 0
alanine aminotransferase level of 66 U/L | 0
fasting triglycerides level of 297 mg/dL | 0
lactate dehydrogenase level of 161 U/L | 0
N-terminal pro-Brain Natriuretic Peptide (NT-pro BNP) level of 10,389 pg/mL | 0
D-dimer level of 3.86 μg/mL | 0
fibrinogen level of 703 mg/dL | 0
ferritin level of 2,350 ng/mL | 0
biopsy of the cervical lymph node | 24
bone marrow aspiration | 24
negative for human immunodeficiency virus (HIV) antibodies | 24
negative for hepatitis B surface antigen and antibody | 24
negative for hepatitis C virus (HCV) antibody | 24
negative for interferon-gamma release assay | 24
negative for rheumatoid factor | 24
negative for antinuclear antibody | 24
tests for Epstein-Barr virus (EBV)-specific antibodies suggested previous infection | 24
tests for Cytomegalo virus (CMV)-specific antibodies suggested previous infection | 24
echocardiography showed diastolic dysfunction | 24
left ventricular ejection fraction (EF) was 62% | 24
E/A ratio was 2.05 | 24
deceleration time was 111 milliseconds | 24
initiated levofloxacin | 24
initiated hydrocortisone 200 mg per day | 24
diuretics | 24
symptoms improved | 48
stopped norepinephrine treatment | 48
laboratory abnormalities improved | 48
IL-6 level of 4.18 pg/mL | 48
soluble interleukin-2 receptor (sIL-2R) level of 7,040 U/m | 48
discharged | 264
histopathological findings of the biopsy specimen of the cervical lymph nodes showed necrotizing lymphadenitis | 264
KFD diagnosed | 264
MIS-A diagnosed | 264