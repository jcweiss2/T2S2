61 years old | 0
male | 0
admitted to hospital | 0
fever | -168
muscle weakness | -168
fatigue | -168
family contacts tested positive for COVID-19 | -168
end-stage renal failure | -0
renal transplant | -0
type 2 diabetes mellitus | -0
cerebrovascular disease | -0
sleep apnea | -0
orthostatic hypotension | -0
benign prostatic hyperplasia | -0
transurethral resection of the prostate | -0
recurrent urinary tract infections | -0
mildly elevated temperature | 0
elevated pulse | 0
elevated blood pressure | 0
urinalysis positive for leucocytes | 0
urinalysis positive for nitrites | 0
urinalysis positive for trace amounts of blood | 0
treated for urosepsis | 0
developed low oxygen saturations | 24
tested positive for COVID-19 | 24
treated with dexamethasone | 24
treated with tocilizumab | 24
transferred to intensive care unit | 168
intubated | 168
hemodialysed | 168
persistent fluctuating low oxygen saturations | 168
computed tomography pulmonary angiogram | 216
saddle pulmonary embolus | 216
bilateral ground-glass attenuation | 216
patchy consolidation | 216
treated with low molecular weight heparin | 216
bilateral edematous eyelids | 264
ophthalmology opinion sought | 264
ocular examination | 264
bilaterally fixed and constricted pupils | 264
asymmetrical right-sided conjunctival injection | 264
chemosis | 264
visual acuity difficult to ascertain | 264
CT head with orbital imaging | 264
expanded and hyperdense right SOV | 264
asymmetrical hyperdensity of the venous structures | 264
swelling of the right pterygoid muscles | 264
effacement of the fat planes | 264
acute thrombosis of the right SOV | 264
acute thrombosis of the right pterygoid venous plexus | 264
dilated left SOV | 264
suspicion of bilateral caroticocavernous fistula | 264
treated with low molecular weight heparin | 264
extubated | 504
repeat interval imaging | 504
complete resolution of the right SOV thrombosis | 504
complete resolution of the pulmonary embolism | 504
marked improvement in lung parenchymal appearances | 504
preserved range of movement in eyes | 720
no diplopia | 720
no deficiency in visual acuity | 720
undergoing speech and language therapy | 720
undergoing physiotherapy | 720
undergoing rehabilitation | 720