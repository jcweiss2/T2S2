76 years old | 0 | 0 
female | 0 | 0 
admitted to the hospital | 0 | 0 
atrial fibrillation | -672 | 0 
rheumatic heart disease | -672 | 0 
congestive heart failure | -672 | 0 
digoxin | -168 | 0 
coumadin | -168 | 0 
generalized malaise | -168 | 0 
shortness of breath | -168 | 0 
lower extremity swelling | -168 | 0 
subjective fever | -168 | 0 
denies chest pain | -168 | 0 
denies orthopnea | -168 | 0 
denies paroxysmal nocturnal dyspnea | -168 | 0 
blood pressure 79/54 mmHg | 0 | 0 
oral temperature 38.3°C | 0 | 0 
heart rate 55 beats/min | 0 | 0 
crackles up to the mid-lung fields bilaterally | 0 | 0 
irregularly irregular heart rhythm | 0 | 0 
2+ pitting edema up to the knees | 0 | 0 
congestion in the bilateral lower lung fields | 0 | 0 
cardiomegaly | 0 | 0 
sodium level 126 | 0 | 0 
potassium 5.2 | 0 | 0 
blood urea nitrogen 33 | 0 | 0 
creatinine 2.77 | 0 | 0 
white blood count 4.9 | 0 | 0 
INR 2.8 | 0 | 0 
signs of digoxin toxicity | 0 | 0 
peak troponin level 0.20 ng/mL | 0 | 0 
digoxin level 3.6 ng/mL | 0 | 0 
given digoxin immune fab | 0 | 1 
ejection fraction 45% to 49% | 1 | 1 
possible vegetation on the mitral valve | 1 | 1 
severe eccentric mitral and tricuspid regurgitation | 1 | 1 
mitral valve vegetation measuring 1.2×0.7 cm | 1 | 1 
severe biatrial enlargement | 1 | 1 
left atrium volume 101.40 mL/m2 | 1 | 1 
right atrium volume 233.80 mL/m2 | 1 | 1 
blood cultures positive for Pasteurella multocida | 1 | 1 
ceftriaxone started | 1 | 432 
septic emboli | 1 | 432 
owned 4 cats | -672 | 0 
evaluated for multi-valve replacement surgery | 24 | 24 
biopsy of the vegetation | 24 | 24 
chose conservative treatment | 24 | 24 
condition stabilized | 168 | 168 
discharged to a skilled nursing facility | 168 | 168 
readmitted for congestive heart failure exacerbation | 720 | 720 
elected for hospice care | 720 | 720