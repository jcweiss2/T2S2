male | 0
newborn | 0
respiratory distress | 0
generalized edema | 0
tachycardia | 0
tachypnea | 0
hypotonia | 0
hypoactivity | 0
facial dysmorphic findings | 0
micropenis | 0
born at 37th gestational week | -168
cesarean section | -168
gestational diabetes | -168
tracheal intubation | 0
mechanical ventilation | 0
surfactant administration | 0
broad-spectrum antibiotics | 0
umbilical catheterization | 0
severe respiratory acidosis | 0
respiratory functions improvement | 72
continuous positive airway pressure | 72
enteral feeding | 72
no hypoglycemic attack | 72
generalized edema persistence | 120
poor feeding | 120
vomiting | 120
hypoactivity | 120
hypotonia | 120
mechanical ventilation | 168
metabolic screening | 168
normal portal | 168
normal splenic | 168
normal renal Doppler | 168
normal echocardiography | 168
central hypothyroidism | 168
low free-thyroxine | 168
elevated thyroid-stimulating hormone | 168
hyponatremia | 168
normal potassium levels | 168
low baseline cortisol | 168
low-dose adrenocorticotropic hormone test | 168
glucocorticoid replacement | 168
thyroid hormone replacement | 168
vomiting cessation | 192
hyponatremia improvement | 192
edema improvement | 192
extubation | 360
no supplemental oxygen | 552
gonadotrophic hormone levels below expected | 360
discharge | 720