28 years old | 0
African woman | 0
gravida 3 | 0
para 0 | 0
past medical history of one miscarriage | 0
past medical history of two abortions | 0
asymptomatic uterine leiomyomas | 0
largest leiomyoma measured 25 cm | 0
spontaneous abortion occurred at 14 weeks and 4 days | -336
referred to the Emergency Department | 0
fever | 0
significant pelvic pain | 0
fourteen days following spontaneous abortion | -336
temperature of 38.3°C | 0
pulse rate of 105/min | 0
blood pressure of 13.3/9.3 kPa | 0
respiratory rate of 16/min | 0
offensive vaginal loss | 0
abdominal tenderness | 0
painful palpation of a large myoma extending to the umbilicus | 0
raised C-reactive protein of 368 mg/L | 0
raised white cell count at 17 × 10⁹/L | 0
anemia with hemoglobin of 95 g/L | 0
platelets at 549 × 10⁹/L | 0
PT time at 68% | 0
blood cultures were negative | 0
ultrasonography demonstrated a significant heterogenous leiomyoma | 0
endometrial thickness of 10 mm | 0
contrast enhanced computed tomography scan | 0
large pelvic mass measuring 16 × 18 × 17 cm | 0
containing air | 0
heterogeneous tissue suggesting necrosis of a uterine fibroid | 0
three additional masses in the right lumbar region and iliac fossa measuring 10 cm, 5 × 3 and 5 × 4 cm diameter | 0
compatible with uncomplicated fibroids | 0
free intraperitoneal fluid in the right lumbar region and right iliac fossa | 0
not associated with any pneumoperitoneum | 0
provisional diagnosis of endometritis | 0
conservative treatment with broad spectrum antibiotics initiated | 0
Amoxicillin/clavulanic acid 1 g three times per day | 0
Ofloxacin 400 mg two times per day | 0
10 days of medical treatment | 240
deterioration of the patient’s clinical status | 240
persistent fever | 240
persistence of biological inflammatory syndrome | 240
C-reactive protein 440 mg/mL | 240
leukocytosis 20 × 10⁹/L | 240
procalcitonin 29 μg/L | 240
occurrence of bleeding disorders with a 49% PT time | 240
cholestasis | 240
PAL 235 UI/L | 240
GGT 307 UI/L | 240
electrolyte disorders | 240
persistent hypokaliemia at 2.35 mmol/L | 240
transferred to the intensive care unit | 240
repeat CT scan | 240
persistence of an aspect of reshapes of the necrobiotic myoma | 240
complicated with an abscess | 240
air fluid level | 240
exploratory laparotomy | 240
surgical exploration | 240
500 mL of a thick reddish-brown fluid | 240
multiple myomas | 240
largest myoma situated in an anterior position and sizing about 20 cm | 240
septic necrobiosis deforming the left side of the uterus | 240
level of the insertion of the left annex | 240
extensive dissection to free the uterus from adhesions | 240
selective myomectomy of a large myoma of 17 × 15 × 11 cm | 240
padding | 240
hemostatic knots using Vicryl suture | 240
extensive lavage of the peritoneal cavity with warm normal saline | 240
decided to preserve the uterus | 240
preserve the other uterine fibroids | 240
postoperative course was favorable | 240
IV antibiotic treatment with Tazocilline | 240
Metronidazole | 240
Amikacin | 240
relayed by Ofloxacin as a monotherapy regimen | 240
culture of the peritoneal fluid yielded no growth of bacteria | 240
histopathologic examination revealed a leiomyoma with advanced ischemic necrosis | 240
inflammation | 240
foci of abscess formation | 240
one month postoperative follow up | 720
resumption of regular and normal menses | 720
pain completely resolved | 720
pelvic ultrasound showed an increased volume of the uterus | 720
largest fibroid measuring 10 cm | 720
two years later | 17520
conceived spontaneously | 17520
fetal growth was normal | 17520
anterior placenta praevia (29 mm from the cervix) | 17520
cesarean section performed | 17520
previous myomectomy | 17520
adhesions on the anterior wall of the uterus | 17520
no signs of uterine rupture | 17520
corporeal hysterotomy performed | 17520
3320 g baby delivered | 17520
Apgar’s of 10 | 17520
post-operative recovery was unremarkable | 17520
