69 years old | 0
    woman | 0
    hypertension | 0
    type 2 diabetes mellitus | 0
    hypersensitivity pneumonitis | 0
    obesity | 0
    gastric band placement | 0
    right breast cancer | 0
    lumpectomy | 0
    chest pain | -12
    shortness of breath | -12
    diaphoresis | -12
    airlifted to emergency department | 0
    ST elevation | 0
    elevated troponin level >10,000 ng/dL | 0
    STEMI | 0
    aspirin | 0
    heparin | 0
    statin therapy | 0
    percutaneous coronary intervention | 0
    cardiac catheterization | 0
    right dominant circulation | 0
    100% occlusion LAD artery | 0
    aspiration thrombectomy | 0
    prasugrel | 0
    dual antiplatelet therapy | 0
    left upper quadrant abdominal pain | 24
    diaphoretic | 24
    short of breath | 24
    fever 103°F | 24
    tachycardia 109 bpm | 24
    hypotension 93/60 mmHg | 24
    leukocytosis WBC 16.5×10³ cells/L | 24
    lactate 1 mmol/L | 24
    CT abdomen | 24
    splenic infarct | 24
    high-grade stenosis celiac artery | 24
    mild thickening splenic flexure | 24
    transthoracic echocardiography | 24
    ejection fraction 40% | 24
    apical wall hypokinesia | 24
    mid/anteroseptal wall hypokinesia | 24
    trace pericardial effusion | 24
    no significant valvular pathology | 24
    distributive shock ruled out | 24
    hypovolemic shock ruled out | 24
    obstructive shock ruled out | 24
    cardiogenic shock | 24
    milrinone | 24
    Swan-Ganz catheter insertion | 24
    blood cultures collected | 24
    cefepime | 24
    metronidazole | 24
    vascular surgery consult | 24
    heparin infusion | 24
    CT angiography | 24
    blood cultures growth gram-positive cocci | 72
    leukocytosis WBC 26×10³ cells/L | 72
    vancomycin | 72
    repeat blood cultures | 72
    E. faecalis identification | 96
    susceptible to ampicillin | 96
    susceptible to gentamicin | 96
    susceptible to penicillin | 96
    ceftriaxone 2g twice daily | 96
    ampicillin every 4 hours | 96
    urinalysis | 96
    urine culture | 96
    afebrile | 120
    WBC count trending downward | 120
    trace leukocytes in urinalysis | 120
    negative nitrites in urinalysis | 120
    urine culture no growth | 120
    repeat blood cultures growth gram-positive cocci | 120
    repeat CT abdomen | 120
    repeat CT thorax | 120
    worsening bilateral pleural effusion | 120
    worsening pericardial effusion | 120
    DENOVA score ≥3 | 144
    TEE performed | 144
    vegetation on mitral valve | 144
    mild mitral regurgitation | 144
    no mitral stenosis | 144
    cardiothoracic surgery consult | 144
    E. faecalis in repeat cultures | 168
    pre-cardiac surgery workup | 168
    head CT subarachnoid hemorrhage | 168
    MRI multiple emboli left frontal lobe | 168
    MRI discitis | 168
    MRI osteomyelitis L1/L2 | 168
    carotid duplex <50% stenosis | 168
    right internal jugular vein thrombus | 168
    heparin withheld | 168
    septic emboli confirmed | 168
    unknown infection source | 168
    GI consult | 168
    general surgery consult | 168
    gastric band fluid aspiration | 168
    esophagogastroduodenoscopy | 168
    gastric mucosal atrophy | 168
    colonoscopy | 168
    rectosigmoid perforation | 168
    endoscopic closure | 168
    hypoxia | 168
    tachycardia | 168
    abdominal pain | 168
    diffuse abdominal tenderness | 168
    guarding | 168
    rebound tenderness | 168
    loss of pulse | 168
    noninvasive positive-pressure ventilation | 168
    epinephrine injection | 168
    exploratory laparotomy | 168
    no intraperitoneal contamination | 168
    extraperitoneal perforation rectum | 168
    end-colostomy | 168
    intensive care transfer | 168
    persistent fever | 168
    peritonitis | 168
    not candidate for mitral valve replacement | 168
    WBC 23×10³ cells/L | 168
    fever 102°F | 168
    hydrocortisone stress dose | 168
    hydrocortisone 100mg TID | 168
    vancomycin | 168
    piperacillin/tazobactam | 168
    no growth in blood cultures | 168
    no growth in tracheal aspirate | 168
    afebrile | 168
    ceftriaxone | 168
    ampicillin | 168
    ventilator-associated pneumonia | 168
    Stenotrophomonas maltophilia | 168
    acute kidney injury | 168
    inpatient rehabilitation | 168
    acute-on-chronic heart failure | 168
    cardiogenic shock | 168
    septic shock | 168
    multiorgan failure | 168
    death | 168

<|end_header_id|>

