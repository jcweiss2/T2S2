63 years old | 0
male | 0
alcoholic cirrhosis | -672
abdominal pain | -72
admitted to the hospital | 0
cachectic | 0
icteric | 0
holosystolic murmur | 0
abdomen diffusely tender | 0
abdomen distended | 0
erythematous macules | 0
purpuric macules | 0
papules | 0
white blood cell count of 16.8 k/uL | 0
hemoglobin of 10 g/dl | 0
platelets of 292 k/uL | 0
prothrombin time 27.8 s | 0
sodium of 125 mEq/L | 0
potassium of 4.8 mmol/L | 0
urea of 54 mg/dL | 0
creatinine 3.3 mg/dL | 0
bilirubin 9.1 mg/dL | 0
alanine transaminase (ALT) of 24 U/L | 0
aspartate transaminase (AST) of 76 U/L | 0
alkaline phosphatase of 93 U/L | 0
lactic acid dehydrogenase (LDH) 829 U/L | 0
total protein of 7.4 g/dL | 0
albumin of 2.6 g/dL | 0
INR of 2.3 | 0
Piperacillin and Tazobactam | 0
Vancomycin | 48
gram-positive cocci in clusters | 48
MSSA | 72
paracentesis | 0
ascitic fluid culture | 0
MSSA in ascitic fluid | 72
echocardiogram | 72
vegetation on the mitral valve | 72
cefazolin | 96
embolic events | 96
high Mayo surgical risk | 96
kidney function deterioration | 96
urine studies | 96
UNa of 79 mEq/L | 96
U creatinine of 50.2 mg/dL | 96
FENa of 4.1% | 96
daily electrocardiography (EKG) | 96
no AV block | 96
no persistent fever | 96
no bacteremia | 96
hepatorenal syndrome (HRS) | 120
octreotide | 120
midodrine | 120
albumin | 120
hemodialysis | 168
discharged to rehab | 336
long-term intravenous antibiotics | 336
repeat echocardiogram | 504
improvement in valve function | 504
clearance of vegetation | 504
refractory symptomatic ascites | 504
hepatic hydrothorax | 504
recurrent pleural effusion | 504
acute liver failure | 504
encephalopathy | 504
palliative peritoneal drainage catheter | 504
transjugular intrahepatic portosystemic shunt (TIPS) | 504
pre-TIPS bilirubin of 2.6 mg/dL | 504