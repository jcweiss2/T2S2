65 years old | 0
male | 0
ischemic cardiomyopathy | -8760
LVAD implantation | -8760
renal insufficiency | -8760
peritoneal dialysis | -8760
septic state | 0
high fever | 0
elevated inflammatory parameters | 0
C-reactive protein 16 mg/dL | 0
leukocytes 17G/L | 0
Staphylococcus aureus in blood cultures | 0
Staphylococcus aureus in peritoneal catheter | 0
right ventricular dysfunction | 0
inotropic support | 0
admission to intensive care unit | 0
driveline infection | 0
massive swelling of subcutaneous tunnel | 0
clean entrance site | 0
surgically opened driveline tunnel | 0
vacuum assisted closure therapy | 0
peritoneal catheter explanted | 0
peritonitis proven laparoscopically | 0
S. aureus identified at surgical site | 0
antibiotic treatment with vancomycin | 0
antibiotic treatment with tigecycline | 0
antibiotic treatment with meropenem | 0
VAC dressing changed every third day | 72
swabs returned sterile | 528
surgical closure of wound | 528
transfer to normal ward | 533
discharged home | 1320
readmitted to hospital | 3528
recurrence of driveline infection | 3528
wound reopened | 3528
debrided | 3528
negative pressure therapy initiated | 3528
VAC Veraflo therapy | 3528
instillation with 0.04% polyhexanide solution | 3528
dressing changed every third day | 3552
local debridement | 3552
surgical closure of wound | 3560
epicutaneous negative pressure wound therapy | 3560
antibiotic treatment with tazobactam/piperacillin | 3528
antibiotic treatment with rifampicin | 3528
discharged | 3864
free from signs of infection | 8760