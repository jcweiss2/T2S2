 \n\n

\boxed{
46 years old | 0 \\
female | 0 \\
decided to undergo elective sleeve gastrectomy | 0 \\
weighed 95 kg | 0 \\
BMI of 38.5 kg/m2 | 0 \\
past medical history of obesity | 0 \\
psoriatic arthritis treated with multiple immunosuppressants | 0 \\
surgical hypoparathyroidism | 0 \\
hypothyroidism following total thyroidectomy for multinodular goitre 20 years previously | -175200 \\
no history of diabetes | 0 \\
no history of dyslipidaemia | 0 \\
no history of hypertension | 0 \\
no history of obstructive sleep apnoea | 0 \\
hypoparathyroidism well managed on long term oral calcium carbonate and calcitriol | 0 \\
planned sleeve gastrectomy | 0 \\
converted to emergency Roux-en-Y gastric bypass surgery due to multiple gastric perforations because of friable mucosa | 96 \\
transferred to intensive care at a tertiary hospital | 96 \\
remained nil orally | 96 \\
calcium level critically low at 0.78 mmol/L | 96 \\
asymptomatic without seizure or arrhythmia | 96 \\
continuous intravenous calcium gluconate infusion required to achieve normocalcaemia | 96 \\
maintenance intermittent IV calcium boluses | 96 \\
prolonged ICU admission of 6 months | 96 \\
required more than 20 abdominal operations | 96 \\
received all medication and nutrition intravenously | 96 \\
lost 14 kg | 96 \\
endocrinology advice required throughout her admission | 96 \\
TSH was 5.83 mU/L | 336 \\
intravenous triiodothyronine (T3) 10 µg BD commenced | 336 \\
euthyroidism achieved after gradual up titration to 40/20/40 µg daily based on TSH levels | 336 \\
high dose intravenous calcium, 4.4 mmol five times daily required through a central line to maintain normocalcaemia | 336 \\
ionised calcium measured daily via routine blood gases | 336 \\
serum phosphate level 1.07 and remained in the normal range throughout the hospital admission | 336 \\
intravenous calcitriol 1 µg alternate daily commenced | 1008 \\
intravenous calcitriol ceased 5 days later due to limited stock and high cost | 1013 \\
150 000 units of intramuscular cholecalciferol trialled | 1344 \\
low 1,25(OH)vitamin D3 level failed to increment | 1344 \\
renal function normal with eGFR > 90 mL/min/1.73 m2 | 1344 \\
intravenous calcium gluconate 4.4 mmol five times daily required to maintain normocalcaemia | 2016 \\
additional intravenous calcitriol obtained and recommenced at a dose of 1 µg alternate daily | 2016 \\
gradually reduced calcium gluconate requirements to 4.4 mmol three times per day | 2016 \\
intramuscular thyroxine 600 µg trialled as a substitute for intravenous triiodothyronine | 2016 \\
patient found the injection painful | 2016 \\
intravenous thyroxine commenced at a dose of 200 µg alternate daily | 2020 \\
maintenance schedule that controlled both the hypocalcaemia and hypothyroidism established | 2020 \\
recommenced oral intake | 5760 \\
discharged on preoperative calcitriol dose (0.75 µg daily) and an increased dose of calcium (1200 mg orally twice daily) | 5760 \\
remained well replaced with normocalcaemia on review 6 weeks after discharge | 5904 \\
remained well replaced with normocalcaemia on review 12 weeks after discharge | 6048 \\
remained well replaced with normocalcaemia on review 4 months after discharge | 6720 \\
weighed 71.8 kg and had a BMI of 29 kg/m2 at 4-month follow up | 6720 \\
} \n\n

Note: The timestamps are calculated based on the provided narrative and the assumption that the admission event is the reference point (0 hours). The timestamps for events occurring before admission are negative, and those occurring after admission are positive. The exact timestamps for some events are approximated based on the context and clinical judgment. \n\n
For example, the event "converted to emergency Roux-en-Y gastric bypass surgery" is assumed to occur 4 days after admission, which is 96 hours. The event "TSH was 5.83 mU/L" is assumed to occur 2 weeks into her admission, which is 336 hours. \n\n
Please let me know if you need further adjustments or additional details. \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n
} \n\n