43 years old | 0
male | 0
admitted to emergency room | 0
history of consuming ALP | -2
abdominal pain | 0
bowel incontinence | 0
breathlessness | 0
heart rate of 113/min | 0
blood pressure of 60 systolic | 0
respiratory rate of 48/min | 0
saturation not recordable | 0
resuscitated with fluid bolus | 0
initiated on dual inotropes | 0
severe left ventricular dysfunction | 0
ejection fraction of 15% | 0
rapid sequence intubation | 0
severe metabolic acidosis | 0
pH of 6.98 | 0
bicarbonate of 8 | 0
lactate levels of 146 | 0
intravenous sodium bicarbonate administered | 0
intravenous magnesium sulfate administered | 0
heart rate dropped to 35/min | 1
intravenous atropine administered | 1
transient variable heart blocks | 1
venoarterial ECMO performed | 2
vitals stabilized | 2
shifted to intensive care unit | 2
decannulated | 72
bilateral cerebral vasculitis | 72
acute kidney injury | 72
renal replacement therapy initiated | 72
coagulopathy | 72
multiple blood transfusions | 72
lower respiratory tract infection | 72
minocycline started | 72
reactive pleural effusion | 72
intercostal drainage placed | 72
intercostal drainage removed | 120
discharged home | 984
no neurological deficits | 984
improving kidney function | 984