76 years old | 0
female | 0
admitted to the hospital | 0
neck pain | -744
productive cough with yellow sputum | -744
denied fever | -744
denied weight loss | -744
thyroid enlargement | -744
indurated texture | -744
no thyroid bruits | -744
lungs clear to auscultation | -744
thyrotropin level of 0.04 µIU/mL | -744
free thyroxine level of 1.64 ng/dL | -744
normal free triiodothyronine level | -744
peripheral blood leukocyte count 11.58 × 10^9/L | -744
erythrocyte sedimentation rate (ESR) 95 mm/hour | -744
solid nodule with intranodular calcifications | -744
subacute thyroiditis | -744
cefixime 0.1 mg | -744
ibuprofen 300 mg | -744
poor treatment response | -720
repeat thyroid function tests | -720
thyrotropin 0.02 µIU/mL | -720
free thyroxine 35.0 pmol/L | -720
free triiodothyronine 5.3 pmol/L | -720
thyroglobulin 78.93 ng/mL | -720
thyroxine receptor antibody 0.46 IU/L | -720
peripheral blood leukocyte count 16.87 × 10^9/L | -720
ESR 86 mm/hour | -720
neuron-specific enolase level 16.6 ng/mL | -720
bone collagen CYFRA21-1 level 11.16 ng/mL | -720
diffuse thyroid disease | -720
hypoechoic solid nodule with calcification | -720
polyglandular lymphadenopathy | -720
Graves’ disease | -8760
hyperthyroidism | -8760
adenomatoid thyroid nodules | -1752
chronic pharyngitis | -8760
type II diabetes mellitus | -8760
hypertension | -8760
cerebral infarction | -8760
pre-excitation syndrome | -8760
radiofrequency ablation | -8760
denied radiation exposure | 0
denied family history of thyroid diseases | 0
hospitalized | 0
oral prednisone acetate 10 mg | 0
rapid-acting insulin | 0
long-acting insulin | 0
oral metformin 0.5 g | 0
irbesartan 150 mg | 0
nifedipine controlled-release tablets 30 mg | 0
bisoprolol 5 mg | 0
rosuvastatin 5 mg | 0
aspirin 100 mg | 0
resolution of neck pain | 384
dysphagia | 384
choking cough | 384
dyspnea | 384
dysphonia | 384
tracheal stenosis | 384
polyglandular lymphadenopathy | 384
stroboscopic laryngoscopy | 384
painless gastroscopy | 384
partial thyroidectomy | 1344
tracheotomy | 1344
postoperative pathological examination | 1344
poorly differentiated malignant tumor | 1344
squamous cell carcinoma | 1344
extensive necrosis | 1344
inflammatory reaction | 1344
invasion of adjacent striated muscle | 1344
invasion of vasculature | 1344
invasion of nerves | 1344
immunohistochemistry | 1344
galectin-3 (+) | 1344
cytokeratin 19 (CK19; +) | 1344
CD56 (−) | 1344
Ki-67 (70% +) | 1344
p53 (−) | 1344
TTF-1 (minority +) | 1344
TG (−) | 1344
calcitonin (−) | 1344
synuclein (−) | 1344
CGA (−) | 1344
Pax8 (+) | 1344
vimentin (scattered +) | 1344
tumor metastasized to lungs | 1680
tumor metastasized to face | 1680
tumor metastasized to other anatomic sites | 1680
surgical site infection | 1680
multiple organ failures | 1680
sepsis | 2184
death | 2184