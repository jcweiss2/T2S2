38 years old | 0
male | 0
admitted to the hospital | 0
HBV-associated PAN | -6 months
medical history of HBV | -6 months
prednisolone | -6 months
cyclophosphamide | -6 months
Tenofovir | -6 months
stopped taking Tenofovir | -2 months
chronic renal failure | 0
diabetes mellitus Type II | 0
acute abdomen | 0
septic shock | 0
free sub diaphragmatic air | 0
peritonitis | 0
three perforations of the small intestine | 0
segmental enterectomy with anastomosis | 0
mechanical ventilation | 0
circulatory support | 0
acute-on-chronic renal failure | 0
weaned off the ventilator | 72
haemodynamically stable | 72
tenofovir orally | 72
IV methylprednisolone | 72
abdominal drain catheter presented enteric content | 168
second explorative laparotomy | 168
two new perforations | 168
multiple areas of patchy necrosis | 168
plasma exchanges | 168
IV cyclophosphamide | 168
IV methylprednisolone | 168
IV prednisone | 168
third laparotomy | 216
three new necrotic lesions | 216
necrotic lesion on the left lobe of the liver | 216
fourth laparotomy | 264
segmental enterectomy with anastomosis | 264
cholecystectomy | 264
anastomotic leak | 264
gangrenous gallbladder | 264
died | 360
septic shock | 360
multiple organ failure | 360
weight loss | -1 year
myalgias | -1 year
fever | -1 year
skin erythema | -1 year
deterioration of renal function | -1 year
new onset of diabetes mellitus Type II | -1 year
hypertension | -1 year
diagnosis of PAN and HBV infection | -6 months
HBsAg | 0
HBeAg | 0
Anti-HBcAb | 0
absence of Anti-HBsAb | 0
absence of Anti-HBeAb | 0