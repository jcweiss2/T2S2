86 years old | 0
male | 0
dementia | 0
hypertension | 0
transferred to the institution | 0
ST-segment elevation myocardial infarction | 0
cough | -168
shortness of breath | -168
no chest pain | -168
presented to outside institution | -168
acute hypoxic respiratory failure | -168
mechanical ventilation initiated | -168
transfer to our institution | -168
anteroseptal ST-segment elevation in precordial leads | -168
confirmed anteroseptal ST-segment elevation | 0
blood pressure 85/57 mmHg | 0
sedated | 0
intubated | 0
cardiopulmonary exam no abnormalities | 0
troponin 4.82 ng/mL | 0
creatinine 1.84 mg/dL | 0
lactate dehydrogenase 496 U/L | 0
C-reactive protein 173 mg/L | 0
chest radiography bilateral infiltrates at the bases | 0
no other abnormalities on chest radiography | 0
ST-segment elevations in leads V2 and V3 | 0
transthoracic echocardiogram ejection fraction 50-55% | 0
no significant regional wall motion abnormalities | 0
no signs of cardiac tamponade | 0
coronary angiography no significant coronary artery disease | 0
admitted to intensive care unit | 0
mechanical ventilation | 0
vasopressor support | 0
troponin increased to 7.84 ng/mL | 24
COVID-19 test positive | 72
respiratory status worsened | 120
required increased oxygen | 120
required positive end-expiratory pressure | 120
improvement with intravenous diuretics | 120
renal function worsened | 120
lymphopenia worsened | 120
inflammatory biomarker abnormalities worsened | 120
required higher amounts of oxygenation | 168
loss of R waves | 168
transient T wave inversions | 168
deepened Q waves | 168
worsening kidney injury | 192
D-dimer level rise | 192
family decided to pursue comfort care measures | 192
patient died | 192
