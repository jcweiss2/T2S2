31 years old | 0
male | 0
admitted to the hospital | 0
fatigue | -160
dizziness | -160
profuse sweating | -160
tremor of hands | -160
tremor of calves | -160
burning sensations in the feet | -160
freezing sensations in the feet | -160
maculopapular rash | -160
elevated liver transaminases | 0
enlarged liver | 0
nonsignificant hyponatremia | 0
diagnosed and treated by a family doctor | -160
diagnosed and treated by an occupational medicine physician | -160
hospitalized for 4 days in a regional hospital | -160
acute mercury vapour poisoning excluded | 0
dizziness | 0
tremor | 0
ataxia | 0
dysarthria | 0
dysphagia | 0
urinary retention | 0
stool retention | 0
diminished deep tendon reflexes | 0
hyponatremia | 0
encephalopathy diagnosed | 0
polyradiculoneuropathy diagnosed | 0
urine sample for mercury test sent | 0
neuro-diagnostic tests performed | 0
brain CT normal | 0
brain MRI abnormal | 0
EEG abnormal | 0
EMG I abnormal | 5
EMG II abnormal | 81
EMG III abnormal | 168
CSF abnormal | 7
antiviral treatment started | 0
antibiotic treatment started | 0
intravenous immunoglobulin treatment started | 0
increased extremity paresthesias | 28
burning sensation of the soles | 28
peripheral facial nerve neuropathy | 28
progressive lower extremity weakness | 28
acute respiratory failure | 28
intubated | 28
mechanical ventilation started | 28
chelation therapy with penicillamine started | 28
transferred to ICU | 28
continuous venovenous hemodiafiltration started | 28
2,3-dimercaptopropane-1-sulfonate treatment started | 28
crackles of subcutaneous emphysema | 28
pneumomediastinum detected | 28
atelectasis detected | 28
consolidation in the lower segments of the left lung | 28
endoscopic examination performed | 28
thick, purulent secretions in the bronchi | 28
mechanical ventilation used for almost 5 months | 28
weaned off the ventilator | 140
control CT scan performed | 140
complete resolution of the air from the mediastinum and neck | 140
progression of pneumonia in the left lung | 140
septic shock developed | 140
multiresistant Acinetobacter baumannii cultured | 140
limb weakness progressed to almost complete tetraplegia | 140
flaccid paralysis | 140
persistent diarrhoea | 140
recurrent Pseudomonas urinary tract infections | 140
formation of multiple urinary calculi | 140
drenching sweats | 140
profound hypovolemia | 140
transient loss of consciousness | 140
intravenous spironolactone added to the penicillamine treatment | 90
tetraplegia began to subside | 113
able to move all extremities | 113
able to stand by the bedside with assistance | 113
weaned off the ventilator | 113
tracheostomy tube removed | 113
EMG showed significant improvement | 113
mercury urine concentration decreased to normal level | 196
return to normal gastrointestinal and urinary functioning | 196
discharged home | 196