35 years old | 0
male | 0
presented to the emergency department | 0
polydipsia | -168
generalized weakness | -168
light headedness | -168
visual disturbances | -168
diabetic ketoacidosis | 0
blood glucose 600 mg/dL | 0
arterial blood pH 7.26 | 0
beta-hydroxybutyrate level greater than 46.8 mg/dL | 0
anion gap 27 mmol/L | 0
hemoglobin A1c 11% | 0
mild leukocytosis 12,250 cells/mcl | 0
admitted to the intensive care unit | 0
intravenous fluids | 0
insulin infusion | 0
transferred to the medical floor | 24
transitioned to subcutaneous insulin | 24
fever 101.6 °F | 24
severely altered mental status | 24
unable to follow multistep commands | 24
unable to tell time on a standard clock | 24
unaware of where he was | 24
unaware of details regarding his hospitalization | 24
unaware of the current President of the United States | 24
auditory hallucinations | 24
visual hallucinations | 24
generalized muscle soreness | 24
neck stiffness | 24
impaired finger to nose testing in both upper extremities | 24
intermittent dysconjugate gaze during extraocular eye movements | 24
no nuchal rigidity | 24
Kernig’s sign negative | 24
Brudzinski’s sign negative | 24
chest radiograph negative for acute cardiopulmonary pathology | 24
computed tomography imaging of the head negative for acute intracranial process | 24
magnetic resonance imaging of the brain negative | 24
lumbar puncture performed | 24
cerebrospinal fluid (CSF) analysis elevated protein 74 mg/dL | 24
CSF normal glucose 95 mg/dL | 24
CSF 14 red blood cells per microliter | 24
CSF 10 white blood cells per microliter | 24
CSF lymphocytes | 24
CSF Gram stain negative for organisms | 24
CSF Herpes virus PCR negative | 24
CSF Enterovirus PCR negative | 24
blood cultures sent | 24
urine cultures sent | 24
urine analysis large blood | 24
urine analysis 2 red blood cells per high power field | 24
possible myoglobinuria | 24
creatine kinase 19,154 U/L | 24
vancomycin started | 24
cefepime started | 24
mental status gradually improved | 96
hallucinations resolved | 96
creatine kinase rose to 118,400 U/L | 96
weakness improved | 96
muscle tenderness mild | 96
muscle tenderness only reproducible with deep palpation | 96
vastus lateralis muscle biopsy obtained | 96
muscle biopsy rare hypotrophic fibers | 96
muscle biopsy no evidence of rhabdomyolysis | 96
muscle biopsy no evidence of myopathy | 96
muscle viral myositis panel sent | 96
paraneoplastic panel sent | 96
CSF culture negative | 96
blood culture negative | 96
urine culture negative | 96
vancomycin stopped | 96
cefepime stopped | 96
continued to improve | 96
fever did not recur | 96
creatine kinase started to decrease | 96
muscle tenderness resolved | 96
discharged home | 264
no neurological deficits | 264
CSF IgM antibodies to West Nile Virus positive | 264
CSF IgG antibodies to West Nile Virus positive | 264
muscle viral panel negative | 264
paraneoplastic panel negative | 264
West Nile Virus encephalitis diagnosis | 264
