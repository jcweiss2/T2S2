71 years old | 0
male | 0
Saudi | 0
rheumatic heart disease | -672
hypertension | -672
chronic kidney disease | -672
admitted to the hospital | 0
anemia | 0
weight loss | 0
gradual decline in vision | -672
no eye redness | -672
no photophobia | -672
no floaters | -672
no flashes | -672
no scotoma | -672
no previous history of eye trauma | -672
no previous history of eye surgery | -672
raw milk ingestion | -672
informed consent | 0
full medical care | 0
treatment | 0
surgical management | 0
chemotherapy treatment | 0
referred to the ophthalmologist | 0
visual acuity 6/200 | 0
visual acuity 20/200 | 0
intraocular pressure 13 mmHg | 0
intraocular pressure 15 mmHg | 0
external examination normal | 0
extra-ocular movements normal | 0
pupils reactive to light | 0
no relative afferent pupillary defect | 0
deep and quite anterior chamber | 0
pinkish hypopyon | 0
iris pigments on the surface of the lens | 0
irregular pupil | 0
posterior synechiae | 0
visually significant nuclear sclerotic cataract | 0
multiple corneal scars | 0
obscuring the dilated fundus exam | 0
extensive systemic work-up | 0
infectious and inflammatory etiologies | 0
three sets of blood culture negative | 0
three sets of sputum culture negative | 0
three sets of urine culture negative | 0
repeated cultures for acid fast bacilli negative | 0
brucella titer negative | 0
B-Scan ultrasonography | 0
flat retina | 0
no vitritis | 0
no subretinal infiltrate | 0
fundus photos | 0
fundus Fluorescein angiography | 0
poor view due to cataract | 0
ultrasound Biomicroscopy | 0
floating cells in the AC | 0
hypopyon | 0
prednisolone acetate 1% drops | 0
cyclopentolate 0.5% drops | 0
left cataract extraction | 24
intraoperative diagnostic paracentesis | 24
atypical small to medium lymphoid cells | 24
blastoid morphology | 24
immunohistochemical staining | 24
T-cell lymphoma | 24
flow cytometry analysis | 24
CD5 positive | 24
CD3 positive | 24
CD2 positive | 24
CD8 positive | 24
CD56 positive | 24
CD4 negative | 24
CD7 negative | 24
CD10 negative | 24
CD34 negative | 24
alpha and beta T-cell receptor positive | 24
gamma T-cell receptor negative | 24
postoperative follow up | 48
visual acuity dropped | 48
counting fingers at 3 feet | 48
intraocular pressure normal | 48
anterior segment examination | 48
reforming pinkish hypopyon | 48
IOL in place | 48
dilated fundus exam | 48
hazy view due to cataract | 48
whitish retinal infiltrate | 48
multiple areas | 48
radiologic investigations | 48
chest x-ray | 48
pulmonary edema | 48
liver ultrasound | 48
heterogeneous liver | 48
no definite mass lesion | 48
computed tomography | 48
large heterogeneous left adrenal mass | 48
suspicious for invasion | 48
consistent with malignancy | 48
no other suspicious lesions | 48
ultrasound guided biopsy | 72
adrenal mass biopsy | 72
infiltration with atypical small to medium lymphoid cells | 72
blastoid features | 72
T-lymphocytes marker CD3 positive | 72
B-lymphocytic marker CD20 negative | 72
haemato-oncology team consultation | 72
chemotherapy regimen | 72
cyclophosphamide | 72
oncovin | 72
prednisolone | 72
lumbar puncture | 96
cerebrospinal fluid negative | 96
bone marrow biopsy | 96
negative for malignancy | 96
PET scan | 96
increase uptake in right nasal and ethmoidal sinuses | 96
lymphoma related | 96
high uptake in scrotum and testicles | 96
metastatic involvement | 96
ultrasonography of scrotum and testicles | 96
local radiotherapy | 120
orbits | 120
testicles | 120
chemotherapy continued | 168
atrial fibrillation | 168
stabilized | 168
transferred to Medical Intensive Care Unit | 168
regular ophthalmic bedside follow up visits | 168
collapsed | 192
unresponsive | 192
impalpable pulse | 192
cardiopulmonary resuscitation | 192
Advanced trauma life support protocols | 192
intubated | 192
deeply comatose | 192
Glasgow Coma scale 6/15 | 192
sepsis | 192
treated with antibiotics | 192
chemotherapy and radiation on hold | 192
Glasgow Coma scale 3/15 | 216
Do not attempt resuscitation | 216
passed away | 216