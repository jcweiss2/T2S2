history of chronic eczema | -720
history of previous alcohol abuse | -720
history of gout | -720
history of hypothyroidism | -720
psychosocial habits included 1 to 2 glasses of wine a day | -720
psychosocial habits included smoking | -720
no significant family history | 0
not on any medications | 0
cutaneous eruption began | -720
desquamation of the hands | -720
desquamation of the feet | -720
desquamation of the perioral skin | -720
desquamation of the perineal skin | -720
associated pain | -720
associated swelling | -720
concurrent hair loss | -720
increasing weakness | -576
fatigue | -576
intermittent diarrhea | -576
unintentional weight loss | -576
admitted to the emergency department | 0
dermatologic examination found erythematous desquamative patches | 0
dermatologic examination found erosions | 0
dermatologic examination found crusted lesions | 0
diffuse nonscarring alopecia of the scalp | 0
scaling patches on the vermillion lips | 0
punch biopsy of the left medial thigh | 0
psoriasiform epidermal spongiosis | 0
superficial perivascular lymphohistiocytic infiltrate | 0
diffuse hypogranulosis | 0
broad overlying parakeratosis | 0
ballooning degeneration of the spinous layer | 0
methicillin-resistant Staphylococcus aureus sepsis | 24
Escherichia coli sepsis | 24
pneumonia | 24
admitted to the intensive care unit | 24
required ventilator respiratory support | 24
systemic antibiotics | 24
laboratory and imaging studies ruled out necrolytic acral erythema | 48
laboratory and imaging studies ruled out pellagra | 48
laboratory and imaging studies ruled out biotin deficiency | 48
low zinc levels | 48
positive antitransglutaminase antibodies | 48
positive antiendomysium antibodies | 48
focal villi blunting | 48
Brunner's gland hyperplasia | 48
treated with a gluten-free diet | 72
treated with zinc sulfate | 72
resolution of gastrointestinal symptoms | 96
resolution of cutaneous symptoms | 96