76 years old | 0
male | 0
admitted to the hospital | 0
history of poorly controlled diabetes | 0
congestive heart failure | 0
hypertension | 0
hyperlipidemia | 0
sore throat | -24
went to a walk-in clinic | -24
negative rapid strep test | -24
prescription for penicillin | -24
became very weak | -12
unable to walk | -12
presented to the emergency room | 0
temperature 102.7°F | 0
pulse 131 | 0
respiration 40 | 0
blood pressure 126/73 | 0
oxygen saturation 96 percent | 0
complained of sore throat | 0
difficulty swallowing | 0
hoarseness | 0
cough | 0
no cervical lymphadenopathy | 0
no tenderness | 0
no pharyngeal erythema | 0
diminished lung sounds at the bases | 0
evaluated by an otolaryngologist | 0
flexible fiber optic laryngoscopy | 0
mild edema and erythema of bilateral aryepiglottic folds | 0
mild post-cricoid edema | 0
bilateral lower extremities edema | 0
treated with Dexamethasone | 0
treated with vancomycin hydrochloride | 0
treated with ceftazidime | 0
treated with Clindamycin | 0
rapid strep test negative | 0
lower respiratory culture grew out beta-hemolytic streptococcus group A | 12
blood culture grew out beta-hemolytic streptococcus group A | 12
Centor score 2 | 0
Centor score modified to 1 | 0
antibiotic regimen narrowed to ceftriaxone | 12
responded well to antibiotic therapy | 24
discharged to a short-term rehabilitation unit | 24
completed treatment course without complications | 168