85 years old | 0
female | 0
spontaneous perforation of the thoracic oesophagus | -168
episode of vomiting | -168
seven days lasting discomfort | -168
moderate fever | -168
clinical conditions progressively deteriorated | -168
CT scan showing lower para-oesophageal pleuro, mediastinal collection with fluid and air | -168
thickened wall of the oesophagus | -168
diagnosed with perforated oesophageal cancer | -168
advised with no treatment except for palliation of symptoms | -168
referred to our hospital | -168
conscious on admission | 0
normal breathing on admission | 0
moderately febrile on admission | 0
normal blood pressure | 0
normal heart rate | 0
white blood cell count of 11,100 cells/μL | 0
C-reactive protein of 243 mg/L | 0
minimal biochemical signs of liver impairment | 0
minimal biochemical signs of renal impairment | 0
accurate anamnesis | 0
episode of vomiting seven days before admission | -168
fever | -168
malaise | -168
continued to feed orally | -168
CT scan showing oral contrast spreading into para-oesophageal mediastinal and left pleural collection | 0
left thoracotomy performed | 0
smelly purulent collection opened and debrided | 0
lower lobe of the lung trapped | 0
necrotic tissues removed | 0
distal third of the oesophagus isolated down to the hiatus | 0
perforation of about 3 cm near gastro-oesophageal junction | 0
muscular layer around perforation diffusely necrotic | 0
necrotic muscular layer removed | 0
mucosal layer exposed | 0
bulging edges of tear inflamed | 0
bulging edges of tear edematous | 0
two stay sutures placed at ends of rupture | 0
mucosal edges grasped with Allis clamp | 0
endoscopic articulating linear cutter placed twice on healthy mucosa | 0
seal tested | 0
nasogastric tube left in stomach | 0
hiatus slightly opened | 0
limited portion of gastric fundus gained | 0
gastric wrap secured over repaired mucosa | 0
lower lobe of the lung decorticated | 0
three chest drainages left in place | 0
Escherichia coli cultured from pleural fluid | 0
Enterococcus faecalis cultured from pleural fluid | 0
postoperative left lower lobe pneumonia | 24
postoperative systemic infection by multidrug-resistant Klebsiella pneumoniae | 24
CT scan on postoperative day 9 confirming seal of repair | 216
excluded residual collections on postoperative day 9 | 216
resumed creamy diet | 216
chest drains removed on postoperative day 11 | 264
discharged home on postoperative day 27 | 648
oesophagogram performed after one month | 648
