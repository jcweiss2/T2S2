66 years old | 0
male | 0
dual-chamber pacemaker | -1296
sick sinus syndrome | -1296
paroxysmal atrial fibrillation | -1296
severe lumbar back pain | 0
mental status changes | 0
hypotension | 0
acute renal failure | 0
hypoxemic respiratory failure | 0
emergent intubation | 0
severe sepsis | 0
hemodynamic support | 0
vasopressin | 0
norepinephrine | 0
blood cultures | 0
methicillin-sensitive Staphylococcus aureus | 0
vancomycin | 0
nafcillin | 0
transthoracic echocardiogram | 0
left ventricular ejection fraction | 0
patent foramen ovale | 0
Doppler of the intra-atrial septum | 0
computed tomography scan | 0
osteomyelitis | 0
magnetic resonance imaging | 0
septic emboli | 0
transesophageal echocardiogram | 0
vegetation | 0
right atrium | 0
pacemaker lead | 0
tricuspid valve | 0
right ventricle | 0
cardiothoracic surgery | 0
surgical intervention | 0
laser lead extraction | 0
Indigo Penumbra system | 0
intracardiac echocardiography | 0
aspiration catheter | 0
vegetation removal | 0
anticoagulation | 0
venovenous bypass | 0
AngioVac system | 0
femoral veins | 0
GORE DrySeal Flex introducer sheath | 0
CARTO SoundStar catheter | 0
Indigo CAT8 XTORQ catheter | 0
aspiration pump | 0
vacuum | 0
blood loss | 72
pathology | 72
gram-positive cocci | 72
methicillin-sensitive Staphylococcus aureus | 72
tissue necrosis | 120
lactic acidosis | 120
worsening renal failure | 120
withdraw care | 120
extubation | 120
death | 120