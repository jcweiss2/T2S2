22 years old | 0
male | 0
admitted to intensive care unit | 0
high-grade fever | -72
hypoxic respiratory failure | -72
ventilatory support | 0
elevated white blood cell count | 0
elevated procalcitonin | 0
elevated troponin | 0
myocarditis | 0
pneumonia | 0
sepsis | 0
fever | -72
sore throat | -72
generalized weakness | -72
myalgia | -72
abdominal pain | -72
treated as outpatient | -72
tachycardia | 0
febrile spikes | 0
tachypnea | 24
tachycardia | 24
chest pain | 24
electrocardiogram showed global ST depression | 24
elevated troponin I | 24
intubated | 24
respiratory distress | 24
2D echo showed new onset global hypokinesia | 24
antimicrobials upgraded | 24
suspecting pneumonia with sepsis and myocarditis | 24
infective causes evaluated | 24
blood cultures negative | 48
throat swab for H1N1 negative | 48
diphtheria negative | 48
febrile spikes persisted | 48
upper abdominal pain | 48
tachycardia | 48
repeat 2D echo normalized | 72
troponin I decreased | 72
hemodynamics maintained | 72
contrast-enhanced computed tomography of the chest and abdomen | 72
bilateral basal consolidation | 72
baseline PCT level elevated | 72
Leptospira negative | 96
dengue negative | 96
malarial parasite negative | 96
HIV negative | 96
hepatitis C virus negative | 96
HbsAg negative | 96
scrub typhus negative | 96
Brucella serology negative | 96
antinuclear antibody negative | 96
ANA profile negative | 96
rheumatoid arthritis negative | 96
C-ANCA negative | 96
P-ANCA negative | 96
antistreptolysin O titers negative | 96
transesophageal echocardiography negative | 96
antibiotics upgraded to colistin | 120
Acinetobacter isolated from bronchoalveolar lavage cultures | 120
febrile spikes continued | 120
episodes of pulmonary edema | 120
serial PCT levels elevated | 120
failed extubation | 168
reintubated | 168
repeat computed tomography chest consistent with prior findings | 168
septic polymerase chain reaction panel negative | 168
bone marrow biopsy and cultures inconclusive | 168
C-reactive protein elevated | 168
serum ferritin levels elevated | 168
initiated on steroids | 192
initiated on nonsteroidal anti-inflammatory drugs | 192
febrile spikes subsided | 192
PCT levels decreased | 192
extubated | 312
steroids tapered | 312
discharged | 480
rheumatic fever | -6048
penicillin prophylaxis | -6048
penicillin prophylaxis stopped | -5040