65 years old | 0 | 0 
female | 0 | 0 
admitted to the hospital | 0 | 0 
fever | 0 | 48 
chills | 0 | 48 
pain in left leg | 0 | 48 
parkinsonism | -8760 | 0 
diabetes mellitus | -8760 | 0 
levodopa / carbidopa | -8760 | 0 
rasagiline | -8760 | 48 
ropinirole | -8760 | 0 
trihexyphenidyl | -8760 | 0 
amantadine | -8760 | 0 
metformin | -8760 | 0 
glipizide | -8760 | 0 
cellulitis | 0 | 0 
intravenous clindamycin | 0 | 48 
intravenous benzylpenicillin | 0 | 48 
high-temperature spikes | 48 | 48 
tachycardia | 48 | 48 
tachypnea | 48 | 48 
hypotensive | 48 | 48 
encephalopathic | 48 | 48 
shifted to ICU | 48 | 48 
intravenous linezolid | 48 | 96 
intravenous piperacillin with tazobactam | 48 | 96 
vancomycin not considered | 48 | 48 
hemodynamics improved | 48 | 48 
inotropic supports | 48 | 96 
oral hypoglycemic agents stopped | 48 | 48 
insulin started | 48 | 240 
confused | 48 | 96 
drowsy | 48 | 96 
disoriented | 48 | 96 
altered sensorium | 48 | 96 
myoclonus | 48 | 96 
tremors | 48 | 96 
jerky movements | 48 | 96 
no neck stiffness | 48 | 48 
computed tomography of the brain | 48 | 48 
cerebrospinal fluid analysis | 48 | 48 
improving white blood cell counts | 48 | 96 
better glycemic control | 48 | 96 
sterile blood and pus cultures | 48 | 96 
serotonin syndrome suspected | 96 | 96 
linezolid and rasagiline stopped | 96 | 96 
temperature settled | 104 | 104 
heart rate normal | 104 | 104 
sensorium improved | 104 | 104 
tremors subsided | 104 | 104 
shifted out of ICU | 192 | 192 
started walking with support | 240 | 240 
discharged from hospital | 240 | 240 
anti-parkinsonism drugs continued | 240 | 0 
rasagiline added | 240 | 0 
regular follow-up with neurologist | 240 | 0 
stable and asymptomatic for serotonin syndrome | 240 | 0