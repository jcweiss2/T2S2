81 years old | 0
    male | 0
    admitted to internal medical department | 0
    longstanding inguinoscrotal hernia | -8760
    upper abdominal pain | 0
    auricular fibrillation | -8760
    chronic heart failure | -8760
    chronic renal dysfunction | -8760
    temperature 36.1°C | 0
    abdominal distention | 0
    epigastric tenderness | 0
    bilateral giant inguinoscrotal hernia | 0
    no tenderness | 0
    no redness | 0
    white blood cell count 4900/mm² | 0
    C-reactive protein 1.2 mg/dl | 0
    creatinin 1.71 mg/dl | 0
    prothrombin time 18.7 s | 0
    PT-INR 1.61 | 0
    computed tomography slightly dilated stomach | 0
    computed tomography slightly dilated jejunum | 0
    bilateral inguinoscrotal hernia containing small bowel | 0
    bilateral inguinoscrotal hernia containing cecum | 0
    bilateral inguinoscrotal hernia containing ascending colon | 0
    bilateral inguinoscrotal hernia containing sigmoid colon | 0
    no remarkable occlusion point | 0
    acute entire abdominal pain | 48
    blood pressure decreased to eighties | 48
    CT scan free air right inguinal hernia sac | 48
    much ascites | 48
    diagnosis acute generalized peritonitis | 48
    diagnosis small bowel perforation in inguinal hernia sac | 48
    emergency operation performed | 48
    mid-lower median abdominal incision | 48
    transverse incision right inguinal area | 48
    dirty ascites inguinal sac | 48
    cecum perforation | 48
    terminal ileum necrotic 100 cm behind Bauhin’s valve | 48
    lateral extension internal hernia ring | 48
    mobilization pancreas head | 48
    mobilization duodenum | 48
    mobilization right side of colon for right hemicolectomy | 48
    substantial amount of bile | 48
    rupture inferior duodenum angle | 48
    right hemicolectomy | 48
    side-to-side anastomosis duodenum and jejunum | 48
    primary closure peritoneum hernia gate | 48
    transferred to intensive care unit | 48
    septic shock | 432
    leakage duodenum–jejunum anastomosis | 432
    use several antibiotic agents | 432
    use vasopressure agent | 432
    continuous hemodiafiltration | 432
    patient passed away | 432
    
    <|eot_id|>
    81 years old|0
    male|0
    admitted to internal medical department|0
    longstanding inguinoscrotal hernia|-8760
    upper abdominal pain|0
    auricular fibrillation|-8760
    chronic heart failure|-8760
    chronic renal dysfunction|-8760
    temperature 36.1°C|0
    abdominal distention|0
    epigastric tenderness|0
    bilateral giant inguinoscrotal hernia|0
    no tenderness|0
    no redness|0
    white blood cell count 4900/mm²|0
    C-reactive protein 1.2 mg/dl|0
    creatinin 1.71 mg/dl|0
    prothrombin time 18.7 s|0
    PT-INR 1.61|0
    computed tomography slightly dilated stomach|0
    computed tomography slightly dilated jejunum|0
    bilateral inguinoscrotal hernia containing small bowel|0
    bilateral inguinoscrotal hernia containing cecum|0
    bilateral inguinoscrotal hernia containing ascending colon|0
    bilateral inguinoscrotal hernia containing sigmoid colon|0
    no remarkable occlusion point|0
    acute entire abdominal pain|48
    blood pressure decreased to eighties|48
    CT scan free air right inguinal hernia sac|48
    much ascites|48
    diagnosis acute generalized peritonitis|48
    diagnosis small bowel perforation in inguinal hernia sac|48
    emergency operation performed|48
    mid-lower median abdominal incision|48
    transverse incision right inguinal area|48
    dirty ascites inguinal sac|48
    cecum perforation|48
    terminal ileum necrotic 100 cm behind Bauhin’s valve|48
    lateral extension internal hernia ring|48
    mobilization pancreas head|48
    mobilization duodenum|48
    mobilization right side of colon for right hemicolectomy|48
    substantial amount of bile|48
    rupture inferior duodenum angle|48
    right hemicolectomy|48
    side-to-side anastomosis duodenum and jejunum|48
    primary closure peritoneum hernia gate|48
    transferred to intensive care unit|48
    septic shock|432
    leakage duodenum–jejunum anastomosis|432
    use several antibiotic agents|432
    use vasopressure agent|432
    continuous hemodiafiltration|432
    patient passed away|432

