35 years old | 0
female | 0
gravida 2 | 0
para 2 | 0
gestational diabetes | 0
admitted to the hospital | 0
excruciating headache | -1
tonic-clonic convulsions | -1
low Glasgow Coma Scores | 0
intubation | 0
CT scan | 0
left frontal hematoma | 0
mild edema | 0
mass effect | 0
midline shift | 0
bleeding | 0
left lateral ventricle | 0
third ventricle | 0
fourth ventricle | 0
left subdural hematoma | 0
basal cisterns | 0
CT angiography | 0
frontal lobe bleeding | 0
carotid bifurcation aneurysm | 0
subarachnoidal bleeding | 0
intraventricular bleeding | 0
hydrocephalus | 0
coiling of the aneurysm | 0
mechanical ventilation | 0
sedated | 0
midposition pupils | 0
sluggish reaction to light | 0
dilatation of the left pupil | 24
sluggish reaction to light | 24
heart rate dropped | 24
hypotension | 24
norepinephrine | 24
crystalloid | 24
colloid therapy | 24
subarachnoidal rebleeding | 48
spastic reaction | 48
ischemia | 48
mesotemporal herniation | 48
third ventricle | 48
aqueduct level | 48
thrombosis | 72
left internal cerebral artery | 72
MCA | 72
partial mechanical thrombectomy | 72
fixed and dilated pupils | 96
decompressive craniotomy | 96
external ventricular drains | 96
ICP monitor | 96
elevated ICP | 120
medical management | 120
muscle relaxants | 120
mannitol | 120
hypertonic saline | 120
thiopental coma | 120
GCS | 216
no gag reflexes | 216
no cough reflexes | 216
apnea test | 216
EEG | 216
ventilatory support | 216
nutritional support | 216
vasoactive drugs | 216
normothermia | 216
hypotension | 216
hypertension | 216
antihypertensives | 216
DDAVP | 216
water flushes | 216
diabetes insipidus | 216
hypernatremia | 216
sepsis | 216
pneumonia | 216
urinary tract infection | 216
line infection | 216
antibiotics | 216
meningitis | 216
meropenem | 216
vancomycin | 216
panhypopituitarism | 216
thyroid hormone replacement | 216
steroids | 216
hypothermia | 216
passive rewarming | 216
blankets | 216
tracheostomy | 432
NG tube | 216
cesarean section | 2640
intrauterine growth retardation | 0
biometry | 0
estimated fetal weight | 0
oligohydramnios | 0
fetal anomalies | 0
ultrasounds | 216
heart rate monitoring | 216
amniocentesis | 216
betamethasone therapy | 216
fetal lung maturity | 216
fetal respiratory distress syndrome | 216
preterm male | 2640
breech presentation | 2640
Apgar score | 2640
NICU | 2640
nasal CPAP | 2640
respiratory distress syndrome | 2640
death | 2640