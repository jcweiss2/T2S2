68 years old | 0
male | 0
admitted to Intensive Care Unit | 0
septic shock | 0
hospital acquired pneumonia | 0
multiple organ dysfunction syndrome | 0
kidney function deteriorated | 0
eGFR 9.8 ml/min/1.73 m2 | 0
blood ureum 221 mg/dl | 0
blood creatinine 5.6 mg/dl | 0
regular hemodialysis | 0
tracheostomy tube placement | -24
prolonged endotracheal tube ventilation | -48
massive bleeding around the tube stoma | -24
arterial bleeding | -24
oxygen saturation 62% | -24
disseminated intravascular coagulation (DIC) | -24
elevated d-dimer | -24
thrombocytopenia | -24
prolonged prothrombin time | -24
flexible bronchoscopy examination | -12
blood clots at larynx and proximal trachea | -12
biopsy forceps extraction | -12
cryoextraction | -6
removal of blood clot | -6
bleeding after removal of blood clot | -6
argon plasma coagulation (APC) | -6
ventilator setting of fraction inspired oxygen (FiO2) 40% | -6
multiple APC | -6
bleeding controlled | -6
oxygen saturation 98% | 0
reevaluation bronchoscopy | 48
no new blood clots | 48
discharged | 1440
regular control at outpatient clinic | 1440