62 years old | 0
    male | 0
    referred to the hospital | 0
    dyspnea | 0
    intermittent chest pain | 0
    end-stage renal disease | -1464
    peritoneal dialysis | -1464
    type 2 diabetes mellitus | -1464
    aortic stenosis | -1464
    transcatheter aortic valve implantation | -1464
    diagnosed with COVID-19 | 0
    anemia | 0
    progressive hypoxia | 0
    intubated | 0
    transferred to tertiary care facility | 0
    treated for cytokine storm | 0
    hypotension | 0
    evaluation of aortic valve prosthesis | 0
    deteriorated rapidly | 0
    hypotensive without palpable pulse | 0
    advanced cardiac life support initiated | 0
    POCUS performed | 0
    large pericardial effusion | 0
    cardiac tamponade | 0
    emergent pericardiocentesis | 0
    serous fluid aspirated | 0
    spontaneous circulation returned | 0
    hemodynamic improvement | 0
    repeat echo performed | 0
    effusion size decreased | 0
    heart expansion | 0
    guide wire advanced | 0
    pigtail placed | 0
    650 mL fluid drained | 0
    resolution of pericardial effusion | 0
    normal LV function | 0
    <|eot_id|>