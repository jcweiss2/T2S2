34 years old | 0
male | 0
primary refractory acute myeloblastic leukemia | -8760
allogeneic bone marrow transplant | -648
delayed engraftment | -648
prolonged severe neutropenia | -648
vancomycin-resistant Enterococcus | -648
Streptococcus viridans | -648
Streptococcus mitis | -648
bacteremia | -648
tedizolid | -648
cefepime | -648
Flagyl | -648
daptomycin | -648
filgrastim | 0
acyclovir | 0
Bactrim | 0
caspofungin | 0
acute abdominal pain | 0
fever | 0
tachycardia | 0
hypotension | 0
tachypnea | 0
distended abdomen | 0
localized peritonitis | 0
white cell count 0.2 x 10^9 /L | 0
absolute neutrophil count (ANC) of zero | 0
anemic | 0
hemoglobin of 7 g/L | 0
thrombocytopenic | 0
platelet count of 10 x 10^9 /L | 0
lactic acid of 3.1 mmol/L | 0
segmental ischemia of the small bowel | 0
exploratory laparotomy | 0
ischemic bowel segment | 0
small bowel resection | 0
primary anastomosis | 0
norepinephrine | 0
vasopressin | 0
transesophageal echo | 0
intensive care unit | 0
pressors weaned | 24
extubated | 24
transferred to the floor | 72
diet advanced | 72
passed flatus | 72
new fevers | 96
increased abdominal pain | 96
lactic acidosis | 96
respiratory decompensation | 96
amphotericin B (AmBisome) | 96
necrotic small bowel | 96
invasive fungal forms | 96
mucormycosis | 96
comfort measures | 120
died | 120