25 years old | 0
G5 now P5 | 0
chronic hypertension | -288
premature prolonged rupture of membranes | -288
latency antibiotics | -288
intravenous ampicillin | -288
oral amoxicillin | -288
single dose azithromycin | -288
completed latency antibiotics | -288
chorioamnionitis | -12
ampicillin for chorioamnionitis | -12
trichomonas infection | -288
negative GBS culture | -288
male infant | 0
preterm | 0
ELBW | 0
26 weeks gestation | 0
birth weight 950 g | 0
spontaneous vaginal delivery | 0
required positive pressure ventilation | 0
required intubation | 0
APGAR scores 6, 3, 4 | 0
admitted to NICU | 0
arterial cord blood pH 6.96 | 0
pCO2 76 mm Hg | 0
base excess -15.9 mmol/L | 0
venous cord blood pH 7.17 | 0
pCO2 42 mm Hg | 0
base excess -12.7 mmol/L | 0
mixed metabolic and respiratory acidosis | 0
required high ventilator support | 0
respiratory acidosis improved | 0
surfactant administration | 0
persistent metabolic acidosis | 0
leukopenia | 0
WBC count 1.5x10^3/mm³ | 0
thrombocytopenia | 0
platelet count 89x10^3/mm³ | 0
CRP 21.1 mg/L | 0
blood culture sent | 0
prescribed ampicillin | 0
prescribed gentamicin | 0
hypotension at 4.5 hours | 4.5
rapid deterioration | 4.5
fluid resuscitation | 4.5
pressors (dopamine, dobutamine) | 4.5
repeat blood culture | 4.5
tracheal aspirate | 4.5
died at 5.5 hours | 5.5
parents declined autopsy | 5.5
blood cultures positive for gram-positive cocci | 12
identified as S. gallolyticus | 12
tracheal aspirate culture negative | 12
placental pathology confirmed chorioamnionitis | 12
fulminant sepsis due to S. gallolyticus | 0
respiratory distress | 0
sepsis | 0
elevated CRP | 0
hypotension | 4.5
death | 5.5
