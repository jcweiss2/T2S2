61 years old | 0
male | 0
admitted to the hospital | 0
left foot and ankle swelling | 0
generalized body aches | 0
intermittent chills | 0
no shortness of breath | 0
no chest pain | 0
no abdominal pain | 0
no urinary symptoms | 0
no diarrhea | 0
no headaches | 0
no runny nose | 0
no sore throat | 0
no tick bites | 0
no skin rashes | 0
cat licks him | -672
healthy cat | -672
cat's immunization status up-to-date | -672
no significant past medical history | 0
outpatient primary care clinic visits up-to-date | 0
not taking any medications at home | 0
tachycardiac | 0
heart rate 128 beats/minute | 0
blood pressure 86/53 mm Hg | 0
saturation 95% on room air | 0
afebrile | 0
alert and oriented to time, place, and person | 0
cardio-pulmonary and gastrointestinal examination unremarkable | 0
left ankle tender | 0
left ankle not erythematous or warm | 0
left foot swollen | 0
good and equal bilateral pulses | 0
white cell count (WBC) 7.5 K/uL | 0
10% bandemia | 0
hemoglobin 13.5 gm/dL | 0
platelets 72 K/mcL | 0
acute kidney injury | 0
creatinine 1.41 mg/dL | 0
glomerular filtration rate 51 mL/min/1.73 m2 | 0
low potassium 3.4 | 0
lactic acidosis 4.1 mmol/L | 0
Red blood cell morphology did not show any schistocytes | 0
urinalysis negative for any infections | 0
high specific gravity of 1.031 | 0
liver function test positive for mildly deranged AST/ALT | 0
AST/ALT 74/72 U/L | 0
total bilirubin 1.4 mg/dL | 0
procalcitonin 29.83 ng/mL | 0
WBC continued to worsen | 24
WBC peaked to 20 K/µL | 144
WBC trended down | 144
hemoglobin remained stable | 24
sepsis-induced thrombocytopenia improved | 192
mild acute kidney injury resolved | 192
liver function tests initially worsened | 24
liver function tests resolved | 192
lactic acidosis resolved | 192
CT chest-abdomen-pelvis did not show any pulmonary consolidations | 24
multiple prominent mesenteric lymph nodes | 24
sizes of lymph nodes improved upon follow-up repeat CT scan | 192
ultrasound of the left lower extremity ruled out deep venous thrombosis | 0
blood cultures drawn | 0
started on broad spectrum intravenous antibiotics | 0
meropenem 500 mg three times a day | 0
vancomycin 1 gm two times a day | 0
admitted to the intensive care unit | 0
MRI of his left ankle-foot showed diffuse soft tissue edema | 48
reticulation around the ankle | 48
trans-thoracic echocardiogram ruled out endocarditis | 48
sent for arthrocentesis | 48
lack of fluid in the ankle joint | 48
blood cultures came back positive for Pasteurella multocida | 48
intravenous antibiotic meropenem continued | 48
ciprofloxacin added | 48
Pasteurella multocida cultures showed good sensitivity to ciprofloxacin | 48
meropenem and piperacillin-tazobactam | 48
worsening left lower extremity edema | 144
ultrasound of the left lower extremity repeated | 144
new partially occlusive deep venous thrombus | 144
left popliteal vein | 144
left posterior tibial vein | 144
started on enoxaparin treatment | 192
sepsis-induced thrombocytopenia resolved | 192
mental status remained stable | 192
purplish discoloration of all finger and toe tips | 192
extensive workup for disseminated intravascular coagulation | 192
vasculitis | 192
hypercoagulable syndrome | 192
autoimmunity | 192
moderately positive lupus anticoagulant antibodies | 192
decreased protein-C activity | 192
positive anti-cardiolipin IgM antibodies | 192
diagnosed with thrombophilia | 192
left lower extremity DVT | 192
secondary to positive anticardiolipin antibodies | 192
low protein-C activity | 192
low-normal complements level | 192
ANA and DsDNA | 192
lupus | 192
vasculitis | 192
connective tissue disease | 192
rheumatoid arthritis | 192
multiple blood cultures negative | 192
discharged to a rehabilitation center | 480
continued to have digital ulcerations | 720
right forefoot turned into wet gangrene | 720
readmitted for right fore-foot amputation | 720
blood cultures sent again | 720
underwent right fore-foot amputation | 720
blood cultures came back positive again for Pasteurella multocida | 720
started on intravenous antibiotic piperacillin-tazobactam | 720
deep tissue cultures and bone biopsy from the gangrenous, infected toes | 720
enterococcus group-D | 720
staphylococcus coagulase negative | 720
started on daptomycin intravenously | 720
left ankle-knee osteomyelitis | 720
underwent below knee amputation | 720
discharged again to a rehabilitation center | 720