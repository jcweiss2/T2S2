history of autoimmune hepatitis | -168
unprotected sexual intercourse | -336
influenza vaccination | -720
COVID-19 vaccination | -720
no recent travel history | 0
admission | 0
bilateral lower extremity pain | 0
edema | 0
ascites | 0
fever | 0
chills | 0
nausea | 0
dizziness | 0
heavy menorrhagia | 0
hemodynamically unstable | 0
blood pressure 67/39 mmHg | 0
heart rate 129 beats per minute | 0
respirations 33 per minute | 0
temperature 35.1 degrees Celsius | 0
jaundice | 0
scleral icterus | 0
abdominal ascites with fluid wave | 0
anasarca | 0
erythematous vaginal vault with minimal discharge | 0
no vesicles, lesions, or retained foreign objects | 0
fine reticular violaceous patches on the right proximal thigh | 0
lactic acidosis | 0
elevated creatinine | 0
elevated aspartate transaminase | 0
elevated alanine transaminase | 0
elevated total bilirubin | 0
elevated direct bilirubin | 0
elevated alkaline phosphatase | 0
low total protein | 0
low albumin | 0
low hemoglobin | 0
low leukocytes | 0
low platelets | 0
elevated prothrombin time | 0
elevated international normalized ratio | 0
negative beta-human chorionic gonadotropin test | 0
occasional schistocytes on peripheral smear | 0
peritoneal fluid analysis with leukocyte count 9821 | 0
CT angiography showing cirrhosis with portal hypertension | 0
large volume abdominal ascites | 0
splenomegaly | 0
generalized edematous wall thickening of the colon and rectum | 0
intubation | 0
intravenous fluids | 0
blood products | 0
vasopressors | 0
broad-spectrum antibiotic therapy | 0
vancomycin | 0
piperacillin-tazobactam | 0
doxycycline | 0
clindamycin | 0
intravenous immunoglobulin | 0
large violaceous non-blanching ecchymoses | 16
flaccid bullae | 16
skin over the entire right leg, as well as the left proximal thigh to mid-shin, was dusky and violaceous | 36
various-sized bullae up to greater than 10 cm filled with red to black-colored fluid | 36
elevated lactate dehydrogenase | 36
low fibrinogen | 36
elevated D-dimer | 36
negative urinalysis | 36
negative salicylate level | 36
negative acetaminophen level | 36
negative Chlamydia trachomatis and Neisseria gonorrhea nucleic acid amplification tests | 36
negative urine toxicology screen | 36
negative peritoneal fluid culture | 36
blood culture grew pan-susceptible Streptococcus pneumoniae | 36
progressive hypoxia | 48
shock | 48
death | 48
autopsy showing cirrhotic liver | 48
diffuse alveolar damage | 48
over five liters of serous fluid in the abdominal compartment | 48