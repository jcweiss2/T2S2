74 years old | 0
white | 0
female | 0
admitted to the hospital | 0
low-grade fever | -48
dry cough | -48
shortness of breath | -48
elective right total knee replacement | -168
post-operative course | -168
pain | -168
redness | -168
swelling | -168
essential hypertension | 0
obesity | 0
myasthenia gravis | 0
osteoarthritis | 0
body temperature 37.3°C | 0
blood pressure 121/82 | 0
pulse 87 beats per minute | 0
respiratory rate 16 breaths per minute | 0
oxygen saturation 87% | 0
bilateral rhonchi | 0
rales | 0
patchy air space opacity | 0
pneumonia | 0
rapid nucleic acid amplification test | 0
nasopharyngeal swab | 0
broad-spectrum antibiotics | 0
cefepime | 0
levofloxacin | 0
supportive care | 0
2 L supplemental oxygen | 0
mild diarrhea | 72
generalized weakness | 72
fatigue | 72
intravenous immunoglobulin | 72
mild MG exacerbation | 72
MG crises | 72
arterial blood gases | 0
complete blood count | 0
basic metabolic profile | 0
mild absolute lymphopenia | 0
anemia | 0
pH 7.46 | 0
pCO2 44.6 mmHg | 0
pO2 94.7 mmHg | 0
bicarbonate 31.4 mmol/L | 0
increasing shortness of breath | 24
oxygen requirements increased | 24
nasopharyngeal swab results | 96
SARS-CoV-2 positive | 96
hydroxychloroquine | 96
azithromycin | 96
zinc sulfate | 96
oral vitamin C | 96
blood and sputum cultures | 96
broad-spectrum antibiotics discontinued | 96
shortness of breath worsened | 144
oxygen requirements increased | 144
drowsy | 144
moderate distress | 144
unable to protect airways | 144
blood pressure 78/56 mmHg | 144
heart rate 112 beats per minute | 144
temperature 38°C | 144
respiratory rate 28 breaths per minute | 144
bilateral alveolar infiltrates | 144
interstitial edema | 144
ARDS | 144
intubated | 144
mechanical ventilation | 144
norepinephrine | 144
septic shock | 144
colchicine | 144
cytokine storm | 144
elevated interleukin-6 | 144
high-dose vitamin C | 168
clinical condition improved | 192
norepinephrine stopped | 192
CXR improved | 240
spontaneous breathing trial | 240
CPAP/PS | 240
ABGs | 240
pH 7.49 mmHg | 240
pCO2 40.2 mmHg | 240
pO2 77.1 mmHg | 240
bicarbonate 30.2 mmol/L | 240
extubated | 240
4 L oxygen | 240
oxygen saturation 92% | 384
CXR nearly complete resolution | 384
discharged | 384
quarantine | 384