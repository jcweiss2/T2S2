73 years old | 0
male | 0
admitted for endoscopic dilatation for achalasia | 0
diabetes mellitus | -8760
Parkinsonism | -8760
trans-urethral resection of the prostate (TURP) | -8760
laparoscopic cholecystectomy | -105120
presented to gastroenterology clinic for dysphagia for solid food | -17520
type II achalasia diagnosis | -17520
manometry confirmed | -17520
water-soluble studies confirmed | -17520
endoscopic pneumatic dilatation | -4320
symptoms free | -4320
symptoms progressively worsened | -4320
scheduled for endoscopic pneumatic dilatation | 0
general anesthesia | 0
endotracheal intubation | 0
placed in left lateral position | 0
Rigiflex dilator introduced | 0
gastroesophageal junction (GEJ) dilated to 35 mm for 60 seconds | 0
GEJ dilated again for 90 seconds | 0
desaturation manifestation | 0
multiple esophageal perforations confirmed | 0
plain chest radiography showed left-sided pneumothorax | 0
minimal pneumomediastinum | 0
chest tube inserted | 0
oxygen saturation improved | 0
thoracic surgical team involved | 0
upper gastrointestinal (GI) surgical team involved | 0
decision for diagnostic laparoscopy | 0
trial of primary esophageal repair | 0
placed in supine position with abducted legs | 0
pneumatic compression devices used | 0
preoperative broad-spectrum antibiotics | 0
pneumoperitoneum created | 0
laparoscope introduced | 0
diagnostic laparoscopy showed no free fluid | 0
left lobe of liver retracted | 0
pars condensa dissected | 0
pars flaccida dissected | 0
hepatic branch of vagus nerve sacrificed | 0
esophago-phrenic ligament dissected | 0
lower esophagus mobilized | 0
umbilical tape applied around GEJ | 0
multiple perforations found in lower esophagus | 0
trial of primary esophageal repair attempted | 0
esophageal mucosa dissected | 0
unhealthy mucosal edges | 0
decision for double-tract reconstruction | 0
distal esophagus transected | 0
anvil introduced through oral cavity | 0
esophagostomy created | 0
proximal gastrectomy | 0
jejunal loop measured 60 cm | 0
camera port extended | 0
Alexis port inserted | 0
jejunal loop delivered | 0
jejuno-jejunostomy created | 0
mesenteric defect closed | 0
circular stapler introduced | 0
esophago-jejunostomy | 0
gastrostomy created | 0
jejunostomy created | 0
gastro-jejunostomy | 0
Blake drain inserted | 0
transferred to ICU | 0
extubated | 24
shifted to regular ward | 24
intravenous fluids | 24
nil per os | 24
empirical antibiotics | 24
antifungal drugs | 24
clear liquid diet | 120
water-soluble study confirmed GI continuity | 120
discharged | 192
followed up | 192
