12 years old | 0
female | 0
admitted to the hospital | 0
fever | 0
shortness of breath | 0
cough | 0
tachycardic | 0
tachypneic | 0
requiring 3 L of supplemental oxygen | 0
given 1 L of normal saline bolus intravenously | 0
bilateral pulmonary edema | 0
sepsis | 0
started on vancomycin | 0
started on cefotaxime | 0
nephrotic syndrome | -2520
renal biopsy | -2160
minimal change disease | -2160
genetic testing | -2160
heterozygous, non-coding mutation in the TRPC6 gene | -2160
cyclophosphamide | -1800
relapse | -1440
tacrolimus | -1080
partial clinical response | -720
repeat biopsy | -240
interstitial nephritis | -240
Acthar | -120
S. pneumoniae | 8
nasopharyngeal swab PCR positive for parainfluenza type 2 | 8
oliguria | 24
creatinine increased | 24
hemoglobin decreased | 24
discontinued Acthar | 24
discontinued tacrolimus | 24
transfused one unit of unwashed packed red blood cells | 24
started on continuous veno-venous hemodiafiltration | 24
respiratory failure | 96
intubation | 96
bilateral patchy consolidation | 96
bilateral pleural effusions | 96
high-dose hydrocortisone | 96
platelet count decreased | 96
intravenous vasoactive support | 96
started plasma exchange | 120
FFP used as replacement fluid | 120
direct Coombs test negative | 120
follow-up direct Coombs test positive | 192
platelet count reached a nadir | 312
slowly improved | 312
discharged home | 936
creatinine returned to baseline level | 936
angiotensin-converting enzyme inhibitor therapy | 936
persistent nephrotic syndrome | 936
PCV7 vaccination | -4320