29 years old | 0
Caucasian | 0
female | 0
diamniotic dichorionic twin pregnancy | 0
admitted to the obstetric unit | 0
preterm premature rupture of membranes | 0
fertilized in-vitro embryo transfer | -280
spontaneous abortion | -728
hyperemesis gravidarum | -196
treated with chlorpromazine | -196
amniocentesis | -168
CGH array | -168
discordant growth between the twins | -112
first fetus small for gestational age | -112
aberrant right subclavian artery | -112
right ventriculum hypertrophy | -112
double left renal artery | -112
corticosteroids | 0
betamethasone | 0
atosiban | 0
prevent very early delivery | 0
magnesium sulfate infusion | 0
twin neuroprotection | 0
cefazoline | 0
bemiparine | 0
prevent thrombosis | 0
inflammatory marker values increased | 96
WBC increased | 96
CPR increased | 96
PCT negative | 96
cefazoline continued | 96
WBC decreased | 264
CPR negative | 264
PCT negative | 264
uterine contractions | 288
substantial discharge of amniotic fluid | 288
counseling on imminent delivery | 288
magnesium sulfate restarted | 288
neuroprotection | 288
biochemical exams | 288
WBC increased | 288
CPR negative | 288
PCT negative | 288
antibiotic therapy continued | 288
first fetus delivered | 336
umbilical cord clamped | 336
kept in uterus | 336
newborn transferred to NICU | 336
newborn died | 432
mother intensively monitored | 336
daily blood exams | 336
ultrasound checks of the second fetus | 336
WBC decreased | 552
tocolysis restarted | 552
atosiban | 552
bemiparine continued | 552
cefazoline continued | 552
ultrasound monitoring | 552
fetus's growth rate slowed | 552
Doppler scans of the umbilical artery | 552
no anomalies | 552
pathological pattern of cardiotocography | 696
low variability | 696
late decelerations | 696
cesarian section | 696
second baby delivered | 696
Apgar score | 696
intubated | 696
admitted to NICU | 696
intubation changed to external pulmonary support | 696
surfactant | 696
blood units | 696
erythropoietin | 696
anemia | 696
clinical condition improved | 696
cardiac ultrasound scans | 696
cerebral ultrasound scans | 696
electroencephalograms | 696
neurophysiological development | 696
urinary functions normal | 696
gastroenterological functions normal | 696
started to eat | 744
parenteral feeding stopped | 744
discharged from hospital | 888
follow-up | 1296
no neurological defects | 1296
no cardiac defects | 1296
no other defects | 1296
antibiotic therapy | 696
ceftriaxone | 696
anti-thrombotic therapy | 696
bemiparine | 696
uterotonic therapy | 696
oxytocine | 696
blood exams returned to normal | 720
discharged | 720
bemiparine prescribed | 720
cefuroxime prescribed | 720