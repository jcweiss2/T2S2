71 years old | 0
female | 0
arthritis | 0
central serous retinopathy | 0
remote deep vein thrombosis | 0
not on anticoagulation | 0
hyperlipidemia | 0
osteoporosis | 0
fatigue | -2160
abdominal pain | -2160
loss of appetite | -2160
referred to emergency room | 0
anemia | 0
hemoglobin 10.7 g/dL | 0
mild thrombocytopenia | 0
abnormal liver function tests | 0
afebrile | 0
pulse 110 beats/minute | 0
blood pressure 115/80 mmHg | 0
O2 saturation 95% | 0
Na+ 128 mmol/L | 0
AST 110 U/L | 0
ALT 73 U/L | 0
GGTP 94 U/L | 0
albumin 2.6 gm/dL | 0
hepatic thrombosis | 0
portal vein thrombosis | 0
hepatitis suspicion | 0
pancreatitis suspicion | 0
colitis suspicion | 0
right hepatic vein thrombosis | 0
pancreatic tail lesion 1.9 × 1.8 cm | 0
pancreatic carcinoma suspicion | 0
pancreatic neuro-endocrine tumor suspicion | 0
multiple foci of large frankly neoplastic cells | 0
infiltrating pancreatic lobules | 0
scant cytoplasm | 0
nuclei with regular contour | 0
prominent nucleoli | 0
mitotic figures | 0
numerous apoptotic bodies | 0
immunohistochemical work-up unrevealing | 0
Ki-67 proliferation index >95% | 0
DLBCL diagnosis | 0
cell block with large atypical cells | 0
CD20 positive | 0
CD79a positive | 0
CD45 positive | 0
PAX-5 focally positive | 0
MUM-1 non-contributory | 0
bone marrow aspirate no involvement | 0
bone marrow biopsy no involvement | 0
Weisella confusa bacteremia | 0
Enterococcus faecalis bacteremia | 0
treated with piperacillin-tazobactam | 0
creatinine up-trending | 0
elevated lactate dehydrogenase | 0
diastolic blood pressure fluctuating | 0
up-trending liver function tests | 0
refractory to intravenous fluid | 0
antibiotic regimen broadened to vancomycin | 0
meropenem | 0
transferred to ICU | 0
septic shock | 0
started on metronidazole | 0
oral vancomycin | 0
fluids and norepinephrine drip | 0
lactic acidosis | 0
intubated | 0
antibiotics broadened to vancomycin | 0
amikacin | 0
micafungin | 0
metronidazole | 0
stress dose steroids | 0
disseminated intravascular coagulopathy | 0
pulmonary emboli | 0
irreversible multi-organ failure | 0
demise | 312
autopsy consent | 312
pancreatic mass 1.9 × 1.8 cm | 312
lymphoma cells in vessels | 312
organizing occlusive thromboemboli in left pulmonary artery | 312
right atrial thrombus | 312
intrahepatic right portal vein thrombus | 312
pancreas mass 2 cm | 312
paraesophageal lymph nodes | 312
perihepatic lymph nodes | 312
hemorrhagic lymph nodes | 312
spleen 350 gm | 312
liver 1520 gm | 312
portal vein thrombosis related to neoplastic involvement | 312
CD5 positive | 312
CD10 negative | 312
MUM1 positive | 312
CD3 negative | 312
Ki-67 >90% | 312
Epstein-Barr encoding region negative | 312
