61 years old | 0
male | 0
admitted to the hospital | 0
T-cell lymphoma | -2160
chemotherapy | -2160
deep venous thrombosis | -672
pulmonary embolism | -672
therapeutic anticoagulation | -672
obtundation | 0
fever | 0
chills | 0
diarrhea | 0
typhlitis of the terminal ileum | -2160
typhlitis of the cecum | -2160
pulmonary involvement | -2160
bilateral pleural effusions | -2160
ground-glass opacification | -2160
alveolar opacities | -2160
respiratory failure | -168
sepsis | -168
acute tubular necrosis | -168
vasogenic edema | -24
agonal breathing | 0
unequal pupils | 0
noncontrast computed tomography | 0
intra-axial lesions | 0
extensive surrounding vasogenic edema | 0
cerebral toxoplasmosis | 0
neurocysticercosis | 0
multiple abscesses | 0
contrast-enhanced MRI | 24
lesions throughout the brain | 24
cervical spine | 24
thoracic spine | 24
lumbar spine | 24
leptomeninges enhancement | 24
osseous hyperdensities | 24
metastases | 24
intradural extramedullary lesion | 24
stereotactic navigation | 48
biopsy | 48
ALK-positive anaplastic large T-cell lymphoma | 48
CD4 | 48
CD45 | 48
CD30 | 48
reactive astrocytosis | 48
cavitation | 48
rarefaction of brain parenchyma | 48
positive IgG antibody against toxoplasmosis | 72
sulfadiazine | 72
pyrimethamine | 72
empiric toxoplasmosis treatment | 72
communicating hydrocephalus | 96
external ventricular catheter | 96
ICP monitoring | 96
therapeutic ventricular drainage | 96
elevated ICP | 120
severe thrombocytopenia | 120
platelet transfusions | 120
hemodynamic instability | 120
norepinephrine | 120
phenylephrine | 120
epinephrine | 120
vasopressin | 120
withdrawal of care | 168
expiration | 168