70 years old | 0
female | 0
Streptococcus pneumoniae aortic valve endocarditis | -120
bioprosthetic porcine aortic valve replacement | -120
recurrent S. pneumoniae endocarditis | -120
aortic root replacement with a homograft | -120
rivaroxaban for atrial fibrillation | -744
pseudomonal bacteremia | -744
cefepime | -744
levofloxacin | -744
admitted with pseudomonal bacteremia | -744
right-sided chest pain | -336
growing pulsatile mass on the right sternal border | -336
computed tomography angiogram (CTA) | 0
2.5 × 2.0-cm proximal thoracic aortic pseudoaneurysm | 0
anterior mediastinal hematoma | 0
labetalol | 0
esmolol | 0
prothrombin complex concentrate | 0
vancomycin | 0
levofloxacin | 0
CTA demonstrated growth of the pseudoaneurysm | 7
3.4 × 2.1-cm pseudoaneurysm | 7
neck 0.6 cm wide | 7
location 1.4 cm superior to the right coronary artery ostium | 7
distance from the right coronary ostium to the innominate artery | 7
60.5 mm | 7
infectious pseudoaneurysm | 0
endovascular stent graft placement | 0
transvenous pacer | 0
right ventricle | 0
right femoral access | 0
left axillary artery | 0
infraclavicular incision | 0
axillary artery punctured | 0
0.035 Glidewire | 0
Terumo Medical | 0
8F sheath | 0
GLIDECATH | 0
left ventricle | 0
double-curved Lunderquist wire | 0
Cook Medical Inc | 0
pigtail catheter | 0
left femoral 5F sheath | 0
36 × 50-mm Zenith abdominal extension stent graft | 0
rapid pacing | 0
device deployed | 0
angiography | 0
continued pseudoaneurysm filling | 0
36 × 50-mm Zenith stent | 0
completion angiography | 0
patency of both coronary arteries | 0
exclusion of the pseudoaneurysm | 0
transferred to the critical care unit | 0
antibiotic therapy changed | 0
tobramycin | 0
meropenem | 0
Pseudomonas aeruginosa | 0
aspirin | 0
prophylactic subcutaneous heparin | 0
rivaroxaban discontinued | 0
heart rate controlled with metoprolol | 0
predischarge computed tomography scan | 240
exclusion of the pseudoaneurysm | 240
discharged to home | 240
postoperative day 10 | 240
home infusions | 240
tobramycin | 240
meropenem | 240
peripherally inserted central catheter | 240
lifelong suppressive therapy with oral levofloxacin | 240
follow-up CTAs | 960
exclusion of the pseudoaneurysm | 960
decreased size of the mediastinal hematoma | 960
stable positioning of the stent grafts | 960
resolution of all symptoms | 960
follow-up CTAs | 1440
exclusion of the pseudoaneurysm | 1440
decreased mediastinal hematoma | 1440
stable stent graft positioning | 1440
no evidence of endoleak | 1440