54 years old|0
    male|0
    admitted to the hospital|0
    malaise|-168
    rigors|-168
    right upper quadrant pain|-168
    flank pain|-168
    septic shock|0
    transferred to tertiary hospital|0
    multi-organ failure|0
    oxygen saturation of 80% on 6L oxygen via Hudson Mask|0
    hemodynamic compromise|0
    systolic blood pressure of 80|0
    sinus tachycardia up to 120 beats per minute|0
    bilateral renal angle tenderness|0
    intubated|0
    transferred to intensive care unit|0
    severe metabolic acidosis|24
    anuric renal failure|24
    thrombocytopenia|24
    dialysis|24
    antibiotics broadened to meropenem|24
    antibiotics broadened to metronidazole|24
    antibiotics broadened to fluconazole|24
    stabilized|24
    CT scan showing bilateral emphysematous pyelonephritis|24
    type 2 diabetes|0
    referral to urology service|24
    discussion with next of kin|24
    decision not to perform bilateral nephrectomies|24
    clinical deterioration|48
    extreme coagulopathy with INR of 16|48
    progressing metabolic acidosis|48
    liver failure|48
    worsening synthetic failure|48
    maximal inotropic support|48
    case conference between next of kin, ICU, and urology team|48
    decision to treat medically|48
    antibiotics rationalized to ceftriaxone|72
    CT scan on day 3 showing no drainable collections|72
    extubated on day 6|144
    ongoing dialysis for acute kidney injury|144
    IV ceftriaxone for 4 weeks|168
    transitioned to oral augmentin duo forte for further 8 weeks|168
    repeat CT after 4 weeks showing no significant change|672
    afebrile|672
    hemodynamically stable|672
    remained on intermittent hemodialysis|672
    creatinine remained 250|672
    required regular hemodialysis|672
    