53 years old | 0
African American | 0
female | 0
admitted to the hospital | 0
altered mental status | -72
feeling unwell | -72
dyspnea | -72
hypertension | -672
diabetes mellitus type 2 | -672
temperature of 36.6 °C | 0
heart rate of 112 beats per minute | 0
blood pressure of 140/72 mm Hg | 0
respiratory rate of 28 breaths per minute | 0
oxygen saturation of 96% on room air | 0
confused | 0
agitated | 0
tachypneic | 0
tachycardic | 0
leukocytosis | 0
white blood cell count of 19.9 × 10^9/L | 0
absolute neutrophils of 89.3% | 0
platelet count of 507 × 10^9/L | 0
sodium level of 131 mmol/L | 0
potassium of 6.2 mmol/L | 0
chloride of 104 mmol/L | 0
total CO2 of 6 | 0
glucose level >38.8 mmol/L | 0
BUN of 25 mmol/L | 0
creatinine of 362.5 µmol/L | 0
high anion gap of 28 | 0
acetone was large | 0
high anion gap metabolic acidosis | 0
compensatory respiratory alkalosis | 0
DKA | 0
acute kidney injury | 0
intravenous fluids | 0
insulin infusion | 0
transferred to the intensive care unit | 0
febrile | 72
Tmax of 39.1 °C | 72
tachycardic | 72
septic workup | 72
empiric broad-spectrum antibiotics | 72
antipyretics | 72
blood cultures grew K pneumoniae | 72
CT scan of the abdomen and pelvis | 96
hypoattenuating hepatic lesions | 96
heterogeneous splenic hyperattenuation | 96
splenic infarcts | 96
magnetic resonance imaging | 120
hepatic abscess | 120
splenic abscesses | 120
piperacillin/tazobactam | 120
ceftriaxone | 120
metronidazole | 120
percutaneous drainage of the left hepatic lobe abscess | 144
pus grew K pneumoniae | 144
repeat blood cultures were negative | 168
renal function stabilized | 168
dialysis was discontinued | 168
worsening of several ill-defined hypoattenuating splenic lesions | 192
percutaneous drainage of the splenic abscesses | 192
acute right femoral vein deep vein thrombosis | 216
popliteal vein deep vein thrombosis | 216
peroneal vein deep vein thrombosis | 216
high-range heparin infusion | 216
inferior vena cava filter | 216
colonoscopy | 240
15-mm polyp in the cecum | 240
nonbleeding hemorrhoids | 240
blood transfusions | 240
discharged | 432
peripherally inserted central catheter line | 432
6-week course of antibiotics | 432