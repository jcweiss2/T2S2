49 years old| 0
female| 0
admitted to the hospital| 0
nausea| -48
vomiting| -48
intermittent fever| -48
unexplained nausea| -72
unexplained vomiting| -72
fever with peak temperature of 38.4°C| -72
diarrhea with watery stools at least twice daily| -72
oliguria| -48
apathy| -48
blood culture| -48
other related tests| -48
transferred to our hospital for further treatment| -48
diagnosed with diarrhea| -48
admitted to the intensive care unit| -48
poor appetite| -48
poor sleep| -48
lost 5 kg of total body weight| -48
history of type 2 diabetes mellitus| -72
oral metformin| -72
unsatisfactory blood sugar control| -72
coma| 0
involuntary movements| 0
temperature: 37.8°C| 0
heart rate: 130 beats/min| 0
respiration: 28 breaths/min| 0
blood pressure: 70/50 mmHg| 0
bowel sounds: 6 beats/min| 0
urine output less than 0.5 mL/kg/min| 0
no swelling of either lower limb| 0
Babinski sign negative| 0
white blood cells (WBC) 9.4 × 109/L| 0
neutral granulocytes 94.5%| 0
platelet count 5.2 × 1010/L| 0
procalcitonin (PCT) 0.4 ng/mL| 0
T-cell subpopulation analysis significant reduction and exhaustion| 0
CD4+ T-cell count 4.4 × 1011/L| 0
CD4+ T-cells 13.89% expressing PD-1| 0
CD8+ T-cell count 1.18 × 1011/L| 0
CD8+ T-cells 26.65% expressing PD-1| 0
liver damage| 0
aspartate aminotransferase 923 U/L| 0
alanine aminotransferase 410 U/L| 0
total bilirubin 27.6 µmol/L| 0
serum creatinine (SCr) 380 µmol/L| 0
metabolic acidosis| 0
respiratory alkalosis| 0
blood gas pH 7.46| 0
partial pressure of carbon dioxide 25 mmHg| 0
bicarbonate level 17.8 mmol/L| 0
base excess -5.0 mmol/L| 0
lactate level 1.2 mmol/L| 0
liver ultrasound multiple mixed-density shadows| 0
NMLA| 0
sepsis| 0
septic encephalopathy| 0
septic shock| 0
SA-AKI| 0
secondary immune deficiency| 0
APACHE II score 18| 0
SOFA score 11| 0
empirical broad-spectrum antibiotic cefoperazone-sulbactam initiated within 1 h| 0
fluid resuscitation for sepsis performed within 3 h with 30 mL/kg crystalloid solution| 0
blood pressure increased to 80/55 mmHg| 0
noradrenaline administered to achieve mean arterial pressure 65 mmHg| 0
antibiotics upgraded to imipenem and linezolid| 0
urine output increased to 1.5–2.0 mL/kg/min| 0
glutathione injection administered| 0
ultrasound-guided puncture and drainage could not be performed| 0
computed tomography confirmed NMLA| 24
sepsis not adequately controlled| 24
lactate rose to 2.9 mmol/L| 24
WBC increased to 1.2 × 1010/L| 48
PCT increased to 200 ng/mL| 48
interleukin-6 (IL-6) 92.5 µmol/L| 48
kidney function deteriorated| 48
SCr increased to 403 µmol/L| 48
proposed performing CRRT combined with HP therapy| 48
family refused treatment due to economic considerations| 48
liver ultrasonography LA still not liquefied| 48
puncture drainage could not be performed| 48
WBC rose to 1.32 × 1010/L| 72
IL-6 increased to 525.2 µmol/L| 72
gram-negative bacterial infection high likelihood| 72
urine output maintained at 2 mL/kg/h| 72
SCr rose to 490 µmol/L| 72
developed septic shock| 72
senescence-associated acute SA-AKI| 72
combination of CRRT and HP performed| 72
PrismaFlex system used for CRRT| 72
M100 filter used for CRRT| 72
HA380 membrane filter used for HP once daily for 6 h| 72
continuous venovenous hemofiltration at 30 mL/kg/h| 72
blood flow rate of 120 mL/h| 72
no adverse effects observed| 72
continuous blood purification therapy terminated on the 7th day| 168
anti-infection and other treatments continued| 168
improvement observed during 5-day CRRT and HP treatment| 120
WBC decreased to 4.0 × 109/L| 168
PCT decreased to 8.43 ng/mL| 168
IL-6 decreased to 82.2| 168
tissue perfusion improved| 168
lactate decreased to 0.9 mmol/L| 168
renal function gradually improved| 168
SCr decreased to 129 µmol/L| 168
immune function improved| 168
CD8+ T-cells rose to 6.71 × 1011/L| 168
LA remained liquefied and could not be drained| 168
APACHE II lowered to 16| 168
SOFA score declined to 3| 168
treated in ICU for 10 days| 240
transferred to gastroenterology department| 240
discharged on the 21st day| 504
recovered after 28 days of follow-up| 672
