55 years old | 0
    male | 0
    simultaneous pancreas-kidney transplantation (SPKT) | 0
    end-stage renal disease due to type 1 diabetes mellitus | 0
    stroke | -14640
    coronary artery disease | -14640
    dialysis | -14640
    started dialysis at age 42 | -14640
    duration of dialysis 1.5 years | -14640
    pancreas and kidney transplantation in 2007 | -17520
    medical history of stroke and coronary artery disease | -17520
    arterial anastomosis of donor-iliac artery graft to recipient common iliac artery | -17520
    portal vein anastomosis to inferior vena cava | -17520
    enteric exocrine drainage via side-to-side duodeno-jejunostomy | -17520
    cold ischemia time pancreas 10 hours 28 minutes | -17520
    warm ischemia time pancreas 30 minutes | -17520
    cold ischemia time kidney 10 hours 28 minutes | -17520
    warm ischemia time kidney 50 minutes | -17520
    tacrolimus | -17520
    mycophenolate mofetil | -17520
    prednisolone | -17520
    anti-thymocyte globulin induction therapy | -17520
    no rejection episodes | -17520
    no infection episodes | -17520
    transferred to our institution in 2019 | -10512
    gastrointestinal bleeding of unknown origin | -10512
    weakness | -10512
    urinary tract infection with Pseudomonas aeruginosa | -10512
    tacrolimus | -10512
    prednisolone | -10512
    azathioprine | -10512
    actively bleeding ulcer at duodenojejunal anastomosis | -10512
    injection of Histoacryl failed | -10512
    recurring hemorrhages | 0
    pancreas graft function normal | 0
    euglycemia (C-peptide 7.9 ng/ml) | 0
    renal allograft function initially impaired (serum creatinine 2.1 mg/dl) | 0
    concomitant urinary tract infection | 0
    anti-infective therapy with imipenem | 0
    renal function normalized | 0
    gastrointestinal bleeding persisted | 0
    esophagogastroduodenoscopy (EGD) repeated | 0
    ulcer at jejuno-duodenal anastomosis | 0
    varicose vessels in the same area | 0
    CT angiography showed no signs of abdominal bleeding | 0
    pantoprazole therapy | 0
    recurring low hemoglobin values (hemoglobin 7.0 g/dl) | 0
    multiple transfusions of RBCs | 0
    double-balloon endoscopy | 0
    colonoscopy | 0
    capsule endoscopy | 0
    negative for acute bleeding focus | 0
    bone marrow biopsy performed for low peripheral leucocyte counts | 0
    no abnormalities in bone marrow biopsy | 0
    recurrent septic episodes | 0
    impairment of renal function | 0
    immunosuppressive medication reduced | 0
    transiently stopped during severe infections | 0
    CD4-positive T lymphocyte count 196/µl | 0
    low-dose hydrocortisone treatment | 0
    elevated liver enzymes (ALAT and ASAT) | 0
    abdominal ultrasound showed no cirrhosis | 0
    hepatitis E infection | 0
    high viral loads | 0
    ascites | 0
    CMV reactivation in blood | 0
    hemorrhagic shock | 1464
    EGD performed during hemorrhagic shock | 1464
    jejunal varices clipped | 1464
    adrenalin injection performed | 1464
    hemorrhage not stopped | 1464
    CT scan showed stenosis of porto-caval anastomosis | 1464
    venous angiography via right superior femoral vein | 1464
    stenosis dilated with balloon catheter | 1464
    partial improvement of stenosis proven by CT scan | 1464
    perfusion of abdominal organs unremarkable | 1464
    recurrent low hemoglobin levels | 1464
    no cardiovascular adverse events | 1464
    normal ejection fraction by echocardiography | 1464
    surgical intervention after 3 months | 2160
    end-to-side anastomosis of splenic vein to right iliac vein | 2160
    pancreas graft unremarkable macroscopically | 2160
    few adhesions | 2160
    tortuous collateral vessels present | 2160
    right internal iliac vein mobilized | 2160
    anastomosis performed with bovine patch | 2160
    color-coded duplex ultrasound verified retrograde perfusion | 2160
    decompression of venous outflow accomplished | 2160
    blood transfusions still needed | 2160
    graft pancreatectomy | 2640
    part of small intestine and donor pancreas resected | 2640
    chronic inflammation of resected tissues | 2640
    intestinal tortuous collateral vessels | 2640
    bleeding stopped | 2640
    over 70 units of RBCs transfused | 2640
    no more blood products needed after pancreatectomy | 2640
    hepatitis E infection no longer detected | 2640
    CMV reactivation treated with ganciclovir | 2640
    CD4 T cell count recovered | 2640
    tacrolimus and prednisolone restarted | 2640
    renal allograft function good (serum creatinine 1.2 mg/dl) | 2640
    no donor-specific HLA antibodies | 2640
    discharged after 180 days | 4320
    patient's health improved over 12 months | 4320