4 years old | 0
male | 0
Progressive symmetrical erythrokeratoderma (PSEK) | 0
Gottron syndrome | 0
hyperkeratotic plaques | 0
peripheral erythema | 0
extensor surfaces | 0
face involvement | 0
trunk involvement | 0
harlequin phenotype | 0
ABCA12 gene mutations | 0
harlequin ichthyosis (HI) | 0
generalized erythroderma | 0
small scales | 0
harlequin-like presentation | 0
amegakaryocytic thrombocytopenia | 0
homozygous variant in KDSR gene | 0
deceased sister | 0
consanguineous parents | 0
born by cesarean section | 0
thick, platelike hyperkeratotic scales | 0
marked ectropion | 0
eclabium | 0
harlequin ichthyosis (HI) diagnosis | 0
admitted to neonatal intensive care unit | 0
transport to tertiary center | 0
severe anemia | 0
thrombocytopenia | 0
multiple transfusions | 0
intravenous antibiotics | 0
recurrent sepsis | 0
skin care | 0
thick scales desquamated | 0
erythematous thick hyperkeratotic plaques | 0
neck involvement | 0
axillae involvement | 0
groin involvement | 0
buttocks involvement | 0
medial aspect of extremities involvement | 0
dorsal aspect of hands and feet involvement | 0
volar aspect of hands and feet involvement | 0
fixed flexion deformity of elbows | 0
fixed flexion deformity of hands | 0
fixed flexion deformity of feet | 0
mitten hand deformity | 0
erythematous scaly plaque on upper face | 0
whole-exome sequencing | 0
inconclusive results | 0
whole-genome sequencing | 0
novel homozygous missense variant in KDSR | 0
skeletal surveys | 0
no evidence of dysplasia | 0
bone marrow biopsy | 0
congenital megakaryocytic aplasia | 0
skin biopsy | 0
hyperkeratosis | 0
acanthosis | 0
papillary dermis fibrosis | 0
discharged in stable condition | 0
admitted for sepsis | 0
epistaxis | 0
mild subdural hematoma | 0
frequent platelet counts below 20 × 109/L | 0
twice-weekly platelet transfusions | 0
monthly intravenous immunoglobulin | 0
packed red blood cells transfusions | 0
acitretin started | 0
remarkable response to acitretin | 0
acitretin replaced by isotretinoin | 0
slow tapering to 0.5 mg/kg/day | 0
good control of skin condition | 0
flareups during febrile episodes | 0
improvement in scales and erythema | 0
lack of availability of acitretin | 0
placed on platelet transfusions | 0
monthly IVIG | 0
packed RBC transfusions | 0
started acitretin | 0
replaced by isotretinoin | 0
slow tapering | 0
elective cesarean section | 0
prior cesarean section | 0
admitted to NICU | 0
spent 2 months in NICU | 0
transfusions for anemia | 0
transfusions for thrombocytopenia | 0
IV antibiotics for sepsis | 0
scales desquamated | 0
flexion deformities | 0
erythematous plaque on upper face | 0
inconclusive exome sequencing | 0
whole-genome sequencing performed | 0
KDSR variant identified | 0
skeletal survey findings | 0
no dysplasia | 0
bone marrow biopsy findings | 0
skin biopsy findings | 0
discharged stable | 0
subsequent admissions for sepsis | 0
admissions for epistaxis | 0
admissions for subdural hematoma | 0
platelet counts below 20 × 109/L | 0
platelet transfusions initiated | 0
IVIG monthly | 0
RBC transfusions | 0
acitretin initiation | 0
acitretin replacement with isotretinoin | 0
tapering of isotretinoin | 0
skin control | 0
flareups during fever | 0
improvement in skin | 0
