59 years old | 0
    female | 0
    referred to hospital | 0
    high temperature | -336
    orthostatic hypotension | 0
    left thigh pain | -336
    back pain | -360
    left hip pain | -360
    thigh pain (persisted) | -360
    fever | -48
    chills | -48
    sweats | -48
    extreme fatigue | -48
    administration of antipyretic agents | -24
    thigh pain (unbearable) | -24
    surgical procedure to the left ilium | -462096
    staphylococcal osteomyelitis | -462096
    smoker | 0
    hypotension (systolic 70 mmHg) | 0
    pulse 90 beats per minute | 0
    normal temperature | 0
    respiratory rate 15 breaths per minute | 0
    oxygen saturation 96% | 0
    chest X-ray normal | 0
    electrocardiogram normal | 0
    left hip pain (exacerbated on movement) | 0
    elevated white blood cell count | 0
    neutrophilic predominance | 0
    elevated erythrocyte sedimentation rate |3D0
    elevated C-reactive protein | 0
    elevated procalcitonin | 0
    mildly elevated liver enzymes | 0
    mildly elevated creatinine kinase | 0
    febrile | 0
    blood cultures obtained | 0
    antipyretics administered | 0
    empirical antibiotics administered | 0
    CT revealed iliopsoas abscess | 0
    MRI confirmed abscesses | 0
    abscess drainage | 0
    pus aspiration for culture | 0
    bilateral pleuritic pain | 0
    difficulty in breathing | 0
    crackles | 0
    diffuse rhonchi | 0
    hypoxia | 0
    chest X-ray bilateral opacities | 0
    CT thorax nodular infiltrates | 0
    differential diagnosis (septic pulmonary emboli) | 0
    differential diagnosis (ARDS) | 0
    transesophageal echocardiogram negative for endocarditis | 0
    thrombosis investigation negative | 0
    health deterioration | 0
    admission to ICU | 0
    acute respiratory failure | 0
    mechanical ventilation | 0
    S. aureus isolated from blood | 120
    S. aureus isolated from pus | 120
    linezolid started | 120
    weaned from ventilator | 168
    CT reduction of abscess | 360
    CT reduction of lung infiltrates | 360
    confirmed septic pulmonary emboli | 360
    intravenous antibiotics continued | 360
    oral antibiotics continued | 864
    CT complete disappearance of abscesses | 2016
    no concomitant diseases | 0
    no skin infection | 0
    no recent trauma | 0
    no bites | 0
    no intramuscular injections | 0
    cultures of skin negative | 0
    cultures of nares negative | 0
    no right-sided endocarditis | 0
    no thrombosis in lower extremities | 0
    no adjacent bone changes | 0
    no osteomyelitis on MRI | 0
    methicillin-susceptible S. aureus | 120