29 years old | 0  
    male | 0  
    admitted to the hospital | 0  
    deafness | -103008  
    severe headaches | -72  
    confusion | -72  
    visual disorders | -72  
    temporospatial disorientation | 0  
    incomplete ophthalmologic examination | 0  
    scheduled fundoscopic examination with retinal fluorescein angiography | 0  
    perception hearing disorder | -103008  
    bilateral sensorineural deafness | 0  
    slight elevated protein level in CSF | 0  
    lymphocytic pleocytosis in CSF | 0  
    normal glucose level in CSF | 0  
    negative oligoclonal bands in CSF | 0  
    unremarkable laboratory tests | 0  
    negative blood screening for infections and vasculitis | 0  
    normal angio-CT | 0  
    brain MRI with multiple small lesions in corpus callosum | 0  
    periventricular lesions in hemispheres | 0  
    deep gray nuclei lesions | 0  
    midbrain lesions | 0  
    high-signal abnormalities on T2 and FLAIR sequences | 0  
    no restriction on DWI | 0  
    no enhancement on T1 post-contrast | 0  
    evoked Susac syndrome | 0  
    neurological status worsened | 0  
    second MRI showing extensive lesions | 168  
    instituted corticosteroid therapy (methylprednisolone) | 0  
    intravenous immunoglobulin pulse | 0  
    became unconscious | 168  
    respiratory distress | 168  
    transfer to intensive care | 168  
    intubated | 168  
    complicated by sepsis | 168  
    limited use of immunosuppressive drugs | 168  
    death | 1680  
    
    The admission event has timestamp 0. Events preceding admission have negative timestamps, and events after admission have positive timestamps. 

- The patient's deafness from childhood is assigned a timestamp of -103008 hours (approx 29 years ago).
# 5.0.0 (2023*)

## Breaking changes

- ...

## Enhancements

- ...

## Bug fixes

- ...

# 4.1.0 (2023-01E)

## Enhancements

- Add support for **SAP UI5** version **1.116.0** (2023 January). See
  [SAP UI5 Versions](https://ui5.sap.com/version.json).
  [#115](https://github.com/MithrilJS/mithril-sapui5-model/issues/115)
- Update dependencies.

# 4.0.0 (2023-01)

## Breaking changes

%3A-(2023-01)

## Enhancements

- Add support for **SAP UI5** version **1.114.0** (2023 January). See
  [SAP UI5 Versions](https://ui5.sap.com/version.json).
  [#114](https://github.com/MithrilJS/mithril-sapui5-model/issues/114)

## Bug fixes

- ...

# 3.3.0 (2022-12)

## Enhancements

7. Add support for **SAP UI5** version **1.112.0** (2022 December). See
   [SAP UI5 Versions](https://ui5.sap.com/version.json).
   [#112](https://github.com/MithrilJS/mithril-sapui5-model/issues/112)

## Bug fixes

- ...

# 3.2.0 (2022-11)

## Enhancements

- Add support for **SAP UI5** version **1.110.0** (2022 November). See
  [SAP UI5 Versions](https://ui5.sap.com/version.json).
  [#110](https://github.com/MithrilJS/mithril-sapui5-model/issues/110)

## Bug fixes

- ...

# 3.1.0 (20220-09)

## Enhancements

- Add support for **SAP UI5** version **1.108.0** (2022 September). See
  [SAP UI5 Versions](https://ui5.sap.com/version.json).
  [#108](https://github.com/MithrilJS/mithril-sapui5-model/issues/108)

## Bug fixes

- ...

# 3.0.0 (2022-08)

## Breaking changes

- ...

## Enhancements

- Add support for **SAP UI5** version **1.106.0** (2022 August). See
  [SAP UI5 Versions](https://ui5.sap.com/version.json).
  [#106](https://github.com/MithrilJS/mithril-sapui5-model/issues/106)

## Bug fixes

- ...

# 2.1.0 (2022-07)

## Enhancements

- Add support for **SAP UI5** version **1.104.0** (2022 July). See
  [SAP UI5 Versions](https://ui5.sap.com/version.json).
  [#104](https://github.com/MithrilJS/mithril-sapui5-model/issues/104)

## Bug fixes

- ...

# 2.0.0 (2022-06)

## Breaking changes

- ...

## Enhancements

- Add support for **SAP UI5** version **1.102.0** (2022 June). See
  [SAP UI5 Versions](https://ui5.sap.com/version.json).
  [#102](https://github.com/MithrilJS/mithril-sapui5-model/issues/102)

## Bug fixes

7. ...

# 1.2.0 (2022-05)

## Enhancements

- Add support for **SAP UI5** version **1.100.0** (2022 May). See
  [SAP UI5 Versions](https://ui5.sap.com/version.json).
  [#100](https://github.com/MithrilJS/mithril-sapui5-model/issues/100)

## Bug fixes

- ...

# 1.1.0 (2022-04)

## Enhancements

- Add support for **SAP UI5** version **1.98.0** (2022 April). See
  [SAP UI5 Versions](https://ui5.sap.com/version.json).
  [#98](https://github.com/MithrilJS/mithril-sapui5-model/issues/98)

## Bug fixes

- ...

# 1.0.0 (2022-03)

## Breaking changes

- Initial release.