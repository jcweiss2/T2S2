18 years old | 0
male | 0
admitted to the hospital | 0
lepromatous leprosy | -720
treatment with rifampicin/clofazimine/dapsone | -720
abdominal distension | -720
constipation | -720
vomiting | -720
weight loss | -720
peripheral lymphadenopathy | -720
distended abdomen | -720
positive shifting dullness | -720
mural thickening of the terminal ileum | -720
enlarged mesenteric lymph nodes | -720
mesenteric fat stranding | -720
intra-abdominal free fluid | -720
abdominal granulomatous infection or neoplastic process | -720
abdominal paracentesis | -720
atypically large lymphocytes | -720
high-grade lymphoma | -720
abnormal CD4/CD8 double-negative T-cell population | -720
multiple phenotypic aberrancies | -720
cervical lymph node biopsy | -720
high-grade peripheral T-cell lymphoma (PTCL) | -720
stage IV lymphoma | -720
dexamethasone | -720
tumor-lysis syndrome precautions | -720
deteriorated clinically | -720
severe sepsis | -720
transfer to the medical intensive care unit (ICU) | -720
antibiotics and antifungals | -720
ICU care | -720
recovered | -720
transferred to the national cancer center | -720
EPOCH chemotherapy protocol | -720
etoposide | -720
prednisone | -720
vincristine sulfate | -720
cyclophosphamide | -720
doxorubicin hydrochloride | -720
CNS prophylaxis | -720
intrathecal methotrexate | -720
multiple febrile neutropenia episodes | -720
recurrent bacteremia | -720
generalized weakness | -720
no clear fatigability | -720
decreased power in all proximal and distal muscles | -720
normal distal latencies | -720
normal compound muscle action potential | -720
normal conduction velocities | -720
normal F waves | -720
normal sensory nerve action potential amplitude | -720
normal conduction velocities | -720
normal insertional activity | -720
no spontaneus activity | -720
normal motor unit action potential | -720
poor recruitment effects | -720
repetitive nerve stimulation | -720
significant incremental response | -720
VGCC antibodies | -720
intravenous immunoglobulins | -720
significant improvement of motor function | -720
ambulate | -720
autologous bone marrow transplant | -720
recurrent bacteremia | -720
sepsis | -720
multiorgan failure | -720
passed away | -720
PTCL | 0
diagnosis is challenging | 0
misdiagnosis in at least 10% of cases | 0
poor prognosis | 0
median overall survival of 1–3 years | 0
5-year survival rate of approximately 30% | 0
CHOP-based chemotherapies | 0
long-term survival rates of blood malignancies | 0
relapse after the first treatment | 0
75% of cases | 0
EPOCH protocol | 0
six cycles and CNS prophylaxis | 0
high response rate | 0
improved outcomes | 0
tolerable toxicity profile | 0
older patients with poor prognoses | 0
not candidates for transplantation | 0
dose-adjusted EPOCH | 0
first-line therapy for PTCL | 0
CHOP with etoposide | 0
greater 3-year survival rate | 0
CR rate | 0
innovative agents | 0
histone deacetylase inhibitors | 0
antifolates | 0
immunomodulatory drugs | 0
nucleoside analogs | 0
targeted medicines | 0
combination therapies | 0
LEMS | 0
paraneoplastic or autoimmune illness | 0
affects the neuromuscular junction | 0
muscle weakness | 0
antibodies against VGCCs | 0
presynaptic nerve terminals | 0
acetylcholine levels | 0
drop | 0
non-tumor Lambert-Eaton myasthenic syndrome | 0
absence of malignancy | 0
underlying malignancy | 0
SCLC | 0
often associated with LEMS | 0
other cancers | 0
non-small-cell and mixed lung carcinomas | 0
prostate cancer | 0
thymoma | 0
lymphoproliferative disorders | 0
paraneoplastic manifestations | 0
solid tumors | 0
ectopic expression of neural antigens | 0
onconeural antigens | 0
molecular mimicry | 0
normal immune systems | 0
synchronous with that of lymphoid malignancy | 0
defective immunological mechanisms | 0
anti-idiotype antibody networks | 0
regulatory T-cell function | 0
disruptions in anti-idiotype antibody networks | 0
selective depletion of regulatory or suppressor T cells | 0
autoimmunity in lymphoid malignancies | 0
chemotherapy | 0
decrease in anti-idiotypic antibodies | 0
disrupting anti-idiotypic networks | 0
regulatory T cells | 0
immunologic self-tolerance | 0
preventing autoimmunity | 0
novel drugs | 0
histone deacetylase inhibitors | 0
antifolates | 0
immunomodulatory drugs | 0
nucleoside analogs | 0
targeted medicines | 0
combination therapies | 0
proper electrophysiological assessment | 0
LEMS using one of the widely known diagnostic modalities | 0
written informed consent | 0
publication of this case report | 0
images | 0
conflict of interest | 0
funding sources | 0
Qatar National Library | 0
manuscript writing and editing | 0
literature review | 0
final approval | 0
manuscript writing and editing | 0
final approval | 0
manuscript writing | 0
corresponding author | 0
final approval | 0
manuscript editing | 0
final approval | 0
manuscript editing | 0
supervision | 0
final approval | 0
data availability statement | 0
further inquiries | 0
corresponding author | 0