30 years old | 0
    gravida 1 | 0
    para 0 | 0
    admitted to a local hospital | 0
    preterm labor | 0
    prenatal laboratories unremarkable | -120
    negative GBS screen | -120
    complete antenatal steroid course | -72
    two doses of betamethasone intramuscular | -72
    latency antibiotics | -72
    ampicillin intravenous | -72
    azithromycin oral | -72
    magnesium for neuroprotection | -48
    preterm labor at 23 weeks | -48
    male neonate | 0
    23 and 4/7 weeks gestational age | 0
    vaginally delivered | 0
    prolonged rupture of membranes | 0
    BW 0.595 kg | 0
    initially vigorous | 0
    intubation | 0
    surfactant for respiratory distress | 0
    APGAR score 5, 6, 8 | 0
    admitted to NICU | 0
    high-frequency oscillator | 0
    respiratory support | 0
    caffeine intravenous | 0
    umbilical catheters inserted | 0
    evaluation for bacterial infection | 0
    empiric therapy with ampicillin and gentamicin | 0
    negative blood culture | 48
    ampicillin and gentamicin discontinued | 48
    nil per os | 0
    total parenteral nutrition | 0
    trialed on conventional mechanical ventilation | 22
    failed mechanical ventilation | 60
    increased oxygen needs | 60
    respiratory acidosis | 60
    transferred to another facility | 72
    leukocytosis | 99
    WBC 19.8K/µL | 99
    bandemia 15% | 99
    septic workup | 99
    blood culture from umbilical arterial catheter | 99
    UVC unable to draw blood culture | 99
    empiric treatment with ampicillin and cefepime | 99
    nationwide shortage of cefotaxime | 99
    abdomen discolored | 99
    abdominal radiograph | 99
    gasless abdomen | 99
    absence of pneumoperitoneum | 99
    absence of portal venous gas | 99
    blood culture positive for gram negative rods | 99
    M. morganii | 99
    umbilical arterial catheter removed | 99
    full sepsis workup | 120
    repeat blood cultures | 120
    peripheral blood culture | 120
    UVC blood culture | 120
    lumbar puncture | 120
    nonsterile urine culture | 120
    antibiotic coverage broadened to meropenem and ampicillin | 120
    speciation pending | 120
    cover for extended spectrum β lactamases | 120
    CSF analysis | 120
    7 red blood cells per µL | 120
    1 WBC per mm³ | 120
    206 mg/dL protein | 120
    78 mg/dL glucose | 120
    CSF culture grew Enterococcus faecalis | 120
    nonsterile urine culture positive for multiple organisms | 120
    Staphylococcus epidermis | 120
    M. morganii | 120
    E. faecalis | 120
    peripheral culture positive for M. morganii | 120
    UVC culture negative | 120
    clinical improvement | 120
    bilious emesis | 192
    increased abdominal discoloration | 192
    never on enteral feeds | 0
    colostrum started | 24
    abdominal radiograph | 192
    free intraperitoneal air | 192
    pneumatosis absent | 192
    SIP | 192
    peritoneal drain placed | 192
    intraoperative peritoneal culture grew M. morganii | 192
    antibiotic coverage changed to vancomycin and fluconazole | 192
    M. morganii sensitivities returned | 192
    meropenem changed back to ampicillin and cefepime | 192
    14-day antibiotic course | 336
    delivery record revisited | 96
    placental maternal culture grew E. coli | 96
    Streptococcus viridans | 96
    coagulase negative Staphylococcus | 96
    Enterococcus | 96
    Bacillus fragilis | 96
    Prevotella species | 96
    M. morganii septicemia | 96
    bacterial translocation from GI tract | 96
    SIP related | 96
    continued clinical improvement | 192
    uncomplicated hospital course | 192
    intestinal perforation healed | 192
    peritoneal drain removal | 192
    enteral feeds advanced | 192
    full enteral feeds | 192
    dexamethasone for chronic lung disease | 240
    extubated | 720
    weaned to room temperature | 2688
    patent ductus arteriosus treated with acetaminophen | 240
    bilateral germinal matrix hemorrhages | 240
    mildly dilated ventricles | 240
    normalized ventricles by discharge | 3024
    corrected full-term cranial ultrasound | 3024
    small left-sided periventricular cyst | 3024
    no ventricular dilation | 3024
    no periventricular white matter changes | 3024
    stage 2 retinopathy of prematurity | 3024
    discharged home | 3024
    corrected GA 41 and 4/7 weeks | 3024
    high-risk infant follow-up clinic | 4032
    corrected GA 6 months | 4032
    feeding therapy | 4032
    infant development services | 4032
    physical therapy | 4032
    normal cognitive skills | 4032
    normal expressive language | 4032
    normal fine motor skills | 4032
    normal gross motor skills | 4032
    normal sensory processing | 4032
    mild delays in receptive language | 4032
    mild delays in social emotional skills | 4032
    outpatient MRI showed no structural abnormality | 4032
    M. morganii sepsis | 99
    LOS | 99
    peritonitis | 192
    SIP | 192
    survived | 3024
    developmental delays | 4032
    maternal antibiotic exposure | -72
    ampicillin resistance | 99
    initial antibiotic therapy with ampicillin and gentamicin | 0
    inadequate coverage | 48
    third-generation cephalosporin and aminoglycoside suggested | 48
    M. morganii bacteremia source GI translocation | 96
    SIP complication | 192
    high mortality in preterm infants | 3024
    survival | 3024
    mild developmental delays | 4032
    negative BCX | 48
    negative UCX | 120
    negative CSF CX | 120
    positive blood cultures | 99
    positive peritoneal culture | 192
    positive peripheral culture | 120
    negative UVC culture | 120
    maternal BCX | 96
    placental cultures | 96
    GI flora contamination | 120
    improved clinical status | 3024
    respiratory distress | 0
    hypotension | 192
    intraventricular hemorrhage | 3024
    NEC | 192
    hydrocephalus | 3024
    VP shunt | 3024
    septic shock | 192
    pulmonary hemorrhage | 192
    stillborn delivery | 96
    apnea of prematurity | 0
    respiratory acidosis | 60
    bilious emesis | 192
    abdominal discoloration | 99
    pneumoperitoneum | 192
    spontaneous intestinal perforation | 192
    peritoneal drain | 192
    ampicillin discontinuation | 48
    gentamicin discontinuation | 48
    cefepime initiation | 99
    meropenem initiation | 120
    vancomycin initiation | 192
    fluconazole initiation | 192
    ciprofloxacin use | 336
    netilmicin use | 336
    amikacin use | 336
    clindamycin use | 192
    cefotaxime shortage | 99
    ELBW program | 72
    APGAR scores improvement | 10
    respiratory distress syndrome | 0
    chronic lung disease | 240
    corrected GA at discharge | 3024
    patent ductus arteriosus treatment | 240
    germinal matrix hemorrhages | 240
    retinopathy of prematurity | 3024
    VP shunt placement | 3024
    psychomotor delay | 4032
    completed antibiotics | 3024
    improved clinical status | 3024
    mortality | 3024
    morbidity | 3024
    gram-negative sepsis | 99
    bacteremia | 99
    facultative anaerobic gram-negative rod | 99
    nosocomial infections | -72
    GI tract infections | 96
    genitourinary tract infections | 96
    neonatal sepsis | 99
    EOS association | 96
    LOS association | 99
    antibiotic resistance | 99
    β-lactamase expression | 99
    maternal ampicillin use | -72
    induced resistance | -72
    neonatal inflammatory markers | 99
    septicemia | 99
    intraabdominal complications | 192
    NEC with perforation | 192
    brain abscess | 3024
    seizures | 3024
    slight psychomotor delay | 4032
    developmental assessment | 4032
    feeding therapy | 4032
    physical therapy | 4032
    outpatient MRI | 4032
    normal structural brain | 4032
    no signal abnormality | 4032
    high-risk follow-up | 4032
    corrected GA 6 months | 4032
    mild delays | 4032
    normal skills | 4032
    literature review | 0
    case reports | 0
    variable clinical presentation | 0
    preterm infants | 0
    EOS cases | 0
    LOS cases | 0
    antibiotic regimens | 0
    complications | 0
    outcomes | 0
    mortality rate | 3024
    morbidity rate | 3024
    hepatobiliary tract infection | 96
    soft tissue infection | 96
    urinary tract infections | 96
    GI translocation | 96
    polymicrobial growth | 120
    contaminated specimen | 120
    adequate antibiotic coverage | 192
    inappropriate antibiotic coverage | 48
    increased mortality risk | 3024
    neonatal literature outcomes | 3024
    extremely premature survival | 3024
    LOS survival | 3024
    SIP survival | 3024
    developmental outcomes | 4032
    conflict of interest | 0
    