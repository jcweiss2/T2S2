50 years old | 0
female | 0
abdominal pain | -240
nausea | -240
vomiting | -240
collapsed | -240
transferred to hospital | -240
acute surgical abdomen | 0
CT scan | 0
appendix with enhanced oedematous wall | 0
retroperitoneal subhepatic air | 0
mild collection | 0
perforated subhepatic appendix | 0
diagnosed as acute abdomen | 0
peritonitis | 0
sepsis | 0
urgent laparotomy | 0
pus evacuated | 0
retrocecal appendix | 0
subhepatic appendix | 0
perforated appendix | 0
retrograde appendectomy | 0
culture and sensitivity swabs | 0
abdomen washed | 0
suction drains secured | 0
admitted to surgical intensive care unit | 0
treated with antimicrobials | 0
estimated recovery and discharge | 0
did not improve as expected | 24
drains continued to drain pus | 24
respiratory distress | 48
intubated | 48
mechanically ventilated | 48
second abdominal CT scan | 72
ill-defined retroperitoneal collection | 72
ultrasound-guided drainage procedure | 96
drained 300 ml of pus | 96
condition improved | 120
extubated | 120
discharged from ICU | 120
accidentally removed drains | 168
repeated CT scan | 168
well-defined enhanced collections | 168
infectious fat necrosis | 168
offered another drain attempt | 168
refused procedure | 168
discharged from hospital | 216
sent home on cefepime | 216
sent home on vancomycin | 216
sent home on metronidazole | 216