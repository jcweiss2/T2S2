9 years old | 0
female | 0
eastern Indian origin | 0
no significant past medical history | 0
admitted to the emergency room | 0
abdominal pain | -72
fever | -72
nausea | -72
vomiting | -72
completed Pfizer-BioNTech COVID-19 immunization series | -744
SARS-CoV-2 PCR test positive | -384
asymptomatic at the time of test | -384
rapid antigen test negative | -384
traveled to US Virgin Islands | -384 to -288
multiple mosquito bites | -384 to -288
persistent fever | -72 to -24
emesis | -72 to -24
nausea (persistent) | -72 to -24
abdominal pain (persistent) | -72 to -24
respiratory viral PCR panel negative | -24
oseltamivir dose | -24
decreased intake | -24
painful area at the tip of the tongue | -24
persistent symptoms leading to emergency department | 0
maximum temperature 40°C | 0
heart rate 124-133 bpm | 0
respiratory rate 20/30 breaths/min | 0
oxygen saturation 96% to 100% | 0
blood pressure 94-102/44-54 mm Hg | 0
mild conjunctival injection | 0
epigastric abdominal tenderness | 0
hyponatremia | 0
leukopenia | 0
thrombocytopenia | 0
lymphopenia | 0
elevated inflammatory markers | 0
SARS-CoV-2 PCR negative | 0
rapid streptococcal antigen test negative | 0
urinalysis abnormalities | 0
IVIG started | 0
ceftriaxone started | 0
doxycycline started | 0
antibiotics discontinued after 72 hours | 72
negative cultures | 72
parasite and viral testing sent | 0
macular nonpruritic nonpetechial rash | 5
rash over neck and hands | 5
sparing of palm and soles | 5
bilateral conjunctival injection | 24
resolved conjunctival injection | 168
afebrile after IVIG completion | 24
prednisone started | 0
confusion episodes | 24
agitation episodes | 24
DVT prophylaxis initiated | 0
anticoagulation discontinued | 0
aspirin not started | 0
unremarkable echocardiogram | 0
inflammatory markers trended downward | 72
pancytopenia persisted | 72
hemoglobin nadir 9.7 g/dL | 72
RBC count nadir 3.61 M/uL | 72
platelet count nadir 30,000/uL | 72
WBC count nadir 2580 cells/uL | 72
absolute lymphocyte count nadir 240 | 72
BNP peak 4114 pg/mL | 72
BNP down trended to 429 pg/mL | 168
normal echocardiography | 0, 72, 168
complement levels normal | 72
ANA positive 1:320 | 72
dsDNA normal | 72
Smith antibodies normal | 72
IL-6 elevated | 72
CXCL-9 elevated | 72
negative DAT | 72
peripheral smear negative for blasts | 72
bone marrow aspiration not performed | 72
thrombocytopenia improved on day 7 | 168
platelet count 104,000/uL at discharge | 168
met criteria for MIS-C | 0
recent positive COVID-19 PCR | -384
fever | -72 to -24
gastrointestinal symptoms | -72 to -24
broad differential diagnosis | 0
negative infectious disease tests | 72
considered HLH | 72
considered ITP | 72
considered DIT | 72
considered MAS | 72
considered sHLH | 72
considered systemic juvenile idiopathic arthritis | 72
considered malignancy | 72
platelet count recovery | 168
ALC recovery | 168
WBC recovery | 168
Hgb recovery | 168
mild persistent fatigue after 2 months | 168
follow-up by specialists | 168
no alternative diagnosis within 4 months | 168
multi-specialty team utilized | 0
IVIG treatment completed | 24
steroids tapered | 72
thrombocytopenia resolution | 168
discharged | 168
