58 years old | 0
male | 0
hypertension | 0
diabetes mellitus | 0
admitted to ICU | 0
septic shock | 0
invasive mechanical ventilation | 0
norepinephrine infusion | 0
febrile | 0
central venous catheter | -144
coronary artery bypass grafting | -312
mitral valve replacement | -312
renal function deteriorated | 0
creatinine clearance higher than 40 ml/min | 0
preserved urine output | 0
CVC removal | 0
blood samples drawn | 0
urine culture | 0
bronchoalveolar lavage | 0
mediastinitis diagnosis improbable | 0
CT scan | 0
transthoracic echocardiography | 0
transesophageal echocardiography | 0
valvular abnormality not shown | 0
empirical antibiotic treatment started | 0
Vancomycin treatment | 0
Imipenem treatment | 0
Colistin treatment | 0
clinical condition worsened | 24
Klebsiella pneumoniae isolated | 24
catheter culture | 24
blood samples culture | 24
Kp intermediate to Amikacin | 24
Kp resistant to Imipenem | 24
Kp resistant to Colistin | 24
Kp resistant to Tigecycline | 24
PCR and sequencing performed | 24
blaOXA-48 gene identified | 24
blaVIM-2 gene identified | 24
blaCMY-2 gene identified | 24
blaSHV-1 gene identified | 24
Vancomycin stopped | 48
Colistin stopped | 48
amikacin treatment started | 48
Imipenem dose increased | 48
CVVHDF started | 49
amikacin dose increased | 72
norepinephrine stopped | 120
CRP decreased | 120
procalcitonin decreased | 120
leukocytes decreased | 120
treatment tolerated | 336
discharged from ICU | 384
serum creatinine values similar to before ICU admission | 384
audiometric test performed | 384
ototoxicity excluded | 384