71 years old | 0
female | 0
hypertension | 0
presented to the emergency department | -4320
dyspnea on exertion | -4320
malaise | -2160
anorexia | -2160
fatigue | -2160
unintentional weight loss | -2160
atrial fibrillation | 0
heart failure | 0
referred to internal medicine service | 0
abdominal ultrasound | 0
pelvic ultrasound | 0
clinical ascites | 0
bilateral adnexal masses | 0
solid and cystic changes | 0
abdominal CT scan | 0
solid peritoneal deposits | 0
moderate ascites | 0
large volume ascites | 0
ovarian malignancy suspected | 0
CA-125 level low | 0
discharged home | 0
urgent follow-up | 0
assessed at gynecology-oncology clinic | 120
paracentesis performed | 120
malignant cells | 120
poorly differentiated carcinoma | 120
sarcoma | 120
epithelioid morphology | 120
planned 3 cycles of Paclitaxel | 120
planned 3 cycles of Carboplatin | 120
interval debulking | 120
presumed epithelial ovarian cancer | 120
received first dose of chemotherapy | 264
presented to emergency department | 384
diarrhea | 384
fatigue | 384
generalized weakness | 384
afebrile | 384
clinically dehydrated | 384
hypotension | 384
pre-renal acute kidney injury | 384
pancytopenic | 384
received volume resuscitation | 384
received PRBC | 384
received GCSF | 384
received prophylactic antibiotics | 384
diagnosis of tumour lysis syndrome | 384
AKI | 384
hyperphosphatemia | 384
hypocalcemia | 384
uric acid elevated | 384
given Rasburicase | 384
transferred to ICU | 384
intubation | 384
hypoxic respiratory failure | 384
volume overload | 384
vasopressor support | 384
septic shock | 384
CRRT initiated | 384
blood cultures grew Group B streptococcus | 384
urine positive for E. coli | 384
continued piperacillin-tazobactam | 384
remained dependant on CRRT | 384
no improvement in haemodynamic state | 384
no improvement in respiratory status | 384
developed fungemia | 384
clinical deterioration | 384
opted for comfort care | 384
life support withdrawn | 384
passed away | 384
autopsy | 384
intramural uterine malignant neoplasm | 384
extensive necrosis | 384
undifferentiated endometrial stromal sarcoma | 384
metastatic involvement | 384
marked autolytic changes | 384
granular casts | 384
- dyspnea on exertion | -480
9malaise | -2640
- anorexia | -2640
: fatigue | -2640
- unintentional weight loss | -2640
