60 years old | 0
female | 0
bipolar disorder | 0
hyperlipidemia | 0
osteoporosis | 0
renal stone | 0
water pipe smoker | 0
electrical burn scar | 0
suicidal behavior | 0
admitted to intensive care unit | 0
dizziness | 0
drowsiness | 0
drug poisoning | 0
amphetamine | 0
benzodiazepine | 0
decreased Glasgow Coma Scale to 9 | 24
decreased Glasgow Coma Scale to 3 | 24
right bundle branch block | 24
complete bundle branch block | 24
therapeutic hemodialysis | 24
severe abdominal distension | 72
lack of defecation | 72
absence of bowel sounds | 72
multiloculated fluid collection | 72
GI perforation | 72
severe peritonitis | 72
transferred to operation room | 72
laparotomy | 72
stomach perforation | 72
acute peritonitis | 72
bowel adhesion repair | 72
stomach perforation repair | 72
retro-gastric fluid collection | 72
sub-diaphragmatic fluid collection | 72
generalized peritonitis | 72
drainage | 72
acute acalculous cholecystitis | 72
chronic acalculous cholecystitis | 72
focal mucosal necrosis | 72
severe constipation | 336
abdominal distention | 336
ascites | 336
edema | 336
multicoated fluid collection | 336
septation | 336
second laparotomy | 336
sepsis | 336
disseminated intravascular coagulation | 336
increased serum BUN | 336
increased serum creatinine | 336
renal failure | 336
cardiorespiratory arrest | 336
death | 336
CMV gastritis | 0
ulceration | 0
foreign body-type giant cell reaction | 0
CMV immunoreactivity | 0
CMV DNA in gall bladder | 0
CMV DNA in gastric wall | 0
