15 years old | 0
female | 0
admitted to the hospital | 0
shortness of breath | -3
chest pain | -3
cough | -24
difficulty breathing | -24
haemoptysis | -3
coryzal symptoms | -168
no cutaneous injury or pathology | -168
no past medical history | 0
no history of immunodeficiency | 0
no drug or food allergies | 0
crackles and reduced air entry in the lower right hemithorax | 0
tachypnoeic | 0
saturating at 92% on room air | 0
heart rate 120 beats/min | 0
blood pressure 105/74 mmHg | 0
afebrile | 0
cold extremities | 0
pH 7.42 | 0
PaCO2 4.0 kPa | 0
PaO2 7.2 kPa | 0
blood lactate 1.7 mmol/L | 0
sodium bicarbonate level 19.5 mmol/L | 0
base excess -5 mmol/L | 0
leukopaenia | 0
neutrophil count 0.8 × 10^9/L | 0
c-reactive protein 3.7 mg/L | 0
full blood count | 0
c-reactive protein results | 0
plain erect radiographs of the chest | 0
rapidly progressive consolidation | 0
four-quadrant opacification | 0
ARDS | 0
diagnostic and therapeutic bronchoscopy | 3
copious yellow, protein-rich plasma-like secretions | 3
bronchial washings | 3
PVL-Staphylococcus aureus | 6
influenza A/H3N2 | 6
surviving sepsis protocols | 1
IV ceftriaxone | 1
enteral azithromycin | 1
enteral oseltamivir | 1
IV linezolid | 6
IV clindamycin | 6
IV ceftriaxone | 6
IV clarithromycin | 6
non-invasive ventilation | 3
emergency intubation | 3
mechanical ventilation | 3
refractory shock | 3
high dose adrenaline | 3
noradrenaline | 3
fluid resuscitation | 3
20% human albumin solution | 3
crystalloids | 3
bedside transthoracic echocardiography | 3
cardiac arrest | 12
ECMO cannulation | 12
venoarterial-ECMO | 12
cardiopulmonary resuscitation | 12
IV corticosteroid | 12
IV immunoglobulin | 12
bronchoalveolar fluid aspiration | 12
VV-ECMO | 18
retained cannula in the left common iliac artery | 18
ischaemia of the distal limbs | 18
disseminated intravascular coagulation | 18
multiple organ failure | 18
conversion of VA-ECMO to VV-ECMO | 24
collateral circulation | 24
adequate lower limb perfusion | 24
extubation | 744
good neurological function | 744
respiratory and functional rehabilitation | 744
renal replacement therapy | 744
transfer to a non-tertiary hospital | 1296
intensive physiotherapy | 1296
mobility improvement | 1296
skin grafting to the left lower leg | 1296
non-healing wounds | 1296
independently mobile | 2592
community rehabilitation services | 2592