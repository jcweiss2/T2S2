63 years old | 0
male | 0
benign prostatic hyperplasia | 0
urinary retention | 0
chronic obstructive pulmonary disease | 0
hypertension | 0
hyperlipidemia | 0
osteoarthritis | 0
foot surgery | -6720
antihypertensives | -672
nebulization | -672
declined history of malignant hyperthermia | 0
declined family history of malignant hyperthermia | 0
elevated baseline creatinine | 0
general anesthesia | 0
induced with lidocaine | 0
induced with propofol | 0
induced with fentanyl | 0
supraglottic laryngeal mask airway | 0
inhaled sevoflurane | 0
spontaneous breathing | 0
stable end tidal CO2 | 0
received fentanyl for analgesia | 0
received ondansetron for antiemesis | 0
surgery uneventful | 0
extubated | 0
transported to recovery unit | 0
alert | 0
awake | 0
non-anxious | 0
comfortable | 0
normothermic | 0
normal oxygen saturation | 0
normotension | 0
normal heart rate | 0
normal respiratory rate | 0
muscle rigidity | 40
elevated temperature | 40
elevated blood pressure | 40
tachypnea | 40
tachycardia | 40
malignant hyperthermia suspected | 40
malignant hyperthermia protocol initiated | 40
malignant hyperthermia hotline contacted | 40
reintubated with propofol | 40
radial artery cannulation | 40
lab studies performed | 40
dantrolene administered | 40
elevated CO2 | 40
elevated white blood cell count | 40
elevated creatine kinase | 40
no more muscle rigidity | 80
normalized blood pressure | 80
normalized CO2 | 120
stable white blood cell count | 120
stable creatine kinase | 120
malignant hyperthermia deemed unlikely | 120
sepsis suspected | 120
blood cultures drawn | 120
clinically stable | 120
hemodynamically stable | 120
extubated | 240
transferred to intensive care unit | 240
elevated temperature improved | 360
white blood cell count improved | 360
creatinine kinase improved | 360
managed for urosepsis | 360
antibiotics administered | 360
discharged home | 720