52 years old | 0
male | 0
diabetes | 0
myelofibrosis | 0
admitted to the hospital | 0
hemorrhagic vesicular eruption | 0
vesiculobullous lesions | 0
necrotic eschar-covered erosive ulcerated lesions | 0
right eye discharge | 0
pale | 0
unwell | 0
severe lower gastrointestinal bleeding | 0
blood pressure 98/54 mmHg | 0
temperature 36.7°C | 0
platelets 396×10^9 | 0
white blood cells 17×10^9/L | 0
hemoglobin 5.7 G/dL | 0
WBC differential 85% neutrophils and 8% lymphocytes | 0
platelet large cell ratio 40% | 0
arterial blood gas analyses pH 7.36 | 0
pCO2 36.9 mmHg | 0
pO2 31 mmHg | 0
aO2 33.4% | 0
urea 39.7 mmol/L | 0
creatinine 290 µmol/L | 0
aspartate transaminase 424 U/L | 0
alanine transaminase 395 U/L | 0
direct bilirubin 20.8 µmol/L | 0
international normalized ratio 3.6% | 0
partial thromboplastin time 45.9 seconds | 0
prothrombin time 46.9 seconds | 0
history of severe beta-lactam-induced allergic reactions | 0
anaphylaxis suspected | 0
septic shock suspected | 0
bacterial culture positive for Pseudomonas aeruginosa | 24
histopathological findings of epidermal necrosis and sloughing | 24
Gram stain preparation of the tissue revealed numerous gram-negative rods | 24
upper and lower gastrointestinal endoscopies performed | 24
no necrotic, inflammatory, or pathologic causes of bleeding found | 24
diagnosis of ecthyma gangrenosum-induced septic shock | 48
levofloxacin initiated | 72
discharged from the intensive care unit | 240
renal and liver functions normal | 1008
coagulation profile normal | 1008
amikacin administered | -72
E. coli-infected amputation stump of the big toe | -72