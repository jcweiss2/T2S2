31 years old | 0
female | 0
SLE | -8760
lupus nephritis | -8760
prior stroke | -8760
intravenous drug use | -8760
admitted to the hospital | 0
cardiogenic shock | 0
mental status changes | 0
elevated jugular venous pressure | 0
prominent v wave | 0
body temperature 36.3°C | 0
blood pressure 95/66 mm Hg | 0
heart rate 94 beats/min | 0
hemoglobin 10.3 g/dL | 0
white blood cell count 18.9 × 10^9/L | 0
platelet count 64 × 10^9/L | 0
international normalized ratio 3.6 | 0
creatinine level 1.7 mg/dL | 0
drug studies positive for narcotics | 0
drug studies positive for cannabis | 0
antiphospholipid serology normal | 0
blood cultures negative | 0
intravenous antibiotics | 0
broad-spectrum intravenous antibiotics | 0
serologic studies | 0
operative cultures | 0
mitral valve prosthesis dehiscence | 0
severe mitral regurgitation | 0
perivalvular regurgitation | 0
annular pseudoaneurysm | 0
transthoracic echocardiography | 0
transesophageal echocardiography | 0
surgical intervention | 0
fourth sternotomy | 24
mitral valve reconstruction | 24
bioprosthesis | 24
bovine pericardium | 24
left atrial dome reconstruction | 24
interatrial septal incision | 24
postbypass TEE | 48
extracorporeal membrane oxygenation | 48
left ventricular ejection fraction 25% | 48
sluggish flow in the left atrium | 48
multiple blood product transfusions | 48
layered thrombus in the left atrium | 120
surgical clot removal | 120
thrombus reaccumulation | 120
extracorporeal membrane oxygenation withdrawn | 144
patient died | 144