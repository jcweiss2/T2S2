26 years old | 0
premenopausal | 0
nulliparous | 0
hypogastric pain | -24
analgesics | -24
uterine myomatosis | -168
pelvic ultrasound | -168
analgesics | -168
abnormal uterine bleeding | 0
abdominal pain | 0
no prior chronic or systemic disease | 0
no prior surgeries | 0
no prior pregnancies or deliveries | 0
regular menstrual cycle | 0
no family history of chronic diseases or cancer | 0
depressible abdomen | 0
tender abdomen | 0
slight increase in hypogastrium volume | 0
normal laboratory findings | 0
negative reverse transcription PCR | 0
MRI mass in posterior uterine wall | 0
T1-weighted hyperintense component | 0
T2-weighted hyperintense component | 0
T1-weighted hyperintense halo | 0
hematic content | 0
liquid content | 0
low ADC value | 0
leiomyoma with red degeneration | 0
pyomyoma differential diagnosis | 0
laparoscopic myomectomy | 0
hypovascularized myoma | 0
friable tissue | 0
postoperative sepsis | 12
hypotension | 12
tachycardia | 12
fever | 12
respiratory distress | 12
drowsiness | 12
intensive care admission | 12
oxygen therapy | 12
fluid resuscitation | 12
empiric antibiotic therapy | 12
anemia | 12
leukocytosis | 12
bandemia | 12
high C-reactive protein | 12
procalcitonin elevation | 12
pCO2 | 12
HCO3 | 12
BEb | 12
lactate | 12
uterine leiomyoma with necrosis | 12
gram-negative cocci bacteria | 12
adjusted antibiotic therapy | 12
normalization of inflammatory markers | 36
clinical improvement | 36
uterine myomatosis with red degeneration | 0
pyomyoma | 0
