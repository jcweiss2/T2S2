65 years old | 0
male | 0
admitted to the hospital | 0
diarrhea | -48
hypotensive | 0
febrile | 0
temperature of 38.4 °C | 0
vomited | -48
brown and green stools | -48
no blood or mucous in stools | -48
contact with granddaughter with diarrheal illness | -72
no significant past medical history | 0
no medication | 0
unvaccinated for rotavirus | 0
distended abdomen | 0
non-tender abdomen | 0
abdomen resonant to percussion | 0
audible bowel sounds | 0
clear chest | 0
equal air entry to both lungs | 0
peripheral limb pulses not palpable | 0
cool peripheries | 0
hemoglobin level 160 g/L | 0
white cell count 18.1×10^9/L | 0
platelet count 128×10^9/L | 0
hypokalemia | 0
potassium level 2.7 mmol/L | 0
raised inflammatory markers | 0
C-reactive protein level 144 mg/L | 0
procalcitonin 235 µg/L | 0
ferritin 2708 µg/L | 0
creatinine level 286 µmol/L | 0
lactate level 6.9 mmol/L | 0
blood cultures sterile | 0
urine cultures sterile | 0
respiratory swabs negative | 0
rotavirus detected in feces | 0
no typing or titer for rotavirus | 0
no other viruses detected | 0
no ova, cysts, and parasites | 0
no bacterial pathogens | 0
cerebrospinal fluid testing negative | 0
high sensitivity troponin level 834 ng/L | 0
type-2 acute myocardial infarction | 0
new anteroinferior T-wave inversion | 0
no ventricular or valvular dysfunction | 0
ischemic liver injury | 0
alanine transaminase 1124 U/L | 0
aspartate transaminase 1101 U/L | 0
hepatitis screen negative | 0
serology testing for hepatitis A, B, and C negative | 0
HIV 1 and 2 negative | 0
urinary albumin/creatinine ratio 112.7 mg/mmol | 0
glomerulonephritis screen negative | 0
acute tubular necrosis | 0
atypical antineutrophil cytoplasmic antibodies pattern | 0
myeloperoxidase and proteinase-3 immunofluorescence negative | 0
CT angiogram of abdomen and pelvis | 0
moderate dilatation of small bowel | 0
entire dilatation of large bowel | 0
no transition point | 0
no clinical evidence of bowel obstruction | 0
resuscitation with intravenous crystalloid rehydration | 0
adrenaline infusion | 0
noradrenaline infusion | 0
potassium infusion | 0
empirical antibiotic cover | 0
vancomycin | 0
piperacillin-tazobactam | 0
intubation | 0
transfer to Intensive Care Unit | 0
continuous renal replacement therapy | 24
intermittent inpatient hemodialysis | 168
transfer to ward | 120
renal function improvement | 720
liver function improvement | 720
amlodipine | 720
aspirin | 720
nosocomial urinary tract infection | 720
pneumonia | 720
urine culture grew Escherichia coli | 720
i.v. meropenem | 720
transfer to subacute facility | 1008
discharged home | 1176