66 years old | 0
female | 0
diffuse pruritus | -168
erythroderma | -168
lymphadenopathy | -168
biopsy | -168
atypical cells with irregular nuclei | -168
abnormal CD3+ CD4+ CD7− CD26− T-cell clone | -168
Sézary cell count of 2312 | -168
positron emission tomography scan | -168
bilateral lymphadenopathy | -168
uncontrolled hypertension | 0
type 2 diabetes | 0
end-stage renal disease | 0
extracorporeal photopheresis | 0
bexarotene | 0
lost to follow-up | -84
pruritus worsened | -84
Sézary count climbed to 11,132 | -84
COVID-19 infection | -56
short of breath | -56
afebrile | -56
recovered fully without medication | -28
Sézary count dropped to 6494 | -28
admitted to the hospital with severe COVID-19 | 0
shortness of breath | 0
chills | 0
fever | 0
hypoxemia | 0
dexamethasone | 0
empiric antibiotics | 0
lymphocyte count began to decrease | 14
discharge from hospital | 25
Sézary count dropped to 936 | 60
romidepsin | 90
pruritus improved | 120
erythroderma resolved | 120
lymphadenopathy resolved | 120
Sézary counts dropped to 389 | 120
admitted to the intensive care unit again | 180
severe COVID-19 | 180
encephalopathy | 180
hypotension | 180
cardiac arrest | 180
death | 180