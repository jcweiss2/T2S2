18 years old | 0  
    Saudi woman | 0  
    presented to the emergency department | -336  
    right lower quadrant (RLQ) abdominal pain | -336  
    nausea | -336  
    vomiting | -336  
    anorexia | -336  
    no fever | -336  
    decayed wheat consumption | -672  
    abdomen distended | 0  
    RLQ tenderness | 0  
    RLQ fullness | 0  
    CT scan of abdomen and pelvis | 0  
    obstructing caecal mass | 0  
    colonoscopy | 0  
    necrotic caecal mass | 0  
    multiple biopsies | 0  
    necrotic tissue | 0  
    decision for surgery | 0  
    laparotomy | 0  
    right hemicolectomy | 0  
    primary anastomosis | 0  
    histopathology negative for malignancy | 0  
    ulcerations | 0  
    necrosis | 0  
    microabscesses | 0  
    multinucleated giant cells | 0  
    fungal hyphae | 0  
    started on amphotericin B | 0  
    postoperative jaundice | 24  
    postoperative high fever | 24  
    postoperative per-rectal bleeding | 24  
    white cell count 33×109/L | 24  
    eosinophilia | 24  
    deranged liver function tests | 24  
    CT scan showing intra-abdominal collection | 24  
    right paracolic gutter collection | 24  
    peritonitis | 24  
    multiple hepatic abscesses | 24  
    exploratory laparotomy | 48  
    ileal perforation | 48  
    white patches over abdominal wall | 48  
    white patches over small bowel | 48  
    white patches over liver | 48  
    bowel resection | 48  
    anastomosis | 48  
    biopsies for histology | 48  
    biopsies for cultures | 48  
    fungal hyphae invading bowel wall | 48  
    Splendore-Hoeppli phenomenon | 48  
    liver biopsies with fungal hyphae | 48  
    Basidiobolus species | 48  
    Candida | 48  
    Klebsiella pneumoniae | 48  
    started on voriconazole | 48  
    started on tigecycline | 48  
    started on meropenem | 48  
    enterocutaneous fistula | 72  
    vacuum-assisted closure | 72  
    total parenteral nutrition (TPN) | 72  
    tapered TPN | 168  
    regular diet | 168  
    inflammatory markers normalized | 168  
    white cell count normalized | 168  
    liver function tests normalized | 168  
    fever spikes to 39°C | 192  
    CT scan showing enlarged paracolic gutter collection | 192  
    common hepatic artery aneurysm | 192  
    porta hepatis/caudate collection | 192  
    large right pleural effusion | 192  
    transferred to tertiary center | 216  
    ultrasound-guided drainage | 216  
    embolisation of aneurysm | 216  
    chest tube insertion | 216  
    follow-up CT scan | 240  
    ruptured liver abscess | 240  
    liver abscess drainage | 240  
    conservative treatment | 240  
    liver abscess cultures Basidiobolus | 240  
    started on liposomal amphotericin B | 240  
    started on posaconazole | 240  
    seizures | 264  
    MRI showing brain edema | 264  
    cortical laminar necrosis | 264  
    meningoencephalitis | 264  
    intubation | 264  
    inotropes | 264  
    CT scan showing lung abscesses | 264  
    expired | 288  

<|eot_id|>