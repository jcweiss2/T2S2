60 years old | 0
male | 0
Asian | 0
hypertensive | 0
diabetic | 0
admitted to the hospital | 0
fever | -72
persistent productive cough | -72
chest pain | -72
myalgias | -72
fatigue | -72
respiratory distress | -72
past history of TB | -10080
unprotected contact with COVID-19 positive individual | -72
decreased breath sounds at the lung bases | 0
saturation of peripheral oxygen (SpO2) 72% | 0
bilateral interstitial infiltrates on portable chest X-ray | 0
lymphocytopenia | 0
increased C-reactive protein | 0
increased lactate dehydrogenase | 0
increased ferritin | 0
diffuse bilateral ground-glass opacities on chest CT scans | 0
COVID-19 confirmed by RT-PCR | 0
admitted to isolation chamber | 0
high flow nasal cannula (HFNC) initiated | 0
awake prone positioning initiated | 0
empiric therapy for COVID-19 started | 0
lopinavir/ritonavir and ribavirin started | 0
dexamethasone started | 0
prophylactic anticoagulation started | 0
nucleic acid amplification test (NAAT) revealed concomitant infection with mycobacterium tuberculosis | 24
isoniazid started | 24
rifampicin started | 24
pyrazinamide started | 24
ethambutol started | 24
HFNC and awake prone positioning discontinued | 288
oxygen therapy administered | 288
oxygen supportive care discontinued | 384
RT-PCR test for COVID-19 negative | 480
microbiology negative | 480
discharged to home isolation | 648