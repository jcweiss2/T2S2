75 years old | 0
woman | 0
brought to the emergency department | 0
unconscious | 0
productive cough | -96
fever | -96
high blood pressure | 0
paroxysmal atrial fibrillation | 0
type 2 diabetes | 0
bisoprolol | 0
propafenone | 0
atorvastatin | 0
metformin | 0
aspirin | 0
nonsmoker | 0
no occupational exposures | 0
tachypnoea | 0
tachycardia | 0
atrial fibrillation | 0
normal blood pressure | 0
transcutaneous arterial oxygen saturation decreased to 86% | 0
auscultation of the lungs | 0
diffuse wheezing | 0
diminished breath sounds | 0
mild dullness at the right base of the lung | 0
severe inflammation | 0
white blood cell count 20.9×109 cells per L | 0
neutrophils 17.2×109 cells per L | 0
C-reactive protein 326.1 mg·L−1 | 0
elevated liver transaminases | 0
alanine aminotransferase 3216 U·L−1 | 0
aspartate aminotransferase 4359 U·L−1 | 0
decreased kidney function | 0
creatinine 313 µmol·L−1 | 0
urea 26.2 mmol·L−1 | 0
severe hypercapnic respiratory failure | 0
carbon dioxide tension (PaCO2) of 107 mmHg | 0
oxygen tension (PaO2) of 63 mmHg | 0
pH 7.04 | 0
HCO3− 28.9 mmol·L−1 | 0
chest CT | 0
pulmonary oedema | 0
right-sided infiltrates | 0
aspiration pneumonia | 0
right-sided aspiration pneumonia | 0
antibiotic therapy with intravenous piperacillin/tazobactam | 0
invasive mechanical ventilation | 0
intubated | 0
transferred to the intensive care unit | 0
regained consciousness | 24
laboratory tests returned to normal | 24
cultures from bronchoalveolar lavage positive for Haemophilus influenzae | 24
persistent hypercapnic respiratory failure | 24
PaCO2 71 mmHg | 24
PaO2 85 mmHg | 24
pH 7.34 | 24
HCO3− 38.3 mmol·L−1 | 24
tracheostomy performed | 24
mechanical ventilation discontinued | 360
breathing spontaneously through the tracheostomy tube | 360
dyspnoea | 360
mild weakness | 360
hypercapnia | 360
pressure support ventilation continued | 360
multiple attempts to evacuate the tracheostomy tube unsuccessful | 360
severe shortness of breath | 360
stridor | 360
acute respiratory insufficiency | 360
bronchoscopy | 360
tracheal dyskinesia | 360
bilateral vocal cord paresis | 360
CT of the head and chest | 360
no major cerebrovascular pathology | 360
no mediastinal pathology | 360
no recent history of surgery | 360
no recent history of trauma | 360
neuromuscular pathology suspected | 360
persistent hypercapnic respiratory failure | 360
dysphagia | 360
slight muscular weakness in the proximal leg muscles | 360
fatigability of the extraocular muscles | 360
myasthenia gravis suspected | 360
critical illness polyneuropathy | 360
Guillain–Barré syndrome | 360
AChR antibodies negative | 360
not tested for MuSK antibodies | 360
RNS studies performed | 360
decremental muscle electrical response up to 20% | 360
myasthenia gravis diagnosed | 360
pyridostigmine 150 mg·day−1 | 360
prednisolone 5 mg·day−1 | 360
dosing gradually increased to 45 mg·day−1 | 360
status greatly improved | 360
dyspnoea disappeared | 360
difficulty breathing disappeared | 360
hypercapnia resolved | 360
PaCO2 returned to normal | 360
active | 360
capable of all self-care | 360
permanent tracheostomy tube placed | 360
discharged | 360
neuromuscular respiratory failure (NRF) | 360
myasthenia gravis | 360
amyotrophic lateral sclerosis | 360
respiratory failure | 360
muscle weakness | 360
neuromuscular disorder | 360
outcomes poor | 360
severe disability | 360
acute NRF | 360
myasthenic crisis | 360
myopathies | 360
disease progression | 360
superimposed respiratory disease | 360
compensatory mechanisms overwhelmed | 360
impaired transmission at the neuromuscular junction | 360
fluctuating weakness | 360
fatigability of the skeletal muscles | 360
ptosis | 360
diplopia | 360
ocular myasthenia gravis | 360
generalised disease | 360
bulbar muscles | 360
facial muscles | 360
neck muscles | 360
limb muscles | 360
proximal weakness | 360
respiratory muscles | 360
advanced disease | 360
serological testing | 360
electrophysiological tests | 360
acetylcholinesterase inhibitor | 360
pyridostigmine | 360
neostigmine | 360
ambenonium chloride | 360
immunosuppressive therapy | 360
prednisone | 360
azathioprine | 360
mycophenolate mofetil | 360
methotrexate | 360
cyclosporine | 360
tacrolimus | 360
rituximab | 360
thymectomy | 360
plasma exchange | 360
intravenous immune globulin | 360
critical illness polyneuropathy (CIP) | 360
neuromuscular weakness | 360
critical illness myopathy | 360
severe sepsis | 360
multiorgan failure | 360
mitochondrial function | 360
stress hormones | 360
cytokines | 360
nitric oxide | 360
ischaemic hypoxia | 360
cytopathic hypoxia | 360
axon degeneration | 360
sodium channels | 360
flaccid and symmetrical weakness | 360
moderate paresis | 360
reduced deep-tendon reflexes | 360
severe quadriplegia | 360
muscle wasting | 360
hypotonia | 360
sensory impairment | 360
distal loss of pain | 360
temperature loss | 360
vibration loss | 360
primary axonal degeneration | 360
reduction in CMAP | 360
sensory nerve action potential amplitudes | 360
no decremental response | 360
supportive treatment | 360
aggressive treatment of sepsis | 360
early rehabilitation | 360
bulbar dysfunction | 360
hypercapnic respiratory failure | 360
persistent bilateral vocal cord paresis | 360
long-term tracheostomy | 360
permanent tracheostomy | 360
CIP | 360
NRF | 360
ICU setting | 360
early recognition | 360
aggressive treatment | 360
outcomes improved | 360
