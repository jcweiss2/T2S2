31-year-old pregnant woman | 0  
    no family history of congenital heart disease | 0  
    referred to centre | -7680  
    foetal aortic valve stenosis | -7680  
    first detected at 18 + 0 weeks of gestation | -7680  
    maternal transabdominal foetal ultrasound imaging at 28 + 4 weeks of gestation | -168  
    severe foetal aortic valve stenosis | -168  
    poorly contracting dilated left ventricle | -168  
    severe mitral valve regurgitation | -168  
    local endocardial fibroelastosis | -168  
    severe mitral regurgitation | -168  
    papillary muscle ischaemia | -168  
    mitral valve inflow biphasic | -168  
    regurgitant velocity exceeded 4 m | -168  
    maximum systolic flow velocity across thickened aortic valve 2 m/s | -168  
    flow across oval foramen left to right | -168  
    retrograde flow inside aortic arch | -168  
    percutaneous ultrasound-guided foetal balloon valvuloplasty attempted at 29 + 4 weeks of gestation | 0  
    general maternofoetal anaesthesia | 0  
    left ventricular function deteriorated further | 0  
    mitral valve flow integral exhibited mostly a-wave filling | 0  
    foetus in dorsoanterior cephalic position | 0  
    left ventricle pointed posteriorly | 0  
    conventional percutaneous ultrasound-guided approach not accessible | 0  
    foetoscopic assistance employed | 0  
    three 11 Fr catheter sheaths percutaneously placed along left flank of foetus | 0  
    amniotic cavity insufflated with carbon dioxide | 0  
    foetoscope introduced through trocars | 0  
    graspers introduced through trocars | 0  
    foetus rotated dorsoposterior position | 0  
    upper extremities postured along foetal sides | 0  
    successful foetoscopic foetal posturing | 0  
    insufflation gas removed | 0  
    18 gauge needle percutaneously advanced into foetal left ventricle | 0  
    needle placed underneath obstructed aortic valve | 0  
    maternal transabdominal foetal echocardiographic guidance | 0  
    successful foetal balloon valvuloplasty achieved via needle shaft | 0  
    3.5 mm coronary angioplasty catheter used | 0  
    mother tolerated procedure well | 0  
    foetus tolerated procedure well | 0  
    no complications observed | 0  
    interventional materials removed | 0  
    maternal skin incisions closed with single stitches | 0  
    marked improvement of flow across aortic valve | 24  
    increase in flow velocity from 1.75 m/s prior to intervention to more than 3 m/s after intervention | 24  
    semi-compliant balloon with inflated diameter 3.5 mm used | 0  
    inflated diameter smaller than aortic annulus | 0  
    decompression observed | 0  
    improved function of left ventricle observed for about 2 weeks | 336  
    further foetal growth | 504  
    fixed stenosis became more effective | 504  
    foetus delivered in third week after prenatal intervention | 504  
    scheduled for postnatal re-valvuloplasty on second day of life | 504  
    infant underwent stent insertions in ductus arteriosus | 504  
    stent insertions in atrial septum | 504  
    insertion of flow occluders into both pulmonary branches | 504  
    two more aortic valvuloplasties carried out | 504  
    left ventricular function improved over time | 504  
    baby died at 6 months of age | 4320  
    Escherichia coli septicaemia | 4320  
    long-standing central venous line | 4320  
    another cardiac surgery addressing mitral valve regurgitation | 4320  
    branch pulmonary artery obstruction | 4320  
    percutaneous ultrasound-guided procedure performed following parental informed consent | 0  
    foetoscopy-assisted procedure performed following parental informed consent | 0  
    ethical standards for human experimentation established by Declaration of Helsinki | 0  
    minimally invasive approach | 0  
    less invasive alternative to maternal laparotomy | 0  
    foetoscopy-assisted foetal transoesophageal echocardiography | 0  
    three-trocar technique combined with insufflation | 0  
    minimally invasive foetoscopic pacemaker insertion | 0  
    techniques developed in foetal sheep models | 0  
    safe anaesthesia protocol for human foetoscopic surgery | 0  
    used for foetal surgery for spina bifida | 0  
    used for haemodynamically compromised foetuses with congenital high airway obstruction syndrome | 0  
    amniotic fluid leakage | 504  
    mean age at delivery 33 weeks of gestation | 504  
    maternal bedrest | 504  
    infection prophylaxis | 504  
    neonatal cardiac intensive care management | 504  
    interventions | 504  
    surgery | 504  
    baby died from Escherichia coli septicaemia | 4320  
    consent obtained from patient | 4320  
    conflict of interest none declared | 4320  
    funding received from Deutsche Forschungsgemeinschaft | 4320  
    development of percutaneous foetoscopic techniques supported by educational and research grants | 4320