43 years old | 0
female | 0
admitted to the hospital | 0
right upper quadrant pain | 0
fevers | 0
vomiting | 0
raised inflammatory markers | 0
raised bilirubin | 0
intravenous antibiotics | 0
abdominal ultrasound demonstrated cholelithiasis | 0
abdominal ultrasound demonstrated choledocholithiasis | 0
no signs of cholecystitis | 0
ERCP | 24
common bile duct cannulated with guidewire | 24
CBD swept via balloon with multiple stones extracted | 24
sphincterotomy performed | 24
CBD stent placed | 24
bile flowed freely through stent | 24
ERCP recovery uneventful | 24
referred to general surgeons | 24
laparoscopic cholecystectomy | 192
surgery uneventful | 192
booked for repeat ERCP and stent removal | 192
appointment postponed due to pandemic | 192
elective ERCP with stent removal | 3504
CBD stent removed | 3504
guidewire passed into biliary tree | 3504
balloon sweep undertaken | 3504
further CBD stones removed | 3504
right shoulder tip pain | 3504
worsening RUQ pain | 3504
pain settled with analgesia | 3504
discharged home | 3504
re-presented with severe RUQ pain | 3528
tachycardic | 3528
CT showed large subcapsular hepatic hematoma | 3528
mass effect on IVC | 3528
advised non-operative management | 3528
repeat hemoglobin testing | 3528
progress CT showed stable hematoma | 3528
pain improved | 3528
discharged | 3600
re-presented with RUQ pain | 4104
shortness of breath | 4104
new fevers | 4104
malaise | 4104
lethargy | 4104
signs of sepsis | 4104
new oxygen requirement | 4104
CT showed continued hematoma | 4104
new right-sided pleural effusion | 4104
admitted under gastroenterology team | 4104
admitted to intensive care | 4104
treated for infected hematoma | 4104
IR guided drainage | 4104
drain did not facilitate resolution | 4104
did not improve sepsis | 4104
consulted UGI surgery team | 4104
laparoscopic washout of infected collection | 4104
right lobe densely adherent to diaphragm | 4104
necrotic capsule present | 4104
partially de-roofed | 4104
drainage of purulent liquid | 4104
necrotic debris suctioned | 4104
old blood suctioned | 4104
required further take back to theater | 4824
on-going fevers | 4824
raised inflammatory markers | 4824
CT showed septated collection | 4824
partial necrosectomy | 4824
cavity irrigated | 4824
no bile leak | 4824
sump drain placed | 4824
Blake drains placed | 4824
continued irrigation of sump drain | 4824
irrigation with normal saline | 4824
IV antibiotics for 40 days | 4824
Klebsiella oxytoca growth | 4824
Escherichia coli growth | 4824
continued drain output monitoring | 4824
no evidence of bile leak | 4824
CT showed reduction of collection | 4824
acute kidney injury | 4824
AKI due to antibiotic toxicity | 4824
acute tubular necrosis | 4824
AKI resolved | 4824
discharged with sump drain | 4824
community nurse reviews | 4824
outpatient clinic reviews | 4824
drain partially removed | 4824
drain completely removed | 4824
no long-term complications | 4824
