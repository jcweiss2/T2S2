69 years old | 0
male | 0
admitted to the hospital | 0
prostate carcinoma | -8760
endoscopic prostatectomy | -8760
adjuvant radiotherapy | -8760
local recurrence of prostate carcinoma | -168
metastatic to bone | -168
docetaxel | -168
tumor induced anemia | -168
Hgb 7.2 g/dL | -168
PSA levels > 200 ng/mL | -168
upper stomach pain | -168
diarrhea | -168
cholecystitis | -168
increased infection parameters | -168
CRP: 280 mg/L | -168
procalcitonin: 6.52 ng/mL | -168
open cholecystectomy | -120
metronidazole | -120
ceftriaxone | -120
blood cultures | -120
purulent gangrenous gallbladder | -120
ileostomy | -120
necrotizing/gangrenous, ulcero-phlegmonous, cholecystitis | -120
fibrinous pericholecystitis | -120
cholecystolithiasis | -120
intraoperative culture | -120
extubated | 24
vasopressor therapy ended | 24
transferred to the ward | 96
discharged | 336
F. plautii detected in blood culture | 96
gram staining | 96
matrix-assisted laser desorption/ionization time of flight (MALDI-TOF) | 96
culture on Columbia agar | 96
16S rRNA sequencing | 120
resistance testing | 120
antimicrobial therapy | 0
improved under treatment | 168
sensitive to metronidazole | 168
sensitive to ceftriaxone | 168
resistant to cotrimoxazole | 168
resistant to fluoroquinolones | 168
intermediate resistance to penicillin | 168
intermediate resistance to linezolid | 168