36 years old | 0
female | 0
admitted to the hospital | 0
fever | -168
hemoptysis | -168
left-sided chest pain | -168
breathlessness | -168
temperature 102°F | 0
respiratory rate 32/min | 0
blood pressure 100/76 mm of Hg | 0
heart rate 108/min | 0
SpO2 of 92% in room air | 0
decreased breath sound on the left side of the chest | 0
crepitation on left infraclavicular, axillary and interscapular area | 0
no significant history of diabetes | 0
no significant history of malignancy | 0
no significant history of drug intake | 0
transferred to Medical Intensive Care Unit | 0
resuscitation of the patient | 0
evaluated for coronary artery diseases | 0
electrocardiography | 0
two-dimensional echo | 0
cardiac markers | 0
normal coronary artery diseases test results | 0
HIV test | 0
HIV test result negative | 0
hepatitis B virus surface antigen test | 0
hepatitis B virus surface antigen test result negative | 0
HCV test | 0
HCV test result negative | 0
autoimmune profile test | 0
autoimmune profile test result negative | 0
Chest X-ray | 0
mass lesion in the left upper and mid-zone of the lung | 0
computed tomography scan thorax with contrast study | 0
large mass-like lesion with contract enhancement | 0
sputum examination | 0
no pathogenic organism in Gram staining | 0
no pathogenic organism in culture reports | 0
fiberoptic bronchoscopy avoided | 0
CT-guided fine-needle aspiration cytology (FNAC) | 0
sample sent for cytological examination | 0
sample sent for Gram staining | 0
sample sent for Ziehl–Neelsen staining | 0
sample sent for aerobic culture | 0
Gram staining showed Gram-positive branching filaments | 0
Gram staining showed coccoid elements | 0
Gram staining suggestive of Nocardia species | 0
conventional Ziehl–Neelsen staining negative | 0
modified Ziehl–Neelsen staining positive | 0
partially acid-fast branching filaments | 0
blood agar plate showed dry whitish-to-tan colonies | 0
colonies showed typical raised, chalky white appearance | 0
colonies showed characteristic earthy odor of Nocardia species | 0
staining of smears from culture showed filamentous bacteria | 0
empirically put on third-generation cephalosporin | 0
empirically put on azithromycin | 0
started cotrimoxazole | 0
rashes all over the body | 24
antibiotic treatment changed to imipenem | 24
imipenem treatment for 10-day duration | 24
started oral linezolid | 240
Chest X-ray showed gradual resolution of pneumonia | 240
Chest X-ray showed cavitation | 240
complete resolution of the left upper lobe lesion | 4320
follow-up chest X-ray | 4320