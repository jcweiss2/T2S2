29 years old | 0 | 0 
male | 0 | 0 
admitted to the hospital | 0 | 0 
biventricular failure | -720 | 0 
ejection fraction 5-10% | -720 | 0 
myopericarditis | -720 | 0 
constrictive physiology | -720 | 0 
peripherally inserted central catheter (PICC) line placed | -720 | 0 
discharged on milrinone | -720 | 0 
fever | -24 | 0 
chills | -24 | 0 
septic shock | 0 | 0 
PICC line removed | 0 | 0 
IV vancomycin | 0 | 24 
piperacillin/tazobactam | 0 | 24 
vasopressor support | 0 | 48 
Chryseobacterium indologenes grew from PICC line | 48 | 48 
Chryseobacterium indologenes grew from peripheral blood cultures | 48 | 48 
antibiotics changed to ciprofloxacin | 48 | 0 
piperacillin/tazobactam | 48 | 336 
weaned off vasopressor support | 48 | 48 
pericardiectomy | 240 | 240 
completed 14 days of antibiotics | 336 | 336 
discharged from the hospital | 336 | 336 
off inotropes | 336 | 336 
stable vital signs | 336 | 336 
stable labs | 336 | 336 
seen in outpatient cardiology clinic | 744 | 744 
remains in good health | 744 | 744 
no evidence of recurrent infection | 744 | 744 
cardiogenic shock | -720 | -720 
atrial flutter | -720 | -720 
radiofrequency ablation | -720 | -720 
inotrope therapy | -720 | 0 
home milrinone infusion | -720 | 0 
elective pericardiectomy | -24 | -24 
fever of 38.7°C | -24 | 0 
tachycardia | -24 | 0 
heart rate in the 110s | -24 | 0 
blood pressure of 96/57 mmHg | -24 | 0 
heart tachycardic | -24 | 0 
normal rhythm | -24 | 0 
no murmurs | -24 | 0 
no rubs | -24 | 0 
no gallops | -24 | 0 
no signs of elevated jugular venous pressure | -24 | 0 
no lower extremity oedema | -24 | 0 
bilateral radial and dorsalis pedis pulses equal | -24 | 0 
lungs clear to auscultation | -24 | 0 
normal work of breathing | -24 | 0 
no redness or drainage around PICC line | -24 | 0 
chest X-ray showed no abnormalities | -24 | 0 
sinus tachycardia | -24 | 0 
normal axis | -24 | 0 
RSR′ pattern in V1 | -24 | 0 
QRS duration of 90 ms | -24 | 0 
non-specific T wave flattening | -24 | 0 
febrile to 39.5°C | 0 | 0 
severe rigours | 0 | 0 
hypotension | 0 | 0 
elevated lactate level of 5.5 mmol/L | 0 | 0 
blood cultures drawn | 0 | 0 
empiric vancomycin | 0 | 24 
piperacillin/tazobactam | 0 | 24 
transferred to cardiac intensive care unit | 0 | 0 
vasopressor support | 0 | 48 
Gram-negative rods | 48 | 48 
Chryseobacterium indologenes | 48 | 48 
ciprofloxacin | 48 | 336 
piperacillin/tazobactam | 48 | 336 
susceptibility testing | 48 | 48 
sensitive to ciprofloxacin | 48 | 48 
sensitive to piperacillin | 48 | 48 
sensitive to trimethoprim/sulfamethoxazole | 48 | 48 
resistant to meropenem | 48 | 48 
improved clinically | 48 | 336 
remained afebrile | 48 | 336 
weaned off vasopressor support | 48 | 48 
follow-up blood cultures remained negative | 168 | 336 
interval echocardiogram | 240 | 240 
dilated and hypertrophied left ventricle | 240 | 240 
diastolic septal bounce | 240 | 240 
constrictive pericarditis | 240 | 240 
ejection fraction of 30-35% | 240 | 240 
right ventricle dilated | 240 | 240 
reduced systolic function | 240 | 240 
no evidence of valvular stenosis | 240 | 240 
no evidence of valvular regurgitation | 240 | 240 
no evidence of vegetations | 240 | 240 
simultaneous right and left heart catheterization | 240 | 240 
discordance of right and left ventricular pressures | 240 | 240 
diastolic equalization of pressures | 240 | 240 
pericardiectomy | 240 | 240 
dense areas of adhesions | 240 | 240 
calcium laterally and towards the apex of the heart | 240 | 240 
adhesions taken down | 240 | 240 
complete removal of pericardium | 240 | 240 
follow-up transthoracic echocardiogram | 288 | 288 
left ventricular ejection fraction increased to 50-55% | 288 | 288 
right ventricular systolic dysfunction improved | 288 | 288 
discharged following completion of antibiotic course | 336 | 336 
inotrope independent | 336 | 336 
guideline-directed medical therapy for heart failure | 336 | 744 
furosemide | 336 | 744 
metoprolol succinate | 336 | 744 
sacubitril-valsartan | 336 | 744 
follow-up with outpatient cardiologist | 744 | 744 
great improvement in functional status | 744 | 744 
denies symptoms of heart failure | 744 | 744 
NYHA Class I | 744 | 744 
no evidence of recurrent infection | 744 | 744