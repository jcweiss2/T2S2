32 years old | 0
female | 0
pregnant | 0
11 weeks pregnant | 0
admitted to the hospital | 0
hyperemesis | 0
sepsis | 0
disseminated intravascular coagulation | 0
admitted to intensive care unit | 0
C. albicans in blood cultures | 0
C. albicans in urine | 0
treatment with L-AMB | 0
treatment with caspofungin | 0
treatment with broad-spectrum antibiotics | 0
lost fetus | -14
discharged from intensive care unit | 18
discharged from hospital | 43
lumbar back pain | 77
pyrexia | 77
CRP 150 mg/l | 77
bone scintigraphy | 85
MRI showed vertebral infection | 90
treatment with caspofungin and fluconazole | 90
biopsy | 91
PCR negative | 91
culture negative | 91
back pain progressed | 104
CRP declined | 104
new MRI showed no regression | 106
treatment failure | 106
treatment changed to L-AMB | 106
slowly improved | 148
discharged | 148
hemodialysis | 148
fluconazole administered after HD | 148
serum fluconazole concentration measured | 148
malaise | 233
vomiting | 233
fluctuating temperature | 233
low back pain | 233
readmitted to hospital | 247
increasing back pain | 247
pyrexia | 247
CRP <8 mg/l | 247
ESR 50 | 247
L-AMB initiated | 252
temporal relief of symptoms | 252
pain returned | 286
L-AMB dose increased | 286
MRI showed progression | 293
L-AMB dose increased to 6 mg/kg | 301
5-FC initiated | 301
PET-CT unchanged | 378
MRI showed minimal regression | 378
bone scintigraphy showed regression | 378
high dose L-AMB continued | 378
leukocyte scintigraphy showed reduced enhancement | 465
MRI showed reduced enhancement | 465
anti-fungal treatment discontinued | 465
ESR remained normal | 538
bone scintigraphy showed minimal activity | 538
no progression on MRI | 538
kidney transplant | 678
gave birth to a healthy child | 1092
no signs of relapse | 1762