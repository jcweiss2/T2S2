26 years old | 0
male | 0
admitted to the hospital | 0
height: 180 cm | 0
weight: 74 kg | 0
kidney transplant | -6048
end-stage kidney disease | -8736
immunosuppression | 0
mycofenolate sodium | 0
methylprednisolone | 0
estimated glomerular filtration rate (eGFR) 35.9 mL/min/1.73 m2 | 0
proteinuria 117 mg/d | 0
chronic kidney transplant disease stage 3bA1 | 0
status post vascular rejection | -6048
chronic calcineurin-inhibitor toxicity | -6048
headache | 0
blurred vision | 0
cranial CT- and MRI scans | 0
methylprednisolone therapy stopped | 0
dexamethasone administered | 0
brain edema | 0
transmitted to the university department of Nephrology | 0
transmitted to the department of Neurosurgery | 0
brain biopsy | 0
diagnosis of cerebral PTLD | 0
diffuse large B-cell lymphoma | 0
positive for Ebstein-Barr virus | 0
CT scan of the thorax | 0
abdomen sonography | 0
bone marrow biopsy | 0
initial chemotherapy regime | 0
high-dose cytarabin | 0
Rituximab | 0
complete remission of PTLD | 24
impairment of the transplant function | 24
eGFR 25.4 mL/min/1.73 m2 | 24
cytomegalovirus (CMV) reactivated | 96
pneumocystis jirovecii pneumonia | 96
chemotherapy changed | 96
Rituximab | 96
antiviral and antibiotic therapy | 96
mycofenolate sodium tapered | 96
generalized seizure | 168
recurrence of PTLD | 168
cerebral MRI scan | 168
HDMTX | 168
Leukovorine | 168
Rituximab | 168
vigorous hydration | 168
HFHD | 192
dialysis procedures | 192
MTX-level measurements | 192
nadir of leucocytes | 216
CMV- and E.coli pneumonia | 240
sepsis | 240
acute kidney transplant failure | 240
transmission to an intensive care unit | 240
invasive ventilation | 240
sepsis managed | 240
discontinuation of mycofenolate sodium | 240
antiviral and antibiotic therapy | 240
follow up cerebral MRI scan | 312
small regredience of PTLD | 312
cerebral radiation | 312
no relevant response of the disease | 312