38 years old | 0
male | 0
admitted to the hospital | 0
abdominal pain | 0
nausea | 0
fever | 0
elevated white cell count | 0
obesity | 0
moderate bilateral symmetrical lower extremity oedema | 0
COVID-19 pneumonia | -336
endotracheal intubation | -336
ventilatory support | -336
CT PE study showed no evidence of PE | -336
pulmonary embolism at the age of 16 | -8032
treated with 6 months of warfarin | -8032
second PE | -2920
chronic thromboembolic pulmonary hypertension | -2920
thromboendarterectomy | -2920
long-term warfarin therapy | -2920
hypercoagulable work-up | -2920
cardiolipin antibody negative | -2920
antithrombin III 92% | -2920
factor V Leiden mutation not identified | -2920
protein C level 147% | -2920
protein S level 58% | -2920
factor II gene mutation not identified | -2920
dilute Russel’s viper venom time 32.9 s | -2920
unremarkable basic metabolic panel | 0
negative high sensitivity troponins | 0
platelets within normal limit | 0
elevated white cell count | 0
INR in therapeutic range | 0
PT elevated to 34.7 s | 0
PTT normal at 37.4 s | 0
CT scan of abdomen showed no abnormalities | 0
incidental finding of a possible filling defect within a partially imaged dilated descending right pulmonary artery | 0
CTPE study showed a large filling defect within the descending right main pulmonary artery | 0
echocardiogram showed a dilated right atrium | 0
bowing of the interatrial septum to the left | 0
severely dilated right ventricle with severely reduced systolic function | 0
diastolic and systolic Left Ventricular septal flattening | 0
dilated inferior vena cava | 0
lower extremity Doppler ultrasounds did not demonstrate a deep vein thrombosis | 0
abdominal infection considered | 0
stress ulcers considered | 0
acute pancreatitis considered | 0
treated with intranasal oxygen | 0
supportive care | 0
transiently on unfractionated intravenous heparin therapy | 0
decision to continue on warfarin with a slightly higher INR target range | 0
advised to follow closely with the haematology department | 0
discharged | 72
follow-up attempts made | 72
patient did not respond to follow-up reminders | 72