24 years old | 0
male | 0
hyperthyroidism | -672
noncompliant with methimazole treatment | -672
MVA | -1
loss of consciousness | -1
self-extricated from the wreckage | -1
ambulatory at the scene | -1
right lower quadrant abdominal pain | -1
right wrist pain | -1
ethanol consumption | -1
heart rate 170 | -1
blood pressure 156/78 | -1
heart rate 163 | 0
blood pressure 153/84 | 0
temperature 37.3°C | 0
Glasgow Coma Score 15 | 0
anxious | 0
fine tremor | 0
hematoma over the left eye | 0
seat belt sign to the left chest | 0
right-sided abdominal tenderness | 0
left hand abrasions | 0
right wrist pain | 0
no neck abrasions or contusions | 0
no goiter | 0
focused abdominal sonography for trauma exam negative | 0
head, maxillofacial, chest, abdomen, and pelvis computed tomography scans negative | 0
plain radiographs of the extremities negative | 0
resuscitated with 2 L of normal saline | 0
IV lorazepam 2 mg | 0
IV fentanyl 50 mcg | 0
laboratory testing | 0
sodium 149 | 0
potassium 3.4 | 0
chloride 108 | 0
carbon dioxide 15 | 0
anion gap 26 | 0
BUN 11 | 0
creatinine 0.51 | 0
AST 43 | 0
ALT 58 | 0
lactic acid 7.6 | 0
free T4 5.61 | 0
thyroid stimulating hormone <0.015 | 0
rapid urine drug screen positive for cannabinoids | 0
ethanol level 101 | 0
serum osmolality 288 | 0
osmolar gap -6 | 0
ethylene glycol negative | 0
methanol negative | 0
hypertensive | 0
tachycardic | 0
TC suspected | 0
methimazole 5 mg | 0
propranolol 1 mg injection | 0
fluid resuscitation continued | 0
admitted to internal medicine service | 0
lactic acidosis improved to 0.8 | 7
sodium 143 | 7
chloride 109 | 7
CO2 21 | 7
anion gap 13 | 7
AST 24 | 7
ALT 50 | 7
blood glucose 102-85 | 7
tachycardia and hypertension resolved | 24
methimazole 5 mg 3 times daily | 24
propranolol 10 mg 3 times daily | 24
blood cultures negative | 24
discharged | 48
follow-up with endocrinology | 48
noncompliant with follow-up | 2160
TC again | 2160
tonsillitis | 2160