69 years old | 0
female | 0
stabbed herself in the abdomen | -1
admitted to the emergency department | 0
blood pressure could not be measured | 0
pulseless electrical activity | 0
body temperature was 35.0 °C | 0
oxygen saturation was 99 % | 0
Glasgow Coma Scale score of 3 | 0
agonal respiration | 0
wound measuring 5 cm on her upper abdomen | 0
intra-abdominal fluid collection | 0
emergency thoracotomy | 0
aortic cross-clamping | 0
open cardiac massage | 0
administration of epinephrine | 0
temporary return of spontaneous circulation | 0
hemodynamically unstable | 0
laparotomy | 0
injuries to the common hepatic and splenic arteries | 0
injuries to the pancreas, spleen, and liver | 0
ligation of the injured arteries | 0
distal pancreatectomy | 0
splenectomy | 0
liver sutured | 0
administration of norepinephrine | 0
second-look surgery | 24
no signs of active bleeding | 24
no ischemic change | 24
no vasopressor requirement | 72
abdominal wall closure | 72
enhanced computed tomography scan | 96
disruption of the celiac artery | 96
gastroduodenal artery arising from superior mesenteric artery | 96
gastroscopy | 216
patchy mucosal necrosis | 216
conservative treatment | 216
fever of 39 °C | 552
pain in the stomach | 552
white blood cell count of 34,000/mm3 | 552
C reactive protein of 13.4 mg/dL | 552
CT scan | 552
air in the gastric wall | 552
intra-abdominal free air | 552
gastric necrosis | 552
emergency surgery | 552
total gastrectomy with Roux-en-Y reconstruction | 552
histological findings of the stomach | 552
diffuse necrotic changes | 552
leakage on the duodenal stump | 696
continuous tube drainage | 696
sepsis due to multidrug-resistant Pseudomonas aeruginosa infection | 1680
disseminated intravascular coagulation | 1680
death | 1680