57 years old | 0
female | 0
visual disturbance | -1440
diplopia | -1440
headaches | -1440
admitted to the hospital | -1440
MRI showed an osteolytic, irregular enhancing lesion occupying the clivus | -1440
TSS | -1440
excisional biopsy was consistent with a chordoma with chondroid differentiation | -1440
tumor not totally removed | -1440
diplopia again | -720
MRI showed that the clival chordoma had increased in size | -720
extended TSS | -720
tumor still remained | -720
postoperative CSF leakage was not observed | -720
tumor had increased again on follow-up MRI | -600
Gamma knife radiosurgery | -600
treatment dose was 18.5 Gy at the tumor margin | -600
proton beam radiotherapy | -420
treatment dose was 6,960 cGy in 29 fractions | -420
unpleasant odor inside her nasal cavity | -120
visited the radiation-oncology department | -120
took antibiotic drugs and steroids | -120
symptoms did not resolve | -120
visited our emergency medical team | 0
copious epistaxis | 0
odor inside her nasal cavity | 0
systemic inflammatory response syndrome | 0
body temperature was 38.2 degrees | 0
WBC was 30,040/mm3 | 0
brain CT scan | 0
comatose mental state | 0
low blood pressure due to septic shock | 0
cardiopulmonary resuscitation | 0
vital signs recovered | 0
CSF examination by lumbar puncture | 0
MRI without enhanced gadolium | 0
exploration inside the nasal cavity with a nasal endoscope | 0
synthetic materials used in the reconstruction of the sellar floor | 0
nasal septum defect due to necrosis | 0
pale and fibrotic mucous membrane | 0
scarring and narrowing of the blood vessels | 0
disruption and necrosis of the membrane | 0
CSF rhinorrhea was not observed | 0
tissue was not biopsied | 0
Enterococcus avium and Escherichia coli were identified on the mucosal culture | 0
CSF examination revealed an increased WBC count | 0
protein level was 345 mg/dL | 0
glucose level was 4 mg/dL | 0
Enterococcus avium and Escherichia coli were identified on the CSF culture and blood culture | 0
diagnosed with bacterial meningitis | 0
administered antibiotic therapy | 0
expired a week later | 168