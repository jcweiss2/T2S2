63 years old | 0
male | 0
admitted to the hospital | 0
respiratory distress | 0
COPD | -672
community-acquired pneumonia | 0
COPD exacerbation | 0
IV moxifloxacin | 0
corticosteroids | 0
intubated | 24
difficult respiratory weaning | 48
widening of the antibiotic spectrum | 48
moxifloxacin ceased | 216
IV ciprofloxacin | 216
piperacillin-tazobactam | 216
hypotensive | 216
feverish | 216
hemocultures negative | 216
cerebral CT scan unremarkable | 216
thoracic CT scan unremarkable | 216
abdominal CT scan unremarkable | 216
cardiac ultrasound unremarkable | 216
sepsis of unknown origin | 216
IV vancomycin | 360
piperacillin-tazobactam substituted to meropenem | 456
fluconazole introduced | 456
oligoanuric acute kidney injury | 360
serum creatinine rising | 360
aggressive fluid administration | 360
IV vitamin C | 456
IV hydrocortisone | 456
IV thiamine | 456
renal replacement therapy | 552
urea elevated | 552
creatinine elevated | 552
estimated GFR decreased | 552
microscopic hematuria | 552
proteinuria | 552
urine sediment revealed calcium oxalate crystals | 552
urinary sodium elevated | 552
urinary creatinine elevated | 552
serum sodium elevated | 552
serum creatinine elevated | 552
serum vitamin C elevated | 552
anti-glomerular basement membrane antibodies negative | 552
perinuclear anti-neutrophil cytoplasmic antibodies negative | 552
proteinase 3 anti-neutrophil cytoplasmic antibodies negative | 552
antibiotics withheld | 552
continuous RRT initiated | 552
renal biopsy performed | 552
acute tubular damage | 552
intratubular translucent crystals | 552
calcium oxalate crystals | 552
glomeruli showed ischemic changes | 552
arterial section revealed discrete intimal fibrosis | 552
immunofluorescence study did not show significant staining | 552
RRT required for several weeks | 600
full renal recovery | 1000
physical rehabilitation | 1000
return home | 1200