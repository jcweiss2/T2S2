40 years old | 0
male | 0
admitted to the hospital | 0
severe left-sided abdominal pain | -120
nausea | -120
vomiting | -120
fevers | -120
rigors | -120
dysuria | -120
dark-colored urine | -120
temperature of 103.3 F | 0
pulse 160 beats/min | 0
blood pressure 102/71 mm Hg | 0
respiratory rate of 28 | 0
92% oxygen saturation | 0
marked tenderness over the left abdomen and flank | 0
left costovertebral angle tenderness | 0
no overlying erythema or warmth of the skin | 0
mildly distended abdomen | 0
no hepatosplenomegaly | 0
no rebound tenderness | 0
no guarding | 0
WBC count of 8,600/µl | 0
serum creatinine of 2.7 mg/dL | 0
total bilirubin of 1.8 mg/dL | 0
alanine aminotransferase 66 U/L | 0
unremarkable urinalysis | 0
blood cultures taken | 0
piperacillin-tazobactam | 0
CT scan | 0
retroperitoneal fluid collection | 0
fascial edema | 0
tachycardia | 24
pain persisted | 24
frequent febrile episodes | 24
WBC increased to over 15,000/µl | 24
hemodynamically stable | 24
breathing comfortably on room air | 24
blood cultures grew group A streptococcus | 24
antibiotic changed to ceftriaxone and clindamycin | 24
abdomen less distended | 48
parasthesia on the left abdomen, flank, and groin | 48
pitting edema of the involved area | 48
no erythema, warmth, or bullae formation | 48
repeat CT scan | 120
persistence of fluid along the left flank musculature and fascial planes | 120
drainage catheter placed | 120
turbid yellow fluid obtained | 120
cell count of 31,400 WBC | 120
gram stain showed many PMNs with no organisms | 120
cultures yielded no growth | 120
immediate pain relief | 120
fever resolution | 120
output from the drain | 120
CT scan showed significant improvement in the amount of fluid | 168
complete renal recovery | 168
bilirubin and alanine aminotransferase normalized | 168
discharged with home infusion of ceftriaxone | 168
elevated ESR | 168
continued on therapy for six weeks | 504
follow-up CT showed near resolution of fascial edema and fluid | 672
full recovery | 672