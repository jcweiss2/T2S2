Here is the table of events and timestamps:

18 years old | 0
male | 0
born | -40
by caesarean section | -40
in the 40th week of gestation | -40
with a birth weight 2100 g | -40
(SDS = –4.86 for gestational age) | -40
birth length 48 cm | -40
(SDS = –1.71 for gestational age) | -40
in good condition (8 points in the Apgar scale) | -40
prominent forehead | -40
relative macrocephaly | -40
limb asymmetry | -40
5th finger clinodactyly of both hands | -40
2/3 toe syndactyly of both legs feet | -40
hypomethylation of the 11p15 region of the paternal chromosome | -17
gene H19 | -17
delayed motor development | -17
walked independently in 16th month of life | -16
hepatic dysfunction | -14
increased concentration of alanine aminotransferase (AlAT 469 U/l) | -14
increased concentration of aspartate aminotransferase (AspAT 439 U/l) | -14
markedly increased creatine kinase level (21 470 U/l) | -14
diagnosis of Duchenne muscular dystrophy | -14
mutation of the maternal DMD gene located on the X chromosome | -14
exon deletion 49–50 | -14
DMD was diagnosed in asymptomatic phase | -14
shortly afterwards health problems typical for DMD appeared | -14
significantly often falling | -14
tiptoed | -14
Achilles tendon contractures | -14
Gover’s syndrome positive | -14
calf enlargement | -14
treated with corticosteroids | -4
prednisone (5 to 6 mg/day) | -4
deflazacort (6 mg/day) | -2
significantly slower height velocity | -2
height velocity 3.3 cm/year | -2
qualified for G-CSF treatment | -6
G-CSF treatment | -6
G-CSF analogue | -6
granulocyte colony stimulating factor (G-CSF) | -6
5 µg/kg/day | -6
5 consecutive days | -6
first, second, third, sixth, and twelfth month | -6
elongation of the distance covered in the 6-minute walk test (6MWT) | -6
334/385 metres to 330/420 metres | -6
sepsis | -6
treatment in the Intensive Care Unit | -6
severe hypoglycaemia | -6
neurological symptoms | -6
glucose level of 14 mg/dl (0.78 mmol/l) | -6
urological care due to hypospadias | -6
cardiological diagnostics | -6
episodes of sinus tachycardia | -6
heart murmur (2/6 degree in Levine scale) | -6
cardiomyopathy excluded | -6
treated with propranolol (15 mg per day in 3 equal doses of 5 mg) | -6
significant deficiency of height and body weight | -6
diagnosed in the Department of Paediatric Endocrinology and Diabetology | -6
growth hormone deficiency excluded | -6
maximum secretion of growth hormone in the sleep test was 31.6 ng/dl | -6
growth hormone deficiency excluded | -6
fulfilled the criteria for treatment with rhGH | -6
treated with rhGH | -6
0.035 mg/kg/per day | -6
improvement of auxological parameters and height velocity | -6
height velocity 6.9 cm/year | -6
IGF-1 increased | -6
exceeding the upper limit of the norm | -6
BMI increased | -6
21.9 kg/m2 (BMI SDS = 1.43) | -6
worsening of glucose metabolism and increasing insulin resistance | -6
HOMA-IR 9.66 | -6
IGT and insulin resistance | -6
distance covered in 6MWT decreased | -6
303/348 m to 315 m | -6
abnormal, weakened gait | -6
rapid weight gain | -6
impaired glucose tolerance | -6
behavioural treatment with lifestyle modification | -6
recommended | -6
rhGH dose reduced to 0.03 mg/kg | -6
2.8 cm growth | -6
rhGH therapy discontinued | -6
auxological and hormonal evaluation | -6
Table II | -6
Patient’s characteristics before the treatment and during the first year of rhGH therapy | -6
Measures | -6
Pre-rhGH | -6
6 months on rhGH | -6
12 months on rhGH | -6
Age (year) | -6
8.9 | -6
9.4 | -6
9.9 | -6
Height (cm) | -6
118.6 | -6
122.0 | -6
125.2 | -6
Height SDS | -6
–2.97 | -6
–2.69 | -6
–2.47 | -6
BMI (kg/m2) | -6
16.6 | -6
18.1 | -6
21.1 | -6
SDS-BMI | -6
–0.2 | -6
0.37 | -6
1.18 | -6
IGF-1 (ng/ml) [normal range] | -6
294 [74–388] | -6
413 [74–388] | -6
457 [88–452] | -6
IGFBP-3 (µg/ml) [normal range] | -6
5.76 [2.1–7.7] | -6
6.83 [2.1–7.7] | -6
7.44 [2.1–7.7] | -6
HbA1c (%) | -6
6.6% [4.5–6.2] | -6
6.4% [4.5–6.2] | -6
6% [4.5–6.2] | -6
densitometry | -6
body mass composition | -6
bioimpedance method | -6
bone density test of the lumbar spine (L1–L4) | -6
Z-score [–] 2.2 | -6
rhGH therapy | 0
improvement of final height | 0
growth retardation | 0
weight gain | 0
insulin resistance | 0
osteoporosis | 0
severe growth failure | 0
glucocorticoids | 0
exaggerated growth retardation | 0
weight gain | 0
insulin resistance | 0
osteoporosis | 0
treatment with rhGH | 0
alleviate or worsen the course of muscular dystrophy | 0
anabolic effect of rhGH | 0
muscle mass and strength | 0
improvement of appetite | 0
increase in lean body (fat free) mass and bone mass | 0
improved mobility | 0
short statured boys | 0
higher strength-to-weight ratio | 0
slower progression of DMD | 0
better prognosis | 0
tall stature | 0
detrimental to muscle function | 0
muscle fibre damage | 0
scoliosis | 0
progression of DMD | 0
muscle strength | 0
muscle weakness | 0
IGF-1 concentrations | 0
elevated levels of IGFBP-3 | 0
lower muscle mass | 0
high content of fat tissue | 0
weight gain | 0
sedentary lifestyle | 0
consumed more food | 0
obesity | 0
harmful to functionality and motility | 0
natural course of muscular dystrophy | 0
progressive muscle weakness | 0
withdrawal from therapy | 0
behavioural therapy | 0
physical rehabilitation | 0
pharmacological treatment | 0
close monitoring of treatment and side effects | 0
immediate decision to withdraw from therapy | 0
alarming symptoms | 0
appropriate behavioural therapy | 0
physical rehabilitation | 0
assumed goal of pharmacological treatment | 0