61 years old | 0
female | 0
diabetes mellitus | -672
admitted to the hospital | 0
fever | 0
headache | 0
anorexia | 0
lethargy | 0
apathetic | 0
poor glycaemic control | 0
dehydration | 0
erythematous patch over the right maxillary bone | 0
tender | 0
neutrophil leukocytosis | 0
high CRP | 0
opacity in her right maxillary sinus | 0
bacterial sinusitis suspected | 0
IV ceftriaxone initiated | 0
blood sugar controlled with insulin | 0
urinary ketone bodies tested | 0
antral washout | 0
antral wash samples sent for bacterial and fungal culture | 0
deteriorated clinically | 0
admitted to the intensive care unit | 0
septic shock | 0
IV fluids and noradrenalin | 0
blood culture grew E. coli | 0
sinus washout culture grew E. coli | 0
antibiotic converted to IV Meropenum | 0
sinus washout fungal culture grew Rhizopus | 24
direct microscopy examination of the natal washout | 24
liposomal amphotericin B administered | 24
necrotic skin over the right maxillary bone | 24
ultrasound scan of the abdomen | 72
chest x-ray | 72
left-sided psoas abscess | 72
CECT of the abdomen | 72
psoas abscess aspirated under USS guidance | 72
samples sent for bacterial culture and AFB | 72
repeat USS of the psoas abscess | 120
recollection of the psoas abscess | 120
aspirated under USS guidance | 120
flexible rhinoscopy repeated | 120
necrotic debris removed | 120
dose of liposomal amphotericin B increased | 120
psoas abscess drained surgically | 168
conscious level deteriorated | 168
metabolic screening normal | 168
NCCT of the brain revealed pneumocephalus | 168
high-flow oxygen | 168
conscious level improved | 192
NCCT brain repeated | 192
pneumocephalus improved | 192
amphotericin B continued | 192
Meropenum continued | 192
flexible rhinoscopy done at the end of the treatment | 336
no necrotic material | 336
referred for facial reconstruction surgery | 336