10 years old | 0
male | 0
admitted to the hospital | -672
born | -8760
birth weight 2100 g | -8760
birth length 48 cm | -8760
prominent forehead | -8760
relative macrocephaly | -8760
limb asymmetry | -8760
5th finger clinodactyly | -8760
2/3 toe syndactyly | -8760
hypomethylation of the 11p15 region | -504
genetic examination | -504
diagnosis of SRS | -504
delayed motor development | -384
walked independently | -384
hepatic dysfunction | -420
increased concentration of alanine aminotransferase | -420
increased concentration of aspartate aminotransferase | -420
increased creatine kinase level | -420
diagnosis of Duchenne muscular dystrophy | -420
genetic test | -384
mutation of the maternal DMD gene | -384
corticosteroids treatment | -192
prednisone treatment | -192
deflazacort treatment | -96
G-CSF treatment | -96
sepsis | -96
hypoglycaemia | -96
neurological symptoms | -96
glucose level of 14 mg/dl | -96
urological care | -96
hypospadias | -96
cardiological diagnostics | -24
episodes of sinus tachycardia | -24
heart murmur | -24
propranolol treatment | -24
growth hormone deficiency | -24
rhGH treatment | 0
growth hormone therapy | 0
height velocity | 0
IGF-1 level | 0
IGFBP-3 level | 0
glucose and insulin levels | 0
HOMA-IR | 0
HbA1c | 0
impaired glucose tolerance | 12
insulin resistance | 12
abnormal gait | 12
weight gain | 12
reduced rhGH dose | 12
discontinuation of rhGH therapy | 18
body mass composition | 12
densitometry | 12
bone density test | 12
scoliosis | 0
BMD assessment | 12