79 years old | 0
female | 0
admitted to ICU | 0
surgical interposition graft | -720
thoracoabdominal aortic aneurysm | -720
hypertension | 0
chronic obstructive pulmonary disease | 0
chronic kidney disease | 0
transcatheter aortic valve implantation | 0
percutaneous coronary intervention | 0
vascular graft of abdominal aorta | 0
acute-on-chronic kidney failure | 0
continuous veno-venous haemofiltration | 0
persistent chylous leakage | 0
re-thoracotomy | 0
third-degree atrioventricular block | 0
pacemaker implanted | 0
surgical tracheostomy | 0
Staphylococcus aureus bacteraemia | -840
infected thoracotomy wound | -840
pleural fluid cultures positive | -840
flucloxacillin treatment started | -840
flucloxacillin 12 g/24 hours | -840
high flucloxacillin blood concentrations | -816
flucloxacillin dose decreased to 3 g/24 hours | -816
flucloxacillin dose changed to 6 g/24 hours | -798
acetaminophen 3 g per day | -840
appendicitis | -720
piperacillin-tazobactam treatment | -720
reduced consciousness | -504
controlled mechanical ventilation | -504
severe respiratory and high anion gap metabolic acidosis | -504
arterial blood gas analysis | -504
acetaminophen prescription stopped | -498
abdominal pain progression | -492
CT scan of abdomen | -492
intra-abdominal abscesses | -492
ICU treatment stopped | -486
patient died | -486
high anion gap metabolic acidosis due to 5-oxoproline accumulation confirmed | -486
urinary analysis | -486
5-oxoproline 1,721 μmol/mmol/creatinine | -486
creatinine 1.69 mmol/l | -486