91 years old | 0
female | 0
mild febrile sensation | -48
general weakness | -48
admitted to the emergency room | 0
hypertension | 0
beta blocker bevantolol | 0
dementia | 0
donepezil | 0
risperidone | 0
ambulate | 0
communicate without assistance | 0
limited ambulation | -336
short-leg splint | -336
undisplaced fractures of the 4th and 5th metatarsal bones of the right foot | -336
no injury with skin defects | 0
no trauma history | 0
no injection history | 0
watery diarrhea | -168
sputum production | -48
abdominal computed tomography scan | 0
fluid retention | 0
gas shadow in the right gluteal area | 0
gas shadow around the greater trochanter of the femur | 0
transferred to our hospital | 0
sepsis following soft tissue infection suspected | 0
systolic blood pressure 149/64 mmHg | 0
pulse rate 74 beats/minute | 0
respiratory rate 17 breaths/minute | 0
body temperature 36.5℃ | 0
physical examination revealed no evidence of skin necrosis | 0
no fluctuation | 0
mild level of heat around the hip and thigh | 0
BP dropped to 81/38 mmHg | 0
body temperature increased to 38.5℃ | 0
chilling sensation | 0
WBC count 14,300/mm3 | 0
neutrophils 95% | 0
erythrocyte sedimentation rate 41 mm/hour | 0
C-reactive protein level 17.46 mg/dL | 0
diagnosis of sepsis | 0
ceftriaxone | 0
clindamycin | 0
gas observed on the right gluteal area on plain radiographs | 0
increased signal intensity along the gluteus fascia to the greater trochanteric area on MRI | 0
abscess formation between the right gluteus maximus and medius | 0
smaller abscess on the left gluteus maximus | 0
air formation on both sides of the hips | 0
cystic shadows in the posterosuperior surface of the uterus | 0
bilateral necrotizing fasciitis confirmed | 0
incisions | 24
debridements | 24
surgery conducted on the right side | 24
posterolateral approach in the right lateral position | 24
no definite skin lesion around the thigh or hip | 24
bacterial cultures | 24
abscess discharged at the time of incision | 24
necrotic tissues observed along the gluteus medius and greater trochanter of the femur | 24
deep muscles invaded | 24
fascia invaded | 24
subcutaneous tissues invaded | 24
removed intraoperatively | 24
debridement | 24
lavage | 24
right hip joint puncture for culture tests | 24
drainage catheter inserted | 24
surgical site sutured | 24
referred to a gynecologist | 24
cystic lesions along the superior surface of the uterus | 24
transvaginal sonography | 24
lithotomy position | 24
puncture and aspiration performed | 24
aspirated fluid clear | 24
lesions non-inflammatory | 24
postoperative intensive care for two days | 24
SBP 132 mmHg | 24
body temperature 36.2℃ | 24
WBC count 9,400/mm3 | 24
neutrophil 95% | 24
ESR 16 mm/hour | 24
CRP level 3.77 mg/dL | 24
Escherichia coli detected | 24
ciprofloxacin | 24
drainage catheter removed | 168
suture removal | 336
ambulation limited | 336
pressure ulcer on the ischial areas | 336
general symptoms not identified | 336
high fever not identified | 336
CRP level elevated to 8.37 mg/dL | 336
body temperature 38.5℃ | 336
pressure ulcer infection | 336
follow-up MRI | 336
increase in the size of the abscess between the left greater trochanter and the gluteus medius | 336
incision | 336
debridement performed on the left aspect | 336
posterolateral incision | 336
no specific pus intraoperatively | 336
bacterial cultures on serosanguinous fluid | 336
drainage catheter inserted | 336
postoperative care in intensive care unit | 336
body temperature not exceeding 36.7℃ | 336
ischial pressure ulcer deterioration | 336
wound dressing | 336
ambulation using a wheelchair | 504
no infection-related complications | 4320
patient conditions improved | 4320
systematic rehabilitation | 4320
no bacteria detected in culture tests from the second operation | 336
body temperature increased to 38.5℃ |A prompt incisions and thorough debridements were performed on the following day. So incisions and debridement happened 24 hours after admission.
