60 years old | 0 | 0 
female | 0 | 0 
admitted to the hospital | 0 | 0 
impaired consciousness | -1 | 0 
atrial fibrillation | -672 | 0 
dilated cardiomyopathy | -672 | 0 
oral warfarin | -672 | 0 
biventricular pacing implantable cardioverter defibrillator | -672 | 0 
found lying at home | -1 | 0 
transported to hospital | -1 | 0 
Japan Coma Scale score was II-10 | 0 | 0 
Glasgow Coma Scale score was 14 | 0 | 0 
no clear neurological deficits | 0 | 0 
non-contrast head CT | 0 | 0 
hemorrhage in the third and fourth ventricles | 0 | 0 
hemorrhage in bilateral lateral ventricles | 0 | 0 
brain 3D-CTA | 0 | 0 
spot enhancement on the lateral wall of the anterior horn of the left lateral ventricle | 0 | 0 
blood pressure control | 0 | 24 
ventricular drainage not performed | 0 | 24 
cerebral angiograph | 72 | 72 
aneurysm at the distal site of the mLSA | 72 | 72 
embolization | 72 | 72 
endovascular treatment | 72 | 72 
N-butyl-2-cyanoacrylate injection | 72 | 72 
aneurysm embolization | 72 | 72 
postoperative head CT | 96 | 96 
no signs of hemorrhagic complications | 96 | 96 
no cerebral infarction | 96 | 96 
no impaired consciousness | 96 | 96 
no paralysis | 96 | 96 
sepsis triggered by pneumonia | 120 | 240 
decrease in muscle strength | 120 | 240 
disuse | 120 | 240 
rehabilitation | 240 | 432 
discharged to home | 432 | 432 
modified Rankin Scale of 1 | 432 | 432 
intraventricular aneurysm | 0 | 0 
distal medial lenticulostriate artery aneurysm | 0 | 0 
primary intraventricular hemorrhage | 0 | 0 
intraventricular hemorrhage | 0 | 0 
DRESS syndrome | 0 | 0 
fever | 0 | 0 
rash | 0 | 0 
acne | 0 | 0 
minocycline | 0 | 0 
increased WBC count | 0 | 0 
eosinophilia | 0 | 0 
systemic involvement | 0 | 0 
diffuse erythematous or maculopapular eruption | 0 | 0 
pruritus | 0 | 0 
DRESS syndrome diagnosis | 0 | 0 
fever persisted | 0 | 24 
rash persisted | 0 | 24 
discharged | 24 | 24 
Note: The events and timestamps are based on the provided case report. The timestamps are in hours, with 0 being the time of admission. Negative timestamps indicate events that occurred before admission, and positive timestamps indicate events that occurred after admission.