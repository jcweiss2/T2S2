85 years old | 0  
    male | 0  
    admitted to the hospital | 0  
    skin ulceration in the left upper limb | -24  
    lethargy | -24  
    fever | -24  
    stabbed in the left upper limb | -48  
    drowsiness | -48  
    fever (maximum body temperature of 38.8°C) | -48  
    skin in the left upper limb ulcerated | -48  
    redness | -48  
    swelling | -48  
    petechiae | -48  
    ecchymosis scattered on the skin of the whole body | -48  
    White blood cell count (WBC) 11.77 × 109/L | 0  
    procalcitonin (PCT) > 100 ng/mL | 0  
    lactate (Lac) 4.28 mmol/L | 0  
    cultures of blood | 0  
    cultures of secretions | 0  
    cultures of fluid seeping from the broken blisters on the skin in the left upper limb | 0  
    antibiotic sensitivity test | 0  
    metagenomic analysis of pathogens in blood sample using next-generation sequencing (NGS) | 0  
    treated with anti-infection (azithromycin and tienam) | 0  
    rehydration | 0  
    pressure promotion | 0  
    anticoagulation | 0  
    blood culture positive for Gram-negative bacilli | 24  
    admitted to emergency intensive care unit (EICU) | 24  
    septic shock | 24  
    history of diabetes for more than 20 years | -17520  
    long-term history of alcoholism | -17520  
    lethargic | 24  
    low spirit | 24  
    left hand and forearm with large areas of fluid exudation | 24  
    local tension blisters | 24  
    dark purple ecchymoses at the base | 24  
    slightly cool ends of the five fingers | 24  
    extensive swelling from the proximal end of the middle segment to the wrist | 24  
    scattered petechiae | 24  
    scattered ecchymosis | 24  
    treated with meropenem | 24  
    treated with levofloxacin | 24  
    norepinephrine | 24  
    vasopressin | 24  
    argatroban | 24  
    ulinastatin | 24  
    multiple incisions to decompress and drain the blisters on the skin in the left upper limb | 24  
    unbroken tension blisters disinfected with iodophor | 24  
    blister fluid aspirated with a syringe | 24  
    wound washed with 3% hydrogen peroxide | 24  
    gentamicin externally applied | 24  
    magnesium sulfate externally applied | 24  
    unstable blood pressure | 24  
    poor oxygenation | 24  
    tracheal intubation | 24  
    ventilator connection | 24  
    fever | 48  
    slight improvement of ulceration in the left limb | 48  
    slight improvement of oedema in the left limb | 48  
    skin on the back of the right hand swollen | 48  
    new petechiae | 48  
    new tension blisters | 48  
    dark purple skin on the neck with patchy ecchymosis | 48  
    PCT high | 48  
    high-sensitivity C-reactive protein (hCRP) levels high | 48  
    stab wound caused by a sea shrimp | -48  
    possibility of V. vulnificus infection considered | 48  
    treated with doxycycline | 48  
    blood culture identification positive for V. vulnificus | 72  
    antibiotic sensitivity test revealed positivity for V. vulnificus | 72  
    V. vulnificus identified as comma-like, flagellate, spore-free, facultative anaerobic bacterium | 72  
    colonies observed on culture medium | 72  
    metagenomic analysis of pathogens in blood sample using NGS indicated V. vulnificus | 72  
    alanine aminotransferase (ALT) level 2295 U/L | 96  
    aspartate aminotransferase (AST) level 1273 U/L | 96  
    liver enzyme levels normal on admission | 0  
    drug-induced liver damage considered | 96  
    doxycycline discontinued | 96  
    body temperature normal | 192  
    significantly alleviated skin ulceration in both upper limbs | 192  
    redness alleviated | 192  
    White blood cell count (WBC) 9.09 × 109/L | 192  
    PCT 2.68 ng/mL | 192  
    Lac 1.74 mmol/L | 192  
    ALT 281 U/L | 192  
    AST 44 U/L | 192  
    sedation stopped | 192  
    conscious | 192  
    passed spontaneous breathing trial (SBT) | 192  
    extubated | 192  
    noninvasive ventilator-assisted ventilation | 192  
    no fever | 408  
    vital signs stable | 408  
    swelling improved | 408  
    ulceration improved | 408  
    granulation tissues at the base of ulcers | 408  
    transferred to general ward | 408  
    history of diabetes | -17520  
    long-term history of alcoholism | -17520  
    stab wound by sea shrimp | -48  
    diabetic | -17520  
    alcohol addiction | -17520  
    immune function low | -17520  
    glucose metabolism disorder | -17520  
    lipid metabolism disorder | -17520  
    reduced protein synthesis | -17520  
    reduced globulin synthesis | -17520  
    decreased immune function | -17520  
    V. vulnificus invasion | -48  
    bacteremia | -48  
    sepsis | -48  
    septic shock | 24  
    MOF | 24  
    V. vulnificus sepsis | 72  
    skin cellulitis in the upper limbs | -48  
    rapid onset | -48  
    rapid progression | -48  
    surgical debridement | 24  
    decompression | 24  
    drainage | 24  
    hydrogen peroxide use | 24  
    gentamicin use | 24  
    magnesium sulfate use | 24  
    antibiotic resistance | 72  
    drug sensitivity test | 72  
    thorough debridement | 24  
    precise antimicrobial therapy | 72  
    improved prognosis | 408  

    