70 years old | 0
male | 0
admitted to the hospital | 0
COVID-19 diagnosis | -96
dyspnea | -96
tachypnea | -96
respiratory symptoms | -96
transferred to ICU | -48
intubation | 48
ventilator care | 48
extubation | 120
re-intubation | 144
tracheostomy planned | 168
preoperative chest X-ray | 170
surgical preparation | 170
thrombocytopenia | 170
platelet transfusion | 170
tracheostomy | 172
surgery | 172
application of PPE | 172
use of portable astral lamp | 172
injection of fentanyl | 172
transverse incision | 172
local injection of lidocaine | 172
repositioning of ET tube | 172
balloon overinflation | 172
attachment of transparent film dressing | 172
tracheostomy tube insertion | 172
ventilator connection | 172
removal of ET tube | 172
maintenance of oxygen saturation | 172
discharge | 105*24
medical staff healthy and asymptomatic | 14*24