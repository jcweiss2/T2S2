space-occupying lesion in the liver | -876 
transarterial embolization | -392 
sorafenib | -274 
dizziness | -182 
skin ulcers | -182 
CT scan | -56 
radiation therapy | -14 
Piggyback LT | 0 
acute renal failure | 0 
hematoma around the liver | 0 
intravenous administration of hepatitis B immunoglobulin | 0 
immunosuppressive drugs | 24 
steroids | 24 
tacrolimus | 24 
continuous hemodialysis | 24 
intermittent infusion of fresh frozen plasma | 24 
leukocyte-depleted red blood cells | 24 
other blood products | 24 
active bleeding in the abdominal cavity ceased | 48 
renal function gradually recovered | 48 
pathological analyses | 240 
HCC | 240 
massive tumor necrosis | 240 
liver function began to improve | 240 
fevers | 240 
procalcitonin levels began to rise | 240 
fever did not subside | 312 
obscure red spots | 312 
no symptoms such as itching | 312 
Nikolsky sign was negative | 312 
tacrolimus administration changed to sirolimus | 408 
mycophenolate mofetil | 408 
sputum culture suggested the presence of Acinetobacter baumannii | 432 
sputum culture suggested the presence of methicillin-resistant Staphylococcus aureus | 432 
rash advanced into erythematous macules and papules | 456 
rash spread to the limbs, palms, neck, and face | 456 
oral examination revealed white ulcers | 456 
severe bone marrow suppression | 456 
white blood cell count dropped | 456 
platelet count dropped | 456 
hemoglobin level dropped | 456 
patient was transferred to the intensive care unit | 456 
dermatologist hypothesized that the rash may be a drug-related adverse reaction | 456 
gamma globulin administration | 456 
skin biopsy | 456 
fluorescence in situ hybridization of the peripheral blood | 456 
abdominal incision split | 696 
abdominal incision sutured again | 696 
bone marrow aspiration | 768 
bone marrow pathology report | 768 
FISH analysis of the peripheral blood | 792 
donor lymphocytes detected | 792 
skin biopsy specimens exhibited epidermal dyskeratosis | 792 
basic vacuolization | 792 
lymphocytic infiltrates | 792 
grade-1 acute lt-GVHD | 792 
multidisciplinary team assembled | 816 
steroids | 816 
tacrolimus | 816 
granulocyte colony-stimulating factor | 816 
meropenem | 816 
voriconazole | 816 
rash was significantly reduced | 816 
patient’s general condition continued to deteriorate | 816 
serum ferritin levels increased | 816 
esophageal and oral ulcers continued to worsen | 816 
patient’s temperature rose | 1128 
hallucinations | 1128 
destruction of the patient’s skin | 1128 
bone marrow | 1128 
mucosal epithelium | 1128 
immunodeficiency | 1128 
multiple infections | 1128 
septic shock | 1320 
multiple organ dysfunction syndrome | 1320 
death | 1320