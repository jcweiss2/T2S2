37 years old | 0
female | 0
OTCD | -25200
seizures | -25200
valproic acid | -25200
hyperammonemia | -25200
liver biopsy | -25200
liver OTC enzyme activity 30% | -25200
hemodialysis | -6840
hemodialysis | -5040
self-restricted protein diet | -25200
L-carnitine treatment | -25200
pregnancy | -280
delivery | 0
male baby | 0
blood ammonia 68 μmol/L | 0
blood ammonia 59 μmol/L | 10
blood ammonia 54 μmol/L | 24
hyperammonemia 194 μmol/L | 96
discharge | 144
consumed hamburger | 144
consumed beef | 144
hospitalized | 168
hyperammonemia 180 μmol/L | 168
impaired consciousness | 168
arginine treatment | 168
blood ammonia 82 μmol/L | 168
hemodialysis | 168
continuous hemodiafiltration | 168
respirator management | 168
high-calorie infusion | 168
arginine | 168
citrulline | 168
sodium benzoate | 168
sodium phenylbutyrate | 168
hyperammonemia improved | 192
extubation | 192
reintubation | 192
sepsis | 192
intensive care unit | 192
maternal milk production | 672
hyperammonemia persisted | 672
brain magnetic resonance imaging | 3024
single-photon emission computed tomography | 3024
atrophy of bilateral frontal and temporal lobes | 3024
decreased blood flow | 3024
discharge | 1008
liver transplantation | -25200
caesarean section | -280
maternal milk production halted | -280
sodium benzoate or sodium phenylbutyrate therapy | -280
blood glutamine levels | -280
liver transplantation | 0