47 years old | 0
male | 0
158 kg | 0
173 cm | 0
diabetes mellitus | -672
hypertension | -672
obstructive sleep apnea | -672
BiPAP ventilation | -672
admitted to intensive care unit | 0
laparoscopic sleeve gastrectomy | -24
anastomotic leak | 0
computed tomography–guided aspiration of abdominal collections | 0
closing gastric fistula and transverse colon | 0
washing abdomen with repeated peritoneal lavage | 0
peritonitis | 0
sepsis | 0
acute kidney injury | 0
sputum cultures positive for coagulase-negative Staphylococcus aureus | 0
vancomycin 1500 mg intravenously twice daily | 0
tigecycline | 0
meropenem | 0
red-man syndrome | -72
peak and trough samples drawn | 144
peak plasma concentration 32.4 mg/L | 144
trough plasma concentration 24.8 mg/L | 144
calculating true elimination rate constant K | 144
calculating true volume of distribution V | 144
recommended dosing interval 36 h | 144
recommended dose 2500 mg | 144
new dose regimen 1500 mg q24 | 168
predicted peak plasma concentration 19 mg/L | 168
actual peak level 22.7 mg/L | 168
trough level 12.5 mg/L | 168
elevated serum creatinine 187 micromole/L | 0
normal baseline serum creatinine 87 micromole/L | -672
discharged | 240