56 years old | 0
    male | 0
    fever | 0
    difficulty breathing | 0
    diabetes | 0
    hypertension | 0
    hyperlipidaemia | 0
    tested positive for COVID-19 | 0
    admitted to the intensive care unit | 0
    intubated | 0
    respiratory deterioration | 0
    ventilation for six weeks | -4032
    brief period of clinical improvement | 0
    developed persistent temperature spikes | 0
    developed fatigue symptoms | 0
    blood culture isolated coagulase-negative Staphylococcus | 0
    echocardiogram showed a 1.4 x 1.5 cm mitral valve vegetation | 0
    received meropenem | 0
    received levofloxacin | 0
    received teicoplanin | 0
    antibiotic combinations for three months | -2592
    no resolution of fever | 0
    no resolution of mitral valve vegetation | 0
    referred to the current centre | 0
    right leg pain | 0
    calf swelling | 0
    pulse of 90 bpm | 0
    blood pressure of 122/77 mmHg | 0
    respiratory rate of 20 breaths/minute | 0
    temperature of 38.5 oC | 0
    pansystolic murmur over the mitral valve area | 0
    bilateral coarse inspiratory crepitations | 0
    right calf swollen | 0
    unable to move ankle due to pain and weakness | 0
    left leg pulses normal | 0
    right foot pulses impalpable | 0
    elevated white blood cell count of 13 x 109/L | 0
    C reactive protein of 341 mg/L | 0
    haemoglobin level of 7.1 g/dL | 0
    antibiotic therapy changed to vancomycin and ceftriaxone | 0
    pre-operative full body computed tomography angiography | 0
    showed right 7 x 7.5 cm tibioperoneal trunk aneurysm | 0
    transoesophageal echocardiogram showed posterior mitral valve leaflet vegetation | 0
    vegetation measured 1.7 x 1.6 cm | 0
    moderate eccentric mitral regurgitation | 0
    no improvement with prolonged antibiotic therapy | 0
    decision for open surgical repair | 0
    underwent lung and cardiac assessment | 0
    considered fit for surgery | 0
    combined one stage operation | 0
    cardiac surgery through median sternotomy | 0
    heparin given | 0
    activated clotting time >400 seconds | 0
    placed on heart-lung machine | 0
    extended vertical transatrial-septal approach | 0
    large amount of vegetation on posterior leaflet | 0
    mitral valve replacement with bioprosthesis | 0
    heparin reversed with protamine | 0
    peripheral aneurysm repaired | 0
    harvest of right saphenous vein | 0
    exposure of distal superficial femoral artery | 0
    posterior tibial artery exposed | 0
    proximal control obtained at distal SFA | 0
    aneurysm approached through medial incision | 0
    aneurysm opened | 0
    organised thrombus without pus observed | 0
    evacuated thrombus | 0
    aneurysm ligated | 0
    distal popliteal artery ligated | 0
    vascular reconstruction with reversed saphenous vein graft | 0
    end to side proximal anastomosis to distal SFA | 0
    vein graft tunnelled anatomically to midcalf | 0
    anastomosed end to side to PTA | 0
    good distal flow along PTA | 0
    no microorganisms recovered from mitral vegetations | 0
    no microorganisms recovered from aneurysm thrombus | 0
    placed on 75 mg aspirin | 0
    placed on 10 mg atorvastatin | 0
    cardiac surgery stage took 3 hours 31 minutes | 0
    vascular surgery took 3 hours 30 minutes | 0
    total blood loss 300 mL | 0
    extubated on post-operative day two | 72
    discharged from ICU on day seven | 168
    discharged from hospital on day 31 | 744
    echocardiography showed normal functioning mitral valve at five months | 3600
    six months follow up free of symptoms | 4320
    palpable right PTA pulse at ankle | 4320
    advised to remain on 75 mg aspirin once daily | 4320
    