18 years old | 0
male | 0
HBV-associated PAN | -720
weight loss | -720
myalgias | -720
fever | -720
skin erythema | -720
deterioration of renal function | -720
new onset of diabetes | -720
hypertension | -720
diagnosed with PAN | -720
diagnosed with HBV | -720
prednisolone | -720
cyclophosphamide | -720
Tenofovir | -720
acute abdomen | 0
septic shock | 0
peritonitis | 0
free sub diaphragmatic air | 0
laparotomy | 0
perforations of the small intestine | 0
segmental enterectomy with anastomosis | 0
mechanical ventilation | 0
circulatory support | 0
acute-on-chronic renal failure | 0
weaned off the ventilator | 24
haemodynamically stable | 24
treatment with tenofovir | 24
IV methylprednisolone | 24
enteric content | 168
second explorative laparotomy | 168
new perforations | 168
patchy necrosis | 168
plasma exchanges | 168
IV cyclophosphamide | 168
IV methylprednisolone | 168
open abdomen | 168
vacuum device | 168
re-laparotomy | 216
third laparotomy | 216
necrotic lesions | 216
IV prednisone | 216
fourth laparotomy | 432
segmental enterectomy with anastomosis | 432
cholecystectomy | 432
gangrenous gallbladder | 432
died | 720