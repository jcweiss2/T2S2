28 years old | 0
female | 0
Japanese | 0
admitted to the hospital | 0
fever | 0
abdominal pain | 0
confusion | 0
blood pressure of 80/50 mm Hg | 0
heart rate of 120 beats/min | 0
respiratory rate of 32 breaths/min | 0
body temperature of 38.3 °C | 0
abdominal tenderness | 0
rebound tenderness | 0
abdominal rigidity | 0
cervical motion tenderness | 0
cervical bleeding | 0
grayish-white and foul-smelling cervical fluids | 0
arterial blood gas pH of 7.35 | 0
HCO3 level of 15.5 mmol/L | 0
lactate level of 6.9 mmol/L | 0
white blood cell count of 0.9 × 10^9/L | 0
C-reactive protein level of 33.98 mg/dL | 0
hepatoportal venous gas | 0
pneumatosis intestinalis | 0
mesenteric emphysema | 0
free air | 0
ascites | 0
small intestinal wall thickening | 0
emergency laparotomy | 0
opaque ascites | 0
inflammatory redness and edema of the uterus and fallopian tubes | 0
adhesion of the right fallopian tube | 0
abdominal cavity washed with physiological saline | 0
abdomen closed | 0
gram-negative cocci | 0
short rods | 0
septic shock | 0
pelvic peritonitis | 0
minocycline | 0
ceftriaxone | 0
metronidazole | 0
negative nucleic acid amplification test for Neisseria gonorrhoeae | 0
negative nucleic acid amplification test for Chlamydia trachomatis | 0
negative nucleic acid amplification test for HIV | 0
Fusobacterium necrophorum in blood culture | 0
Fusobacterium necrophorum in ascites culture | 0
Gardnerella vaginalis in ascites culture | 0
Gardnerella vaginalis in vaginal fluid culture | 0
Mobiluncus species in vaginal fluid culture | 0
resolution of hepatoportal venous gas | 72
resolution of pneumatosis intestinalis | 72
left the ICU | 288
postcoital bleeding | -504
dyspareunia | -504
cloudy and odorous vaginal fluid | -504
multiple sexual partners | -504
receptive oral sex | -504
no intrauterine device | -504
no condom | -504
no upper respiratory symptoms | -504
no antibiotics | -504
bacterial vaginosis | -504