81 years old | 0
    woman | 0
    admitted to the hospital | 0
    fatigue | -72
    lethargy | -72
    fever | -72
    chills | -72
    phlegm | -72
    wheezing | -72
    coma | 0
    oxygen saturation dropped to 70%-80% | 0
    admitted to the intensive care units | 0
    progressive drop in blood pressure | 0
    norepinephrine | 0
    chronic obstructive pulmonary disease | -131328
    bronchial asthma | -131328
    long-term home oxygen therapy | -131328
    chronic heart insufficiency | -131328
    bisoprolol | -131328
    no history of abdominal pain | 0
    no history of chronic renal failure | 0
    no smoking history | 0
    no alcohol consumption | 0
    body temperature 36 °C | 0
    pulse 85 beats/min | 0
    respiratory rate 18 breaths/min | 0
    blood pressure 105/45 mmHg | 0
    decreased breath sounds in both lungs | 0
    wet rales at the bottom of both lungs | 0
    unremarkable cardiac examination | 0
    unremarkable abdominal examination | 0
    troponin level increased from 0.05 ng/mL to 3.92 ng/mL | 0
    B-type natriuretic peptide 4164 pg/mL | 0
    carbon dioxide partial pressure 58.7 mmHg | 0
    oxygen partial pressure 86.5 mmHg | 0
    oxygenation index 172.97 mmHg | 0
    white blood cell 8.12 × 109/L | 0
    neutrophil percentage 93.2% | 0
    C-reactive protein 298.38 mg/L | 0
    procalcitonin 6.26 ng/mL | 0
    interleukin-6 > 5000 pg/mL | 0
    negative PCR-SARS-CoV-2 test | 0
    negative multiple blood cultures | 0
    normal fecal examinations | 0
    normal coagulation function | 0
    sinus rhythm | 0
    T wave high and sharp | 0
    R wave V1-V4 progression poor | 0
    V1 Qr type | 0
    ST-segment elevation (> 0.05 mv) | 0
    left atrial enlargement | 0
    segmental abnormal motion of the left ventricular wall | 0
    left ventricular apical bulge | 0
    decreased left ventricular diastolic function | 0
    LVEF 51% | 0
    chronic bronchitis | 0
    emphysema | 0
    multiple infections in both lungs | 0
    right pleural cavity small effusion | 0
    aortic arch calcification | 0
    coronary artery calcification | 0
    abdominal aorta calcification | 0
    assisted ventilation | 0
    vasoactive drugs | 0
    milrinone | 0
    amiodarone | 0
    anti-infection treatment | 0
    PCI via left femoral artery approach | 24
    no significant abnormalities in left and right coronary arteries | 24
    abdominal distension | 48
    decreased bowel sounds (1-2/min) | 48
    glycerin enema | 48
    sudden loss of consciousness | 96
    blood pressure dropped | 96
    abdominal wall swelling | 96
    increased abdominal wall tension | 96
    bowel sounds disappeared | 96
    extensive pneumatosis intestinalis | 96
    hepatic portal system gas | 96
    intestinal wall necrosis | 96
    mesenteric artery involvement | 96
    AMI | 96
    septic shock | 96
    refractory shock | 120
    death | 120

<|eot_id|>
