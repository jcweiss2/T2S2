43 years old | 0
female | 0
Chron’s disease | 0
infliximab | 0
azathioprine | 0
admitted to the hospital | 0
fever | -72
thoracic pain | -72
elevated inflammatory parameters | -72
nasopharyngeal swab for SARS-CoV-2 negative | -72
bilateral community-acquired pneumonia (CAP) | -72
cefuroxime | -72
returned to the hospital | -48
Streptococcus pneumoniae urinary antigen test negative | -48
Legionella pneumophila urinary antigen test negative | -48
nasopharyngeal swab for SARS-COV-2 negative | -48
piperacillin-tazobactam | -48
admitted to the hospital | -48
acute rapidly progressive respiratory failure | -24
invasive mechanical ventilation | -24
admitted to the intensive care unit (ICU) | -24
vancomycin | -24
methylprednisolone | -24
mixed acidaemia | -12
refractory hypoxemia | -12
extracorporeal membrane oxygenation (ECMO) | -12
transferred to Infectious Diseases ICU | 0
meropenem | 0
liposomal amphotericin | 0
cardiovascular failure | 12
hypoperfusion | 12
hypotension | 12
anasarca | 12
hyperlacticaemia | 12
anuric acute kidney injury | 12
liver failure | 12
worsening pancytopenia | 12
multiple blood transfusions | 12
vasopressor therapy | 12
continuous renal replacement therapy | 12
sodium bicarbonate supplementation | 12
albumin supplementation | 12
plasmapheresis | 12
Saprochaete clavata in blood culture | 24
identified as Saprochaete clavata by MALDI-TOF technology | 48
died | 120
Legionella pneumophila in bronchoalveolar lavage | 120