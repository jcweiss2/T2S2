right-sided abdominal pain | -48
vomiting | -48
fever | -48
presentation to emergency department | 0
conscious | 0
alert | 0
oriented | 0
pale | 0
sick | 0
temperature of 37.8°C | 0
blood pressure of 150/90 mmHg | 0
oxygen saturation of 95% on room air | 0
abdomen distended | 0
tympanic | 0
right upper quadrant tenderness | 0
right flank tenderness | 0
total leukocyte count was 20 × 10^3 | 0
hemoglobin 10.7 gm% | 0
acidotic with pH 7.33 | 0
laboratory evidence of end-stage renal disease | 0
chest X-ray demonstrated air under the right hemi-diaphragm | 0
evaluated by the general surgeon | 0
impression of perforated viscous | 0
computed tomography (CT) scan with contrast | 0
right perinephric collection with extension into the right sub-phrenic region | 0
gas in the right collecting system and urinary bladder | 0
no gas in the renal parenchyma | 0
incidental finding of the right atrial thrombus | 0
started on parenteral antibiotics | 0
admitted to intensive care unit | 0
trial of percutaneous drainage | 12
percutaneous drainage failed | 12
evaluated by the anesthetist | 12
not fit for general anesthesia | 12
open drainage of a very thick, foul smelly, loculated perinephric and sub-phrenic collection | 24
cystoscopy | 24
abnormal bladder mucosa with multiple cystic lesions with air “bubbles” all over the bladder | 24
ureteric Double J stent inserted in the right ureter | 24
urethral catheter to drain the bladder | 24
reasonably well during the procedure | 24
condition started to deteriorate | 48
culture of the collection showed Klebsiella pneumonia extended-spectrum β-lactamase | 48
condition continued to deteriorate | 72
died | 72
severe sepsis | 72
multiple organ failure | 72
history of diabetes mellitus | -1000
history of end-stage renal disease | -1000
history of peripheral vascular disease | -1000
left below knee amputation | -1000
right above knee amputation | -1000
right extra anatomical axillobifemoral bypass graft | -1000
known case of adult polycystic kidney disease | -1000 
no shortness of breath | 0
denies chest pain | 0