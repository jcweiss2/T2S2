35 years old | 0
female | 0
admitted to the hospital | 0
dyspnea | -72
loss of consciousness | -72
hyaluronic acid injection | -72
confused mental state | 0
petechial rash | 0
body temperature 36.8 | 0
blood pressure 150/110 mm Hg | 0
pulse rate 127/min | 0
respiratory rate 28/min | 0
crackles in both lower lung fields | 0
liver function test normal | 0
renal function test normal | 0
white blood cells 21,080/µL | 0
hemoglobin 11 g/dL | 0
platelets 240,000/µL | 0
troponin I 0.16 ng/mL | 0
CK-MB 0.6 ng/mL | 0
C-reactive protein 5.307 mg/dL | 0
D-dimer 1.278 µg/mL | 0
N-terminal of the prohormone brain natriuretic peptide 9,177 pg/mL | 0
arterial blood gas analysis | 0
pH 7.505 | 0
PCO2 28.6 mm Hg | 0
PO2 66.1 mm Hg | 0
HCO3- 22.4 mmol/L | 0
plain chest radiography showed ground glass opacity and consolidation | 0
contrast-enhanced chest CT showed diffuse ground glass opacity | 0
mechanical ventilation | 0
hemorrhagic eruptions | 72
antibiotics | 0
corticosteroids | 0
diuretics | 0
hypoxemia improved | 120
blood culture showed no growth | 120
discontinued antibiotics | 120
weaned from mechanical ventilation | 120
discharged | 192
follow-up chest CT showed improvement | 720
no fibrosis | 720