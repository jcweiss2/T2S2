66 years old | 0
male | 0
Billroth II gastrectomy | -8400
peptic ulcer disease | -8400
open cholecystectomy | -240
diffuse abdominal pain | 0
vomiting | 0
diarrhea | 0
nonsteroidal anti-inflammatory drugs | -72
colchicine | -72
gout crisis | -72
diffuse articular pain | -72
mild tenderness to deep palpation | 0
enlarged prostate | 0
leukocytosis | 0
INR of 2.5 | 0
C-reactive protein of 48 mg/l | 0
pH of 7.21 | 0
base excess of 13.6 mEq/l | 0
pCO2 of 33 mmHg | 0
no acute abdominal disease | 0
plain abdominal X-ray | 0
simple left renal cyst | 0
dilatation and edema of the jejunal loops | 0
minimal quantity of free fluid in the peritoneal space | 0
possible localized peritonitis | 0
respiratory failure | 2
intubation | 2
mechanical ventilation | 2
severely hypotensive | 2
oliguric | 2
inotropic support | 2
macroscopic hematuria | 2
emergency explorative laparotomy | 2
no anastomotic leak | 4
no source of abdominal sepsis | 4
multiorgan failure | 16
death | 16
colchicine overdose | 16
autopsy not performed | 16