54 years old | 0
male | 0
obese | 0
Caucasian | 0
admitted to hospital | 0
fever | -120
rigors | -120
persistent cough | -120
myalgia | -120
shortness of breath | -120
no chest pain | -120
no palpitation | -120
no hemoptysis | -120
non-smoker | 0
does not drink alcohol | 0
no history of liver disease | 0
no co-morbidities | 0
temperature of 39.5 °C | 0
low O2 saturation at 88% | 0
blood pressure of 140/82 mm Hg | 0
heart rate of 95/min | 0
respiratory rate of 22/min | 0
bibasilar crackles | 0
no pleural rub | 0
no pericardial rub | 0
no deep vein thrombosis | 0
lymphopenia | 0
high CRP | 0
high ferritin | 0
elevated LDH | 0
normal clotting | 0
normal liver function | 0
normal renal function | 0
atypical pneumonia screen negative | 0
blood cultures negative | 0
type 1 respiratory failure | 0
bilateral patchy consolidation on CXR | 0
diagnosed with COVID-19 pneumonia | 0
O2 therapy | 0
intravenous antibiotics | 0
dexamethasone | 0
remdesivir | 0
high-flow O2 | 24
tocilizumab | 24
good recovery | 120
discharged home | 120
readmitted | 336
generally unwell | 336
extreme fatigue | 336
poor appetite | 336
reduced oral intake | 336
high temperature | 336
heart rate of 132/min | 336
hypotensive | 336
tachypnea | 336
Glasgow Coma Scale of 14/15 | 336
icterus positive | 336
peripherally cyanosed | 336
flapping tremors | 336
encephalopathic | 336
distended tender abdomen | 336
severe type 1 respiratory failure | 336
severe metabolic acidosis | 336
severe acute kidney injury | 336
hyperkalemia | 336
high creatinine | 336
low GFR | 336
acute hepatic injury | 336
high ALT | 336
high AST | 336
high bilirubin | 336
high amylase | 336
high ALP | 336
high GGT | 336
low albumin | 336
undetectable paracetamol | 336
coagulopathy | 336
high INR | 336
high aPTT | 336
high D-dimer | 336
thrombocytopenia | 336
high CRP | 336
extremely high ferritin | 336
admitted to ICU | 336
central venous catheter inserted | 336
high-flow oxygen | 336
potential for intubation and ventilation | 336
intravenous piperacillin/tazobactam | 336
intravenous fluids | 336
human albumin serum | 336
fresh frozen plasma | 336
dexamethasone | 336
proton pump inhibitors | 336
bicarbonate | 336
CXR done | 336
CT of abdomen and pelvis done | 336
discussed with hepatology and liver transplant unit | 336
best supportive care | 336
GCS dropped | 339
hypotensive | 339
intubated and ventilated | 339
cardiac arrest | 339
died | 339