24 years old | 0
female | 0
pregnant | 0
admitted to the hospital | 0
abdominal pain | -120
abdominal distension | -120
constipation | -120
increasing severity of pain | -120
no significant past medical history | 0
no significant past surgical history | 0
uneventful menstrual history | 0
uneventful antenatal history | 0
dehydrated | 0
hypotension | 0
tachycardia | 0
tachypnea | 0
asymmetrically distended abdomen | 0
tenderness all over abdomen | 0
empty rectum on digital examination | 0
vaginal examination not suggestive of threatened preterm labour | 0
elevated white cell count | 0
clear urine analysis | 0
distended bowel loop on ultrasound | 0
moderate amount of free fluid in peritoneal cavity | 0
single viable fetus | 0
clinical diagnosis of intestinal obstruction | 0
abdominal X-ray | 0
dilated large bowel on X-ray | 0
abnormal gas pattern on X-ray | 0
coffee bean appearance on X-ray | 0
sigmoidoscopy | 0
twisted sigmoid colon | 0
failure to negotiate obstruction | 0
foetal distress | 0
deceleration in heart rate | 0
concomitant caesarean section | 0
premature fetus | 0
male preterm infant | 0
weight 750g | 0
mechanical ventilation | 0
lung immaturity | 0
enormously distended sigmoid loop | 0
ischemic and gangrenous changes | 0
no signs of perforation | 0
necrotic colon | 0
posteriorly displaced by pregnant uterus | 0
lower segment caesarean section | 0
delivery of preterm infant | 0
admitted to neonatal ICU | 0
resection of sigmoid colon | 0
Hartmann’s procedure | 0
end colostomy | 0
closure of rectal stump | 0
post-operative course uneventful | 0
discharged home on 9th post-operative day | 216
child discharged home after 10 weeks in neonatal ICU | 720
reversal of Hartmann’s | 4320
bowel continuity restored through colo-rectal anastomosis | 4320