27 years old | 0
female | 0
fell from a bicycle | -2
landed on the handlebar | -2
pancreatic contusion | -2
trauma CT scan | -2
referred to a level 1 trauma center | -2
grade III lesion of the pancreas | -2
rupture of the pancreatic neck | -2
retroperitoneal hematoma | -2
admitted to the hospital | 0
nasogastric tube | 0
intravenous proton pump inhibitor | 0
subcutaneous octreotide | 0
intravenous cefuroxime | 0
metronidazole | 0
parenteral nutrition | 0
ERCP | 72
papillotomy of the pancreatic duct | 72
diastasis of the duct ends | 72
large hematoma | 72
displacement of the fractured parts | 72
attempt to insert a bridge prosthesis | 72
abdominal pain | 96
inflammatory parameters | 96
free intraperitoneal fluid | 96
ultrasonography | 96
laparotomy | 96
removal of 2000 ml ascites | 96
external 18 Fr tubes | 96
abdomen closed | 96
general condition improved | 120
no need for pain killers | 120
systemic inflammatory response decreased | 120
started eating regular food | 120
one abdominal tube discontinued | 120
decreasing amount of fluid | 120
stable level of liquid | 120
amylase of 10,000 U/l | 120
discharged | 384
followed up at the outpatient clinic | 384
intermittent retraction of the drain | 384
fistula to the skin formed | 672
drain removed | 672
discharge ceased from the fistula | 784
increasing discomfort | 784
abdominal pain | 784
CT scan | 784
pseudocyst | 784
MRCP | 784
MR angiography | 784
severed pancreatic duct | 784
arterial perfusion | 784
endoscopic ultrasonography | 784
HOT AXIOSTM stent | 784
insertion of the stent | 784
collection punctured | 784
distal flange deployed | 784
proximal flange deployed | 784
patient could eat normally | 808
abdominal pain ceased | 808
discharged | 808
CT scan | 952
collapsed cyst | 952
stent removed | 1008
CT scan | 1056
no recurrence of the cyst | 1056
pancreatic duct measured 6 mm | 1056
blood supply | 1056
patient doing well | 1056
no signs of malabsorption | 1056
no diabetes | 1056
follow-ups terminated | 1056