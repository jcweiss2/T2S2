42 years old | 0
male | 0
chronic alcohol abuse | 0
cocaine abuse | 0
admitted to the medical floors for altered mental status secondary to alcohol intoxication with impending withdrawal | 0
elevated heart rate (115 bpm) | 0
elevated blood pressure (168/111 mmHg) | 0
hypoxia (O2 saturation 70% on room air) | 0
agitation | 0
altered mental status | 0
expiratory wheezes | 0
white blood cell count 14,500/μL | 0
Hb 15.2 g/dL | 0
platelet count 380,000/μl | 0
elevated serum creatinine (1.27 mg/dL) | 0
urine drug screen positive for cocaine | 0
blood alcohol level elevated (34) | 0
normal CT scan of the head | 0
chest X-ray showing possible right small pleural effusion | 0
CT pulmonary angiogram showing moderate hiatal hernia | 0
moderate distention of the esophagus | 0
mild debris in the left main stem bronchus concerning aspiration | 0
patchy subsegmental bibasilar opacities | 0
mild nonspecific ground-glass opacities | 0
started on CIWA protocol for alcohol withdrawal | 0
started on antibiotics (Piperacillin-Tazobactam) for aspiration pneumonia | 0
oxygen supplementation with nasal cannula | 0
COVID-19 test negative | 0
episode of coffee ground vomitus | 0
started on IV Protonix | 0
consultation with gastroenterology department | 0
no further active bleeding | 0
hemoglobin value within normal range | 0
worsening mental status on the 2nd day | 48
transferred to the intensive care unit for worsening delirium tremens and respiratory distress | 48
increasingly hypoxic | 48
decreased breath sounds on the right side of the chest | 48
repeat CXR showing large right-sided pleural effusion | 48
thoracic surgery consultation obtained | 48
insertion of right inferior chest thoracostomy tube | 48
draining 2 L of dark fluid | 48
pleural fluid analysis suggestive of exudative effusion (WBC 82831, Polys 92%, fluid glucose <10, LDH 1459, protein 2.1, PH 6) | 48
fluid cultures positive for Candida Albicans | 48
infectious diseases consultation | 48
antibiotics switched to meropenem and vancomycin | 48
addition of antifungal agent micafungin | 48
transferred to the medical floor | 72
worsening agitation | 96
readmitted to the ICU | 96
treated with lorazepam infusion | 96
persistently febrile (T max 101.7 °F) | 96
leukocytosis (WBC count up to 24,000) | 96
repeat CT scan of the chest showing multiple right-sided loculated pleural effusions with air-fluid levels | 96
blood cultures no growth | 96
thoracic surgery consultation indicating patient was a poor surgical candidate | 96
insertion of two chest tubes by interventional radiology department | 96
superiorly inserted chest tube draining 300 mL of pus | 96
inferior chest tube draining 50 mL of purulent fluid and air | 96
pleural fluid cultures showing candida and staphylococcus epidermidis growths in superior chest tube | 96
candida in inferior chest tube | 96
antibiotic regimen changed to meropenem, vancomycin, and fluconazole | 96
3rd chest tube placed inferiorly following repeat CT chest | 144
increased effusion size in basilar portion of the right lung | 144
two upper chest tubes removed later | 168
meropenem switched to ampicillin-sulbactam | 168
mental status improved after about 15 days of hospitalization | 360
oral feeding started | 360
repeat CT chest demonstrating empyema on the right side with slight decrease in size | 360
moderate left pleural effusion | 360
food contents coming out from the chest tube | 360
chest tube output high at 1.5–2 L per day | 360
contrast esophagogram demonstrating leak from the right side of the distal esophagus | 504
discussion with gastroenterology and thoracic surgery departments | 504
feeding tube placement with esophageal stent insertion | 504
percutaneous endoscopic gastrostomy (PEG) | 672
endoscopic findings confirming esophageal defect | 672
endoscopic esophageal stent placement | 672
vancomycin stopped | 672
switched to ampicillin-sulbactam | 672
completed additional month of fluconazole treatment after discharge | 1344
diagnosed with esophagopleural fistula | 672
candida empyema | 672
esophageal perforation | 672
esophageal stent placement | 672
discharge | 1344
