61 years old | 0
female | 0
hypertension | 0
chronic cough | 0
dyspnea | 0
50-pound weight loss | 0
nausea | -504
vomiting | -504
cachexia | 0
scleral icterus | 0
jaundice | 0
dry mucous membranes | 0
decreased breath sounds in the left lower lung fields | 0
tachycardia | 0
hypotension | 0
hyponatremia | 0
sodium level of 131 mEq/L | 0
bicarbonate level of 32 mEq/L | 0
elevated alkaline phosphatase level of 215 u/L | 0
total bilirubin level of 5.8 mg/dL | 0
aspartate aminotransferase level of 58 u/L | 0
alanine aminotransferase level of 36 u/L | 0
innumerable pulmonary parenchymal nodules throughout both lungs | 0
large mass extending into the lingula | 0
large mass extending into the superior segment of the left lower lobe | 0
pleural effusion | 0
severely dilated common bile duct | 0
moderately distended gall bladder | 0
large heterogeneous mass in the pancreatic head | 0
grossly dilated common bile duct | 0
enlarged retroperitoneal lymph nodes | 0
lung mass biopsy | 0
emergent biliary stenting via endoscopic retrograde cholangiopancreatography | 0
high nuclear pleomorphism | 0
prominent nuclei | 0
immunohistological staining positive for thyroid transcription factor−1 (TTF-1) | 0
cytokeratin-7 (CK-7) staining | 0
absence of tumor protein 63 (p63) expression | 0
metastases to the brain | 0
radiation therapy | 0
adjunctive chemotherapy | 0
metastases to the pancreas | 0
metastases to the retroperitoneum | 0
severe pneumonia | 0
sepsis | 0
female |[![Build Status](https://travis-ci.org/microsoft/vstest.svg?branch=master)](https://travis-ci.org/microsoft/vstest)
