39 years old | 0  
    Thai | 0  
    man | 0  
    street vendor | 0  
    lives in Bangkok | 0  
    presented to the emergency department | 0  
    fever | -120  
    myalgia | -120  
    breathlessness | -6  
    haemoptysis | -6  
    no medical history | 0  
    20-pack-year smoking | 0  
    high body temperature | 0  
    39.8°C | 0  
    tachypnea | 0  
    respiratory distress | 0  
    no conjunctival suffusion | 0  
    no icteric sclera | 0  
    chest radiography bilateral diffuse opacification pattern | 0  
    arterial blood gas pH 7.42 | 0  
    pCO2 35.7 mm Hg | 0  
    pO2 55 mm Hg | 0  
    SpO2 89% | 0  
    lactate 1.2 | 0  
    FiO2 1.0 | 0  
    haemoglobin 108 g/L | 0  
    mean corpuscular volume 93 fL | 0  
    platelet 117,000 | 0  
    white blood cell count 10,250 | 0  
    neutrophil 89.9% | 0  
    lymphocyte 5.4% | 0  
    monocyte 4.4% | 0  
    eosinophil 0% | 0  
    basophil 0.3% | 0  
    prothrombin time 13.7 | 0  
    INR 1.23 | 0  
    aPTT 29.3 | 0  
    total bilirubin 1.51 mg/dL | 0  
    alanine aminotransferase 48 U/L | 0  
    creatinine 0.93 mg/dL | 0  
    albumin 3.4 g/dL | 0  
    urinalysis mild proteinuria | 0  
    microscopic haematuria | 0  
    Thai-Lepto score 8.5 | 0  
    intubation | 0  
    fresh blood suctioned | 0  
    admitted to intensive care unit | 0  
    APACHE II score 17 | 0  
    respiratory distress | 0  
    oxygen desaturation | 0  
    diffuse alveolar haemorrhage | 0  
    severe ARDS | 0  
    ventilator support | 0  
    lung-protective strategy | 0  
    sedation cisatracurium | 0  
    propofol | 0  
    midazolam | 0  
    fentanyl | 0  
    ceftriaxone | 0  
    levofloxacin | 0  
    plasmapheresis | 2  
    IVMP 250 mg | 2  
    ANCA negative | 0  
    anti-MPO negative | 0  
    anti-PR3 negative | 0  
    anti-GBM negative | 0  
    severe hypoxaemia | 12  
    hypercapnia | 12  
    mechanical ventilator PCV mode | 12  
    VV$ECMO started | 12  
    leptospirosis diagnosis confirmed | 24  
    anti-Leptospira IgM negative | 24  
    anti-Leptospira IgM positive | 192  
    transthoracic echocardiography normal | 0  
    LVEF 60% | 0  
    haemoculture negative | 0  
    sputum culture negative | 0  
    sputum acid-fast bacilli negative | 0  
    modified acid-fast bacilli negative | 0  
    anti-HIV negative | 0  
    anti-HCV negative | 0  
    HBsAg negative | 0  
    anti-HBs negative | 0  
    anti-HBc negative | 0  
    Weil-Felix test negative | 0  
    OX 19 titre negative | 0  
    OX K titre negative | 0  
    OX 2 titre negative | 0  
    scrub typhus Ab negative | 0  
    murine typhus Ab negative | 0  
    dengue NS1 antigen negative | 0  
    dengue IgM negative | 0  
    dengue IgG positive | 0  
    influenza A/B/RSV rapid test negative | 0  
    RT-PCR negative | 0  
    respiratory virus 19 subtypes negative | 0  
    thin blood film negative | 0  
    thick blood film negative | 0  
    ANA negative | 0  
    CH50 44.9 U/mL | 0  
    C3 138 mg/dL | 0  
    C4 53.4 mg/dL | 0  
    renal function slightly impaired | 96  
    renal function returned to normal | 96  
    liver function test normal | 0  
    condition improved | 120  
    weaned off VV$ECMO | 120  
    withdrawal of VV$ECMO | 192  
    endotracheal tube removed | 240  
    discharged from intensive care unit | 240  
    stable condition | 240  
    good consciousness | 240  
    no dyspnoea | 240  
    discharged home | 336  
    recovered | 336  
    healthy after 1 year | 8760  
<|eot_id|>
    