71 years old | 0
female | 0
admitted to the hospital | 0
unconscious state | 0
history of hypertension | 0
history of ischaemic heart disease | 0
history of peripheral vascular disease | 0
stroke | 0
head computed tomographic scan | 0
inotropic support | 24
septic shock | 24
elevated levels of inflammatory markers | 24
erythrocyte sedimentation rate | 24
C-reactive protein | 24
blood culture | 24
yeast in blood culture | 24
caspofungin treatment | 24
died | 72
Lodderomyces elongisporus | 48
identification by VITEK 2 yeast identification system | 48
identification by PCR sequencing of ITS region of rDNA | 48
turquoise blue colonies on CHROMagar Candida | 48
long ellipsoidal-shaped ascospores | 48
antifungal susceptibility testing | 48
amphotericin B | 48
fluconazole | 48
voriconazole | 48
posaconazole | 48
itraconazole | 48
flucytosine | 48
caspofungin | 48
micafungin | 48
hospitalization for lower limb ischaemia | -336
discharge from hospital | -336
fungaemia | 24
primary fungaemia | 24
Lodderomyces elongisporus fungaemia | 24
catheter tip culture | 24
caspofungin treatment | 24
death | 72
treatment outcome | 72
antifungal therapy | 72
echinocandins | 72
caspofungin | 72
micafungin | 72
antifungal susceptibility | 48
in vitro MIC values | 48
Infectious Disease Society of America guidelines | 72
therapeutic use of echinocandins | 72
treatment of candidaemia | 72
Candida parapsilosis | 48
Candida parapsilosis complex | 48
Candida orthopsilosis | 48
Candida metapsilosis | 48
matrix-assisted laser desorption/ionization time-of-flight mass spectrometry | 48
rare yeast species | 72
reduced susceptibility to antifungal agents | 72
prolonged survival of seriously ill patients | 72
administration of multiple broad-spectrum antibiotics | 72
dependence on life support systems | 72
extended use of intravascular catheters | 72
prophylactic and therapeutic use of antifungal agents | 72
selection pressure | 72
increased colonization and invasive infection | 72
delay in accurate identification | 72
lack of experience in management of rare yeast infections | 72
diagnostic and therapeutic challenges | 72
higher mortality rates | 72