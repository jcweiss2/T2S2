49 years old | 0
    female | 0
    generalized weakness | -720
    abdominal pain | 0
    back pain | 0
    onset of weakness 1 month prior | -720
    abdominal fullness for a year | -8760
    marked splenomegaly | 0
    hemoglobin 9 | 0
    platelet count 40 | 0
    WBC count 45 | 0
    17% blasts | 0
    bone marrow core biopsy 100% cellular | 0
    marked myeloid predominance | 0
    30% to 40% blasts | 0
    chromosome analysis identified 2 related abnormal clones | 0
    complex 4-way rearrangement between chromosomes 1, 11, 9, and 22 | 0
    BCR:ABL rearrangement | 0
    deletion in chromosome 14 | 0
    translocation between chromosomes 7 and 12 | 0
    FISH confirmed BCR-ABL1 gene rearrangement 62% | 0
    next-generation sequencing negative for multiple genes | 0
    bone marrow biopsy and cytogenetic studies suggested de novo BCR-ABL positive AML or CML-BC | 0
    diagnosis of CML-BC | 0
    treated with induction chemotherapy (cytarabine plus daunorubicin) | 0
    started on dasatinib 140 mg twice daily | 0
    follow-up bone marrow biopsy confirmed complete morphologic remission | 24
    chromosomal analysis showed normal female karyotype | 24
    FISH negative for BCR-ABL translocation | 24
    referred for allogeneic hematopoietic stem cell transplant | 24
    underwent matched related donor SCT | 24
    received myeloablative conditioning with fludarabine and busulfan | 24
    stable course until day +81 | 1944
    new leukocytosis | 1944
    increased blast count | 1944
    hemoglobin 11.7 | 0
    platelet count 20 | 0
    WBC 39 | 0
    10% peripheral blasts | 0
    PT 18 | 0
    INR 1.6 | 0
    aPTT 26 | 0
    fibrinogen 456 | 0
    negative soluble fibrin monomers | 0
    fever 38.4°C | 24
    hypotension | 24
    sepsis | 24
    blood cultures showed no growth | 24
    CT scan of abdomen and pelvis showed colitis | 24
    stool testing positive for Clostridioides difficile | 24
    peripheral blast count increased from 10% to 41% | 96
    bone marrow aspirate and core biopsy on day 3 | 72
    100% cellular marrow | 72
    absent erythroids | 72
    absent megakaryocytes | 72
    85% to 90% blasts | 72
    relapse of CML-BC | 72
    FISH analysis confirmed BCR-ABL1 fusion 54% | 72
    worsening coagulopathy | 0
    worsening anemia | 0
    worsening thrombocytopenia | 0
    hemoglobin 6.4 | 0
    hematocrit 19.2 | 0
    platelet count 9 | 0
    INR increased to 4.1 | 48
    peripheral blast count increased | 48
    PT 52.7 seconds | 48
    factor deficiency or weak inhibitor | 48
    FVII activity 3% | 48
    Factor II 55% | 48
    Factor X 57% | 48
    Factor V 77% | 48
    oral vitamin K 5 mg administered | 48
    no improvement in INR | 48
    no improvement in factor levels | 48
    decreased level of responsiveness | 48
    transfer to ICU | 48
    CT scan of head ruled out intracranial hemorrhage | 48
    no further evidence of bleeding | 48
    started on chemotherapy (cladribine, cytarabine, venetoclax) | 120
    clinical improvement | 120
    transferred back to hematology ward | 168
    regained consciousness | 168
    vision loss | 168
    dilated fundus exam showed severe bilateral retinal hemorrhages | 168
    coagulopathy improved | 168
    peripheral blast count declined | 168
    FVII activity improved to 63% | 336
    improvement of blurry vision | 336
    hospital discharge | 336
    two months later | 1488
    bone marrow aspirate and biopsy showed persistent disease 70% blasts | 1488
    FVII activity 14% | 1488
    INR 2.2 | 1488
    started on decitabine and venetoclax | 1488
    FVII level 15% 10 days later | 1536
    no bleeding | 1536
    achieved remission after 1 cycle | 1488
    not candidate for second SCT | 1488

<|eot_id|>