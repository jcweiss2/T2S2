6 years old | 0
male | 0
admitted to the hospital | 0
seizure | -24
hypertensive encephalopathy | -24
posterior reversible encephalopathy syndrome | -24
abdominal mass | -24
adrenal mass | -24
pheochromocytoma | -24
nifedipine | -24
labetalol | -24
dexamethasone | -24
weight gain | -720
moon face | 0
central obesity | 0
Buffalo hump | 0
abdominal striae | 0
hirsutism | 0
hypertension | 0
elevated blood pressure | 0
tachycardia | 0
abdominal pain | 48
hematuria | 48
anuria | 48
bilateral ureteral stones | 48
acute kidney injury | 48
fever | 48
elevated C-reactive protein | 48
broad-spectrum antibiotics | 48
etomidate | 48
hydrocortisone | 72
ureteral stent indwelling | 72
continuous renal replacement therapy | 48
discontinuation of losartan | 96
discontinuation of minoxidil | 96
discontinuation of nicardipine | 96
improvement of oliguria | 96
improvement of renal function | 96
discontinuation of CRRT | 96
adrenal mass resection | 120
histologically confirmed adrenocortical adenoma | 120
ureteral stones removal | 120
calcium carbonate apatite | 120
discharge | 168
replacement therapy of hydrocortisone | 168