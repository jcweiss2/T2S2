63 years old | 0
male | 0
achalasia | -6720
dyspepsia | -6720
admitted to the hospital | 0
severe right chest pain | 0
epigastric pain | 0
chest retrosternal pain | 0
respiratory distress | 0
tachycardic | 0
normal arterial pressure | 0
no fever | 0
diminished breath sounds | 0
pain and tenderness of epigastric | 0
O2 saturation 88% | 0
pneumomediastinum | 0
pleural effusion | 0
collapsed right lobe of the lung | 0
esophageal rupture | 0
Candida albicans in the pleural space | 0
intubated | 24
antibiotics | 24
chest physical therapy | 24
adequate intravenous fluids | 24
nasogastric tube feeding | 24
elevated WBC count | 72
elevated BUN | 72
elevated potassium | 72
tachyarrhythmia | 72
multiple organ failures | 96
hemodialysis | 96
thoracotomy | 96
debridement | 96
drainage of the mediastinum and pleural space | 96
6-cm longitudinal rupture in the upper esophagus | 96
noradrenaline and vasopressin support | 96
T-tube implanted | 96
sutures to anchor fistula | 96
two chest tubes inserted | 96
ventilator support | 96
broad-spectrum IV piperacillin/tazobactam antibiotic therapy | 96
two stents placed in the esophagus | 120
oral liquid feeding started | 120
discharged from the ICU | 936
discharged from the hospital | 944
tracheostomy | 960
good condition at 2-month follow-up | 1488