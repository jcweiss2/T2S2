55 years old | 0
man | 0
admitted to the hospital | 0
pulled into a cement mixer | -60
right lower limb completely torn off | -60
conscious | -60
drowsy | -60
patent airway | -60
injury severity score of 75 | -60
blood pressure 70 to 85/40 to 50 mmHg | -60
pulse 120 beats per minute | -60
bandaging applied with strong mechanical pressure | -60
intravenous rehydration treatment | -60
oxygen inhalation | -60
open wound over the right costal arch | 0
perineum extension | 0
ending near the right sacroiliac joint | 0
entire area stripped of skin | 0
peritoneum holding in abdominal contents | 0
cement and other foreign matters covering the wound | 0
displaced extremity cold | 0
extensively crushed | 0
pulseless | 0
fluid resuscitation through central venous line | 0
fluid resuscitation through peripheral lines | 0
tetanus prophylaxis | 0
broad-spectrum antibiotics | 0
computed tomography (CT) imaging | 0
loss of the right lower limb | 0
loss of the right lower abdominal wall | 0
no intra-abdominal injury | 0
bladder intact | 0
rectum intact | 0
CT angiography | 0
transection of the right common iliac vessels | 0
general anesthesia | 0
systemic exploration of the pelvic wound | 0
gross loss of skin from the right lower abdomen | 0
severely contaminated peritoneum | 0
bowel peristalsis observed | 0
right scrotum avulsed | 0
exposed testis | 0
spermatic cord extravasation | 0
missing soft tissue around anus | 0
missing soft tissue around right ilium | 0
exposed sacrum | 0
arterial bleeding in the pelvic cavity | 0
right external iliac vessels transected | 0
right internal iliac vessels transected | 0
thrombosed vessels | 0
ligation of main vessels | 0
sutured to stop pelvic hemorrhage | 0
wound washed with saline | 0
wound washed with hydrogen peroxide | 0
wound washed with iodophor diluent | 0
extensive skin loss | 0
wound left open | 0
vacuum-sealing drainage (VSD) device | 0
rectal tube for bowel integrity | 0
packed red blood cells (800 mL) | 0
crystalloids (1000 mL) | 0
colloids (1500 mL) | 0
transferred to ICU | 0
mechanical ventilation support | 0
blood transfusion (600 mL) | 0
aggressive fluid resuscitation | 0
preventive broad-spectrum antibiotics | 0
imipenem (0.5 g, q6h) | 0
metronidazole (1 g, q8h) | 0
antifungal medication | 0
linezolid (0.6 g, q12h) | 0
fever persisted in ICU | 24
white blood cell count peak of 16.95 × 10^9/L | 120
closed drainage | 120
pneumothorax in the right lung | 120
pneumonia in the left lung | 120
no localized pelvic abscess | 120
second operation for debridement | 144
granulation tissue observed | 144
devitalized tissue removed | 144
pus samples collected for culture | 144
repetitive irrigation | 144
repetitive debridement | 144
VSD therapy continued | 144
presence of Proteus mirabilis | 144
presence of Providencia alcalifaciens | 144
blood sample showing Pseudomonas aeruginosa | 216
antibiotic regimen changed | 216
meropenem (1 g, q8h) | 216
levofloxacin (0.5 g, qd) | 216
tigecycline (0.1 g, q12h) | 216
fluconazole (0.4 g, qd) | 216
diverting colostomy | 336
body temperature remained high | 336
temperature fluctuations | 336
body temperature dropping to baseline | 600
skin defect of 28 × 21 cm² | 504
psychiatric management | 504
nutritional management | 504
chronic pain management | 504
skin regeneration | 2016
skin defect decreased 50% | 2016
VSD therapy discontinued | 2016
split-skin graft from left thigh | 2016
able to walk with crutches | 1680
squatting maneuvers performed | 1680
semi-laparotomy prosthesis | 5280
healed wound | 8760
phantom pain | 8760
prescribed pain medicine | 8760
no symptoms of depression | 8760
