35 years old | 0
female | 0
newly diagnosed diabetes | -672
persistent generalized headache | -168
non-productive cough | -96
sore throat | -96
altered mental status | 0
lethargic | 0
confused | 0
unresponsive | 0
random rhythmic movements of bilateral upper and lower extremities | 0
no tongue biting | 0
no fecal or urinary incontinence | 0
taking food to a COVID-19 positive family member | -336
no close contact | -336
no history of substance use | 0
no smoking | 0
no recent travel | 0
Glasgow Coma Scale of 9 | 0
afebrile | 0
temperature 36.6 | 0
heart rate 93 | 0
blood pressure 133/70 | 0
no nuchal rigidity | 0
Brudzinski and Kernig’s signs were negative | 0
agitation | 0
vomiting | 0
endotracheal intubation | 0
white blood cell count of 6900/μL | 0
lactate of 1.1 mmol/L | 0
head CT without contrast showed no abnormalities | 0
urinalysis was negative | 0
chest x-ray showed bilateral patchy infiltrates | 0
nasopharyngeal SARS-CoV-2 PCR resulted positive | 0
pharyngeal swab for rapid Streptococcus test was positive for Streptococcus pyogenes | 0
blood cultures were drawn | 0
vancomycin | 0
ceftriaxone | 0
acyclovir | 0
admitted to the intensive care unit | 0
fluoroscopy-guided lumbar puncture | 48
cerebrospinal fluid analysis showed glucose of 109 mg/dL | 48
cerebrospinal fluid analysis showed protein of 250 mg/dL | 48
cerebrospinal fluid analysis showed RBC of 231/mm3 | 48
cerebrospinal fluid analysis showed WBC of 42/mm3 | 48
infectious workup of the CSF resulted negative | 48
elevated C-reactive protein | 0
elevated erythrocyte sedimentation rate | 0
elevated D-dimer | 0
normal ferritin | 0
normal lactate dehydrogenase | 0
normal interleukin-6 levels | 0
blood and CSF cultures finalized negative | 120
vancomycin was discontinued | 48
ceftriaxone was continued | 48
acyclovir was continued | 48
mental status markedly improved | 96
extubated | 96
discharged home | 216
PO penicillin V | 216
PO valacyclovir | 216