30 years old | 0
female | 0
pregnancy | 0
G1P0 | 0
27 weeks of gestation | 0
admitted to the emergency department | 0
progressive dyspnea | -120
lethargy | -120
fever | -120
bacterial pneumonia | 0
Amoxicillin | 0
Clavulanate | 0
Clarithromycin | 0
Oseltamivir | 0
consolidation in the base of the left hemithorax | 0
no auscultatory findings | 0
hospitalization | 0
worsening dyspnea | 4
increased demand of supplemental oxygen | 4
transferred to ICU | 4
continuous non-invasive ventilation (NIV) | 4
full-face mask (10 L/min O2) | 4
unsatisfactory clinical response | 7
unsatisfactory laboratorial response | 7
elective endotracheal intubation | 7
severe hypoxemia | 16
PaO2/FiO2 <80 | 16
ARDS | 16
neuromuscular blockade | 16
alveolar recruitment | 16
no adequate response | 16
semi-pronation position (900) to the left | 16
new alveolar recruitment | 16
no satisfactory improvement in oxygenation | 16
veno&shy;venous ECMO installation | 24
cannulation of the right internal jugular vein | 24
cannulation of the right femoral vein | 24
preserved cardiac function | 24
decision not to interrupt the gestation | 24
fetus viability monitoring | 24
daily cardiac rhythm evaluation | 24
bedside ultrasound | 24
betamethasone administration | 24
increased white blood cell count | 96
new culture samples obtained | 96
Piperacillin-Tazobactam | 96
Oseltamivir continued | 96
Amoxicillin and Clavulanate resistant Enterobacter | 96
important impairment of lung function | 168
Methylprednisolone (2mg/kg) | 168
mechanical ventilation | 168
ECMO cessation | 264
extubation | 312
intermittent NIV requirement | 312
ICU discharge | 360
discharge after 21 days of hospitalization | 504
current pregnancy (30 weeks) | 504
normodramnia | 504
fetal biometry compatible with gestational age | 504
antenatal evaluation | 504
Caesarean section at 38 weeks of gestation | 504
delivery of a healthy male infant | 504
H1N1 infection | -120
ARDS secondary to H1N1 infection | 16
refractory hypoxemia | 24
ECMO use | 24
ECMO circuit-related complications | 24
systemic anticoagulation | 24
heparin use | 24
corticosteroid administration | 168
lung-protective mechanical ventilation | 24
no fetal distress | 24
delayed antiviral therapy institution | 0
antiviral therapy with Oseltamivir | 0
increased risk factors (pregnancy) | 0
physiological and anatomical changes during pregnancy | 0
respiratory signs and symptoms | 0
masking the adequate diagnosis | 0
delaying the treatment | 0
increased risk of severe influenza-associated complications | 0
need for mechanical ventilation | 16
severe pneumonia | 16
refractory hypoxemia resistant to conventional ventilation | 24
improved lung function | 264
significant improvement in lung function | 264
lung recruitment maneuvers | 16
prone positioning | 16
inhaled nitric oxide | 16
high-frequency oscillatory ventilation | 16
ECMO as salvage therapy | 24
successful use of ECMO | 24
ECMO feasibility during pregnancy | 24
hemorrhagic complications | 24
fetal survival rate | 504
maternal survival rate | 504
increased ICU admission rate for ARDS | 0
mortality rate for ARDS | 0
fetal loss rate | 0
preterm deliveries | 0
neonatal ICU admission rate | 0
cesarean section | 504
neonatal morbidity | 504
neonatal mortality | 504
safety of Oseltamivir during pregnancy | 0
no competing interests | 0
no specific funding | 0
30 years old|0
female|0
pregnancy|0
G1P0|0
27 weeks of gestation|0
admitted to the emergency department|0
progressive dyspnea|-120
lethargy|-120
fever|-120
bacterial pneumonia|0
Amoxicillin|0
Clavulanate|0
Clarithromycin|0
Oseltamivir|0
consolidation in the base of the left hemithorax|0
no auscultatory findings|0
hospitalization|0
worsening dyspnea|4
increased demand of supplemental oxygen|4
transferred to ICU|4
continuous non-invasive ventilation (NIV)|4
full-face mask (10 L/min O2)|4
unsatisfactory clinical response|7
unsatisfactory laboratorial response|7
elective endotracheal intubation|7
severe hypoxemia|16
PaO2/FiO2 <80|16
ARDS|16
neuromuscular blockade|16
alveolar recruitment|16
no adequate response|16
semi-pronation position (900) to the left|16
new alveolar recruitment|16
no satisfactory improvement in oxygenation|16
veno-venous ECMO installation|24
cannulation of the right internal jugular vein|24
cannulation of the right femoral vein|24
preserved cardiac function|24
decision not to interrupt the gestation|24
fetus viability monitoring|24
daily cardiac rhythm evaluation|24
bedside ultrasound|24
betamethasone administration|24
increased white blood cell count|96
new culture samples obtained|96
Piperacillin-Tazobactam|96
Oseltamivir continued|96
Amoxicillin and Clavulanate resistant Enterobacter|96
important impairment of lung function|168
Methylprednisolone (2mg/kg)|168
mechanical ventilation|168
ECMO cessation|264
extubation|312
intermittent NIV requirement|312
ICU discharge|360
discharge after 21 days of hospitalization|504
current pregnancy (30 weeks)|504
normodramnia|504
fetal biometry compatible with gestational age|504
antenatal evaluation|504
Caesarean section at 38 weeks of gestation|504
delivery of a healthy male infant|504
H1N1 infection|-120
ARDS secondary to H1N1 infection|16
refractory hypoxemia|24
ECMO use|24
ECMO circuit-related complications|24
systemic anticoagulation|24
heparin use|24
corticosteroid administration|168
lung-protective mechanical ventilation|24
no fetal distress|24
delayed antiviral therapy institution|0
antiviral therapy with Oseltamivir|0
increased risk factors (pregnancy)|0
physiological and anatomical changes during pregnancy|0
respiratory signs and symptoms|0
masking the adequate diagnosis|0
delaying the treatment|0
increased risk of severe influenza-associated complications|0
need for mechanical ventilation|16
severe pneumonia|16
refractory hypoxemia resistant to conventional ventilation|24
improved lung function|264
significant improvement in lung function|264
lung recruitment maneuvers|16
prone positioning|16
inhaled nitric oxide|16
high-frequency oscillatory ventilation|16
ECMO as salvage therapy|24
successful use of ECMO|24
ECMO feasibility during pregnancy|24
hemorrhagic complications|24
fetal survival rate|504
maternal survival rate|504
increased ICU admission rate for ARDS|0
mortality rate for ARDS|0
fetal loss rate|0
preterm deliveries|0
neonatal ICU admission rate|0
cesarean section|504
neonatal morbidity|504
neonatal mortality|504
safety of Oseltamivir during pregnancy|0
no competing interests|0
no specific funding|0
