76 years old | 0
    male | 0
    admitted to the hospital | 0
    diabetes | 0
    hypertension | 0
    post-coronary artery bypass graft surgery | 0
    magnetic resonance imaging-compatible ICD implantation | -26280
    secondary prevention of ventricular tachycardia | -26280
    low left ventricular ejection fraction of 30% | -26280
    computerized tomography coronary angiography | -4392
    atypical chest pain | -4392
    patent grafts | -4392
    metoprolol XL | 0
    telmisartan | 0
    spironolactone | 0
    multiple ICD shocks | -6
    fever | -120
    myalgia | -120
    tested positive for SARS-CoV-2 infection | -120
    clinical examination unremarkable | 0
    stable vital signs | 0
    oxygen saturation of 97% on room air | 0
    electrocardiogram: normal sinus rhythm | 0
    electrocardiogram: no ST-T changes | 0
    electrocardiogram: QTc interval of 464 milliseconds | 0
    echocardiogram: global hypokinesia | 0
    echocardiogram: left ventricular ejection fraction of 30% | 0
    serum potassium within normal limits | 0
    serum magnesium within normal limits | 0
    elevated C-reactive protein | 0
    elevated ferritin | 0
    elevated creatine kinase | 0
    elevated troponin T | 0
    elevated NT-proBNP | 0
    ICD interrogation: multiple episodes of monomorphic ventricular tachycardias | 0
    ICD interrogation: ventricular ectopic | 0
    tachycardia persisted despite anti-tachycardia pacing | 0
    terminated by 38 shocks of 35 J each | 0
    amiodarone infusion | 0
    increased metoprolol doses | 0
    VT storm controlled | 24
    symptomatic treatment for COVID-19 infection | 0
    recovered in 10 days | 240
    discharged | 240
    amiodarone | 240
    metoprolol XL | 240
    telmisartan | 240
    torsemide-spironolactone | 240
    aspirin | 240
    statins | 240
    oral hypoglycemics | 240
    no episodes of VT at 3-month follow-up | 2184
    asymptomatic at 3-month follow-up | 2184