67 years old | 0
male | 0
multiple cerebrovascular events | 0
myocardial infarction | 0
hypertension | 0
30 pack-year smoking history | 0
dull 5/10 sacral pain | 0
pelvic magnetic resonance imaging (MRI) examination | 0
large, well circumscribed, heterogeneously enhancing mass through the mid body of the sacrum | 0
core biopsy | 0
sacral chordoma | 0
preoperative external beam radiation | -72
sacrectomy | -72
abdominoperineal resection | -72
colostomy exteriorized through the left rectus abdominus muscle | -72
pelvic defect | -72
perineal defect | -72
reconstructed using a right VRAM flap | -72
postoperative admission to the intensive care unit | 0
transferred to the orthopedic surgery unit | 120
regular flap checks | 120
flap consistently well perfused | 120
postoperative day 13 | 312
fever | 312
tachycardia | 312
significant abdominal discomfort | 312
increase in white blood cell count | 312
septic workup initiated | 312
flap demonstrated signs of venous insufficiency | 312
flap demonstrated signs of arterial insufficiency | 312
computed tomography of the pelvis | 312
markedly distended bladder | 312
bilateral hydronephrosis | 312
deep inferior epigastric pedicle visualized | 312
pedicle occluded by the distended bladder | 312
bladder decompressed | 312
improvement in clinical status | 312
perfusion to the flap did not improve | 312
total flap loss | 312
debridement of the VRAM flap | 504
significant thrombosis of the deep inferior epigastric pedicle | 504
necrotic flap | 504
bilateral advancement flaps elevated for closure | 504
discharged from hospital | 960
wound completely healed | 1440
