34 years old| 0
    African-American woman| 0
    gravida 3| 0
    para 1| 0
    presented with left uterine mass| 0
    menorrhagia| -8760
    pelvic pain| -8760
    newly developed left uterine mass| 0
    multiple small myomas| 0
    diagnostic laparoscopy| 0
    possible myomectomy| 0
    laparotomy with left oophorectomy| -8760
    ovarian cysts| -8760
    elective terminations of pregnancy| -8760
    inflammatory process| -8760
    asthma| 0
    use of nonsteroidal anti-inflammatory drugs| 0
    bradycardia| 0
    small thyroid nodule| 0
    mild iron deficiency anemia| 0
    hemoglobin 11.6 g/dL| 0
    hematocrit 35.3%| 0
    inconclusive thyroid studies| 0
    clinically euthyroid| 0
    open entry method| 0
    adherent small bowel loops| 0
    careful dissection| 0
    establishment of pneumoperitoneum at 15 mm Hg| 0
    extensive adhesions| 0
    careful port placement| 0
    adhesiolysis using disposable scissors| 0
    uterus adherent to sigmoid colon| 0
    uterine bulges consistent with myoma or adenomyoma| 0
    myolysis| 0
    serial bipolar needle punctures| 0
    abdomen lavaged with saline| 0
    generous amount of saline left to minimize adhesion reformation| 0
    operative time 75 minutes| 0
    anesthetic inhalation agents: sevoflurane and nitrous oxide| 0
    estimated blood loss <30 mL| 0
    discharged on same day of surgery| 0
    postoperative recovery uneventful for first 3 days| 0
    afebrile| 0
    voiding well| 0
    tolerating oral intake| 0
    passed flatus on second day| 48
    small bowel movement on third day| 72
    bloody drainage from incision attributed to hydroflation| 24
    black and blue mark around umbilicus| 48
    abdominal pain| 0
    abdominal distention| 0
    vomited| 96
    presented to emergency room| 96
    acute abdomen diagnosed| 96
    sudden onset of atrial fibrillation| 96
    hypotension| 96
    triple lumen catheter placed| 96
    exploratory laparotomy| 96
    enteric fluid exit from umbilical port site| 96
    midline laparotomy performed| 96
    gross spillage of enteric fluid| 96
    extremely dense adhesions between bowel and anterior abdominal wall| 96
    extensive mobilization of small bowel| 96
    perforated bowel seeping fluid| 96
    incidental enterotomy during adhesiolysis| 96
    affected bowel resected| 96
    Prasad double barrel ileostomy done| 96
    foreshortening of mesentery| 96
    3-cm defect in resected bowel| 96
    ischemic necrosis| 96
    bowel mucosa slightly edematous| 96
    transferred to ICU| 96
    treated with broad-spectrum antibiotics| 96
    activated protein C (Xigris)| 96
    2-month ICU course| 1680
    candidemia| 1680
    unsuccessful extubation trials| 1680
    profound multiple neuropathy| 1680
    nosocomial pneumonia| 1680
    pressure ulcer| 1680
    drug-induced thrombocytopenia| 1680
    gastrointestinal bleeding| 1680
    shock| 1680
    2 cardiopulmonary arrests| 1680
    gastrostomy tube placed| 1680
    tracheostomy tube placed| 1680
    inferior vena cava filter placed| 1680
    deep-vein thrombosis| 1680
    currently in rehabilitation| 4320