45 years old | 0
male | 0
admitted to the emergency department | 0
cough | -216
sore throat | -216
oxygen saturation of 88% on room air | 0
heart rate of 104 beats per minute | 0
blood pressure of 105/75 mmHg | 0
temperature 38.5 °C | 0
SARS-CoV-2 infection | -216
COVID-19 pneumonia | -216
BMI of 22.7 kg/m2 | 0
no significant medical history | 0
no known drug allergies | 0
no history of smoking or drinking alcohol | 0
no regular medications | 0
antiviral treatment with favipiravir | 0
dexamethasone | 0
LMWH with 1 × 40 mg enoxaparin | 0
3/L oxygen support | 0
d-dimer level of 660 μg/L | 0
oxygen support gradually decreased | 0
antiviral treatment completed | 0
discharged with LMWH | 168
left upper quadrant and left flank pain | 168
physical examination normal | 168
mild tenderness without peritonitis findings | 168
leukocytosis of 17.2 × 10∧3/μL | 168
D-dimer of 310 μg/L | 168
troponin of 0.001 | 168
abdominal CT showed noncontrast hypodense area | 168
thorax CT showed subpleural dominant irregular ground-glass opacities | 168
oral intake stopped | 168
intravenous hydration started | 168
nonopioid analgesics started | 168
anticoagulant treatment increased to 2 × 0,6 mL | 168
sudden onset chest pain | 192
ST segment elevation in the limb leads | 192
acute inferior MI | 192
emergency coronary angiography | 192
stent placed in the RCA | 192
transferred to the general surgery clinic | 216
regressive abdominal pain | 216
oral intake increased | 216
abdominal findings regressed | 216
discharged with 100 mg acetylsalicylic acid and ticagrelor | 240
genetic hypercoagulant tests negative | 720
control abdominal ultrasonography normal | 720
no intra-abdominal fluid or abscess collection | 720
meningococcal and Haemophilus influenza vaccines not necessary | 720
follow-up imaging not indicated | 720