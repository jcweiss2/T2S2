45 years old | 0
male | 0
high-speed motor vehicle accident | -6120
BTAI with near aortic transection | -6120
exploratory laparotomy | -6120
splenectomy | -6120
repair of a bladder injury | -6120
TEVAR with Gore TAG Endoprosthesis | -6120
thrombosis of the left subclavian artery | -3600
stent graft at the origin of the left subclavian artery | -3600
lost to follow-up | -1092
evaluated at an outside hospital for fever, chills, and malaise | -192
completed an outpatient course of antibiotics for pneumonia | -192
presented again with prolonged fevers and chills | -128
Streptococcus viridans and Mycoplasma bacteremia | -128
treated with an inpatient course of parenteral antibiotics | -128
intermittent fevers | -128
30-pound weight loss | -128
presented to our institution with high fevers and sepsis | 0
Staphylococcus capitis bacteremia | 0
admitted to the intensive care unit | 0
tranthoracic echocardiography | 0
freely mobile pedunculated vegetations within the thoracic aortic endograft | 0
computed tomography angiography of the chest | 0
right lower lobe consolidation with collapse and bilateral pleural effusions | 0
open surgical explantation of the aortic endograft and left subclavian artery stent graft | 24
aortic débridement | 24
inline reconstruction with a rifampin antibiotic-soaked prefabricated Dacron graft | 24
wedge resection of the portion of involved lung | 24
hypothermic circulatory arrest | 24
excision of the aortic endograft, left subclavian artery stent graft, and proximal descending thoracic aorta | 24
inline anatomic reconstruction of the aorta | 24
intraoperative cultures from the endograft, aortic wall, and vegetations grew Candida | 24
initiated on lifelong oral antifungal therapy | 24
short course of broad-spectrum antibiotics | 24
postoperative course complicated by a chylothorax | 48
treated with total parenteral nutrition | 48
coil embolization and Onyx glue obliteration of the thoracic duct | 72
discharged home | 264
computed tomography angiography demonstrated a patent repair and no evidence of infection | 1440
doing well at 6-month postoperative check | 4320