46 years old | 0 | 0 | Factual
Asian-Indian | 0 | 0 | Factual
male | 0 | 0 | Factual
tropical chronic pancreatitis | -8760 | 0 | Factual
oral pancreatic enzyme therapy | -8760 | 0 | Factual
exocrine pancreatic insufficiency | -8760 | 0 | Factual
non-insulin-dependent diabetes mellitus | -2190 | 0 | Factual
glucotrol | -2190 | 0 | Factual
midepigastric pain | -6 | 0 | Factual
pain control with narcotics | -6 | 0 | Factual
nausea | 48 | 48 | Factual
vomiting | 48 | 48 | Factual
no fever | 48 | 48 | Negated
CT scan | 48 | 48 | Factual
fatty atrophy of pancreatic head and uncinate process | 48 | 48 | Factual
pancreatic duct filled with large calcifications | 48 | 48 | Factual
possible obstruction at the level of the neck | 48 | 48 | Possible
marked upstream ductal dilatation | 48 | 48 | Factual
admitted for management of pain | 48 | 48 | Factual
previous CT scan | -144 | -144 | Factual
chronic atrophic calcific pancreatitis | -144 | -144 | Factual
dilated pancreatic duct | -144 | -144 | Factual
intraductal calculi | -144 | -144 | Factual
ERCP | -144 | -144 | Factual
pancreatography | -144 | -144 | Factual
medically managed | -144 | -144 | Factual
discharged | -144 | -144 | Factual
fever | 48 | 48 | Factual
chills | 48 | 48 | Factual
rigors | 48 | 48 | Factual
severe sepsis | 48 | 48 | Factual
septic shock | 48 | 48 | Factual
intubated | 48 | 48 | Factual
hypoxemic respiratory failure | 48 | 48 | Factual
acute respiratory distress syndrome | 48 | 48 | Factual
multiorgan failure | 48 | 48 | Factual
broad-spectrum antibiotics | 48 | 240 | Factual
vasopressor support | 48 | 240 | Factual
activated recombinant human protein C | 48 | 240 | Factual
ultrasound of abdomen | 48 | 48 | Factual
markedly dilated pancreatic duct | 48 | 48 | Factual
calculus within the duct | 48 | 48 | Factual
diffusely echogenic pancreas | 48 | 48 | Factual
prominent common bile duct | 48 | 48 | Factual
no obvious obstructing calculi | 48 | 48 | Negated
bedside emergency ERCP | 72 | 72 | Factual
frank pus expelling spontaneously | 72 | 72 | Factual
no evidence of papillitis | 72 | 72 | Negated
no evidence of tumor | 72 | 72 | Negated
no previous sphincterotomy | 72 | 72 | Negated
evacuation of pus | 72 | 72 | Factual
cholangiogram | 72 | 72 | Factual
normal biliary tree | 72 | 72 | Factual
no stones | 72 | 72 | Negated
pancreatogram | 72 | 72 | Factual
marked dilatation of main pancreatic duct | 72 | 72 | Factual
single distal calculus | 72 | 72 | Factual
guide wire introduced | 72 | 72 | Factual
evacuation of pus | 72 | 72 | Factual
5-cm-long 5 F stent placed | 72 | 72 | Factual
no more pus draining | 72 | 72 | Negated
ASPD | 72 | 240 | Factual
reevaluation of pancreas | 144 | 144 | Factual
inflammatory changes | 144 | 144 | Factual
edema | 144 | 144 | Factual
diminished ductal dilatation | 144 | 144 | Factual
distal migration of calculus | 144 | 144 | Factual
no evidence of pancreatic necrosis | 144 | 144 | Negated
no fluid collection | 144 | 144 | Negated
bilateral moderate pleural effusions | 144 | 144 | Factual
dramatic signs of clinical improvement | 168 | 168 | Factual
stabilization of hemodynamic parameters | 168 | 168 | Factual
blood cultures grew Klebsiella ornithinolytica | 168 | 168 | Factual
sensitive to antibiotics | 168 | 168 | Factual
extubated | 240 | 240 | Factual
transferred from intensive care unit | 240 | 240 | Factual
completed antibiotic course | 240 | 240 | Factual
discharged home | 240 | 240 | Factual
follow-up examinations | 720 | 2160 | Factual
no further complications | 720 | 2160 | Negated