87 years old | 0
white | 0
male | 0
end-stage renal disease | 0
atrial fibrillation | 0
warfarin | -672
maintenance HHD | -672
NxStage machine | -672
laparoscopic appendicectomy | -24
intra-abdominal abscess | -24
sepsis | -24
tamponade | -24
bloody pericardial effusion | -24
therapeutic pericardiocentesis | -24
warfarin discontinued | -24
heparin-free HHD | 0
intermittent heparin-free hemodialysis | 0
Fresenius machine | 0
Optiflux 160 NR dialyzers | 0
normal saline flushes | 0
extracorporeal circuits clotting | 0
high venous pressures | 0
compromised HHD | 0
heparin anticoagulation contraindicated | 0
normal saline flushes failed | 0
clotting problem | 0
Locke-Onuigbo Maneuver | 0
CAR-170-C NXSTAGE Chronic cartridge | 0
rotating filter | 0
clockwise rotation | 0
counterclockwise rotation | 0
clotting resolved | 0
smooth heparin-free HHD | 24
no normal saline flushes | 24
stable HHD treatments | 24
discharged home | 0
home hemodialysis | 0
 NxStage machine | 0
CAR-170-C NXSTAGE Chronic cartridge | 0
heparin-free HHD | 0
normal saline-flush-free HHD | 0
patient satisfied | 168
wife satisfied | 168
daily diary | 0
December 2019 | -720
January 2020 | 0
Locke-Onuigbo Maneuver | 0
repeated rotational manipulations | 0
antigravity effect | 0
thrombogenesis prevention | 0
sustainable HHD | 0
fluidity maintenance | 0
extracorporeal circuit | 0
adequate hemodialysis | 0
further study | 168
biomedical engineers | 168
repeatability | 168
reproducibility | 168
electric motor | 168
commercially successful method | 168