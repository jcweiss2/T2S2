78 years old | 0
female | 0
admitted to the hospital | 0
acute non-ST segment elevation myocardial infarction | -240
chest pain | -240
shortness of breath | -240
dyspnea | -240
tracheal intubation | -240
ventilator-assisted ventilation | -240
vasodilation | -240
transferred to the ICU | -240
hypertension | -3600
coronary heart disease | -3600
cerebral infarction | -3600
anterior wall myocardial infarction | -3600
decreased blood pressure | 0
increased heart rate | 0
fever | 0
septic shock | 0
cardiogenic shock | 0
blood oxygen saturation (SpO2) fluctuations above 97% | 0
thick breath sounds in lungs | 0
slight moist rale in lower lungs |-0
heart rate of 100 bpm | 0
low and blunt heart sound | 0
no noise in each valve area | 0
dry necrosis of the right lower foot | 0
scattered ecchymoses | 0
serum creatine kinase-MB concentration of 25.8 ng/mL | 0
white blood cell count of 24.25 × 109/L | 0
double lung infection | 0
moderate mitral regurgitation | 0
mild aortic regurgitation | 0
right leg gangrene | 0
right leg peripheral arterial occlusive disease | 0
imipenem | 0
cilastatin sodium | 0
dopamine | 0
norepinephrine | 0
percutaneous coronary intervention (PCI) | -72
coronary angiography | -72
right coronary artery stent implantation | -72
70%-80% stenosis in the anterior descending artery | 0
80% stenosis in the circumflex artery | 0
90% stenosis in the right coronary artery | 0
right coronary artery dominant type | 0
three-vessel coronary lesions | 0
increased body temperature (38.5-39 ºC) | -72
white blood cell count of 33.74 × 109/L | -72
dry skin necrosis of the right lower extremity | -72
scattered ecchymoses | -72
right middle iliac artery occlusion | -72
endotracheal tube in place | -72
fever | -72
SpO2 over 97% with medium flow oxygen inhalation | -72
mid-thigh amputation | 0
tracheal catheter in place | 0
dopamine infusion at 5 µg/kg/min | 0
norepinephrine infusion at 0.06 µg/kg/min | 0
non-invasive blood pressure of 95/45 mmHg | 0
heart rate of 98 bpm | 0
SpO2 of 99% | 0
left radial artery puncture catheter | 0
anesthesia system connected to tracheal catheter | 0
ultrasound-guided fascia iliaca compartment block | 0
ropivacaine hydrochloride injection | 0
midazolam | 0
sufentanil | 0
cisatracurium | 0
etomidate | 0
sevoflurane inhalation anesthesia | 0
operation duration of 65 min | 0
bispectral index maintained between 45 and 60 | 0
vasoactive drugs used | 0
stable vital signs during perioperative period | 0
CPOT score of 2 at 6 h after surgery | +6
Ramsay sedation score of 3 | +6
improved inflammatory indicators two days after operation | +48
tracheal intubation removed | +48
discharged | +48
