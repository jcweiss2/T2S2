75 years old | 0
male | 0
hypertension | 0
sequelae of ischemic stroke | 0
mild right hemiplegia | 0
accidentally fell into a creek | -1
submerged in the water | -1
rescued | -1
Glasgow Coma Scale was E3V3M6 | 0
body temperature was 33.4°C | 0
heart rate was 88 beats/min | 0
blood pressure was 120/60 mmHg | 0
respiratory rate was 26 breaths/min | 0
oxygen saturation was 92% | 0
bilateral coarse crackles | 0
hypothermia | 0
rewarming using a warming blanket | 0
antibiotic therapy (ampicillin and sulbactam) | 0
non-invasive ventilation | 0
oxygenation steadily deteriorated | 0
intubated and mechanically ventilated | 0
transferred to the emergency department | 0
sedated with propofol | 0
body temperature was 36.4°C | 0
heart rate was 104 beats/min | 0
blood pressure was 123/84 mmHg | 0
respiratory rate was 30 breaths/min | 0
oxygen saturation level was 91% | 0
bilateral diminished breath sounds | 0
arterial blood gas analysis | 0
pH of 7.34 | 0
PaCO2 of 42 mmHg | 0
PaO2 of 199 mmHg | 0
HCO3 of 21.9 mmol/L | 0
white blood cell count of 2980/μL | 0
neutrophils 63.5% | 0
hemoglobin level of 15.3 g/dL | 0
platelet level of 159,000/μL | 0
C-reactive protein level of 0.6 mg/dL | 0
procalcitonin level of 59.37 ng/mL | 0
ultrasonographic examination of the heart | 0
normal ejection fraction | 0
no valvular disease | 0
chest radiography | 0
computed tomography (CT) of the lung | 0
diffuse infiltrates bilaterally | 0
no pleural effusion | 0
diagnosis of acute respiratory distress syndrome (ARDS) | 0
diagnosis of septic shock | 0
treated with isotonic crystalloids | 0
intravenous broad-spectrum antibiotic (meropenem) | 0
vasopressors | 0
protective ventilation | 0
methylprednisolone 80 mg daily | 24
beta-D-glucan assay | 72
elevated at 37.6 pg/mL | 72
tracheal aspirate culture was found positive for Aeromonas hydrophila | 120
blood culture was negative | 120
switched to piperacillin/tazobactam | 120
hypoxia continued to worsen | 120
died | 168
CT scans obtained at autopsy | 168
no focal lesion in the brain | 168
both lungs were completely infiltrated with effusion | 168
severely congested | 168
each weighed over 1000 g | 168
embolus was detected in the right pulmonary artery | 168
microscopic analysis with Grocott staining | 168
diffuse filamentous fungi throughout the lungs | 168
within necrotizing tissue and intravascular lesions | 168
in the heart, stomach, and thyroid gland | 168
pulmonary embolus contained filamentous fungi | 168
cultured biopsies from both lungs | 168
identified as Aspergillus fumigatus | 168
diagnosed as invasive aspergillosis complicated by pulmonary embolism | 168