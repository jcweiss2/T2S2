56 years old | 0
male | 0
admitted to the hospital | 0
multiply recurrent ventral hernia | -672
open recurrent umbilical hernia repair | -672
Atrium C-QUR mesh | -672
seroma formation | -672
open wound | -672
wound vacuum therapy | -672
multiple washouts | -672
mesh excision | -672
repeat ventral hernia repair | -672
Alloderm mesh | -672
medial component separation | -672
recurrence | -672
significant pain | -672
discomfort | -672
large ventral hernia defect | -672
preoperative body mass index | -24
tobacco chewer | -24
hypertension | -24
multiply operated abdomen | -24
combined endoscopic bilateral component separation | 0
open recurrent giant ventral incisional hernia repair | 0
underlay biologic mesh | 0
extensive open lysis of adhesions | 0
dermatolipectomy | 0
hernia defect | 0
estimated blood loss | 0
peak airway pressures | 0
extubation | 0
transferred to the medical-surgical ward | 0
oliguric | 4
elevated creatinine level | 4
hyperkalemia | 4
intubation | 4
paralysis | 4
nasogastric tube decompression | 4
intraabdominal pressures | 4
diagnosis of ACS | 4
urine output | 6
creatinine level | 12
potassium level | 12
bladder pressures | 12
peak airway pressures | 12
paralytic medication discontinued | 48
bladder pressures monitored | 48
peak airway pressures monitored | 48
urine output monitored | 48
creatinine level monitored | 48
continuous positive airway pressure trials | 72
extubated | 96
trickle-tube feeds | 96
ambulatory | 96
abdominal binder | 96
clear liquid diet | 120
regular diet | 144
transferred to the floor | 120
discharged | 192
home oxygen | 192