75 years old | 0
male | 0
admitted to the hospital | 0
arterial hypertension | -8760
chronic atrial fibrillation | -8760
type 2 diabetes | -8760
moderate chronic renal failure | -8760
myocardial infarction | -7920
coronary artery bypass grafting | -7920
implantable defibrillator | -7920
low left ventricle ejection fraction | -7920
ramipril | -8760
cardensiel | -8760
aldactone | -8760
fluindione | -8760
metformin | -8760
furosemide | -8760
anasarca | -144
exertional dyspnea | -144
diuretic treatment | -144
furosemide | -144
spironolactone | -144
indwelling urinary catheterization | -144
acute renal failure | -144
dobutamine | -144
arterial hypotension | -144
increased inflammatory syndrome | -144
oliguria | -144
persistent hypotension | -144
confused | 0
hypothermic | 0
atrial tachycardia | 0
capillary blood glucose level | 0
mottling | 0
deep hypotension | 0
cloudy and foul-smelling urinary residues | 0
thrombocytopenia | 0
hyperleukocytosis | 0
inflammatory syndrome | 0
C-reactive protein | 0
procalcitonin | 0
acute renal failure | 0
creatinine | 0
urea | 0
liver function tests | 0
troponins | 0
hyperlactatemia | 0
glycated hemoglobin | -72
vasoplegic hemodynamic profile | 0
mixed cardiogenic and septic shock | 0
thoraco-abdomino-pelvic computed tomography | 2
bilateral pleural effusions | 2
cardiomegaly | 2
intra- and peri-bladder air | 2
emphysematous cystitis | 2
central venous line | 2
noradrenaline | 2
mineralocorticoids | 2
intravenous insulin therapy | 2
microbiological sampling | 2
probabilistic antibiotic therapy | 2
piperacillin/tazobactam | 2
amikacin | 2
hemodynamic monitoring | 2
cardiorespiratory arrest | 3
ventricular tachycardia | 3
external cardiac massage | 3
adrenalin | 3
internal electric shock | 3
intubated | 3
sedated | 3
series of cardiorespiratory arrest | 6
shockable rhythm | 6
electromechanical dissociation | 6
no flow | 6
low flow | 6
refractory shock | 9
multivisceral failure | 9
cytobacteriological examination of urine | 9
Enterobacter cloacae | 9
methicillin Staphylococcus aureus | 9
blood cultures | 9
death | 9