66 years old | 0
female | 0
morbid obesity | 0
hypertension | 0
hyperlipidemia | 0
non-insulin dependent diabetes mellitus | 0
coronary artery disease | 0
admitted to the hospital | 0
sepsis | 0
lower extremity ulceration | 0
osteomyelitis | 0
immobilized in the collapsed floor of her mobile home | -336
without access to hydration for long time | -336
contacted family members for assistance | -336
refused outside assistance | -336
requested medical attention | -336
transported by emergency medical services to the emergency department | -24
anxious | 0
temperature 99.8o F | 0
pulse 109 beats per minute | 0
blood pressure 128/60 mm Hg | 0
respiratory rate 18 breaths per minute | 0
multiple necrotic ulcers with brown discharge | 0
bilateral lower extremities | 0
left heel | 0
sacral decubitus area | 0
atrial fibrillation with rapid ventricular response | 0
computed tomography of the thorax and abdomen | 0
no acute abnormalities | 0
vancomycin | 0
piperacillin-tazobactam | 0
empiric coverage of common pathogens | 0
white cell count of 23.6k per mm3 | 0
hemoglobin 9.7 g/dL | 0
platelet count of 601k per mm3 | 0
sodium 128 mEq/L | 0
bicarbonate 18 mEq/L | 0
urea nitrogen 46 mg/dL | 0
creatinine 2.03 mg/dL | 0
lactic acid 2.76 mmol/L | 0
cultures of urine and blood | 0
orthopedic and infectious disease services were consulted | 0
blood cultures grew Clostridium sporogenes | 24
urine cultures grew Enterococcus spp. | 24
daptomycin | 24
ertapenem | 24
clindamycin | 24
repeat blood cultures were negative | 120
clinical gas gangrene | 120
severe destruction to the subcutaneous tissue | 120
whole planter surface of the left foot | 120
parts of the right foot | 120
general surgery was consulted | 120
below knee amputation of the left leg | 120
right foot disarticulation | 120
patient refused the amputations | 120
treatment with antimicrobial agents | 120
patient clinical conditions continued to deteriorate | 168
patient refused all medical management | 168
placed on comfort measures | 168
expired | 192