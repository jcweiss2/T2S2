90 years old | 0
male | 0
admitted to the hospital | 0
severe abdominal pain | 0
nausea | 0
vomiting | 0
inability to defecate or pass gas | 0
abdominal pain and constipation | -4380
lost weight | -8760
hypertension | -8760
cachectic | 0
abdomen distended | 0
mucosae dry | 0
blood pressure 90/50 mmHg | 0
pulse rate 95 bpm | 0
body temperature 37.9°C | 0
rebound tenderness | 0
guarding | 0
WBC 8.890 | 0
neutrophil 86.1% | 0
Hemoglobin 14 gr/dL | 0
BUN 38 mg/dL | 0
creatinine 0.8 mg/dL | 0
diffuse air-fluid levels | 0
intestinal obstruction | 0
tumoral obstruction | 0
viscus perforation | 0
laparotomy | 0
encapsulation of small intestine | 0
fibrocollagenous membrane | 0
abdominal cocoon syndrome | 0
loop ileostomy | 0
intensive care unit | 0
septic shock | 72
multiorgan failure | 72
WBC 1880/µL | 72
BUN 123 mg/dL | 72
creatinine 2.92 mg/dL | 72
albumin 2.4 gr/dL | 72
died | 72