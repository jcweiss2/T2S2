low-grade fever | -48
dry cough | -48
shortness of breath | -48
admission | 0
elective right total knee replacement | -168
pain in the right knee | 0
redness in the right knee | 0
swelling in the right knee | 0
essential hypertension | 0
obesity | 0
myasthenia gravis in remission | 0
osteoarthritis | 0
body temperature of 37.3°C | 0
blood pressure of 121/82 | 0
pulse of 87 beats per minute | 0
respiratory rate of 16 breaths per minute | 0
oxygen saturation of 87% | 0
bilateral rhonchi with rales | 0
patchy air space opacity in the right upper lobe suspicious for pneumonia | 0
rapid nucleic acid amplification test for influenza A and B negative | 0
nasopharyngeal swab specimen obtained | 0
broad-spectrum antibiotics with cefepime and levofloxacin started | 0
supportive care with 2 L of supplemental oxygen started | 0
mild diarrhea | 72
generalized weakness | 72
fatigue | 72
evaluation by Neurology | 72
intravenous immunoglobulin started | 72
mild MG exacerbation | 72
pending MG crises | 72
arterial blood gases monitored | 0
complete blood count monitored | 0
basic metabolic profile studies monitored | 0
mild absolute lymphopenia | 0
anemia | 0
pH of 7.46 | 0
pCO2 of 44.6 mmHg | 0
pO2 of 94.7 mmHg | 0
bicarbonate of 31.4 mmol/L | 0
creatinine kinase normal | 144
lactic acid normal | 144
lactate dehydrogenase elevated | 144
ferritin elevated | 144
interleukin-6 elevated | 144
progressively increasing shortness of breath | 24
oxygen requirements increased | 24
nasopharyngeal swab results positive for SARS-CoV-2 | 96
hydroxychloroquine started | 96
azithromycin started | 96
zinc sulfate started | 96
oral vitamin C started | 96
blood and sputum cultures did not grow any organisms | 96
broad-spectrum antibiotics discontinued | 96
shortness of breath worsened | 144
oxygen requirements increased | 144
drowsy | 144
moderate distress | 144
unable to protect the airways | 144
blood pressure of 78/56 mmHg | 144
heart rate of 112 beats per minute | 144
temperature of 38°C | 144
respiratory rate of 28 breaths per minute | 144
bilateral alveolar infiltrates due to pneumonia and interstitial edema | 144
intubated | 144
mechanical ventilation started | 144
norepinephrine started | 144
colchicine started | 144
high-dose vitamin C infusion started | 168
clinical condition improved | 192
norepinephrine support stopped | 192
CXR showed significant improvement | 240
spontaneous breathing trial tolerated | 240
pH of 7.49 mmHg | 240
pCO2 of 40.2 mmHg | 240
pO2 of 77.1 mmHg | 240
bicarbonate of 30.2 mmol/L | 240
extubated | 240
oxygen saturation of 92% | 384
CXR revealed almost complete resolution of the infiltrates | 384
discharged from the hospital | 384
hydroxychloroquine treatment completed | 120
azithromycin treatment completed | 120
colchicine treatment completed | 120
high-dose vitamin C infusion completed | 240
oral zinc sulfate completed | 240