67 years old | 0
    man | 0
    hospitalized with severe acute pancreatitis | 0
    transferred to our hospital | 72
    past medical history of chronic pancreatitis | -72
    past medical history of diabetes | -72
    consumed 5 liters of beer every day for 47 years | -72
    body temperature 36.6℃ | 0
    blood pressure 172/94 mmHg | 0
    heart rate 96 beats/min | 0
    respiratory rate 21 breaths/min | 0
    abdomen hard and flat | 0
    tenderness | 0
    defensiveness | 0
    increased white blood cell count (20,000 /μL) | 0
    increased serum CRP (31.03 mg/dL) | 0
    increased serum amylase (280 IU/L) | 0
    increased serum lipase (254 U/L) | 0
    HbA1c 9.6% | 0
    CE-CT revealed low enhancement of pancreatic parenchyma | 0
    CE-CT revealed surrounding fluid collection | 0
    prognostic factor score 2 points (CRP >15 mg/dL and SIRS) | 0
    diagnosed with severe acute pancreatitis | 0
    fluid resuscitation (100 mL/kg daily) started | 0
    treated with nafamostat mesylate (240 mg daily) for 5 days | 0
    treated with antibiotics (meropenem 1.5 g daily) for 10 days | 0
    stayed in ICU for 12 days | 0
    abdominal pain improved | 0
    inflammation improved | 0
    developed high fever | 384
    no urinary tract infection | 384
    no pneumonia | 384
    no infected pancreatic fluid | 384
    Candida albicans detected in blood cultures | 384
    Candida albicans detected in central venous catheter cultures | 384
    blood β-D glucan 47.4 pg/mL | 384
    diagnosed with candidemia | 384
    ophthalmologic examinations performed | 384
    exudative plaques consistent with fungal infection observed | 384
    diagnosed with candida endophthalmitis | 384
    no visual disturbance | 384
    administered micafungin (150 mg daily) | 384
    administered caspofungin (75 mg daily) | 384
    administered fluconazole (800 mg daily) | 384
    intravenous fluids administered for 59 days | 384
    blood cultures evaluated weekly | 384
    disappearance of C. albicans from blood stream | 456
    exudative plaques disappeared | 456
    blood β-D glucan negative (19.8 pg/mL) | 1200
    discharged | 2280
    