20 years old | 0
pregnant | 0
26-weeks of gestation | 0
anti-epileptic therapy with carbamazepine | 0
consumption of 4000 mg of carbamazepine | -4
denied concomitant overdose with other medications | -4
gastric lavage | -4
transferred to hospital | 0
Glasgow coma score (GCS) was 3/15 | 0
pulse rate was 138/min | 0
blood pressure 110/70 mmHg | 0
respiratory rate 25/min | 0
capillary blood glucose level was 109 mg/dl | 0
pupils were dilated 6 mm bilaterally | 0
pupils reacting to light | 0
deep tendon reflexes were sluggish | 0
Babinski sign was negative | 0
intubated for low sensorium | 0
multi-dose activated charcoal therapy | 0
shifted to ICU | 0
serum carbamazepine level was > 20 μg/ml | 0
hemoglobin was 8 g/dl | 0
white count 15,200/cumm | 0
renal function was normal | 0
liver function test was normal | 0
coagulation profile was normal | 0
circulatory shock | 6
fluid resuscitation | 6
low dose vasopressors | 6
empiric antibiotic therapy | 6
negative cultures | 6
low procalcitonin (0.34) | 6
absence of a definite focus of infection | 6
discontinued antibiotic therapy | 12
hypoglycemia | 48
bolus doses of 50% dextrose | 48
infusion of 25% dextrose | 48
infusion given for 60 hours | 108
no further episodes of hypoglycemia | 108
serum carbamazepine level on the third day was 17.3 μg/ml | 72
serum carbamazepine level decreased to sub therapeutic range | 168
extubated | 168
vasoactive agents were weaned | 168
serum carbamazepine level normalized | 168
no further hypoglycemic episodes at 2-months follow-up | 720