4 months old| 0
mulatto | 0
boy | 0
admitted to the service | 0
miliaria rubra-like lesions on the neck | -2928
miliaria rubra-like lesions on the upper limb folds | -2928
miliaria rubra-like lesions on the lower limb folds | -2928
referred to a pediatrician | -2928
prescription of powder with bismuth subgallate and zinc oxide | -2928
prescription of cream with ketoconazole, betamethasone dipropionate, and neomycin sulfate | -2928
application of cream for one month | -2928
no improvement | -2232
prescription of prednisolone 0.8mg/kg/day for seven days | -2232
prescription of potassium permanganate topical solution | -2232
refractoriness of the condition | -2232
prescription of single-dose ampoule of betamethasone intramuscularly | -2232
lesions spread to trunk | -2232
lesions spread to face | -2232
lesions spread to scalp | -2232
lesions became crusty | -2232
referred to dermatology clinic | -2232
diagnosis of severe seborrheic dermatitis | -2232
mother followed throughout pregnancy | -2232
negative serological tests (VDRL, hepatitis B, toxoplasmosis, HIV) | -2232
denied intercurrence except topical treatment for scabies during pregnancy | -2232
child born healthy | -2232
multiple erythematous papules | 0
crusted lesions | 0
erythematous lesions | 0
disseminated lesions on body | 0
lesions mainly affecting trunk | 0
lesions mainly affecting scalp | 0
nail dystrophy | 0
abdominal fissures | 0
hypoactive | 0
tachycardic | 0
febrile | 0
cushingoid facies | 0
anasarca | 0
diagnostic hypothesis of crusted scabies | 0
diagnostic hypothesis of Norwegian scabies | 0
secondary infection | 0
sepsis | 0
mother complained of pruritus | 0
grandparents complained of pruritus | 0
nocturnal pruritus | 0
mother's erythematous hyperchromic papules on abdomen | 0
mother's erythematous hyperchromic papules on back | 0
compatible with scabies | 0
dermoscopy showing triangular structures | 0
dermoscopy showing millipede-like structures | 0
skin biopsy conducted | 0
laboratory tests requested | 0
hospitalized in pediatric hospital | 0
histopathology revealing tunnels in stratum corneum | 0
presence of parasite | 0
significant leukocytosis | 0
left shift | 0
thrombocytopenia | 0
increased inflammatory markers | 0
intravenous antibiotic therapy | 0
topical permethrin lotion 1% once daily | 0
contact isolation | 0
family treated with oral ivermectin | 0
family treated with topical permethrin lotion 5% | 0
improvement of cutaneous lesions on day 10 | 240
septic shock | 240
treatment in intensive care unit | 240
cardiac arrest | 240
death | 240
