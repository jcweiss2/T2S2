42 years old| 0
    woman | 0
    admitted | 0
    dyspnea | 0
    enduring cough | 0
    several days | 0
    no underlying illness | 0
    oseltamivir | -96
    influenza A (H1N1) | -96
    PCR | -96
    blood pressure 90/60 mm Hg | 0
    pulse rate 100 beats per minute | 0
    respiratory rate 22 breaths per minute | 0
    body temperature 36.3℃ | 0
    oxygen saturation 93.3% | 0
    2 L/min oxygen via nasal cannula | 0
    coarse breathing sounds in both lung fields | 0
    chest X-ray peribronchial consolidations | 0
    multifocal ground glass opacities in both hilar areas | 0
    arterial blood gas analysis pH 7.390 | 0
    PCO2 27.9 mm Hg | 0
    PO2 67.9 mm Hg | 0
    bicarbonate 17.0 mmol/L | 0
    hemoglobin 13.8 g/dL | 0
    white blood cell count 4,640 cells/mm3 | 0
    neutrophils 77.4% | 0
    platelet count 161,000 cells/mm3 | 0
    C-reactive protein 30.24 mg/dL |*0
    serum albumin 3.7 g/dL | 0
    aspartate aminotransferase 35 U/L | 0
    alanine aminotransferase 27 U/L | 0
    total bilirubin 0.9 mg/dL | 0
    serum creatinine 1.8 mg/dL | 0
    chest CT tracheobronchial wall thickening | 0
    multifocal patchy consolidations | 0
    nodular opacities with cavitations on both lungs | 0
    bronchoscopy severe mucosal inflammation | 0
    sloughing | 0
    diffuse cobblestone-like multiple mucus swelling of exudates | 0
    partial obstruction of airways | 0
    pseudomembranous tracheobronchitis | 0
    no bronchoscopic biopsy | 0
    respiratory failure | 0
    transferred to ICU | 0
    mechanical ventilation | 0
    MSSA isolated from bronchial washing fluid | 0
    acid fast bacillus stain negative | 0
    PCR for Mycobacterium tuberculosis negative | 0
    serum galactomannan test negative | 0
    pseudomembranous tracheobronchitis following influenza | 0
    changed antibiotics to ciprofloxacin and amoxicillin/clavulanate | 0
    required tube thoracotomy for bilateral pneumothoraces | 0
    infected pneumatoceles | 0
    drained fluid from infected pneumatocele | 0
    changed antibiotics to colistin | 0
    multi-drug resistant Acinetobacter baumannii isolated | 0
    improvement of dyspnea | 0
    improvement of chest X-ray | 0
    remove pigtail catheter | 0
    follow-up bronchoscopy improvement | 0
    discharged | 1248
    <|eot_id|>
