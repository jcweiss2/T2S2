79 years old | 0
female | 0
myalgias | -672
spontaneous bowel diverticula perforation | -672
resection | -672
ileostomy | -672
polyarteritis nodosa | -672
corticosteroids | -672
immunosuppressants | -672
admitted to the medical Intensive Care Unit | 0
severe acute on chronic abdominal pain | 0
sepsis | 0
abdominal computed tomography | 0
gallbladder fundus wall thickening | 0
pericholecystic edema | 0
dependent cholelithiasis | 0
right posteroinferior hepatic abscess | 0
hepatobiliary scan | 24
Tc-99m diisopropyliminodiacetic acid | 24
incomplete gallbladder filling | 24
no radiotracer filling of the distal gallbladder fundus | 24
catheter intervention for the hepatic abscess | 48
Escherichia coli | 48
metastatic septic arthritis | 72
osteomyelitis | 72
persistent bacteremia | 96
second Tc-99m DISIDA hepatobiliary scan | 120
nonfilling of the gallbladder | 120
acute cholecystitis | 120
surgical and medical management | 144
improvement in the patient's condition | 168
partial gallbladder stricture | -672
dumbbell-shaped gallbladder | -672
percutaneous cholangiogram | 192
focal inflammation of the distal end of the dumbbell gallbladder | 192
dumbbell gallbladder cholecystitis | 192
focal gallbladder wall thickening | 0
focal pericholecystic edema | 0
layering cholelithiasis | 24
biliary sludge | 24
retained bile | 24
mass effect from tumor | 24
hepatic abscess adjacent to the distal end of the dumbbell gallbladder | 0
acute on chronic upper abdominal pain | 0