70 years old | 0
    male | 0
    type 2 diabetes mellitus | 0
    previous kidney transplantation in 2007 | -105216
    previous kidney transplantation in 2017 | -57600
    end-stage renal disease | -105216
    focal segmental glomerulosclerosis | -105216
    chronic antibody-mediated rejection | -57600
    presented to intensive care unit | 0
    distributive shock | 0
    requiring vasopressor support | 0
    empirically started on piperacillin-tazobactam | 0
    blood cultures grew non-lactose fermenting gram-negative bacillus | 19
    underwent cystoscopy for microscopic hematuria | -96
    no peri-procedural antimicrobials | -96
    bilobar prostatic hypertrophy | -96
    no significant macroscopic bladder abnormalities | -96
    blood culture isolate identified as Pseudomonas aeruginosa | 19
    susceptible to all anti-pseudomonal antimicrobials | 19
    appropriate piperacillin-tazobactam dosing | 19
    rapid defervescence | 19
    normalized hemodynamic parameters | 19
    transferred to ward | 19
    transitioned to oral ciprofloxacin | 19
    persistent P. aeruginosa bacteremia | 19
    high-dose ceftazidime added | 19
    persistent bacteremia for 7 days | 168
    no indwelling catheters or prosthetic devices | 168
    no perinephric abscess | 168
    no hydronephrosis | 168
    no clinical evidence of pneumonia | 168
    no radiographic evidence of pneumonia | 168
    no known cardiac valvulopathy | 168
    no arterial aneurysms | 168
    ongoing delirium | 168
    reported rectal pain | 168
    digital rectal examination revealed enlarged and tender prostate | 168
    endorectal ultrasound confirmed prostatomegaly | 168
    increased vascularity | 168
    multiple prostatic abscesses | 168
    largest abscess 3.4 cm | 168
    ultrasound-guided transrectal needle aspirate | 168
    drained small amounts of thick purulent fluid | 168
    cultures grew P. aeruginosa | 168
    underwent transurethral resection of prostate | 168
    unroofing of prostatic abscess | 168
    surgical pathology revealed foamy histiocytes | 168
    abundant necrotic debris | 168
    rare hemosiderin deposition | 168
    Auramine-rhodamine stain negative for acid-fast bacilli | 168
    Grocott-Gomori’s methamine silver stain negative for fungi | 168
    histiocytes did not express cytokeratin AE1/AE3 | 168
    excluded epithelial neoplasm | 168
    diagnostic of XG prostatitis | 168
    completed 10 days of oral ciprofloxacin | 408
    surveillance urine cultures grew P. aeruginosa | 408
    new lower urinary tract symptoms | 408
    decision for 6 additional weeks of ciprofloxacin | 408
    completed without adverse events | 1272
    follow-up assessment one month after discontinuing antimicrobials | 1704
    clinically doing very well | 1704
    no infectious symptoms | 1704
    no urinary tract symptoms | 1704
    prior urological instrumentation | -96
    microscopic hematuria | -96
    chronic urinary tract infections | -96
    immune dysregulation | -96
    bacterial sepsis triggered by cystoscopy | -96
    abnormal immune response | -96
    recurrent or chronic subclinical infection | -96
    chronic allograft dysfunction | -96
    chronic rejection | -96
    chronic kidney disease | 0
    immunosuppression | 0
    diabetes mellitus | 0
    prostatic abscesses | 168
    gram-negative bacilli bloodstream infections | 168
    persistent P. aeruginosa bacteremia | 168
    XG prostatitis | 168
    transurethral resection of the prostate | 168
    surgical resection | 168
    histopathology diagnosis | 168
    no significant adverse events | 1272