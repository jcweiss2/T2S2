69 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
stabbed herself in the abdomen | -1 | -1 | Factual
admitted to emergency department | 0 | 0 | Factual
blood pressure could not be measured | 0 | 0 | Factual
pulseless electrical activity | 0 | 0 | Factual
body temperature 35.0 °C | 0 | 0 | Factual
oxygen saturation 99 % | 0 | 0 | Factual
Glasgow Coma Scale score 3 | 0 | 0 | Factual
agonal respiration | 0 | 0 | Factual
wound 5 cm on upper abdomen | 0 | 0 | Factual
intra-abdominal fluid collection | 0 | 0 | Factual
emergency thoracotomy | 0 | 1 | Factual
aortic cross-clamping | 0 | 15 | Factual
open cardiac massage | 0 | 15 | Factual
epinephrine administration | 0 | 15 | Factual
temporary return of spontaneous circulation | 15 | 15 | Factual
hemodynamically unstable | 15 | 24 | Factual
laparotomy | 15 | 24 | Factual
injuries to common hepatic and splenic arteries | 15 | 24 | Factual
injuries to pancreas, spleen, and liver | 15 | 24 | Factual
ligation of injured arteries | 15 | 24 | Factual
distal pancreatectomy | 24 | 24 | Factual
splenectomy | 24 | 24 | Factual
liver sutured | 24 | 24 | Factual
norepinephrine administration | 24 | 48 | Factual
second-look surgery | 24 | 24 | Factual
no active bleeding or ischemic change | 24 | 24 | Factual
abdominal wall closure | 72 | 72 | Factual
regular examinations for ischemic changes | 72 | 168 | Factual
enhanced CT scan | 96 | 96 | Factual
disruption of celiac artery | 96 | 96 | Factual
gastroduodenal artery arising from superior mesenteric artery | 96 | 96 | Factual
gastroscopy | 216 | 216 | Factual
patchy mucosal necrosis | 216 | 216 | Factual
conservative treatment | 216 | 552 | Factual
fever 39 °C | 552 | 552 | Factual
pain in stomach | 552 | 552 | Factual
white blood cell count 34,000/mm3 | 552 | 552 | Factual
C reactive protein 13.4 mg/dL | 552 | 552 | Factual
CT scan | 552 | 552 | Factual
air in gastric wall | 552 | 552 | Factual
intra-abdominal free air | 552 | 552 | Factual
gastric necrosis suspected | 552 | 552 | Factual
gastroscopy | 552 | 552 | Factual
extensive mucosal necrosis | 552 | 552 | Factual
emergency surgery | 552 | 552 | Factual
total gastrectomy with Roux-en-Y reconstruction | 552 | 552 | Factual
histological findings of stomach | 552 | 552 | Factual
diffuse necrotic changes | 552 | 552 | Factual
inflammatory cell infiltrations | 552 | 552 | Factual
no invasive fungal infection | 552 | 552 | Factual
leakage on duodenal stump | 696 | 696 | Factual
continuous tube drainage | 696 | 696 | Factual
consciousness clear | 696 | 696 | Factual
rehabilitation in bed | 696 | 1680 | Factual
sepsis due to multidrug-resistant Pseudomonas aeruginosa | 1680 | 1680 | Factual
disseminated intravascular coagulation | 1680 | 1680 | Factual
general condition deteriorated | 1680 | 1680 | Factual
death | 1680 | 1680 | Factual