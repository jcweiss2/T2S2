45 years old | 0
female | 0
American Society of Anesthesiologists Grade I | 0
right sided hemi-arthroplasty | -1304
subcapitate fracture of neck of femur | -1304
infected implant | -728
implant removal | -728
antibiotic coated spacer insertion | -728
wound debridement | -728
regional anesthesia | -1304
perioperative period uneventful | -1304
injection teicoplanin | -24
injection amikacin | -24
raised total leucocyte count | -24
raised erythrocyte sedimentation rate (ESR) | -24
raised C-reactive protein (CRP) | -24
capsule pregabalin 150 mg | -24
capsule pregabalin 150 mg | -2
noninvasive blood pressure 100/70 mmHg | 0
SpO2 99% | 0
coarse AF | 0
heart rate 150-160 beats/min | 0
irregularly irregular rhythm | 0
drowsy | 0
arousable | 0
responding to verbal commands | 0
denied anxiety | 0
denied headache | 0
denied nausea | 0
denied chest pain | 0
denied palpitation | 0
denied difficulty in breathing | 0
defibrillator ready | 0
resuscitative drugs and equipments ready | 0
injection metoprolol | 0
12-lead ECG | 0
cardiology opinion sought | 0
surgery postponed | 0
cardiologist confirmed AF | 0
amiodarone infusion advised | 0
systolic blood pressure above 90 mmHg | 0
intravenous amiodarone 150 mg bolus | 1
amiodarone infusion at 1 mg/min | 1
heart rate reduced to 90/min | 20
systolic blood pressure increased to 120 mmHg | 20
AF reverted to sinus rhythm | 20
arterial blood gas within normal limits | 20
serum electrolytes within normal limits | 20
shifted to intensive care unit (ICU) | 20
troponin T within normal limits | 24
creatine phosphokinase-myoglobin within normal limits | 24
serum electrolytes within normal limits | 24
transthoracic echocardiography within normal limits | 24
amiodarone infusion continued | 24
aspirin 75 mg once daily started | 24
transferred to ward | 48
CRP decreasing trend | 336
right sided hemiarthroplasty | 336
surgery conducted successfully | 336
no perioperative ECG changes | 336