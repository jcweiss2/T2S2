Here is the extracted table of clinical events and timestamps:

pneumonia | -672
SARS-CoV-2 | -672
COVID-19 | -672
fever | -672
cough | -672
fatigue | -672
dyspnea | -672
anorexia | -672
diarrhea | -672
vomiting | -672
abdominal pain | -672
ACE II receptor expression | -672
abdominal imaging | 0
CT scan | 0
abdominal CT | 0
ultrasonography | 0
bowel wall thickening | 0
fluid-filled colon | 0
intestinal distention | 0
mucosal hyperenhancement | 0
peri enteric fat stranding | 0
mesenteric inflammation | 0
vascular engorgement | 0
pneumatosis | 0
portal venous gas | 0
ileus | 0
GI bleeding | 0
abdominal pain | 0
sepsis | 0
nausea | 0
vomiting | 0
abdominal distention | 0
GI perforation | 0
ascites | 0
intussusception | 0
contrast-enhanced CT | 0
ischemic bowel disease | 0
hypercoagulable state | 0
mesenteric ischemia | 0
pneumoperitoneum | 0
acute diverticulitis | 0
ileocolic intussusception | 0
perforated jejunal diverticulitis | 0
periportal edema | 0
hematomas | 0
retroperitoneum | 0
abdominal wall | 0
rectosigmoid | 0
small bowel obstruction | 0
cecal wall thickening | 0
ileocolonic intussusception | 0
MIS-C | 0
appendicitis | 0
Kawasaki-like presentations | 0
mucocutaneous symptoms | 0
non-compressible appendix | 0
dilated appendix | 0
mural hyperemia | 0
periappendiceal mesenteric fat stranding | 0
edema | 0
ascites | 0
thickened terminal ileum | 0
luminal dilatation | 0
wall thickening of the appendix | 0
calcified deposit within the appendix | 0
pelvic free fluid | 0
enlarged lymph nodes | 0
perforation | 0
adjacent small rim-enhancing fluid collections | 0
thromboembolic complications | 0
coagulation dysfunction | 0
endothelial damage | 0
complement proteins | 0
acute stroke | 0
acute myocardial infarction | 0
extracorporeal membrane oxygenation circuit thrombosis | 0
multiple organ failure | 0
death | 0
microvascular involvement | 0
end-organ ischemia | 0
bowel loops | 0
spleen | 0
kidneys | 0
liver infarctions | 0
SMA thrombotic occlusion | 0
intestinal gangrene | 0
dilated ileal loops | 0
non-enhancing barely discernible walls | 0
direct viral infection | 0
small vessel thrombosis | 0
non-occlusive mesenteric ischemia | 0
deep venous thrombosis | 0
acute pulmonary thromboembolism | 0
AMI | 0
CT angiography | 0
emboli | 0
SMA | 0
celiac | 0
inferior mesenteric arteries | 0
intramural bowel gas | 0
absence of bowel wall enhancement | 0
hepatic portal venous gas | 0
ischemia of other organs | 0
SMV thrombosis | 0
filling defect in the SMV | 0
diffuse small bowel wall thickening | 0
mesenteric fat stranding | 0
mesenteric venous congestion | 0
non-occlusive AMI | 0
thrombosis of distal SMA branches | 0
thromboembolic occlusion of SMA | 0
decreased peristalsis | 0
interloop fluid | 0
increased intraluminal contents | 0
stasis | 0
intra-abdominal hemorrhage | 0
extraperitoneal hemorrhage | 0
intramuscular hematomas | 0
iliopsoas | 0
rectus sheath | 0
active bleeding | 0
hyperdense fresh hematoma | 0
vascular abnormalities | 0
fat stranding surrounding the mesenteric vessels | 0
hypoperfused distal SMA1 branches | 0
SMA thrombosis | 0
mesenteric congestion | 0
gas in the transverse mesocolon vasculature | 0
significant filling defect in the superior mesenteric vein | 0
psoas muscle hemorrhage | 0
contrast extravasation | 0
pelvic extraperitoneal hemorrhage | 0
active bleeding | 0
massive right iliopsoas muscle hematoma | 0
extravasation extending to the retroperitoneal area | 0
small low-density area in the left iliopsoas muscle | 0
hematoma | 0
spontaneous iliopsoas muscle hematoma | 0