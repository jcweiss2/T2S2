55 years old | 0
woman | 0
presented with chest pain | -72
presented with palpitations | -72
presented with shortness of breath | -72
presented with nausea | -72
blood pressure of 182/87 mmHg | 0
heart rate of 74 bpm | 0
temperature of 98.3°F | 0
oxygen saturation of 94% | 0
troponin elevation of 0.26 ng/mL | 0
creatinine elevation of 1.5 mg/dL | 0
white blood cell count elevation of 21.6 K/uL | 0
blood glucose elevation of 497 mg/dL | 0
AST elevation of 110 U/L | 0
ALT elevation of 133 U/L | 0
lactic acid elevation of 6.9 mmol/L | 0
pro-BNP elevation of 926 pg/mL | 0
EKG showing ST segment elevations in leads V1 and V2 | 0
CTPA negative for pulmonary embolism | 0
incidental finding of right adrenal mass | 0
admitted to ICU | 0
STEMI | 0
hyperglycemia | 0
sepsis | 0
heparin drip started | 0
metoprolol started | 0
cefepime started | 0
lactated ringers bolus administered | 0
insulin drip started | 0
worsening chest pain | 24
worsening palpitations | 24
troponin rise to 1.00 ng/mL | 24
echocardiogram showing 40-45% ejection fraction | 24
septal hypokinesis | 24
lateral hypokinesis | 24
anteroseptal hypokinesis | 24
posterolateral hypokinesis | 24
cardiac angiography showing normal coronary vessels | 24
myocarditis considered | 24
erythrocyte sedimentation rate of 0 mm/hr | 24
chest pain improvement | 48
oxygen requirement decreased to room air | 48
lactic acid decrease to 2.0 mmol/L | 48
blood glucose decrease to 179 mg/dL | 48
AST improvement to 39 U/L | 48
ALT improvement to 41 U/L | 48
diagnostic work-up for pheochromocytoma | 48
plasma metanephrine elevation of 2.13 nmol/L | 48
normetanephrine elevation of 4.15 nmol/L | 48
doxazosin started | 48
carvedilol started | 48
CT Adrenal showing right adrenal mass | 48
robotic assisted laparoscopic right adrenalectomy | 120
resolution of cardiomyopathy | 2880
cardiomyopathy | 0
pulmonary edema | 0
acute kidney injury | 0
acute liver injury | 0
hyperglycemia without diabetes | 0
elevated lactic acid | 0
normal coronary vessels | 24
unexpected improvement in clinical symptoms | 48
pheochromocytoma diagnosis | 48
