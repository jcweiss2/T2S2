39 years old | 0  
male | 0  
admitted to the hospital | 0  
intermittent fever | -1440  
moderate exertion dyspnoea | -168  
orthopnoea | -24  
systolic murmurs in aortic and pulmonary areas | 0  
high C-reactive protein | 0  
leucocytosis | 0  
neutrophilia | 0  
empiric antibiotic therapy started | 0  
transoesophageal echocardiography | 24  
5 mm vegetation attached to the non-coronary cusp of the aortic valve | 24  
severe aortic regurgitation | 24  
aortic root abscess | 24  
left ventricle-to-right atrium fistula | 24  
blood cultures | 24  
Ceftriaxone started | 48  
surgery | 72  
aortic valve replacement with a biological prosthesis | 72  
closure of the fistula | 72  
worsening of patient's general condition | 360  
computed tomography | 360  
transthoracic echocardiography | 360  
acute mediastinitis | 360  
pericardial abscess | 360  
cardiac tamponade | 360  
emergency surgery | 360  
patient exits intensive care unit after second surgery | 480  
Pericardial abscess culture | 480  
Enterococcus faecalis | 480  
Ampicillin added to therapy | 480  
patient discharged | 912  
36 days of ceftriaxone | 912  
24 days of metronidazole | 912  
19 days of ampicillin | 912  
antibiotic therapy to be finished under outpatient regimen | 912  
occasional smoking | 0  
alcohol consumption | 0  
no lower limb swelling | 0  
no palpitations | 0  
no dizziness | 0  
no syncope | 0  
no weight loss | 0  
no symptoms suggestive of constitutional syndrome | 0  
mild tachypnoea at rest | 0  
temperature of 36.9°C | 0  
blood pressure of 129/40 mmHg | 0  
heart rate of 105 b.p.m. | 0  
blood oxygen saturation 96% | 0  
diastolic murmurs in both aortic and pulmonary areas | 0  
slight crackles in both lung bases | 0  
no skin alterations | 0  
normal oropharyngeal cavity | 0  
abdomen soft and depressible | 0  
no pain on palpation | 0  
no masses | 0  
no megalia | 0  
no oedema in the lower limbs | 0  
anaemia | 0  
haemoglobin 10.8 g/dL | 0  
no significant electrocardiogram findings | 0  
mild bilateral pleural effusion | 0  
right basal atelectasis | 0  
admitted to Internal Medicine department | 0  
unknown origin fever | 0  
first episode of heart failure | 0  
suspicion of infective endocarditis | 0  
blood cultures extracted | 0  
piperacillin-tazobactam started | 0  
transthoracic echocardiography | 0  
moderately dilated left ventricle | 0  
biplane end-diastolic volume 252 mL | 0  
preserved ejection fraction 62% | 0  
normal size right atrium and right ventricle | 0  
normal right ventricle function | 0  
tricuspid annular plane systolic excursion 24 mm | 0  
tricuspid annulus S' wave 14 cm/s | 0  
mild tricuspid regurgitation | 0  
peak velocity 297 cm/s | 0  
estimated systolic pulmonary artery pressure 40 mmHg | 0  
severe aortic regurgitation | 0  
wide central jet exceeding anterior mitral valve plane | 0  
pressure half-time 117 ms | 0  
vegetation in non-coronary cusp of aortic valve | 0  
aortic root pseudoaneurysm | 0  
left ventricle-to-right atrium fistula | 0  
transoesophageal echocardiography confirmed 5 mm vegetation | 24  
18 x 7 mm periannular pseudoaneurysm | 24  
subaortic left ventricle-to-right atrium fistula | 24  
Gerbode defect | 24  
Gram-negative bacilli in blood cultures | 24  
identified as C. canimorsus | 24  
dog bite 4 months earlier | -2880  
owned a pet dog | 0  
antibiotic therapy switched to ceftriaxone | 48  
metronidazole added | 336  
persistent fever | 336  
sensitivity to metronidazole demonstrated | 336  
urgent surgical treatment decided | 72  
10 mm defect next to non-coronary cusp | 72  
aortic root diameter 18 mm | 72  
aortic root enlargement via Nicks procedure | 72  
bovine pericardial patch used for aortic defect | 72  
fistula repaired with bovine pericardial patch | 72  
native aortic valve replaced | 72  
significant bleeding detected | 72  
revision and reinforcement of sutures | 72  
admission to intensive care unit | 72  
post-operative echocardiogram normal function | 72  
persistence of left ventricle-to-right atrium fistula | 72  
dehiscence of pericardial patch | 72  
peak velocity 4.7 m/s | 72  
peak gradient 89 mmHg | 72  
Qp/Qs ratio 1.2 | 72  
post-operative day +12 worsening | 360  
low-grade fever | 360  
profuse sweating | 360  
purulent secretion in pacemaker leads | 360  
thoracic computed tomography | 360  
acute mediastinitis | 360  
pericardial abscess | 360  
cardiac tamponade | 360  
emergency surgery | 360  
Enterococcus faecalis in culture | 480  
ampicillin added | 480  
progressive clinical improvement | 480  
resolution of mediastinitis | 480  
no residual pericardial effusion | 480  
discharged with oral antibiotics | 912  
metronidazole continued | 912  
linezolid started | 912  
subsequent check-ups showed improvement | 912  
no fever | 912  
no heart failure symptoms | 912  
normal physical activity | 912  