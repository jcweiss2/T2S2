47 years old | 0
female | 0
admitted to the hospital | 0
skin ecchymosis | 0
vaginal bleeding | 0
WBC count 7.91×10^9/l | 0
hemoglobin 84 g/l | 0
platelet count 14×10^9/l | 0
prothrombin time 16.9 s | 0
activated partial thromboplastin time 40.7 s | 0
fibrinogen level 1.66 g/l | 0
d-dimer level 20 μg/mL | 0
bone marrow smear showed hypercellularity | 0
abnormal promyelocytic granulocytes 96.5% | 0
Auer bodies observed | 0
peroxidase staining positive | 0
immunophenotype analysis showed positivity for myeloperoxidase | 0
immunophenotype analysis showed positivity for CD13 | 0
immunophenotype analysis showed positivity for CD33 | 0
immunophenotype analysis showed positivity for human leukocyte antigen-DR | 0
immunophenotype analysis showed positivity for CD56 | 0
treated with ATRA | 0
treated with ATO | 0
chest tightness | 14
dyspnea | 14
systemic edema | 14
pleural effusion | 14
differentiation syndrome | 14
WBC count 9.4×10^9/l | 14
hemoglobin 59 g/l | 14
platelet count 38×10^9/l | 14
prothrombin time 18.3 s | 14
fibrinogen level 0.91 g/l | 14
d-dimer level 20 μg/mL | 14
karyotype 45, X, –X, del(9)(q13q22), t(11;12)(p15;q13) | 14
PML–RARA fusion transcript negative | 14
mutations detected in IDH2 | 14
mutations detected in TET2 | 14
mutations detected in ASXL1 | 14
mutations detected in TP53 | 14
mutations detected in WT1-exon7 | 14
mutations detected in WT1-exon9 | 14
treatment with ATRA and ATO discontinued | 14
diuretic detumescence | 14
ventilator-assisted respiratory therapy | 14
second bone marrow smear showed 95.5% abnormal promyelocytic granulocytes | 20
Auer body in the form of an Auer bundle | 20
peroxidase staining positive rate 100% | 20
treated with idarubicin | 20
treated with cytarabine | 20
severe pulmonary infection | 27
antibiotics | 27
WBC and platelet counts remained low | 27
third bone marrow smear showed 10.5% blasts | 34
treated with homoharringtonine | 34
treated with idarubicin | 34
treated with cytarabine | 34
treated with GCSF | 34
bone marrow examination showed 0.5% blasts | 41
complete remission | 41
consolidation therapy with HIAG regimen | 41
severe pulmonary infection | 41
septic shock | 41
metabolic acidosis | 41
heart failure | 41
admitted to intensive care unit | 41
recovered after 1 month | 71
refused allogeneic hematopoietic stem cell transplantation | 71
received CAG regimen | 71
received HA regimen | 71
minimal residual disease detected by flow cytometry negative | 71
alive and leukemia-free at 24-month follow-up | 720
NUP98–RARG fusion gene detected | -672
RT-PCR analysis | 0
FISH analysis | 0
cytogenetic analysis | 0
fluorescence in situ hybridization | 0