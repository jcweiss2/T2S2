50 years old | 0
woman | 0
presented to the hospital | 0
abdominal pain for 10 days | -240
mild abdominal pain | -240
colicky abdominal pain | -240
right flank pain | -240
nausea | -240
vomiting | -240
pain worsened | 0
collapsed while walking | 0
transferred to the hospital | 0
acute surgical abdomen | 0
CT scan revealed enhanced oedematous appendiceal wall | 0
retroperitoneal subhepatic air | 0
mild collection indicative of perforated subhepatic appendix | 0
diagnosed with acute abdomen | 0
perforated appendix | 0
peritonitis | 0
sepsis | 0
underwent urgent laparotomy | 0
pus evacuated | 0
retrocecal appendix | 0
subhepatic appendix | 0
retrograde appendectomy | 0
culture and sensitivity swabs taken | 0
abdomen washed extensively | 0
suction drains secured to the right abdomen | 0
surgery not complicated | 0
admitted to surgical intensive care unit | 0
managed accordingly | 0
estimate of recovery and discharge within 10 days | 0
treated with antimicrobials based on culture and sensitivity report | 0
did not improve as expected | 0
drains continued to drain 200 ml pus daily | 0
appropriate antimicrobial coverage | 0
developed respiratory distress | 0
intubated | 0
mechanically ventilated | 0
second abdominal CT scan | 0
ill-defined retroperitoneal collection on right side | 0
two pockets of retroperitoneal collection | 0
first pocket under abdominal muscles and peripherally | 0
second pocket anterior to Gerota's fascia of right kidney |
