74 years old | 0
    male | 0
    admitted to the hospital | 0
    obstructive sleep apnea | 0
    interstitial lung disease | 0
    morbid obesity | 0
    hypertension | 0
    atrial fibrillation | 0
    diabetes mellitus | 0
    epigastric abdominal pain | -24
    chest pain | -24
    progressive abdominal distension | -24
    poor appetite | -24
    nausea | -24
    belching | -24
    constipation | -24
    cardiac workup negative for acute coronary syndrome | -24
    computed tomography abdomen and pelvis | -24
    moderate colonic stool | -24
    enlarged pelvic lymph nodes | -24
    enlarged mediastinal lymph nodes | -24
    enlarged retroperitoneal lymph nodes | -24
    mild increase in lymph node size since 2018 | -24
    bronchoscopy | -2016
    fine-needle aspiration of level 7 lymph node | -2016
    flow cytometry analysis | -2016
    no specific pathology | -2016
    laboratory examination unremarkable | -24
    discharged | -24
    aggressive bowel regimen | -24
    emergency department presentation | -24
    no improvement in pain | 0
    worsening abdominal distension | 0
    baseline oxygen use | 0
    normal vital signs | 0
    soft abdomen | 0
    mildly distended abdomen | 0
    non-tender abdomen | 0
    no rebound tenderness | 0
    no guarding | 0
    admission laboratory values | 0
    repeat CT chest | 0
    repeat CT abdomen | 0
    repeat CT pelvis | 0
    chest adenopathy | 0
    abdominal adenopathy | 0
    pelvic adenopathy | 0
    aortoiliac atherosclerotic disease | 0
    right upper-quadrant ultrasound | 0
    heterogeneous hepatic parenchyma | 0
    coarsened echotexture of hepatic parenchyma | 0
    no biliary tree disease | 0
    no gallbladder disease | 0
    concern for acute mesenteric ischemia | 0
    CT angiography abdomen | 0
    extensive atherosclerosis of superior mesenteric artery | 0
    moderate stenosis at ostium | 0
    endoscopy | 0
    non-obstructing Schatzki ring | 0
    gastric ulcer | 0
    oozing hemorrhage | 0
    bipolar cautery | 0
    serum immunofixation | 0
    M spike 0.2 g/dL | 0
    polyclonal gammopathy | 0
    IgM kappa | 0
    quantitative IgM 233 mg/dL | 0
    normal free light chain ratio | 0
    flow cytometry peripheral blood | 0
    no increased blast proliferation | 0
    no lymphoproliferative disease | 0
    declined bone marrow biopsy | 0
    worsening abdominal pain | 192
    altered mental status | 192
    asterixis | 192
    afebrile | 192
    normal vitals | 192
    oxygen saturation 94% | 192
    white blood cell count 16.4×109/L | 192
    platelets 89×109/L | 192
    ALT 101 U/L | 192
    AST 328 U/L | 192
    lactic acid 4.2 mmol/L | 192
    total bilirubin 2.5 mg/dL | 192
    direct bilirubin 1.9 mg/dL | 192
    INR 6.35 | 192
    ammonia level 117 µmol/L | 192
    repeat CT abdomen and pelvis | 192
    no acute findings | 192
    worsening abdominal pain | 192
    encephalopathy | 192
    elevated transaminases | 192
    lactic acidosis | 192
    coagulopathy | 192
    transferred to PCU | 192
    acute liver failure | 192
    IV N-acetylcysteine | 192
    lactulose | 192
    IV vitamin K | 192
    acute encephalopathy | 192
    CT head | 192
    no acute abnormalities | 192
    EEG diffuse slowing | 192
    serology negative for HAV | 192
    serology negative for HBV | 192
    serology negative for HCV | 192
    serology negative for HIV | 192
    serology negative for EBV | 192
    serology negative for CMV | 192
    tick panel negative | 192
    anti-smooth muscle antibodies negative | 192
    continued clinical worsening | 192
    respiratory status decompensation | 192
    CXR bilateral ground-glass opacities | 192
    concern for pneumonia | 192
    broad-spectrum antibiotics | 192
    lethargy | 216
    tachypnea | 216
    ABG pH 7.46 | 216
    ABG pCO2 34 mmHg | 216
    ABG HCO3 24 mEq/L | 216
    BiPAP | 216
    ICU admission | 240
    unresponsive | 240
    comatose | 240
    hypotensive | 240
    worsening septic shock markers | 240
    lactic acidosis 7.3 mmol/L | 240
    total bilirubin 7.9 mg/dL | 240
    direct bilirubin 5.3 mg/dL | 240
    ALT 174 U/L | 240
    AST 396 U/L | 240
    hemoglobin 6.6 g/dL | 240
    thrombocytopenia 29×109/L | 240
    INR 7.04 | 240
    intubation | 240
    gram-negative bacteremia | 240
    septic shock | 240
    IV fluids | 240
    vasopressors | 240
    ventricular tachycardia | 240
    defibrillation | 240
    atrial fibrillation with rapid ventricular response | 240
    ARDS | 240
    continued deterioration | 240
    comfort care | 240
    palliative extubation | 240
    death | 336
    autopsy diffuse large B-cell lymphoma | 336
    liver involvement | 336
    lung involvement | 336
    bone marrow involvement | 336
    lymph node involvement | 336
    extensive lymphadenopathy | 336
    right cervical lymphadenopathy | 336
    peri-bronchial lymphadenopathy | 336
    subcarinal lymphadenopathy | 336
    pelvic lymphadenopathy | 336
    large hilar mass | 336
    matted lymph nodes | 336
    enlarged liver | 336
    pale-yellow nodules | 336
    infiltration of atypical lymphoid cells | 336
    CD20 positive | 336
    CD10 positive | 336
    BCL-2 positive | 336
    cyclin D1 negative | 336
    CD5 negative | 336
    CD138 negative | 336
    MUM1 negative | 336
    CD21 negative | 336
    CD3 negative | 336
    BCL6 negative | 336
    hepatic necrosis | 336
    nodular infiltrate | 336
    diffuse infiltrate | 336
    bone marrow involvement >90% | 336
    acute liver failure | 192
    transaminitis | 192
    jaundice | 192
    abnormal coagulation profile | 192
    INR >1.5 | 192
    hepatic encephalopathy | 192
    persistent lymphadenopathy | 192
    refused bone marrow biopsy | 192
    gram-negative bacteremia | 240
    septic shock | 240
    ventricular tachycardia | 240
    ARDS | 240
    comfort care | 240
    palliative extubation | 240
    death | 336
    autopsy findings | 336
    acute liver failure due to DLBCL | 336
    <|eot_id|>
    