48 years old | 0
male | 0
admitted to the Emergency Department (ED) | 0
chest pain | 0
shortness of breath | 0
stabilized in the ED | 0
transferred to the intermediate general ward | 0
drug optimization | 0
hemodialysis | 0
coronary angiography | 0
3-vessel CAD (3VD) | 0
61% ejection fraction (EF) | 0
body mass index 28.7 kg/m2 (overweight) | 0
history of CKD | 0
stroke | 0
angina | 0
diabetes | 0
dyslipidemia | 0
smoking | 0
scheduled for urgent CABG surgery | 0
anemia (8.4 g/dL) | 0
leukocytosis (11,100/µL) | 0
increased cardiac enzymes | 0
CKMB (30 U/L) | 0
decreased pCO2 (27.9 mmHg) | 0
increased pO2 (170.5 mmHg) | 0
decreased HCO3 (19.6 mmol/L) | 0
thorax X-ray showed cardiomegaly | 0
normal appearance of both lungs before surgery | 0
CABG surgery | 192
LIMA-LAD | 192
SVG-OM1 | 192
SVG-PDA | 192
transferred to the Intensive Care Unit (ICU) | 192
extubated | 212
treated in the ICU for 21 hours | 192
transferred to the intermediate ward | 216
transferred to the ward | 336
increased difficulty in breathing | 432
decreased saturation | 432
low PO2 | 432
fever | 432
transferred to the isolation ICU room | 432
reintubated | 432
COVID-19 RT-PCR test | 432
positive for COVID-19 | 432
neutrophil-to-lymphocyte ratio (NLR) 14.03 | 312
thorax X-rays showed consolidation of both lungs | 216
pneumonia | 216
hemodynamically unstable due to sepsis | 432
deterioration of urea and creatinine levels | 432
considered for continuous renal replacement therapy (CRRT) | 432
respiratory failure | 528
pO2 low | 528
saturation low | 528
high fiO2 | 528
died | 528
respiratory distress caused by COVID-19 infection | 528
