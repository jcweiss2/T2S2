58 years old | 0
female | 0
history of Hodgkin lymphoma | 0
status post radiation therapy | 0
hypertension | 0
diabetes mellitus | 0
hypothyroidism | 0
dyspnea on exertion | -336
metformin | 0
aspirin | 0
levothyroxine | 0
metoprolol | 0
blood pressure 96/60 mmHg | 0
heart rate 110 beats per minute | 0
oxygen saturation 96% | 0
elevated jugular venous pressure | 0
faint and distant heart sounds | 0
weak peripheral pulses | 0
low voltage on 12-lead electrocardiogram | 0
sinus tachycardia | 0
cardiomegaly on chest X-ray | 0
large circumferential pericardial effusion | 0
end diastolic right ventricular compression | 0
swing sign | 0
left ventricular ejection fraction 60%-65% | 0
pericardiocentesis | 0
rapid drainage of 2200 mL of serous fluid | 1
minimal improvement in hemodynamics | 1
worsening dyspnea | 1
hypotension | 1
labored breathing | 1
pulmonary edema | 1
intubation | 1
hemodynamic support with dobutamine and norepinephrine | 1
low-normal left ventricular ejection fraction | 1
mild to moderately dilated right ventricle | 1
mild right ventricular hypokinesis | 1
septal shift towards the left ventricle | 1
intravenous saline bolus | 1
hemodynamic support with intravenous vasopressors | 1
inotropes | 1
diuresed with intravenous lasix | 2
vasopressor-inotropic support weaned off | 48
CT-chest angiography | 48
no evidence of pulmonary embolism | 48
improvement in pulmonary edema | 48
extubation | 72
normalized ventricular function | 120
trivial/minimal pericardial effusion | 120
discharged | 144