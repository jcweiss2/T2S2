55 years old | 0
    man | 0
    nonalcoholic steatohepatitis | -15120
    alpha 1 antitrypsin deficiency | -15120
    orthotopic liver transplant | -15120
    incarcerated inguinal hernia | -15120
    repaired inguinal hernia | -15120
    cytomegalovirus viremia | -15120
    treated with valganciclovir | -15120
    discharged | -15120
    maintenance immunosuppression | -15120
    mycophenolate mofetil | -15120
    tacrolimus | -15120
    prednisone | -15120
    presented 5 weeks post-transplant | 0
    encephalopathy | -48
    increasing home oxygen requirements | -48
    arrival | 0
    required 4L nasal cannula | 0
    maintain oxygen saturation >92% | 0
    encephalopathy characterized by sparse speech | 0
    encephalopathy characterized by disorientation | 0
    nonfocal neurologic examination | 0
    vital signs within normal limits | 0
    physical examination within normal limits | 0
    white blood cell count 9.3 × 109/L | 0
    creatinine 2.12 mg/dL | 0
    blood urea nitrogen 53 mg/dL | 0
    synthetic liver function within normal limits | 0
    international normalized ratio within normal limits | 0
    alanine aminotransferase within normal limits | 0
    aspartate aminotransferase within normal limits | 0
    bilirubin within normal limits | 0
    arterial ammonia 204 µmol/L | 0
    intensive care unit admission | 0
    induction dosing of intravenous ganciclovir | 0
    elevated CMV titers | 0
    started on empiric antibiotic coverage | 0
    vancomycin | 0
    meropenem | 0
    micafungin | 0
    blood cultures drawn | 0
    intravenous micronutrient supplementation | 0
    B1 | 0
    B6 | 0
    levocarnitine | 0
    lumbar puncture | 0
    opening pressure 8 cmH2O | 0
    Gram stain revealed encapsulated yeast | 0
    suspicious for Cryptococcus | 0
    started on liposomal amphotericin B | 0
    flucytosine | 0
    hyperammonemia | 0
    started on continuous renal replacement therapy | 0
    rifaximin | 0
    zinc | 0
    lactulose | 0
    ammonia climbed to 692 µmol/L | 24
    neurological deterioration | 24
    mechanical ventilation | 24
    empiric intravenous doxycycline | 24
    urine obtained for Mycoplasma PCR | 24
    bronchial aspirate obtained for Mycoplasma PCR | 24
    urine obtained for Ureaplasma PCR | 24
    bronchial aspirate obtained for Ureaplasma PCR | 24
    48 hours after antifungal induction | 48
    48 hours after CRRT | 48
    ammonia levels <100 µmol/L | 48
    Cryptococcal serum antigen positive | 48
    cerebrospinal fluid antigen positive | 48
    cultures from bronchoalveolar lavage revealed cryptococcal growth | 48
    CSF cultures revealed cryptococcal growth | 48
    blood cultures revealed cryptococcal growth | 48
    disseminated disease | 48
    repeat lumbar punctures | 72
    opening pressures >45 cmH2O | 72
    large volume drainage every 48 hours | 72
    permanent CSF diversion not possible | 72
    persistent thrombocytopenia | 72
    thrombocytopenia nadir 16 × 103/µL | 72
    mental status transiently improved | 72
    unable to wean from mechanical ventilation | 72
    tracheostomy | 72
    continued complications of cryptococcal infection | 120
    sludging | 120
    obstruction of microvascular structures | 120
    persistent hydrocephalus | 120
    oliguric renal failure | 120
    progressive splenic infarcts | 120
    necrosis requiring splenectomy | 120
    magnetic resonance imaging of the brain | 120
    no cytotoxic edema | 120
    rapid correction of ammonia levels | 120
    hospital course complicated by sepsis | 120
    duodenal leak | 120
    persisting renal failure | 120
    failure to thrive | 120
    poor quality of life | 120
    multiple unresolved end-organ problems | 120
    family decided on comfort care in hospice | 120
    urea cycle disorder screening studies | 120
    low urine orotic level | 120
    normal serum citrulline | 120
    normal serum arginine | 120
    urea cycle disorder unlikely | 120
    