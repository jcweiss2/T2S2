22 years old | 0
female | 0
admitted to hospital | 0
headache | -48
neck pain | -48
vomiting | -48
diarrhea | -48
abdominal pain | -48
photophobia | -48
malaise | -48
tachycardic | 0
pyrexial | 0
normal blood pressure | 0
suspected meningitis | 0
treated with ceftriaxone | 0
treated with acyclovir | 0
CSF sampling | 0
CSF sampling unremarkable | 0
managed on the ward | 0
deteriorated on Day 3 | 72
persistent fever | 72
severe hypoxia | 72
lactatemia | 72
hypotension | 72
unresponsive to IV fluids | 72
admitted to ITU | 72
high-flow nasal oxygen | 72
vasopressors | 72
intubated | 72
ventilated | 72
multisystem failure | 90
hypotension | 90
hypoxia | 90
azotemia | 90
oliguria | 90
nonabsorption of feeds | 90
diarrhea | 90
focused intensive care echocardiogram | 90
poorly contracting right and left ventricles | 90
dobutamine | 90
renal dysfunction | 90
severe metabolic acidosis | 90
hemofiltration | 90
CT chest/abdomen | 90
multiple enlarged mesenteric lymph nodes | 90
diagnostic laparoscopy | 108
multiple mesenteric lymph node enlargement | 108
minimal ascites | 108
small left ovarian cyst | 108
lymph node biopsy | 108
ascitic sampling | 108
no source of sepsis | 108
broad-spectrum antibiotics | 108
ciprofloxacin | 108
vancomycin | 108
meropenem | 108
no clinical improvement | 108
MIS-A diagnosis | 108
IV immunoglobulin | 108
methylprednisolone | 108
rapid improvement | 144
resolution of hyperpyrexia | 144
cardiovascular instability | 144
decreasing oxygen requirements | 144
extubated | 168
normal ventricular function | 168
discharged | 312
raised white cell count | 0
CRP | 0
clear CSF | 0
no cells in CSF | 0
no organisms in CSF | 0
normal chest X-ray | 0
normal CT head | 0
mesenteric lymphadenopathy | 72
negative microbiology | 0
negative virology | 0
negative vasculitis | 0
negative autoimmune screen | 0
biventricular dysfunction | 0
resolved biventricular dysfunction | 168
lymph node biopsy | 108
marked suppurative inflammation | 108
acute vasculitic changes | 108
negative SARS-CoV-2 PCR | 0
positive COVID-19 antibodies | 0
mildly elevated ferritin | 0
no hypofibrinogenemia | 0
no cytopenias | 0