35-year-old pregnant woman | 0
    34 + 4 wk pregnancy | 0
    fever | -240
    cough | -240
    aggravated dyspnoea | -120
    admitted to the hospital | 0
    body temperature of 36.4 ℃ | 0
    blood pressure of 117/87 mmHg | 0
    heart rate of 130 beats/min | 0
    respiratory rate of 20 times/min | 0
    cyanosis of the lip | 0
    thick breathing sounds in both lungs | 0
    dry and wet rales in the right lower lung | 0
    gestational and symmetric abdominal type | 0
    height of 166 cm | 0
    pre-pregnancy weight of 46.5 kg | 0
    body mass index of 16.87 | 0
    weight gain of 8.8 kg during pregnancy | 0
    uterine height was 34 cm | 0
    abdominal circumference was 89 cm | 0
    sporadic and weak contractions | 0
    head presentation | 0
    foetal heart sounds of 142 beats/min | 0
    normal intrapelvic and extrapelvic measurements | 0
    arterial blood gas pH 7.472 | 0
    partial pressure of carbon dioxide 34.0 mmHg | 0
    partial pressure of oxygen 56 mmHg | 0
    sulfur dioxide 88.6% | 0
    C-reactive protein 186.33 mg/L | 0
    erythrocyte sedimentation rate 69.00 mm/h | 0
    procalcitonin 2.24 ng/mL |: 0
    white blood cell 18.29 × 109/L | 0
    neutrophil 90.10% | 0
    lymphocyte 0.97 × 109/L | 0
    alkaline phosphatase 232 U/L | 0
    total bilirubin 23.1 μmol/L | 0
    albumin 33.9 g/L | 0
    K+ 2.93 mmol/L | 0
    sodium 129 mmol/L | 0
    chloride 89 mmol/L | 0
    normal cardiac markers | 0
    D-dimer 3.50 mg/L | 0
    chest CT multiple plaques | 0
    miliary foci | 0
    nodular foci with partial consolidation and cavities | 0
    obstetric ultrasound single viable foetus | 0
    head presentation | 0
    oligohydramnios | 0
    no significant cardiac ultrasound findings | 0
    no significant lower extremity vascular ultrasound findings | 0
    first menarche at 15 years | 0
    menstrual cycle regular every 30 d | 0
    menstruation lasting 3-4 d | 0
    last menstruation on May 2, 2022 | 0
    moderate menstrual volume | 0
    normal menstrual color | 0
    no blood clots | 0
    no painful menstruation | 0
    married at appropriate age | 0
    healthy spouse | 0
    G2P1 | 0
    full-term normal delivery in 2006 | 0
    female infant weighing 3500 g | 0
    good health of infant | 0
    pregnancy combined with severe pneumonia | 0
    novel coronavirus infection | 0
    S. aureus infection | 0
    respiratory failure | 0
    late pregnancy 34 + 4 wk G2P1 left occiput anterior | 0
    elderly second parturient women | 0
    maternal lower weight | 0
    oligohydramnion | 0
    premature live baby | 0
    electrolyte disturbance | 0
    hypoproteinaemia | 0
    cefoperazone sodium and sulbactam sodium treatment | 0
    dexamethasone 10 mg | 0
    oxyhemoglobin saturation decline | 0
    foetal heart sounds 146 beats/min | 0
    caesarean section of the lower uterus | 0
    high-flow nasal cannula oxygen therapy | 0
    fraction of inspired oxygen 100% | 0
    flow rate 50 L/min | 0
    cyanosis improvement | 0
    oxyhemoglobin saturation 95%-98% | 0
    oxyhemoglobin saturation measured on 2nd day | 48
    foetus transferred to neonatal ICU | 0
    puerperant woman transferred to respiratory ICU | 0
    assisted ventilation by endotracheal intubation | 0
    empirical antibiotic therapy | 0
    meropenem | 0
    vancomycin | 0
    fluid infusion | 0
    albumin infusion | 0
    tracheoscopy irrigation solution tested with mNGS | 0
    S. aureus detection | 0
    novel coronavirus detection | 0
    no acid-fast bacilli in sputum | 0
    TB-PCR negative | 0
    nontuberculosis mycobacterium-PCR negative | 0
    normal galactomannan experiments | 0
    continued vancomycin 1 g q12h | 0
    meropenem 1 g q8h | 0
    anticoagulant therapy | 0
    cough relief treatment | 0
    sputum reduction treatment | 0
    transition to nasal tube oxygen on 2nd day | 48
    flow rate 3-4 L/min | 48
    chest CT on 4th day post-surgery | 96
    multiple areas of inflammation in both lungs | 96
    mildly enlarged mediastinal lymph nodes | 96
    small amount of bilateral pleural effusion | 96
    CRP 38.54 mg/L | 96
    WBC 8.25 × 109/L | 96
    PCT 0.129 ng/mL | 96
    potassium 4.04 mmol/L | 96
    D-dimer 2.44 mg/L | 96
    TB-PCR negative | 96
    chest CT on 9th day post-surgery | 216
    inflammatory lesions | 216
    absorbed pleural effusion | 216
    antibiotics adjusted to sitafloxacin 50 mg twice daily | 216
    stable condition on 11th day post-surgery | 264
    discharged from hospital | 264
    chest CT one week post-discharge | 432
    multiple lung inflammation absorbed slightly | 432
    chest CT one month post-discharge | 720
    multiple lung inflammation apparently absorbed | 720
    S. aureus sequence number 43700 | 0
    S. aureus coverage 93.1785% | 0
    2019-nCoV sequence number 10 | 0
    2019-nCoV coverage 5.8690% | 0
    S. aureus resistant to macrolides and lincosamides | 0
    chest CT inflammatory lesions improved | 216
    <|eot_id|>
    