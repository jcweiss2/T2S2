48 years old | 0
    male | 0
    referred to urology by renal physicians | 0
    possible Fournier's gangrene | 0
    necrotic lesion on glans penis | 0
    broad spectrum antibiotics for sepsis | 0
    infected calciphylaxis-related ulcer on thigh | 0
    no suprapubic pain | 0
    clinical anuria | 0
    increasing bladder volumes on ultrasound | 0
    UTI posited as alternative sepsis source | 0
    infrequent urinary incontinence | -24
    end-stage renal failure (ESRF) | 0
    transitioned from peritoneal dialysis to haemodialysis | -2928
    calciphylaxis | -2928
    type 2 diabetes | 0
    previous cerebrovascular accident due to AF | 0
    palpable bladder | 0
    tender necrotic lesion over glans tip | 0
    involvement of urethral meatus | 0
    penile shaft oedema | 0
    ultrasound showing 400ml urine | -336
    bladder scan showing 600ml | 0
    ultrasound-guided bladder aspiration | 0
    continued medical treatment for infected ulcers | 0
    protracted admission | 24
    slow resolution of infected ulcer | 24
    physical deconditioning | 24
    further bladder aspiration 3 months later | 2160
    1300mL urine drained | 2160
    stable glans lesion at 3 months | 2160
    stable glans lesion at 5 months | 3600
    no urethral voiding | 0
    discharged to nursing home | 3600
    increasing physical care needs | 3600
    urinary retention | 0
    meatal obstruction | 0
    penile calciphylaxis | 0
    risk of complications from indwelling suprapubic catheter | 0
    anticipated need for aspiration | 0
    plan to review in 4 months | 2880
    calciphylaxis diagnosis | 0
    ESRF | 0
    hyperphosphataemia | 0
    hypercalcaemia | 0
    hyperparathyroidism | 0
    vitamin K deficiency | 0
    diabetes mellitus | 0
    wound care | 0
    analgesia | 0
    infection prevention | 0
    serum vitamin D regulation | 0
    calcium regulation | 0
    phosphate regulation | 0
    diet modification | 0
    calcium chelating agents | 0
    phosphate chelating agents | 0
    Cinacalcet use | 0
    sodium thiosulfate with haemodialysis | 0
    surgical intervention consideration | 0
    intractable pain | 0
    unresolving infection | 0
    progressive gangrene | 0
    debridement | 0
    partial penectomy | 0
    total penectomy | 0
    urinary diversion | 0
    parathyroidectomy consideration | 0
    sepsis due to UTI | 0
    catheter-associated UTI risk | 0
    aspiration on triannual basis | 0
    life expectancy less than one year | 0
    sepsis mortality risk | 0
    sterile ultrasound-guided aspiration | 0
    informed consent obtained | 0
    funding declaration | 0
    author contributions | 0
    declaration of competing interests | 0