69 years old| 0
male | 0
admitted to the hospital | 0
worsening abdominal pain | -48
nausea | -48
atrial fibrillation | 0
diabetes | 0
chronic kidney disease | 0
left thoracotomy for lung cancer resection | 0
presented to a urology clinic | -336
micropenis | -336
microhematuria | -336
cystoscopy | -336
negative cystoscopy | -336
CT scan | -336
left perinephric mass | -336
enlarged peri-renal lymph nodes | -336
enlarged para-aortic lymph nodes | -336
retroperitoneal streaky changes | -336
CT-guided peri-renal lesion biopsy | -336
atypical cellular proliferation | -336
no clear pathological diagnosis | -336
elected surveillance | -336
hospital admission | 0
increasing abdominal pain | 0
tachycardia | 0
distended abdomen | 0
tender abdomen | 0
positive fluid wave | 0
no rebound tenderness | 0
no guarding | 0
clean biopsy site | 0
no evidence of hematoma | 0
leukocytosis | 0
normal hematological profile | 0
normal biochemical profile | 0
normal coagulation profile | 0
ascites | 0
ultrasound-guided paracentesis | 0
extracted 6 L bloody fluid | 0
CT imaging | 0
concern for urine extravasation | 0
fluid analysis not consistent with urinary ascites | 0
SAAG <1.1 g/dL | 0
paracentesis | 72
extracted 8 L bloody fluid | 72
cytology negative for malignant cells | 72
consulted Urology | 0
retrograde pyelogram | 0
extravasation at proximal ureter | 0
left ureteral stent | 0
left nephrostomy tube | 0
discharged home | 0
readmitted | 24
syncopal event | 24
painful abdominal distention | 24
ascites requiring frequent paracenteses | 24
withdrew 23 L hemorrhagic ascites | 24
consulted Surgical Oncology | 24
malignancy workup | 24
negative tumor markers | 24
AFP negative | 24
CEA negative | 24
CA 19-9 negative | 24
diagnostic laparoscopy | 24
purplish discoloration of omentum | 24
thickening of omentum | 24
inflammatory reaction on parietal peritoneum | 24
viable small bowel | 24
no evidence of enteric leakage | 24
biopsy of omentum | 24
frozen section analysis | 24
atypical cellular proliferation | 24
extensive areas of necrosis | 24
aspirated 12 L bloody peritoneal fluid | 24
systemic inflammatory response | 24
intensive care unit admission | 24
exploratory laparotomy | 48
omentectomy | 48
continued sepsis | 48
ongoing tissue necrosis | 48
normal liver | 48
normal gallbladder | 48
normal pancreas | 48
serositis of small bowel | 48
no necrosis in small bowel | 48
necrotic greater omentum | 48
purplish discoloration of greater omentum | 48
resected greater omentum | 48
retroperitoneal peri-renal mass | 48
involving Gerota’s fascia | 48
normal kidney | 48
aspirated 9 L bloody ascites fluid | 48
high-grade angiosarcoma | 48
not candidate for palliative chemotherapy | 48
clinical status decline | 48
died | 168
