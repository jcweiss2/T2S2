19 years old | 0
male | 0
admitted to the hospital | 0
trauma | 0
shock state | 0
motor vehicle accident | -72
resuscitation | -24
crystalloid infusion | -24
intra-abdominal complications ruled out | -24
bilateral epidural hematoma | 0
tachycardic | 0
blood pressure 110/65 mmHg | 0
premedication with fentanyl | 0
anesthesia induction with sevoflurane | 0
endotracheal tube placement | 0
cisatracurium use | 0
cranial decompressive surgery | 24
large intravenous lines malfunctioning | 24
preparation of large bore peripheral IV line | 24
failed trials | 24
hemodynamically unstable | 24
femoral artery pulsation not palpable | 24
femoral vein catheterization decision | 24
introducer catheter insertion | 24
central vein catheterization | 24
aspiration of catheter lumens | 24
retrograde flow confirmation | 24
catheter fixation | 24
packed RBCs infusion | 48
crystalloid infusion | 48
norepinephrine infusion | 48
blood loss | 48
transfer to ICU | 72
intubated | 72
stable hemodynamic status | 72
abdominal distension | 96
ultrasound findings of fluid | 96
laparotomy | 96
femoral catheter misplacement | 96
catheter extraction | 96
right inguinal hernia | 96
retroperitoneal fluid | 96
no intestinal perforation | 96
iliac vein perforation bleeding | 96
