60 years old | 0
male | 0
hypothyroidism | -672
alcohol abuse | -672
admitted to the hospital | 0
unresponsive | 0
subacute cognitive decline | -720
sepsis | 0
aspiration pneumonia | 0
opioid and benzodiazepine overdose | 0
acute respiratory failure | 0
intubation | 0
ICU | 0
rehabilitation | 96
discharged home | 168
behavioral changes | 168
re-admitted to the hospital | 192
progressive neuropsychiatric decline | 192
decrease in awareness | 192
decrease in engagement | 192
near akinetic mutism | 192
extensive workup | 192
laboratory testing | 192
paraneoplastic panel | 192
lumbar puncture | 192
CT of the head | 192
MRI of the brain | 192
MRA of the head and neck | 192
cerebral angiogram | 192
T2-weighted image hyperintensities | 192
elevated protein | 192
EEG | 192
lacosamide | 192
IVMP | 192
transferred to Tampa General Hospital | 216
awake and alert | 216
non-verbal | 216
unable to follow commands | 216
required assistance with daily living | 216
extensive workup | 216
serum laboratory testing | 216
autoimmune workup | 216
infectious workup | 216
paraneoplastic panel | 216
elevated CRP | 216
elevated ESR | 216
lumbar puncture | 216
elevated protein | 216
MRI brain | 216
diffuse slowing on EEG | 216
CT of the chest, abdomen, and pelvis | 216
IVIG | 216
brain biopsy | 240
white matter spongiform changes | 240
reactive gliosis | 240
absence of inflammation | 240
discharged to rehabilitation facility | 264
slow clinical improvement | 4320
alert and attentive | 8760
non-dysarthric speech | 8760
normal speech content | 8760
following commands | 8760
mild expressive aphasia | 8760
fully ambulatory | 8760
MMSE examination | 8760
genetic evaluation | 8760
no inheritable metabolic defect | 8760
continued clinical improvement | 10920
insecticides | -720
non-FDA approved anabolic steroids | -720
opioids | -720
benzodiazepines | -720
rodent-repellents | -720