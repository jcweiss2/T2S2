47 years old | 0
    male | 0
    admitted to the hospital | 0
    primary school director | 0
    goiter in euthyroidism | 0
    renovation work one month before | -672
    onset one week ago | -168
    high fever | -168
    repeated chills | -168
    diffuse myalgias | -168
    onset 4 days later | -96
    mucocutaneous jaundice | -96
    yellowish diarrhea | -96
    more than 4 stools/day | -96
    abdominal pain | -96
    right hypochondrium pain | -96
    patient altered | 0
    dehydrated | 0
    conscious | 0
    temperature 38°C | 0
    blood pressure 90/70 mm Hg | 0
    oxygen saturation 98% | 0
    jaundice | 0
    liver normal size | 0
    spleen normal size | 0
    white blood cells 29,000/mm3 | 0
    neutrophils 91% | 0
    hemoglobin 8.7 g/dL | 0
    platelet counts 30,000/mm3 | 0
    serum creatinine 76 mg/L | 0
    urea 1.38 g/L | 0
    alanine aminotransferase 140 IU/L | 0
    aspartate aminotransferases 180 IU/L | 0
    alkaline phosphatase 194 IU/L | 0
    total bilirubin 425 mg/L | 0
    conjugated bilirubin 80% | 0
    prothrombin level 95% | 0
    clear cerebrospinal fluid | 0
    cytochemical normal | 0
    chest radiograph unremarkable | 0
    abdominopelvic ultrasound normal-sized liver | 0
    non-dilated bile ducts | 0
    low abundance fluid effusion | 0
    treated with ceftriaxone | 0
    treated with ciprofloxacin | 0
    treated with metronidazole | 0
    parenteral rehydration | 0
    3rd day | 72
    blood pressure 60/40 mm Hg | 72
    moderate hematemesis | 72
    unable to eat | 72
    abdominal pain | 72
    nausea | 72
    abdomen tense | 72
    abdomen bloated | 72
    depressible to palpation | 72
    transit preserved | 72
    diuresis null | 72
    worsening renal insufficiency | 72
    urea 3.31 g/L | 72
    creatinine 106 mg/L | 72
    hyponatremia 115 mEq/L | 72
    hemoglobin 6.7 g/dL | 72
    procalcitonin 111 ng/mL | 72
    creatine phosphokinase 833 IU/L | 72
    lactate dehydrogenase 955 IU/L | 72
    lipaemia 273 IU/L | 72
    amylasemia 429 IU/L | 72
    electrocardiography normal | 72
    echocardiography normal | 72
    abdominal CT angiography enlarged pancreas | 72
    caudal part losing lobulated aspect | 72
    slight densification peri-caudal fat | 72
    necrosis flow back cavity omentums | 72
    liquid digestive distension | 72
    hydro-aeric level 38 mm | 72
    densification mesenteric fat | 72
    intraperitoneal effusion medium abundance | 72
    transferred to medical resuscitation service | 72
    noradrenaline | 72
    vascular filling | 72
    blood transfusions | 72
    extrarenal purification sessions | 72
    Inexium | 72
    antibiotic therapy maintained | 72
    gradual improvement clinical | 72
    gradual improvement biological | 72
    initiated diuresis | 72
    colors return | 72
    17th day | 408
    kidney tests correct | 408
    liver tests correct | 408
    blood cultures negative | 408
    HBsAg negative | 408
    anti-HAV IgM negative | 408
    anti-HCV antibodies negative | 408
    HIV serology negative | 408
    SARS-CoV-2 PCR negative | 408
    MAT serology positive Leptospira biflexa | 408
    discharged from the hospital | 408
    followed up several times | 408
    no complication | 408
    