65 years old | 0
female | 0
Guatemalan | 0
admitted to the hospital | 0
nausea | -48
vomiting | -48
diarrhea | -48
CIDP | -7200
prednisone 40-60 mg daily | -7200
emigrated from Guatemala | -7200
visited Guatemala annually | -7200
prior positive Strongyloides serology | -7200
peripheral eosinophilia | -7200
no prior anti-helminthic treatment | -7200
blood pressure 94/72 mmHg | 0
heart rate 158 beats/min | 0
respiratory rate 26 breaths/min | 0
oxygen saturation 94% | 0
temperature 37.0 °C | 0
rigors | 0
dry mucous membranes | 0
clear lung fields | 0
suprapubic tenderness | 0
WBC count 22,000/mm3 | 0
19% bands | 0
0% eosinophils | 0
urinalysis 22 WBC/high powered field | 0
IV fluids | 0
ciprofloxacin | 0
metronidazole | 0
methylprednisolone 100 mg IV | 0
admitted to ICU | 0
piperacillin-tazobactam | 0
methylprednisolone discontinued | 0
prednisone 30 mg twice daily | 0
admission blood cultures grew Escherichia coli | 24
admission urine cultures grew Escherichia coli | 24
stool studies negative for enteric pathogens | 24
hemodynamic status improved | 48
transferred to medical ward | 48
progressive hypoxemia | 120
contrast-enhanced chest CT | 120
small bilateral pleural effusions | 120
diffuse perihilar and peripheral air space opacities | 120
chest X-ray | 192
progressive bilateral infiltrates | 192
bronchoscopy | 192
blood throughout the tracheobronchial tree | 192
serial aliquots of bronchoalveolar lavage fluid | 192
persistently hemorrhagic fluid | 192
intubated | 192
transferred to ICU | 192
WBC count 24,000/mm3 | 192
7% bands | 192
13% eosinophils | 192
platelets 348,000/mm3 | 192
prothrombin time 13.9 s | 192
DAH | 192
methylprednisolone 1 g daily | 192
oral ivermectin | 192
BAL fluid positive for Strongyloides stercoralis | 216
corticosteroids discontinued | 216
subcutaneous ivermectin | 216
repeat bronchoscopy | 216
resolving hemorrhage | 216
serologies negative for ANCA | 216
serologies negative for anti-GBM | 216
serologies negative for ANA | 216
serologies negative for HIV | 216
serologies negative for HTLV-1 | 216
stool studies monitored | 216
discharged | 240
completed 4 weeks of daily oral ivermectin therapy | 672