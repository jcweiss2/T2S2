59 years old | 0
male | 0
chronic obstructive pulmonary disease | -672
generalized fatigue | -24
dyspnea | -24
oliguria | -24
blood pressure 70/40 mmHg | 0
pulse rate 122 bpm | 0
temperature 36.4°C | 0
peripheral oxygen saturation 88% | 0
decreased breath sounds in the lower right lung fields | 0
pretibial edema | 0
hepatomegaly | 0
serum potassium 6.0 mEq/dL | 0
phosphorus 5.2 mg/dL | 0
alanine aminotransferase 672 U/L | 0
alkaline phosphatase 489 U/L | 0
total bilirubin 1.6 mg/dL | 0
direct bilirubin 0.87 mg/dL | 0
lactate dehydrogenase 2954 U/L | 0
creatinine 2.15 mg/dL | 0
uric acid 20.32 mg/dL | 0
serum calcium level 10.2 mg/dL | 0
albumin 3.0 g/dL | 0
C-reactive protein 115 mg/L | 0
pulmonary medicine department suspected cancer | -168
thoracoabdominal computed tomography scan | -168
11 cm × 9 cm × 8 cm solid mass | -168
surrounding atelectasis | -168
mediastinal lymphadenopathies | -168
multiple liver metastases | -168
biopsy conducted with bronchoscopy | -72
admitted to the intensive care unit | 0
diagnosis of TLS | 0
intravenous fluid hydration | 0
antipotassium treatment | 0
allopurinol | 0
blood and urine cultures | 0
meropenem | 0
serial laboratory examinations | 0
increases in the levels of Cr | 24
increases in the levels of potassium | 24
increases in the levels of phosphorus | 24
hemodialysis | 24
official pathology reports confirmed SCLS | 24
death | 72
urea 215 mg/dL | 0
urea 202 mg/dL | 24
urea 241 mg/dL | 48
creatinine 2.02 mg/dL | 24
creatinine 2.19 mg/dL | 48
uric acid 19.2 mg/dL | 24
uric acid 17.6 mg/dL | 48
potassium 6.8 mmol/L | 24
potassium 7.1 mmol/L | 48
phosphorus 6.2 mg/dL | 24
phosphorus 7.2 mg/dL | 48
calcium 9.8 mg/dL | 24
calcium 9.6 mg/dL | 48
ALT 824 U/L | 24
ALT 986 U/L | 48
LDH 3277 U/L | 24
LDH 5450 U/L | 48
total bilirubin 1.5 mg/dL | 24
total bilirubin 1.63 mg/dL | 48
C-reactive protein 115 mg/L | 24
C-reactive protein 139 mg/L | 48
venous blood pH 7.21 | 0
venous blood pH 7.23 | 24
venous blood pH 6.82 | 48
sodium bicarbonate 14.7 mEq/L | 0
sodium bicarbonate 15.4 mEq/L | 24
sodium bicarbonate 4.9 mEq/L | 48
lactic acid 7.3 mmol/L | 0
lactic acid 7.2 mmol/L | 24
lactic acid 9.1 mmol/L | 48