17 years old | 0
female | 0
admitted to the hospital | 0
headache | -744
occupying lesion located in bilateral and third ventricles | 0
neuronavigation-assisted IVT tumor excision | 0
external ventricular drainage (EVD, right side) | 0
cefazolin | 0
vancomycin | 48
ceftriaxone | 144
leucocytosis | 48
abnormal CSF laboratory examination | 48
fever | 408
nausea | 408
emesis | 408
apathy | 408
carbapenem-resistant Enterobacter cloacae infection | 480
MIC to imipenem ≥16 mg/mL | 480
blood culture positive | 480
tigecycline | 480
amikacin | 480
cardiac and respiratory arrest | 480
herniation of the brain | 480
EVD (right side) | 480
meropenem | 528
cotrimoxazole | 528
allergic to cotrimoxazole | 528
fever persisted | 528
lethargy | 528
CSF cultures still showed carbapenem-resistant Enterobacter cloacae infection | 528
IVT amikacin | 576
informed consent | 576
amikacin administered IVT | 576
CSF drainage tube temporarily closed | 576
elevated WBC count | 624
CSF culture persistently positive | 624
EVD (left side) | 696
hydrocephalus | 768
EVD (right side) | 768
CSF culture negative | 864
IVT treatment well tolerated | 864
ventricular drainages removed | 960
IVT amikacin discontinued | 1104
meropenem and amikacin stopped | 1696
CSF culture continuously negative | 1696
mental status improved | 1696
fever subsided | 1696
no nephrotoxicity or seizures | 1696
no focal deficits | 1696
central neurocytoma | 1696
radiotherapy and rehabilitation | 1696
third ventriculostomy and septostomy | 1696
full recovery | 1696