baby boy | 0 | 0 
born by emergency cesarean section | 0 | 0 
severe preeclampsia in the mother | -672 | 0 
gestational week 25 6/7 | 0 | 0 
birthweight 665 g | 0 | 0 
intubated in the delivery room | 0 | 0 
transferred to the neonatal intensive care unit | 0 | 0 
mechanical ventilation | 0 | 0 
total parenteral nutrition | 24 | 0 
minimal enteral nutrition with breast milk | 24 | 0 
delayed meconium passage | 48 | 0 
abdominal distension | 48 | 0 
increased gastric residuals | 48 | 0 
necrotizing enterocolitis | 48 | 0 
gastric free drainage | 144 | 0 
broad-spectrum antibiotic therapy | 144 | 0 
perforated NEC | 144 | 0 
surgery | 144 | 0 
short bowel syndrome | 144 | 0 
thyroid screening tests | 336 | 0 
low circulating free and total throxine | 336 | 0 
low TSH | 336 | 0 
cortisol 5.75 µg/dL | 336 | 0 
serum total bilirubin level 12.12 mg/dL | 336 | 0 
direct reacting bilirubin 11.48 mg/dL | 336 | 0 
enteral levothyroxine 5 µg/kg/day | 336 | 504 
increased enteral levothyroxine 10 µg/kg/day | 504 | 576 
rectal levothyroxine 10 µg/kg/day | 576 | 1824 
increased fT4 levels | 1584 | 0 
decreased bilirubin levels | 1584 | 0 
severe bronchopulmonary dysplasia | 1824 | 0 
surgical NEC | 1824 | 0 
sepsis | 1824 | 0 
death | 1824 | 1824 
written informed consent | 0 | 0 
publication | 0 | 0