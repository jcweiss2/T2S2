65 years old | 0
male | 0
admitted to the hospital | 0
multiple blisters | -432
erosions | -432
oral mucosa | -432
scalp | -432
superadded maggot infection | -432
previous episodes of lesions | -720
treatment with steroids | -720
unknown generic medications | -720
lesions all over the body | -216
febrile | 0
flaccid blisters | 0
erosions | 0
Nikolsky sign positive | 0
diagnosis of PV | 0
skin biopsy | 0
tzanck smear | 0
intravenous dexamethasone pulse | 0
supportive care | 0
intravenous antibiotics | 0
isolation intensive care unit | 0
oozing from skin ulcerations | 0
hemorrhagic excoriation | 0
peeling of skin | 0
oral methyl prednisolone | 0
hypoproteinemia | 72
pleural effusion | 72
blood culture showed enterobacter | 72
pus culture showed Staphylococcus aureus | 72
pus culture showed Proteus mirabilis | 72
intravenous Tigecycline | 72
intravenous vancomycin | 72
sepsis | 72
high grade fever | 72
albumin levels fell | 72
TPE cycle | 72
TPE performed | 96
anticoagulation with citrate | 96
replacement of plasma | 96
monitoring of hemodynamic parameters | 96
complications during procedure | 96
Nikolsky sign negative | 168
no new lesions | 168
exudation from lesions reduced | 168
dressings dry | 168
lesions showed re-epithelization | 168
lesions showed healing | 240
oral lesions healed | 240
IV methyl prednisolone pulse | 240
cyclophosphamide | 240
discharged | 360
monthly IV dexamethasone pulse | 360
daily oral prednisolone | 360