8 years old | 0
male | 0
admitted to the hospital | 0
severe abdominal pain | 0
diagnosed with ALL | -3456
first relapse | -1095
bone marrow transplant | -1095
second relapse | -672
last chemotherapy | -72
high dose of methotraxate | -72
no vaccination against chickenpox | -1095
normal body temperature | 0
hepatosplenomegaly | 0
tenderness in the periumbilical area | 0
hemoglobin of 12.1 g/dL | 0
WBCs count of 3,490/mm3 | 0
segmented neutrophils of 80.0% | 0
platelet count of 135,000/mm3 | 0
slightly increased levels of AST | 0
slightly increased levels of ALT | 0
fever | 24
empirical intravenous antibiotics | 24
abdominal pain remained constant | 24
multiple erythematous vesicles | 48
acyclovir | 48
vesicles developed across the whole body | 96
dyspnea | 96
varicella pneumonia | 96
WBCs of 5,090/mm3 | 96
platelet count of 32,000/mm3 | 96
AST of 931 U/L | 96
ALT of 788 U/L | 96
LDH of 3,196 U/L | 96
DIC profile was positive | 96
intravenous immunoglobulin | 96
single donor platelets | 96
fresh frozen plasma | 96
antithrombin III | 96
transferred to the ICU | 96
drowsy mental state | 108
dyspnea was aggravated | 108
total haziness and ARDS | 108
intubation | 108
mechanical respiratory support | 108
increased dose of IVIG | 108
cardiomegaly | 144
platelet count was 69,000/mm3 | 144
AST and ALT were 224 U/L and 280 U/L | 144
recovered from DIC | 144
fever persisted | 144
vesicular skin lesions showed no change | 144
VZV was detected in patient serum | 168
increased blood pressure | 168
intravenous labetarol | 168
generalized tonic-clonic seizure | 204
hypertensive crisis | 204
VZV involvement in central nerve system | 204
intravenous nitroprusside | 204
cerebrospinal fluid tapping | 204
normal CSF results | 204
VZV antibody and PCR in CSF were negative | 204
increased antihypertensives dose | 204
intravenous phenytoin | 204
no more seizures | 204
pulmonary condition was stable | 240
taken off the ventilator | 240
no fever | 240
all skin lesions reached the scarring stage | 240
transferred from the ICU to the general ward | 312
vital signs were stable | 312
all laboratory data showed improvements | 312
lymphocyte subset showed CD3 of 87.0% | 312
lymphocyte subset showed CD4 of 14.8% | 312
lymphocyte subset showed CD8 of 70.6% | 312
lymphocyte subset showed CD19 of 9.6% | 312
lymphocyte subset showed CD56 of 3.0% | 312
brain MRI showed multiple patchy high-signal-intensity lesions | 312
EEG looked normal | 312
phenytoin was stopped | 312
ceased administration of intravenous antibiotics | 360
ceased administration of acyclovir | 360
discharged | 360
chemotherapy was resumed | 720
follow-up brain MRI was done | 2160
multiple high-signal-intensity lesions due to VZV-induced encephalitis were disappeared | 2160