59 years old | 0
    woman | 0
    advanced lung cancer | 0
    pulmonary hypertension | 0
    cirrhosis of the liver | 0
    hepatitis C positivity | 0
    history of alcohol abuse | 0
    consumed raw oysters | -24
    generalized lower abdominal pain | -12
    non-radiating dull abdominal ache | 0
    denied fever | 0
    denied chills | 0
    no nausea | 0
    no vomiting | 0
    blood pressure 75/50 mm Hg | 0
    pulse rate 100 beats/min | 0
    respiratory rate 22 breaths/min | 0
    temperature 36.7°C | 0
    no signs of distress | 0
    nontoxic appearance | 0
    lungs clear | 0
    lower abdominal tenderness | 0
    no peritoneal signs | 0
    WBC count 0.7 K/uL | 0
    hemoglobin 12.5 g/dL | 0
    platelet count 32 K/uL | 0
    sodium 144 mEq/L | 0
    potassium 3.6 mEq/L | 0
    creatinine 1.75 mg/dL | 0
    BUN 16 mg/dL | 0
    glucose 71 mg/dL | 0
    albumin 1.9 g/L | 0
    urinalysis +1 protein | 0
    urinalysis +1 blood | 0
    urinalysis +4 urobilinogen | 0
    2.5 hyaline casts per high power field | 0
    51 to 100 WBCs with clumps | 0
    CT scan right colon wall thickening | 0
    inflammation terminal ileum and appendix | 0
    portal venous congestion | 0
    cirrhosis of the liver confirmed | 0
    right lower lobe infiltrate | 0
    no splenomegaly | 0
    admitted to ICU | 0
    sepsis with shock | 0
    colitis | 0
    right lower lobe pneumonia | 0
    urinary tract infection | 0
    IV fluid boluses | 0
    remained hypotensive | 0
    norepinephrine initiated | 0
    broad-spectrum antibiotics initiated | 0
    cefepime | 0
    metronidazole | 0
    levofloxacin | 0
    no pharmacologic DVT prophylaxis | 0
    Granix administered | 0
    radiation 2 months prior | -1440
    dyspnea treated with albuterol/ipratropium | 0
    oxygen saturation above 93% | 0
    acute hypoxic respiratory failure | 24
    progressive encephalopathy | 24
    endotracheal intubation | 24
    mechanical ventilation | 24
    orogastric tube placed | 24
    septic shock persisted | 24
    hypotension persisted | 24
    albumin administered | 24
    sodium bicarbonate infusion | 24
    vitamin C sepsis protocol initiated | 24
    vitamin C 500 mg IV | 24
    hydrocortisone 100 mg IV | 24
    thiamine 200 mg IV | 24
    gram-negative bacteremia | 24
    doxycycline added | 24
    blisters and boils forming | 34
    E. tarda bacteremia | 34
    died | 34
