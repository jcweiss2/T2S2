\
\boxed{
65 years old | 0
female | 0
admitted to the hospital | 0
fever | 0
chills | 0
pain in left leg | 0
known case of parkinsonism | 0
diabetes mellitus | 0
levodopa / carbidopa | 0
rasagiline | 0
ropinirole | 0
trihexyphenidyl | 0
amantadine | 0
metformin | 0
glipizide | 0
multiple hospital and ICU admissions | 0
worsening parkinsonism | 0
admitted to the ward for cellulitis | 0
intravenous clindamycin | 0
intravenous benzylpenicillin | 0
anti-parkinsonism and diabetic medications continued | 0
persistently high-temperature spikes | 72
tachycardia | 72
tachypnea | 72
hypotensive | 72
encephalopathic | 72
shifted to ICU | 72
sepsis with multi-organ dysfunction syndrome | 72
intravenous linezolid | 72
intravenous piperacillin with tazobactam | 72
vancomycin not considered | 72
hemodynamics improved | 72
minimal inotropic supports | 72
anti-parkinsonism drugs continued | 72
oral hypoglycemic agents stopped | 72
switched to insulin | 72
confused | 72
drowsy | 72
disoriented | 72
altered sensorium | 72
myoclonus | 72
tremors | 72
jerky movements | 72
no neck stiffness | 72
computed tomography of the brain not significant | 72
cerebrospinal fluid analysis not significant | 72
improving white blood cell counts | 72
better glycemic control | 72
blood and pus cultures sterile | 72
high temperature | 168
altered mental status | 168
myoclonus | 168
jerky movements | 168
tremors | 168
serotonin syndrome suspected | 168
linezolid and rasagiline stopped | 168
temperature settled | 176
heart rate normal | 192
sensorium improved | 192
tremors completely subsided | 192
shifted out of the ICU | 192
started walking with support | 264
discharged from the hospital | 264
discharged with anti-parkinsonism drugs | 264
rasagiline added | 264
regular follow-up with the neurologist | 264
stable and remained asymptomatic for serotonin syndrome | 264
}
\boxed{
65 years old | 0
female | 0
admitted to the hospital | 0
fever | 0
chills | 0
pain in left leg | 0
known case of parkinsonism | 0
diabetes mellitus | 0
levodopa / carbidopa | 0
rasagiline | 0
ropinirole | 0
trihexyphenidyl | 0
amantadine | 0
metformin | 0
glipizide | 0
multiple hospital and ICU admissions | 0
worsening parkinsonism | 0
admitted to the ward for cellulitis | 0
intravenous clindamycin | 0
intravenous benzylpenicillin | 0
anti-parkinsonism and diabetic medications continued | 0
persistently high-temperature spikes | 72
tachycardia | 72
tachypnea | 72
hypotensive | 72
encephalopathic | 72
shifted to ICU | 72
sepsis with multi-organ dysfunction syndrome | 72
intravenous linezolid | 72
intravenous piperacillin with tazobactam | 72
vancomycin not considered | 72
hemodynamics improved | 72
minimal inotropic supports | 72
anti-parkinsonism drugs continued | 72
oral hypoglycemic agents stopped | 72
switched to insulin | 72
confused | 72
drowsy | 72
disoriented | 72
altered sensorium | 72
myoclonus | 72
tremors | 72
jerky movements | 72
no neck stiffness | 72
computed tomography of the brain not significant | 72
cerebrospinal fluid analysis not significant | 72
improving white blood cell counts | 72
better glycemic control | 72
blood and pus cultures sterile | 72
high temperature | 168
altered mental status | 168
myoclonus | 168
jerky movements | 168
tremors | 168
serotonin syndrome suspected | 168
linezolid and rasagiline stopped | 168
temperature settled | 176
heart rate normal | 192
sensorium improved | 192
tremors completely subsided | 192
shifted out of the ICU | 192
started walking with support | 264
discharged from the hospital | 264
discharged with anti-parkinsonism drugs | 264
rasagiline added | 264
regular follow-up with the neurologist | 264
stable and remained asymptomatic for serotonin syndrome | 264
} \n
\boxed{
65 years old | 0
female | 0
admitted to the hospital | 0
fever | 0
chills | 0
pain in left leg | 0
known case of parkinsonism | 0
diabetes mellitus | 0
levodopa / carbidopa | 0
rasagiline | 0
ropinirole | 0
trihexyphenidyl | 0
amantadine | 0
metformin | 0
glipizide | 0
multiple hospital and ICU admissions | 0
worsening parkinsonism | 0
admitted to the ward for cellulitis | 0
intravenous clindamycin | 0
intravenous benzylpenicillin | 0
anti-parkinsonism and diabetic medications continued | 0
persistently high-temperature spikes | 72
tachycardia | 72
tachypnea | 72
hypotensive | 72
encephalopathic | 72
shifted to ICU | 72
sepsis with multi-organ dysfunction syndrome | 72
intravenous linezolid | 72
intravenous piperacillin with tazobactam | 72
vancomycin not considered | 72
hemodynamics improved | 72
minimal inotropic supports | 72
anti-parkinsonism drugs continued | 72
oral hypoglycemic agents stopped | 72
switched to insulin | 72
confused | 72
drowsy | 72
disoriented | 72
altered sensorium | 72
myoclonus | 72
tremors | 72
jerky movements | 72
no neck stiffness | 72
computed tomography of the brain not significant | 72
cerebrospinal fluid analysis not significant | 72
improving white blood cell counts | 72
better glycemic control | 72
blood and pus cultures sterile | 72
high temperature | 168
altered mental status | 168
myoclonus | 168
jerky movements | 168
tremors | 168
serotonin syndrome suspected | 168
linezolid and rasagiline stopped | 168
temperature settled | 176
heart rate normal | 192
sensorium improved | 192
tremors completely subsided | 192
shifted out of the ICU | 192
started walking with support | 264
discharged from the hospital | 264
discharged with anti-parkinsonism drugs | 264
rasagiline added | 264
regular follow-up with the neurologist | 264
stable and remained asymptomatic for serotonin syndrome | 264
} \n
\boxed{
65 years old | 0
female | 0
admitted to the hospital | 0
fever | 0
chills | 0
pain in left leg | 0
known case of parkinsonism | 0
diabetes mellitus | 0
levodopa / carbidopa | 0
rasagiline | 0
ropinirole | 0
trihexyphenidyl | 0
amantadine | 0
metformin | 0
glipizide | 0
multiple hospital and ICU admissions | 0
worsening parkinsonism | 0
admitted to the ward for cellulitis | 0
intravenous clindamycin | 0
intravenous benzylpenicillin | 0
anti-parkinsonism and diabetic medications continued | 0
persistently high-temperature spikes | 72
tachycardia | 72
tachypnea | 72
hypotensive | 72
encephalopathic | 72
shifted to ICU | 72
sepsis with multi-organ dysfunction syndrome | 72
intravenous linezolid | 72
intravenous piperacillin with tazobactam | 72
vancomycin not considered | 72
hemodynamics improved | 72
minimal inotropic supports | 72
anti-parkinsonism drugs continued | 72
oral hypoglycemic agents stopped | 72
switched to insulin | 72
confused | 72
drowsy | 72
disoriented | 72
altered sensorium | 72
myoclonus | 72
tremors | 72
jerky movements | 72
no neck stiffness | 72
computed tomography of the brain not significant | 72
cerebrospinal fluid analysis not significant | 72
improving white blood cell counts | 72
better glycemic control | 72
blood and pus cultures sterile | 72
high temperature | 168
altered mental status | 168
myoclonus | 168
jerky movements | 168
tremors | 168
serotonin syndrome suspected | 168
linezolid and rasagiline stopped | 168
temperature settled | 176
heart rate normal | 192
sensorium improved | 192
tremors completely subsided | 192
shifted out of the ICU | 192
started walking with support | 264
discharged from the hospital | 264
discharged with anti-parkinsonism drugs | 264
rasagiline added | 264
regular follow-up with the neurologist | 264
stable and remained asymptomatic for serotonin syndrome | 264
} \n
\boxed{
65 years old | 0
female | 0
admitted to the hospital | 0
fever | 0
chills | 0
pain in left leg | 0
known case of parkinsonism | 0
diabetes mellitus | 0
levodopa / carbidopa | 0
rasagiline | 0
ropinirole | 0
trihexyphenidyl | 0
amantadine | 0
metformin | 0
glipizide | 0
multiple hospital and ICU admissions | 0
worsening parkinsonism | 0
admitted to the ward for cellulitis | 0
intravenous clindamycin | 0
intravenous benzylpenicillin | 0
anti-parkinsonism and diabetic medications continued | 0
persistently high-temperature spikes | 72
tachycardia | 72
tachypnea | 72
hypotensive | 72
encephalopathic | 72
shifted to ICU | 72
sepsis with multi-organ dysfunction syndrome | 72
intravenous linezolid | 72
intravenous piperacillin with tazobactam | 72
vancomycin not considered | 72
hemodynamics improved | 72
minimal inotropic supports | 72
anti-parkinsonism drugs continued | 72
oral hypoglycemic agents stopped | 72
switched to insulin | 72
confused | 72
drowsy | 72
disoriented | 72
altered sensorium | 72
myoclonus | 72
tremors | 72
jerky movements | 72
no neck stiffness | 72
computed tomography of the brain not significant | 72
cerebrospinal fluid analysis not significant | 72
improving white blood cell counts | 72
better glycemic control | 72
blood and pus cultures sterile | 72
high temperature | 168
altered mental status | 168
myoclonus | 168
jerky movements | 168
tremors | 168
serotonin syndrome suspected | 168
linezolid and rasagiline stopped | 168
temperature settled | 176
heart rate normal | 192
sensorium improved | 192
tremors completely subsided | 192
shifted out of the ICU | 192
started walking with support | 264
discharged from the hospital | 264
discharged with anti-parkinsonism drugs | 264
rasagiline added | 264
regular follow-up with the neurologist | 264
stable and remained asymptomatic for serotonin syndrome | 264
} \n
\boxed{
65 years old | 0
female | 0
admitted to the hospital | 0
fever | 0
chills | 0
pain in left leg | 0
known case of parkinsonism | 0
diabetes mellitus | 0
levodopa / carbidopa | 0
rasagiline | 0
ropinirole | 0
trihexyphenidyl | 0
amantadine | 0
metformin | 0
glipizide | 0
multiple hospital and ICU admissions | 0
worsening parkinsonism | 0
admitted to the ward for cellulitis | 0
intravenous clindamycin | 0
intravenous benzylpenicillin | 0
anti-parkinsonism and diabetic medications continued | 0
persistently high-temperature spikes | 72
tachycardia | 72
tachypnea | 72
hypotensive | 72
encephalopathic | 72
shifted to ICU | 72
sepsis with multi-organ dysfunction syndrome | 72
intravenous linezolid | 72
intravenous piperacillin with tazobactam | 72
vancomycin not considered | 72
hemodynamics improved | 72
minimal inotropic supports | 72
anti-parkinsonism drugs continued | 72
oral hypoglycemic agents stopped | 72
switched to insulin | 72
confused | 72
drowsy | 72
disoriented | 72
altered sensorium | 72
myoclonus | 72
tremors | 72
jerky movements | 72
no neck stiffness | 72
computed tomography of the brain not significant | 72
cerebrospinal fluid analysis not significant | 72
improving white blood cell counts | 72
better glycemic control | 72
blood and pus cultures sterile | 72
high temperature | 168
altered mental status | 168
myoclonus | 168
jerky movements | 168
tremors | 168
serotonin syndrome suspected | 168
linezolid and rasagiline stopped | 168
temperature settled | 176
heart rate normal | 192
sensorium improved | 192
tremors completely subsided | 192
shifted out of the ICU | 192
started walking with support | 264
discharged from the hospital | 264
discharged with anti-parkinsonism drugs | 264
rasagiline added | 264
regular follow-up with the neurologist | 264
stable and remained asymptomatic for serotonin syndrome | 264
} \n
\boxed{
65 years old | 0
female | 0
admitted to the hospital | 0
fever | 0
chills | 0
pain in left leg | 0
known case of parkinsonism | 0
diabetes mellitus | 0
levodopa / carbidopa | 0
rasagiline | 0
ropinirole | 0
trihexyphenidyl | 0
amantadine | 0
met