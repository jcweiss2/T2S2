52 years old | 0
    woman | 0
    history of bipolar disorder | -87600
    treated with lithium (1650 mg/day) | -87600
    treated with risperidone (2.5 mg/day) | -87600
    presented to general practitioner | -168
    dry cough | -48
    sweats | -48
    feeling feverish | -48
    upper respiratory tract infection | -168
    symptoms persisted | 0
    addressed to emergency department | 0
    delirium | 0
    pain in upper right abdominal quadrant | 0
    fever (39°C) | 0
    tachycardia | 0
    irregular heart rhythm | 0
    blood pressure 149/87 mm Hg | 0
    tenderness of upper right abdominal quadrant | 0
    normal white blood cell count | 0
    elevated CRP (43.5 mg/dL) | 0
    hyponatraemia (129 mmol/L) | 0
    corrected calcium (2.61 mmol/L) | 0
    potassium level (3.5 mmol/L) | 0
    acute kidney injury | 0
    creatinine (120 µmol/L) | 0
    urine culture positive for Escherichia coli | 0
    serum lithium concentration elevated (2.0 mmol/L) | 0
    ECG atrial fibrillation | 0
    wide QRS complex (160 ms) | 0
    ST-segment elevation in V1 and V2 | 0
    previous ECG sinus rhythm | 0
    narrow QRS | 0
    abdominal CT scan confirmed pyelonephritis | 0
    ruled out cholecystitis | 0
    delirium complicating symptoms assessment | 0
    ECG alterations | 0
    possibility of acute coronary syndrome | 0
    ST elevation limited to V1 and V2 | 0
    no reciprocal changes | 0
    high-sensitivity troponin slightly elevated (20 ng/L) | 0
    no dynamic change | 0
    acute kidney injury | 0
    focused transthoracic echocardiography no wall-motion abnormality | 0
    full TTE confirmed normal biventricular function | 72
    no wall-motion abnormality | 72
    normal filling pressures | 72
    absence of left atrial enlargement | 72
    no valvular disease | 72
    AF multifactorial | 0
    sepsis | 0
    electrolyte imbalance | 0
    lithium intoxication | 0
    diagnosis of Brugada syndrome not immediately evoked | 0
    admitted to intensive care unit | 0
    continuous cardiac monitoring | 0
    lithium suspended | 0
    normal saline infusion initiated | 0
    empirical ceftriaxone | 0
    switched to ciprofloxacin | 48
    continued for seven days | 48
    blood cultures sterile | 0
    rapid clinical improvement | 0
    heart rate 100-110 bpm | 0
    no rate or rhythm control for AF | 0
    complete resolution of delirium | 168
    complete resolution of fever | 168
    complete resolution of abdominal pain | 168
    discharge | 168
    correction of renal function | 0
    lithium concentration 0.68 mmol/L | 48
    electrolyte levels normalized | 48
    spontaneous cardioversion of AF | 24
    ECG sinus rhythm | 48
    first-degree atrioventricular block | 48
    narrow QRS (120 ms) | 48
    ST-segment elevation less than 1 mm in V1 and V2 | 48
    final diagnosis conduction abnormalities | 0
    acute-on-chronic lithium intoxication | 0
    sepsis | 0
    acute renal failure | 0
    reduced lithium posology (1320 mg/day) | 168
    discharge | 168
    Brugada pattern suspected | 720
    ECG Brugada type 1 pattern | 720
    episodes of near-syncope | -87600
    vasovagal origin | -87600
    ECG 3 years earlier slightly convex ST segment elevation in V2 | -26280
    type 2 Brugada pattern | -26280
    hospitalised again | 720
    lithium withdrawal | 720
    valproic acid replacement | 720
    ECG no persistent Brugada pattern | 720
    declined genetic testing | 720
    brother's ECG discrete alterations | 720
    ajmaline provocation test positive | 720
    SCN5A mutation confirmed (c.3840+1G>A) | 720
    no implantable cardioverter-defibrillator | 720
    clinical follow-up | 720
