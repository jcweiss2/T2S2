56 years old | 0
female | 0
admitted to the hospital | 0
neck swelling | -144
tenderness | -144
diagnosed with hypertension | -4380
blood pressure well controlled via medication | -4380
Mallampatti class IV | 0
mouth opening of less than three finger widths | 0
neck computed tomography (CT) findings | 0
right side retropharyngeal abscess | 0
anterior and posterior cervical space and carotid space | 0
preoperative airway evaluation | 0
vital signs | 0
blood pressure 140/83 mmHg | 0
heart rate 110 beats/min | 0
saturation of percutaneous oxygen (SpO2) 97% | 0
arterial blood gas analysis | 0
mild respiratory alkalosis | 0
tachypnea | 0
respiration rate 25 breaths/min | 0
pH 7.50 | 0
partial pressure of CO2 34.1 mmHg | 0
partial pressure of O2 124.6 mmHg | 0
O2 saturation 99% | 0
preoxygenation | 0
facial mask with 100% oxygen | 0
indirect videolaryngoscope | 0
endotracheal tubes (ETTs) of various diameters | 0
lidocaine spray | 0
topicalization of the airway | 0
epiglottis visible | 0
glottis not visible | 0
Cormack and Lehane grade 3 | 0
intubation using indirect videolaryngoscope | 0
general anesthesia | 0
propofol 120 mg | 0
rocuronium 60 mg | 0
mask ventilation | 0
tidal volume 300 mL | 0
peak airway pressure 20 cmH2O | 0
intubation with an ETT with an internal diameter (ID) of 7.0 mm | 0
intubation with an ETT with an internal diameter (ID) of 6.5 mm | 0
oxygen saturation maintained above 97% | 0
anesthesia maintained | 0
sevoflurane 1.7 volume % | 0
remifentanil | 0
air 2 L/min | 0
O2 2 L/min | 0
pressure-controlled ventilation mode | 0
end-tidal CO2 28-30 mmHg | 0
pulse oximetry 100% | 0
surgery | 0
incision and retropharyngeal abscess drainage | 0
transcervical approach | 0
wound closure delayed | 0
transferred to the intensive care unit (ICU) | 24
mechanical ventilator | 24
saturation above 95% | 24
pressure-controlled ventilation | 24
tidal volume 450 mL | 24
respiration rate 12 breaths/min | 24
PEEP 5 cmH2O | 24
FiO2 0.4 | 24
recommenced spontaneous breathing | 48
extubated | 48
wound closure | 72
packing gauze removal | 72
monitored anesthesia care | 72
noninvasive blood pressure monitoring | 72
electrocardiography | 72
pulse oximetry | 72
end-tidal CO2 measurement | 72
nasal cannula with 100% O2 at 3 L/min | 72
dexmedetomidine 6 µg/kg/hr | 72
SpO2 decreased to 95% | 72
reservoir mask with 100% O2 at 6 L/min | 72
SpO2 dropped to 94% | 72
high-flow nasal cannula | 72
humidified oxygen flow 30 L/min | 72
fractional inspired oxygen 1.0 | 72
SpO2 maintained at 100% | 72
dexmedetomidine 0.6 µg/kg/hr | 82
fentanyl 50 µg | 82
midazolam 1 mg | 82
dexmedetomidine increased to 0.7-1.0 µg/kg/hr | 82
vital signs stable | 82
no signs of bradycardia | 82
no discomfort | 82
OAA/S score 2 | 82
recovery room | 120
100% O2 at 3 L/min via a nasal cannula | 120
O2 saturation 96-100% | 120
transported to a general hospital room | 120
discharged | 288