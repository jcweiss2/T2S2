66 years old|0
female|0
maintenance hemodialysis|0
COVID-19 infection|0
mild cough|0
sore throat|0
asthma|0
no personal travel history|0
attended extended family gathering|-120
family members with respiratory symptoms|0
fever of 38°C|0
placed on droplet and isolation precautions|0
nasopharyngeal swab ordered|0
discharged in stable condition|0
instructed to self-isolate|0
positive COVID-19 NP swab|0
admitted to hospital|24
private room|24
denied dyspnea|24
productive cough|24
blood pressure 113/65 mm Hg|24
oxygen saturation 91%|24
low-grade fever 38°C|24
bibasilar crackles|24
chest X-ray diffuse patchy infiltrates bilaterally|24
lymphopenia|24
progressive anemia|24
normal lactate|24
ferritin 275 μg/L|24
elevated partial thromboplastin time 39.4 seconds|24
D-dimer not performed|24
normal biventricular function|24
hypoxia|48
oxygen saturation 86%|48
improved with oxygen 2 L/min|48
dyspneic|48
respiratory deterioration|72
FiO2 50%|72
nonrebreather mask|72
intubated|72
transferred to ICU|72
septic shock|96
ceftriaxone|96
ciprofloxacin|96
hydroxychloroquine 400 mg|96
hydroxychloroquine 200 mg daily|96
negative influenza swab|96
salmeterol use|96
hemodynamic instability|96
continuous renal replacement therapy|96
regional citrate anticoagulation|96
vasopressors|96
prefilter replacement fluid|96
postfilter replacement fluid|96
no bleeding|96
no thrombosis|96
additional PPE training|96
care bundle approach|96
CRRT dosing reduced|96
CRRT for 13 days|240
transitioned to intermittent hemodialysis|240
PPE education|240
safety leader implemented|240
practice standards established|240
extubated|456
discharged home|600
droplet and contact precautions|600
surveillance COVID-19 swabs|600
persistently detectable PCR|600
laboratory abnormalities|600
readmitted|888
sinus tachycardia|888
biliary obstruction|888
endoscopic retrograde cholangiopancreatographies|888
secondary sclerosing cholangitis|888
infected liver abscesses|888
fluconazole|888
moxifloxacin|888
contact tracing|0
self-isolation of staff|0
self-isolation of patients|0
asymptomatic staff return to work|0
universal PPE precautions|0
no nosocomial spread|0
detectable viral PCR for 42 days|1008
two negative COVID# swabs|1008
elevated transaminases|600
synthetic liver function tests elevated|600
readmissions|888
antimicrobial therapy|888
clear to return to work|336
cleared by IP & C|1008
