68 years old | 0
male | 0
admitted to the hospital | 0
superficial bite wound | -24
bite delivered by 3-year-old child | -24
limb appeared swollen and cyanotic | -4
general discomfort | -4
swelling and pain in the distal right upper extremity | -16
visited a local clinic | -16
diagnosed with gout arthritis | -16
given nonsteroidal anti-inflammatory treatment | -16
worsening of the swelling and pain of the limb | -8
purpura around the wound and right hand | -8
systemic symptoms including weakness, palpitation, and cold sweats | -8
visited the emergency department | 0
acute pain | 0
in shock | 0
hypotension | 0
rapid pulse | 0
cold sweats | 0
flaky plaques | 0
swelling | 0
weak iliac artery pulsation | 0
dopamine administered | 0
laboratory and imaging examinations conducted | 0
swelling and ecchymosis of the patient’s limb continued to expand | 0
crepitus of the subcutaneous soft tissue | 0
gas bubbles in the subcutaneous tissue with edema | 0
anti-infection treatment administered | 0
condition did not alleviate | 0
limb lesions continued to expand | 0
deterioration of consciousness | 0
white blood cell count, 4.85 × 109/L | 0
hemoglobin concentration, 70 g/L | 0
platelet count, 36 × 109/L | 0
C-reactive protein concentration, 68.35 mg/L | 0
procalcitonin concentration, 48.960 ng/mL | 0
blood coagulation normal | 0
X-ray and computed tomography examinations revealed a large volume of gas in the soft tissue | 0
smear examination of the bite wound showed a large number of Gram-negative bacilli | 0
gas gangrene-like infection | 0
open amputation | 3
fish mouth incision in the skin | 3
entered the limb layer by layer | 3
revealed important vascular nerves and disconnected them | 3
ligated the blood vessels | 3
cut the bone at the upper part of the humerus | 3
trimmed the stump | 3
muscle sutured to cover the end of the bone | 3
wound not sutured but wrapped in a large amount of sterile wound dressing | 3
sent to the ICU for isolation treatment | 3
endotracheal intubation | 3
dissection of the amputated limb caused a large amount of malodorous gas to escape | 3
lesions were necrotic and dark purple | 3
some tissues had dissolved | 3
combination of penicillin, meropenem, and clindamycin for infection | 3
vasoactive drugs to maintain blood pressure | 3
intermittent fever after the operation | 12
infection index, procalcitonin concentration, and C-reactive protein concentration still elevated for 3 days postoperatively | 72
HGB concentration and PLT count remained at low levels during ICU treatment | 72
multi-point bacteriological culture revealed Aeromonas hydrophila | 72
postoperative pathologic examination revealed a large amount of necrotic tissue and inflammatory cell infiltration | 72
bone marrow smear revealed mild myeloid hyperplasia with decreased megakaryocytes | 72
bone marrow biopsy revealed interstitial edema and megakaryocyte reduction | 72
diagnosis of acute myeloid leukemia (AML) | 72
surgeons replaced the wound dressing daily | 72
exposed stump tissue emitted a foul odor and exudate | 96
local muscle tissue necrosis and a small number of ecchymoses around the wound | 96
stump trimmed to remove the necrotic tissue | 168
6 cm of the humerus removed from the proximal end | 168
wound sutured layer by layer and covered with a vacuum sponge | 168
vacuum sponge removed 1 week after stump revision surgery | 336
vital signs gradually recovered and stabilized | 240
laboratory indicators gradually recovered to near normal levels | 240
extubated on the 11th day after amputation | 264
resumed spontaneous breathing | 264
state of consciousness remained clear | 264
wound healed | 336
discharged | 336
died of blood system disease 2 years later | 17520