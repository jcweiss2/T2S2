73 years old | 0
    woman | 0
    duodenal switch surgery | 0
    pancreatic head adenocarcinoma | 0
    obstructive jaundice | 0
    DBE-ERCP attempted | 0
    unsuccessful DBE