39 years old | 0
male | 0
caucasian | 0
non-verbal | 0
stimulant abuse | -8760
traumatic anoxic brain injury | -8760
quadriplegia | -8760
reversed tracheostomy stoma | -8760
percutaneous gastrostomy tube dependence | -8760
PEG tube replaced | -432
high grade fever | 0
coffee ground emesis | 0
intubated | 0
aspiration pneumonia | 0
diffused crackles throughout the lung fields | 0
mild epigastric distention | 0
left lower quadrant tenderness | 0
PEG tube in place | 0
loose external bumper | 0
inability to twirl, retract or advance the tube | 0
normal bowel sounds | 0
normal sphincter tone | 0
hemoccult negative stool | 0
hemodynamically unstable | 0
low blood pressure | 0
norepinephrine | 0
mechanical ventilation | 0
100% fraction of inspired oxygen | 0
white blood cells 26,000 k/ul | 0
hemoglobin 12.9 g/dl | 0
granulocyte 80.1% | 0
sodium 157 mmol/l | 0
potassium 2.9 mmol/L | 0
chloride 116 mmol/L | 0
bicarbonate 31 mmol/l | 0
BUN 50 mg/dl | 0
glucose 212 mg/dl | 0
Lactic Acid 1.8 mmol/L | 0
AST 45 U/L | 0
bilateral infiltrations | 0
thickening at the distal end of stomach wall | 0
thickening at the proximal duodenum | 0
gastric tube retention of the balloon in the third part of duodenum | 0
PEG tube removal | 0
broad spectrum antibiotics | 0
vancomycin | 0
cefepime | 0
tapered off the norepinephrine | 24
new PEG tube insertion | 24
balloon inflated with 20cc of water | 24
external bumper fixed at 4 cm to skin level | 24
distance to the skin 1 cm | 24
significant improvement | 48
tolerating tube feeds again | 48
discharged to nursing home | 72