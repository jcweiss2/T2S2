85 years old | 0
    male | 0
    admitted to the hospital (initial clinic presentation) | -4320
    prior total hip arthroplasty (1997) | -17520
    head and liner exchange (2014) | -76800
    atrial fibrillation | -76800
    congestive heart failure | -76800
    peripheral vascular disease | -76800
    abdominal aortic aneurysm | -76800
    renal artery stenosis | -76800
    chronic kidney disease | -76800
    hypertension | -76800
    chronic obstructive pulmonary disease | -76800
    prostate cancer | -76800
    anticoagulated with rivaroxaban | -76800
    abdominal aortic aneurysm repair | -76800
    aortobifemoral bypass | -76800
    hospitalized for Escherichia coli sepsis (6 months before clinic) | -4320
    right hip pain (during sepsis hospitalization) | -4320
    readmitted with worsening right hip pain and swelling (2 months after sepsis hospitalization) | -2016
    transferred to institution | -2016
    serum laboratory work | -2016
    fluoroscopically guided hip joint aspiration | -2016
    diagnosed with periprosthetic joint infection | -2016
    cultures grew Escherichia coli | -2016
    plain radiographs at admission | -2016
    irrigation and debridement | -1920
    removal of total hip arthroplasty | -1920
    extended trochanteric osteotomy | -1920
    placement of antibiotic-impregnated cement spacer | -1920
    postoperative radiographs | -1920
    treated with 6 weeks intravenous antibiotics | -1920
    further 6 weeks oral antibiotics | -1920
    2-week antibiotic holiday | -1920
    fluoroscopically guided aspiration | -1920
    serologic markers normalized | -1920
    synovial fluid cell count normalized | -1920
    alpha defensin testing negative | -1920
    bacterial cultures negative | -1920
    infection cleared | -1920
    scheduled second-stage reimplantation | -1920
    physical examination (pre-second-stage surgery) | -1920
    well-healed posterolateral scar | -1920
    no signs of infection | -1920
    passive range of motion | -1920
    flex to 110° | -1920
    20° internal rotation | -1920
    40° external rotation | -1920
    no leg length discrepancy | -1920
    palpable dorsalis pedis pulses | -1920
    palpable posterior tibial pulses | -1920
    radiographs (pre-second-stage surgery) | -1920
    cement spacer in appropriate position | -1920
    fracture of greater trochanter | -1920
    evaluated by vascular surgeon | -1920
    evaluated by cardiologist | -1920
    rivaroxaban discontinued 72 hours pre-surgery | -72
    revision right total hip arthroplasty | 0
    posterior approach | 0
    irrigation and debridement (second surgery) | 0
    removal of antibiotic spacer | 0
    reimplantation of right total hip arthroplasty | 0
    noncemented acetabular component | 0
    2 screws for secondary fixation | 0
    proximal femoral replacement | 0
    estimated blood loss 500 cc | 0
    postanesthesia care unit | 0
    palpable dorsalis pedis pulses (postoperative) | 0
    palpable posterior tibial pulses (postoperative) | 0
    postoperative hemoglobin 7.4 | 0
    preoperative hemoglobin 9.7 | 0
    rivaroxaban reinitiated (postoperative day 1) | 24
    postoperative day 1 hemoglobin 5.8 | 24
    transfused 2 units packed red blood cells | 24
    white blood cell count increased from 15 to 25 | 24
    loose bowel movements | 24
    Clostridioides difficile positive | 24
    started on oral vancomycin | 24
    right lower extremity cool to touch | 24
    no palpable distal pulses | 24
    denied pain | 24
    denied weakness | 24
    denied changes in sensation | 24
    computed tomography angiography | 24
    occlusion of right limb aortobifemoral graft | 24
    emergency thrombectomy | 24
    arterial injury (brachial artery) | 24
    open repair left brachial artery | 24
    open balloon thrombectomy | 24
    intraoperative angiogram confirmed restored blood flow | 24
    extubated | 24
    intensive care unit admission | 24
    heparin drip started | 24
    rivaroxaban held | 24
    heparin stopped | 24
    rivaroxaban restarted | 24
    vascular examination stable | 24
    compartments soft | 24
    discharged to skilled nursing facility | 336
    ambulating with walker | 5760
    ankle-foot orthosis use | 5760
    residual right foot weakness | 5760
    no recurrent infection | 5760
    no compromised blood flow | 5760
    chronic anticoagulation with warfarin | 5760
    