64 years old | 0
male | 0
end-stage liver disease | -672
secondary biliary cirrhosis | -672
non-alcoholic steatohepatitis | -672
robotic cholecystectomy | -1344
hepatic duct leak | -1344
open choledochojejunostomy | -1344
persistently elevated liver function tests | -672
magnetic resonance cholangiopancreatography | -672
choledochojejunostomy stricture | -672
intrahepatic biliary tree dilation | -672
liver biopsy | -672
cirrhosis | -672
chronic biliary obstruction | -672
superimposed non-alcoholic steatohepatitis | -672
liver transplantation | 0
extended two-hepatic vein piggy-back technique | 0
portal vein to portal vein anastomosis | 0
common HA to common HA anastomosis | 0
reconstruction of a small accessory right HA | 0
biliary reconstruction | 0
steroid taper | 0
Myfortic | 0
Tacrolimus | 0
Micafungin | 0
Valcyte | 0
Bactrim | 0
thrombus of the accessory right HA | 24
computed tomography angiography | 24
therapeutic low molecular weight heparin | 24
perihepatic hematoma | 48
percutaneous drain | 48
drain fluid cultures | 48
negative drain output | 48
nonbilious drain output | 48
Apixaban | 192
perihepatic drain removal | 240
sudden onset right upper quadrant abdominal pain | 528
lightheadedness | 528
hemodynamically unstable | 528
tachycardic | 528
hypotensive | 528
abdominal distension | 528
massive transfusion protocol | 528
resuscitation | 528
sepsis protocol | 528
severe lactic acidosis | 528
acute blood loss anemia | 528
acute kidney injury | 528
worsening liver function tests | 528
computed tomography | 528
main HA pseudoaneurysm | 528
active extravasation | 528
hemoperitoneum | 528
endovascular therapy | 528
acute decompensation | 528
pulseless electrical activity | 528
advanced cardiac life support | 528
intubation | 528
right femoral arterial line | 528
REBOA sheath | 528
inflation at zone 1 | 528
MTP resuscitation | 528
cardiopulmonary resuscitation | 528
REBOA inflated | 528
spontaneous cardiac activity | 528
emergency transport | 528
operating room | 528
rapid laparotomy | 528
open abdominal opening | 528
fresh blood clot | 528
hematoma | 528
hepatic hilum | 528
no biloma formation | 528
no bile leak | 528
no enteric leak | 528
no abscess formation | 528
ischemic hepatic allograft | 528
cessation of abdominal aortic perfusion | 528
REBOA deflation | 528
intraabdominal aorta re-perfuse | 528
severe reperfusion injury | 528
recurrent PEA | 528
REBOA re-inflated | 528
ACLS | 528
pulse | 528
donor proper HA thrombosed | 528
damaged | 528
anterior wall of the donor HA ruptured | 528
disintegrated | 528
mycotic change | 528
recipient HA stump ligated | 528
open abdomen negative pressure therapy | 528
surgical intensive care unit | 528
continuous renal replacement therapy | 528
goal directed resuscitation | 528
refractory septic shock | 528
severe acidosis | 528
electrolyte abnormalities | 528
coagulopathy | 528
hepatic ischemic | 528
hemorrhagic insult | 528
Streptococcus Constellatus bacteremia | 528
Klebsiella Pneumoniae colonization | 528
evacuated hematoma | 528
condition decline | 552
refractory septic shock | 552
multiorgan failure | 552
allograft non-function | 552
bradycardic | 542
pulseless | 542
further resuscitative efforts discontinued | 542
pronounced deceased | 542
postmortem preoperative microbiology results | 542
Streptococcus Constellatus bacteremia | 542
Strep Constellatus | 542
Klebsiella Pneumoniae colonization | 542
evacuated hematoma | 542