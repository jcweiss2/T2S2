60 years old | 0
male | 0
admitted to the hospital | 0
biopsy proven PAN | -8760
on prednisone | -8760
on cyclophosphamide | -8760
prior failure on cyclophosphamide alone | -8760
paroxysmal atrial fibrillation | 0
hypertension | 0
not on calcium channels blocker | 0
dyslipidemia | 0
non-insulin dependent diabetes mellitus | 0
multiple prior admissions for PAN flares | -8760
history of an admission for septic shock | -17520
scrotal pain | 0
fever of 103°F | 0
fatigue | 0
tachycardic to 130 beats per minute | 0
hypotensive to 103/40 mm Hg | 0
broad-spectrum antibiotics | 0
vancomycin | 0
Zosyn (piperacillin/tazobactam) | 0
kidney function worsened | 24
switch in antibiotics to meropenem | 24
creatinine level continued to rise | 48
suspicion of acute interstitial nephritis less likely | 48
continued to spike fevers | 48
no specific source of an infection found | 48
no focus found on the CT chest, abdomen, and pelvis | 48
stopping all antibiotics | 48
macular rash | 168
rash progressed slowly | 168
involved axillary area | 168
involved chest, head, neck, and abdomen | 168
decline of mental status | 168
worsening of skin lesions | 168
element of bullae and vesicles | 168
dermatology team involved | 240
biopsy obtained | 240
initiating local steroid cream | 240
diagnosis of AGEP | 240
kidney injury | 240
neutrophilia | 240
cyclic fevers | 240
rash became pustular | 312
high grade fever of 109°F | 312
transfer to the intensive care unit | 312
protocol of cooling | 312
pulse steroids | 312
fever subsided | 336
improvement of the initial rash | 336
decreased progression of sloughing | 336
complete resolution of acute kidney injury | 336
taper in steroids | 336
skin biopsy | 0
urine analysis | 0
CT chest/abdomen/pelvis | 0
CBC/BMP/coagulation | 0
differential diagnosis | 0
Generalized acute pustular psoriasis (von Zumbusch type) | 0
Acute generalized exanthematous pustulosis (AGEP) | 0
Drug reaction with eosinophilia and systemic manifestation (DRESS) | 0
Steven Johnson syndrome | 0
Leukocytoclastic vasculitis | 0
Subcorneal pustular dermatosis (Sneddon–Wilkinson disease) | 0
Cutaneous candidiasis | 0
intra- and subcorneal spongiform | 240
superficial, interstitial, mid-dermal infiltrate rich in neutrophils | 240
dermal edema | 240
tender erythematous nodules | -8760
purpura | -8760
livedo reticularis | -8760
ulcers | -8760
bullous or vesicular eruption | -8760
systemic corticosteroids | 312
withdrawal of the offending drug | 48
supportive care | 0
symptomatic treatment of pruritus and skin inflammation | 0
immunosuppressive management | 336
abstain from using penicillin antibiotics | 336