31 years old | 0
male | 0
asymptomatic | 0
exposure to COVID-19-positive colleague | -336
nasal swab positive for COVID-19 | -336
home quarantine/isolation | -336
admitted to hospital | 0
acute severe left flank pain | 0
mild shortness of breath | 0
nausea | 0
occasional cough | 0
no fever | 0
no dehydration | 0
no vomiting | 0
no change in urinary/bowel habits | 0
mild tenderness in left lumbar region | 0
vital signs stable | 0
elevated inflammatory markers | 0
mild leukocytosis | 0
mildly deranged D-dimer | 0
mildly deranged PT | 0
mildly deranged INR | 0
normal renal functions | 0
no proteinuria | 0
thrombophilia work up negative | 0
hypothyroidism | -672
dyslipidemia | -672
levothyroxine treatment | -672
atorvastatin treatment | -672
sinus tachycardia | 0
rare premature atrial contractions | 0
rare premature ventricular contractions | 0
no intra-cardiac shunt | 0
multiple infarctions at mid and lower poles of left kidney | 0
patent main renal vessels | 0
subpleural patchy ground glass | 0
reticular opacities in lung bases | 0
COVID-19 pneumonia | 0
therapeutic enoxaparin | 0
injectable acetaminophen | 0
no specific treatment for COVID-19-related pulmonary findings | 0
no intubation | 0
no ICU admission | 0
no supplementary oxygen | 0
discharged | 120
follow-up CT abdomen | 432
focal scaring at lower pole of left kidney | 432
warfarin treatment | 120
poor compliance to medical treatment | 432
sub-therapeutic INR | 432
advised to continue warfarin for life-long | 432
no complications reported | 432