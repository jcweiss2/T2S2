22 years old | 0
gravid woman | 0
admitted to the hospital | 0
dysuria | -168
febrile | 0
tachycardia | 0
suprapubic and left-sided costovertebral angle tenderness | 0
sepsis | 0
acute pyelonephritis | 0
leukocytosis | 0
urinalysis was positive for nitrites and leucocytes esterase | 0
urine squamous cell was 4.8/UL | 0
urine WBC was 566.8/UL | 0
urine bacteria was >10000/UL | 0
urinary tract infection [UTI] | 0
urine culture was positive for Escherichia coli [E. coli] | 0
renal ultrasound revealed hyperechoic kidneys | 0
started on intravenous [IV] antibiotics | 0
started on intravenous fluid | 0
blood culture was positive for bacteremia with E. coli | 24
septic shock | 48
hypotension | 48
hypoxic | 48
diffused crackles | 48
intubated | 48
started on norepinephrine infusion | 48
ABG showed PH 7.41/PCO2 33mmHg/PO2 60 mmHg | 48
fetal heart tracings were reassuring | 48
chest x-ray revealed bilateral lung consolidation | 48
severe ARDS | 48
initiate V-V ECMO | 72
pre-ECMO vital signs were blood pressure of 103/72mmHg | 72
oxygen saturation of 75% | 72
respiratory rate [RR] of 18 | 72
body temp of 99.3°F | 72
pulse rate of 102 bpm | 72
right femoral and a right internal jugular vein were placed | 72
cannulas were passed over an Amplatz wire | 72
fetal distress | 75
emergency cesarean section | 75
delivery of a viable neonate | 75
newborn was admitted to the Neonatal Intensive Care Unit | 75
given broad-spectrum antibiotics | 75
mechanical ventilation was reduced to FiO2 of 0.4 | 75
ECMO circuit consisted of a Maquet Rotaflow centrifugal pump | 75
ECMO circuit consisted of a Maquet oxygenator | 75
initial ECMO settings were: pump speed initially was at 1500 revolution per minute [RPM] | 75
flow rate was 4 L per min [LPM] | 75
sweep of 5.5 LPM | 75
patient’s saturation was 96% | 75
monitored for ECMO “chatter” | 75
cannula site was examined daily for migration | 75
anticoagulation for ECMO circuit was performed | 75
hemoglobin level was maintained above 10 g/dl | 75
received a total of 4 units of PRBC while on ECMO | 96
initial ECHO showed an ejection fraction [EF] of 38% | 96
mild left ventricular [LV] dilatation | 96
moderate global and diffuse LV hypokinesis | 96
mild RV dilatation | 96
mild RV dysfunction | 96
no pericardial effusion | 96
successfully weaned off ECMO support | 120
de-cannulated | 120
extubated | 144
chest x-ray showed marked improvement in lung fields | 144
repeat ECHO showed an ejection fraction of 53% | 144
no evidence of hemodynamically significant valve disease | 144
no wall motion abnormality was detected | 144
discharged | 312
no oxygen requirement | 312