73 years old | 0
male | 0
admitted to the hospital | 0
signs of infection at the surgical site on his left hip | 0
avascular necrosis | -175200
staged bilateral total hip arthroplasty | -175200
empty sella syndrome | 0
multiple complications from neurosurgical bleeding | 0
penicillin allergy | 0
adrenal insufficiency | 0
prolonged hospitalization due to drug addiction | 0
aseptic loosening of his left hip | -105120
one-stage revision | -105120
white cell count 5560/mm3 | -105120
erythrosedimentation 43 mm/hr | -105120
ultrasensitive C-reactive protein 10 mg/L | -105120
purulent wound drainage | -105000
elevation of ESR to 33 mm/hr | -105000
elevation of CRP to 20 mg/L | -105000
deep THA infection | -105000
WBC in normal range | -105000
blood glucose levels in normal range | -105000
joint aspiration | -105000
Escherichia coli with resistance to ampicillin | -105000
open debridement and irrigation with prosthetic retention | -105000
administration of antibiotic therapy | -105000
DAIR performed | -105000
deep tissue samples sent for culture | -105000
broad-spectrum antibiotics initiated with intravenous ciprofloxacin | -105000
same germ isolated from intraoperative cultures | -105000
persistent signs of infection | -105000
two DAIR performed | -105000
three weeks postoperatively | -104400
six weeks postoperatively | -103680
Staphylococcus epidermidis cultured in all samples | -103680
six-week course of IV antibiotic therapy with vancomycin and rifampicin | -103680
asymptomatic with no signs of infection | -103680
two episodes of prosthetic dislocation | -105120
WBC 13700/mm3 | -105120
ESR 35 mm/hr | -105120
CRP 108 mg/dL | -105120
instability | -105120
chronic wound infection | -105120
two-stage revision performed | -105120
placement of a cement spacer with antibiotics | -105120
empirical IV meropenem and trimethoprim/sulfamethoxazole administered | -105120
S. epidermidis detected in intraoperative cultures | -105120
six-week course of teicoplanin and ciprofloxacin | -105120
hospitalized for fever | -105120
persistent wound drainage | -105120
WBC 11240/mm3 | -105120
ESR 25 mm/hr | -105120
CRP 137 mg/dL | -105120
new surgical debridement performed | -105120
spacer kept in place | -105120
E. coli detected in intraoperative cultures | -105120
deep vein thrombosis | -105120
intestinal ischemia | -105120
resection of the transverse and small colon | -105120
transferred to the ICU | -105120
persistent signs of infection | -105120
additional surgical debridements performed | -105120
revision of the spacer | -105120
Candida parapsilosis detected in intraoperative samples | -105120
treatment adjusted to include antifungals | -105120
patient's condition improved | -105120
discharged from the hospital | -105120
reactivation of chronic wound infection | -105120
fever | -105120
fistulous lesions | -105120
purulent spontaneous drainage | -105120
WBC 7611/mm3 | -105120
ESR 47 mm/hr | -105120
CRP 36 mg/dL | -105120
revision of the cement spacer | -105120
antibiotic-loaded with vancomycin and liposomal amphotericin B | -105120
methicillin-sensitive S. aureus detected | -105120
E. coli detected | -105120
Acinetobacter baumannii detected | -105120
markers of inflammation normalized | -105120
absence of clinical signs of infection | -105120
second stage of re-implantation arthroplasty performed | -105120
femoral tumor stem | -105120
uncemented porous tantalum cup created with 3D printing | -105120
acetabular defect addressed | -105120
episode of dislocation | -105120
reactivation of chronic infection | -105120
WBC 8455/mm3 | -105120
ESR 32 mm/hr | -105120
CRP 57 mg/dL | -105120
DAIR performed again | -105120
wide resection of necrotic tissue | -105120
retention of all components | -105120
large number of WBC by microscopic analysis | -105120
no microorganisms isolated | -105120
conduct of an overseeding sample resulted in identification of S. maltophilia | -105120
suppressive antibiotic therapy with levofloxacin | -105120
new prosthesis dislocation | -105120
chronically dislocated hip revision prosthesis | -105120
taking suppressive antibiotics for one year | -105120
no signs of reactivation of the chronic infection | -105120
plan on discontinuing suppressive antibiotic therapy | -105120
latest laboratory results showed WBC 7430/mm3 | -105120
ESR 36 mm/hr | -105120
CRP 47 mg/dL | -105120
patient and family decided not to undergo another revision surgery | -105120
