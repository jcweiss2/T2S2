56 years old | 0
female | 0
presented to the ER | 0
fever | 0
painful rash on the hands | 0
abnormal blood culture report indicating growth of yeast | -48
shortness of breath | 0
progressively worsening cough | -336
non-bloody white sputum | -336
subjective fever | -336
chills | -336
hemodialysis through a left-arm arteriovenous graft | 0
hypertension | 0
diabetes mellitus | 0
referred to the hospital | -48
yeast identified in blood cultures | -48
candida zeylanoides identified | -48
obese | 0
alert | 0
comfortable | 0
febrile at 102 °F | 0
blood pressure 156/86 mmHg | 0
oxygen saturation 98% on room air | 0
left-arm arteriovenous graft with good thrill | 0
1-mm violaceous macular lesions on the palm and ventral aspects of 4th and 5th fingers of left hand | 0
basilar crackles | 0
normal heart sounds | 0
no murmurs | 0
hypertensive retinopathy | 0
white hypo-pigmented inferotemporal lesion suggestive of fungal chorioretinitis | 0
leukocytosis with WBC count 1.34 × 104/μL | 0
WBC count increased to 1.82 × 104/μL on day 3 | 72
blood cultures positive for yeast | -48
ultrasound showing fluid collection around arteriovenous graft | 0
fine needle aspiration | 0
culture grew candida zeylanoides | 0
excision of infected arteriovenous graft | 0
temporary Shiley catheter placed for hemodialysis | 0
permanent permacath placed | 0
transesophageal echocardiogram negative for vegetation | 0
chest CT showed peripheral nodular lesions suggestive of infective emboli | 0
bronchoscopy with bronchoalveolar lavage | 0
white exudate | 0
transbronchial biopsy | 0
tissue cultures yielded Candida zeylanoides | 0
negative serum precipitins to Aspergillus fumigatus and Aspergillus niger | 0
started on caspofungin | 0
fluconazole replacement per Infectious disease team recommendations | 0
repeat blood cultures negative for fungal growth | 0
discharged from the hospital | 0
orders to complete 6 weeks of parenteral fluconazole during hemodialysis | 0
completed antifungal therapy as outpatient | 0
followed in dialysis center | 0
