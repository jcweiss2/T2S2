54 years old | 0
female | 0
admitted to the Emergency Department | 0
syncope | 0
hematemesis | 0
smoking habit | -6720
alcohol consumption | -6720
hemodynamically stable | 0
asymptomatic | 0
physical examination anodyne | 0
hemoglobin 10.2 mg/dl | 0
coagulation parameters normal | 0
cranial computed tomography scan | 0
no pathological findings | 0
esophagogastroduodenoscopy | 0
traces of blood in the stomach | 0
uncomplicated hiatal hernia | 0
no active bleeding | 0
in-hospital observation | 0
no hemodynamic instability | 72
several stools compatible with melenae | 72
hemoglobin level stable | 72
esophagogastroduodenoscopy | 48
no traces of blood | 48
no pathological features | 48
discharged | 72
readmitted | 96
syncope | 96
hypotension | 96
heart rate 92 bpm | 96
fluid replacement | 96
hemodynamic stability | 96
hemoglobin 8.4 mg/dl | 96
transfusion of 2 units of packed red blood cells | 96
new episode of melenae | 96
esophagogastroduodenoscopy | 96
pulsatile vessel in the second portion of the duodenum | 96
no active bleeding | 96
irregular fusiform aortic aneurysm | 96
CT scan imaging | 96
aneurysm contacted with the third duodenal portion | 96
extended itself toward the iliac bifurcation | 96
1 cm mural thrombus in the right iliac artery | 96
duodenal AEF originating from the aneurysm | 96
urgent laparotomy | 96
inflammatory infrarenal aortic aneurysm | 96
ligation of both common iliac arteries and infrarenal aorta | 96
vascular perfusion with an axilo-bifemoral bypass | 96
resection of the aortic-jejunal fistula | 96
primary suture repair of the defect | 96
low dose vasoactive drugs | 96
transfusion of 5 additional units of packed red blood cells | 96
admitted to the Intensive Care Unit | 96
favorable evolution | 102
transferred to the ward | 150
discharged | 264
no signs of active bleeding | 264
stable hemoglobin analysis | 264
pathology report of the surgical specimen | 264
AEF with no presence of pathogens | 264
culture positive for gram positive aerobic flora | 264
Streptococcus viridians | 264
coagulase-negative Staphyloccocus | 264
treated with Piperacillin/Tazobactam | 264
follow-up CT scan | 2160
no evidence of recurrent AEF | 2160
good condition | 2160
no further gastrointestinal bleeding | 2160