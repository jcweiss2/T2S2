29 years old | 0
female | 0
Crohn’s disease | -8760
perianal fistula | -8760
Infliximab monotherapy | -8760
peri-anal abscess drainage | -8760
Certolizumab Pegol | -8760
pregnancy | -840
mild peri-anal pain | -120
discharged | -120
worsening pain | -96
admitted | -96
fetal monitoring | -96
colorectal evaluation | -96
anal stricture | -96
white blood cell count of 13 500 | -96
C-reactive protein of 115 mg/L | -96
perineal ultrasound | -96
intravenous ceftriaxone | -96
metronidazole | -96
emergency cesarean section | -72
fetal distress | -72
tachycardia | -60
hypo-tension | -60
perianal pain progressed | -60
diffuse hyperemia | -60
swelling of the vulva | -60
purple discoloration of the skin | -60
Fournier’s gangrene suspected | -60
wide drainage and debridement | -60
necrosis of the ischiorectal fat | -60
foul-smelling purulent discharge | -60
anoscopy | -60
rectal ulcers | -60
fistulous opening | -60
purulent discharge | -60
laparoscopic loop ileostomy | -60
intraoperative colonic lavage | -60
vacuum-assisted therapy | -60
hydrocolloid paste | -60
cultures revealed polymicrobial infection | -48
Eschericia Coli | -48
Citrobacter freundii complex | -48
Candida albicans | -48
antibiotics adjusted | -48
discharged from the Intensive Care Unit | 72
debridements | 72
vacuum-therapy exchanges | 72
perineal defect closed | 336
unilateral medial thigh advancement flap | 336
draining seton | 336
discharged | 672
medial thigh flap completely healed | 1008
Infliximab monotherapy resumed | 1008
ileostomy reversal planned | 1008
baby recovered well | 1008