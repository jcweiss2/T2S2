84 years old | 0
female | 0
admitted to the hospital | -936
Alzheimer's dementia | 0
fever | 0
pulmonary thromboembolism | -936
deep vein thrombosis | -936
blood pressure 87/44 mm Hg | 0
heart rate 105 bpm | 0
body temperature 38.2° | 0
leukocytosis | 0
elevated C-reactive protein | 0
serum lactate level 3.57 mmoL/L | 0
septic shock | 0
methicillin-resistant Staphylococcus aureus bacteremia | 0
contrast-enhanced chest CT | 4
contrast-enhanced abdominal CT | 4
multiple peripheral nodules in both lungs | 4
septic embolism | 4
mild swelling of the thyroid gland | 4
heterogeneous enhancement of the thyroid gland | 4
perithyroidal fluid collection | 4
shock thyroid | 4
admitted to the intensive care unit | 4
glycopeptide antibiotic administered | 4
fluid resuscitation administered | 4
diluted norepinephrine administered | 4
hemodynamically stable | 4
follow-up neck CT | 26
thyroid function tests | 26
normalization of thyroid gland size | 26
normalization of thyroid gland enhancement pattern | 26
resolution of perithyroidal fluid collection | 26
normal serum free thyroxine (T4, 1.23 ng/dL) | 26
normal serum thyroid-stimulating hormone (0.53 mIU/L) | 26
low serum triiodothyronine (T3, 58.5 ng/dL) | 26
moved to the general ward | 96
discharged | 96
