19 years old | 0
male | 0
admitted to the hospital | 0
motor vehicle accident | -2
trauma | -2
shock state | -2
resuscitated | -2
infusion of crystalloids | -2
intra-abdominal complications ruled out | -2
physical exam | -2
ultrasound studies | -2
bilateral epidural hematoma | -1
tachycardic | -1
acceptable blood pressure | -1
premedication with fentanyl | -1
induction of anesthesia | -1
sevoflurane | -1
cisatracurium | -1
cranial decompressive surgery | 0
large intravenous lines malfunctioning | 1
planning for central intravenous catheter | 1
femoral vein catheterization | 2
insertion of introducer catheter | 2
aspiration of catheter lumens | 2
visualization of retrograde flow | 2
infusion of packed RBCs | 2
infusion of crystalloid | 2
infusion of norepinephrine | 2
stable hemodynamic status | 4
transferred to intensive care unit | 4
intubated | 4
abdominal distension | 24
ultrasound findings of fluid in abdominal cavity | 24
laparotomy | 24
misplacement of femoral catheter | 24
extraction of femoral catheter | 24
right inguinal hernia | 24
retroperitoneal blood | 24
iliac vein perforation | 24
bleeding | 24
removal of catheter | 24
patient care at ICU | 48