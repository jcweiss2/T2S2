50 years old | 0
female | 0
relapsing idiopathic membranous nephropathy | -192 months
maculopapular rash | -168 hours
rituximab | -168 hours
complete remission | -192 months
cyclophosphamide | -192 months
prednisolone | -192 months
methotrexate | -192 months
cyclosporine | -192 months
nephrotic syndrome | -28 days
renal biopsy | -28 days
diabetic nephropathy | -28 days
serum antiphospholipase-A2 receptor antibody negative | -28 days
trimethoprim-sulfamethoxazole | -168 hours
metformin | -168 hours
admission to hospital | 0
widespread maculopapular rash | 0
haemodynamically stable | 0
allergic urticaria | 0
prednisolone | 0
cetirizine | 0
promethazine | 0
hypotensive | 24
febrile | 24
tachycardic | 24
generalized myalgias | 24
arthralgias | 24
cervical lymphadenopathy | 24
inotropic support | 24
empirical antibiotics | 24
intravenous hydrocortisone | 24
leucocytosis | 24
lymphocytosis | 24
normal serum eosinophils | 24
normal neutrophils | 24
non-specific reactive leucocytosis | 24
elevated C-reactive protein | 24
low C3 | 24
normal C4 | 24
lactic acidosis | 24
acute kidney injury | 24
urine microscopy | 24
procalcitonin not tested | 24
symptoms resolved | 48
inotropic support weaned | 24
renal function normalized | 48
rituximab-induced serum sickness | 48
antibiotics ceased | 48
hydrocortisone changed to prednisolone | 48
trimethoprim-sulfamethoxazole rechallenged | 48
no issues | 48
outpatient skin allergen testing | 48
discharged home | 72
no recurrence of symptoms | 2160