30 years old | 0
female | 0
pregnant | 0
27 weeks of gestation | 0
admitted to the hospital | 0
5-day history of progressive dyspnea | -120
5-day history of lethargy | -120
5-day history of fever | -120
gravid uterus | 0
treated as bacterial pneumonia | 0
Amoxicillin plus Clavulanate | 0
Clarithromycin | 0
Oseltamivir | 0
no auscultatory findings | 0
chest X-ray showed consolidation | 0
fetal ultrasound had no alteration | 0
transferred to the ICU | 4
started continuous non-invasive ventilation | 4
unsatisfactory clinical and laboratorial response | 7
elective endotracheal intubation | 7
severe hypoxemia | 12
ARDS criteria | 12
neuromuscular blockade | 12
alveolar recruitment | 12
semi-pronation position | 12
veno-venous ECMO installation | 24
preserved cardiac function | 24
echocardiogram | 24
cannulation of the right internal jugular vein | 24
cannulation of the right femoral vein | 24
decision not to interrupt the gestation | 24
fetus viability monitored | 24
betamethasone administered | 24
increased white blood cell count | 96
new culture samples obtained | 96
Piperacillin-Tazobactam | 96
Oseltamivir continued | 96
tracheal aspirates showed Amoxicillin and Clavulanate resistant Enterobacter | 96
Methylprednisolone | 168
significant improvement in lung function | 216
ECMO cessation | 216
extubated | 264
intermittent NIV | 264
ICU discharge | 312
hospital discharge | 504
antenatal evaluation performed regularly | 504
Caesarean section | 1008
delivery of a healthy male infant | 1008