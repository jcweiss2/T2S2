21 years old | 0
female | 0
presented to a tertiary care hospital | 0
history of on and off low-grade fever | -2160
abdominal pain | -168
no history of cough | -2160
no weight loss | -2160
no facial rashes | -2160
conscious | 0
anxious | 0
pale | 0
blood pressure on the lower side of normal | 0
distended abdomen | 0
tuberculosis ruled out | 0
vasculitis like systemic lupus erythematosus ruled out | 0
anti-dsDNA negative | 0
anti-sm-RNA negative | 0
erect X-ray | 0
abdomen ultrasonography | 0
developed septic shock | 72
mean blood pressure <65 mmHg | 72
altered sensorium | 72
intubated | 72
transferred to the intensive care unit | 72
magnetic resonance imaging of head | 72
cerebrospinal fluid study | 72
serum sodium level 137 mmol/L | 72
leukocytosis 21000/cmm | 72
anemia 5 gm/dL | 72
thrombocytopenia 20000/cmm | 72
deranged liver function tests | 72
prothrombin time 6 s prolonged | 72
echocardiography showed mild diastolic dysfunction | 72
ejection fraction >60% | 72
managed conservatively with fluids | 72
sedation | 72
noradrenaline 0.5–3 μg/kg/min | 72
vasopressin 0.01 U/min infusion | 72
broad-spectrum antibiotics | 72
platelet transfusion | 72
packed cell transfusion | 72
blood cultures sterile | 72
endotracheal tube aspirate cultures sterile | 72
repeat ultrasonography of the abdomen | 120
thickened bowel loops | 120
dilated nonobstructed bowel loops | 120
coarse hepatic echo-texture | 120
refused active management | 120
high nasogastric aspirates | 96
feed intolerance | 96
prokinetics use | 96
started accepting nasogastric feeds | 144
enteral feed | 144
developed rapidly rising intraabdominal pressure >18 mmHg | 144
sudden deterioration in hemodynamics | 144
increasing metabolic academia | 144
hyponatremia serum sodium 124 mmol/L | 144
passed large amounts of fresh blood-mixed loose stools | 144
Clostridium difficile negative | 144
bedside abdominal ultrasonography suspected air shadows within the hepatic portal vein | 144
urgent computed tomography scan abdomen | 144
pneumatosis intestinalis of the small bowel | 144
dilated bowel loops | 144
gas in portal venous system | 144
prolonged septic shock | 144
vasopressor support | 144
metabolic acidosis | 144
exploratory laparotomy | 144
multiple areas of gangrenous patches | 144
dusky discoloration of the jejunum | 144
air bubbles in the subserosa | 144
major mesenteric vessels pulsating | 144
no evidence of thrombus | 144
no atherosclerosis | 144
no visible occlusion | 144
no bowel perforation | 144
surgical incisions in the wall of the jejunum | 144
succumbed | 148
postmortem examination not conducted | 148
nonocclusive mesenteric ischemia | 144
