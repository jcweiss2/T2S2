57 years old | 0
female | 0
alpha-1 antitrypsin deficiency | 0
chronic obstructive pulmonary disease | 0
home oxygen | 0
polysubstance use disorder | 0
buprenorphine | 0
severe malnutrition | 0
hemicolectomy | 0
colostomy | -17520
large bowel obstruction | -17520
acute abdominal pain | -96
vomiting | -96
constipation | -96
generalized weakness | -96
slurred speech | -96
black stools | -672
tobacco use | 0
assistance with activities of daily living | 0
clonidine | 0
paroxetine | 0
buprenorphine/naloxone | 0
albuterol/ipratropium inhaler | 0
temperature 36.6°C | 0
heart rate 122 bpm | 0
respiratory rate 22 breaths per minute | 0
blood pressure 155/109 mmHg | 0
oxygen saturation 100% | 0
severe cachectic | 0
BMI 14 kg/m² | 0
abdomen tender to light palpation | 0
ostomy output black | 0
WBC count 27.1 ×10⁹ cells/L | 0
lactate 3.7 mmol/L | 0
urine toxicology positive for cocaine | 0
urine toxicology positive for buprenorphine | 0
fecal occult blood test negative | 0
CT abdomen/pelvis with contrast | 0
small bowel dilatation | 0
small bowel obstruction (SBO) | 0
admitted to surgery service | 0
managed non-operatively | 0
initial improvement | 72
WBC decreased to 13.6 ×10⁹ cells/L | 72
clinical deterioration | 96
WBC increased to 22.4 ×10⁹ cells/L | 120
repeat CT abdomen/pelvis with contrast | 120
pelvic abscess 8.2 ×14.0 ×16.3 cm | 120
persistent SBO | 120
percutaneous transgluteal pigtail catheter placed | 120
purulent, malodorous fluid removed | 120
abscess cultures grew mixed flora | 120
Enterococcus faecium | 120
Candida dubliniensis | 120
ampicillin/sulbactam 3g IV q6h | 120
micafungin 100mg IV q24h | 120
repeat CT abdomen/pelvis | 192
drainage catheter within abscess | 192
bowel rupture | 192
poor surgical candidate | 192
transgluteal drain upsized | 192
confusion | 192
hypothermic | 192
tachycardic | 192
tachypneic | 192
transferred to ICU | 192
sepsis | 192
blood cultures positive for Dietzia cinnamea | 192
antimicrobials continued | 192
improved | 240
repeat blood cultures negative | 240
taken to OR | 336
jejunal enterotomy | 336
jejunojejunal anastomosis | 336
ileocolic anastomosis | 336
abdominal washout | 336
removal of transgluteal drain | 336
cultures of soft tissue | 336
abscess cultures | 336
post-operative confusion | 336
deconditioning | 336
ongoing malnutrition | 336
imaging showed resolution of abscess | 672
antimicrobials completed | 672
discharged | 1344
