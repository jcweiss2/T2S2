75 years old | 0
man | 0
body mass index 24.49 kg·m⁻² | 0
presents to the emergency department | 0
fever | -96
myalgia | -96
dyspnoea | -96
quit smoking | -131040
40 pack-years | -131040
hypertension | -131040
valsartan | -131040
amlodipine | -131040
travelled recently | 0
stayed in a motel | 0
temperature 38.7°C | 0
blood pressure 132/67 mmHg | 0
heart rate 102 beats per min | 0
respiratory rate 24 breaths per min | 0
arterial blood gases analysis | 0
severe hypoxaemia | 0
arterial oxygen tension 47.1 mmHg | 0
arterial carbon dioxide tension 40.9 mmHg | 0
pH 7.464 | 0
HCO3⁻ 28.4 mmol·L⁻¹ | 0
arterial oxygen saturation 84.2% | 0
anaemia | 0
haemoglobin 10.7 g·dL⁻¹ | 0
elevated white blood cells | 0
11420 per μL | 0
92.0% neutrophils | 0
4.6% lymphocytes | 0
elevated C-reactive protein | 0
19.97 mg·dL⁻¹ | 0
hyponatraemia | 0
serum Na+ 127 mmol·L⁻¹ | 0
normal laboratory tests | 0
chest radiograph infiltrates in both lungs | 0
antibiotic therapy with intravenous ampicillin/sulbactam | 0
3 g per 6 h | 0
antiviral therapy with oral oseltamivir | 0
75 mg per 12 h | 0
Legionella urinary antigen test positive | 0
antibiotic therapy changed to moxifloxacin | 0
400 mg per 24 h | 0
haemoptysis | 24
haemodynamic instability | 24
type I respiratory failure | 24
noninvasive ventilation | 24
ABGs PaO2 41.7 mmHg | 24
ABGs PaCO2 40.6 mmHg | 24
ABGs pH 7.427 | 24
ABGs HCO3⁻ 25.9 mmol·L⁻¹ | 24
ABGs SaO2 77.1% | 24
intubated | 24
transferred to respiratory failure unit | 24
chest computed tomography | 24
extensive bilateral infiltrates | 24
blood in bronchial secretions | 24
high oxygenation index 51.3 | 24
increased need for haemodynamic support | 24
renal function deteriorated | 24
creatinine 4.75 mg·dL⁻¹ | 24
haemoglobin 6.7 g·dL⁻¹ | 24
urine sample many red blood cells | 24
160–170 per optical field | 24
severe morphological deterioration indicating glomerular origin | 24
bronchoscopy performed | 24
bronchoalveolar lavage | 24
iron-laden macrophages | 24
microbiology results negative for bacteria | 24
mycobacteria negative | 24
fungi negative | 24
cytology negative for malignancy | 24
transfused with fresh frozen plasma | 24
red blood cells | 24
positive C+ANCA | 24
proteinase+3 150.46 EU·mL⁻¹ | 24
anti+GBM 0.54 U·mL⁻¹ | 24
methylprednisolone 1 g per 24 h i.v. | 24
cyclophosphamide 15 mg·kg⁻¹ | 24
severe diffuse alveolar haemorrhage | 24
respiratory instability | 24
adjustment of mechanical ventilation | 24
plasma | 24
blood transfusion | 24
vasopressor therapy | 24
acute renal failure | 24
Legionella infection | 24
vasculitis | 24
positive C-ANCA | 24
proteinase-3 150.46 EU·mL⁻¹ | 24
anti-GBM 0.54 U·mL⁻¹ | 24
