54 years old | 0
male | 0
shortness of breath | -168
seizure | -168
right lung non-small cell lung cancer | -168
brain metastasis | -168
superior vena caval syndrome | -168
stage IV | -168
phenytoin | -168
dexamethasone | -168
palliative radiotherapy | -168
radiotherapy to the mediastinum | -168
radiotherapy to the whole brain | -168
20 Gray in 5 fractions | -168
Co-60 gamma rays | -168
general condition improved | -14
paclitaxel-carboplatin combination | -14
painful erythematous lesions | -7
afebrile | -7
pulse rate 98/min | -7
respiratory rate 28/min | -7
blood pressure 109/83 mm Hg | -7
mild dehydration | -7
erythematous tender macules | -7
confluent epidermal detachment | -7
blistering | -7
conjunctivitis | -7
hemorrhagic crusting on lips | -7
erosions over buccal and nasal mucosa | -7
erosions over glans penis | -7
hyponatremia | -7
phenytoin discontinued | 0
intravenous fluid replacement | 0
electrolyte correction | 0
systemic antibiotics | 0
dexamethasone 16 mg/day | 0
local skin care | 0
condition worsened | 7
septicemia | 7
death | 7