62 years old | 0
woman | 0
congestive heart failure | 0
type 1 diabetes | 0
hypertension | 0
progressive dysphagia | 0
encephalopathy | 0
acute respiratory failure | 0
admitted to the intensive care unit | 0
intubated | 0
influenza A | 0
bacterial pneumonia | 0
acute respiratory distress syndrome | 48
septic shock | 48
broad-spectrum antibiotics | 48
vasopressors | 48
ejection fraction of 20% | 0
cardiogenic shock | 0
Impella device placed | 0
extracorporeal membranous oxygenation initiated | 0
systemic heparin started | 0
transferred to the cardiac intensive care unit | 0
continuous renal replacement therapy started | 192
anasarca | 192
oliguria | 192
hemodynamic status improved | 288
Impella support weaned off | 288
vasopressors weaned off | 288
hematochezia | 288
hemoglobin level 6.4 g/dL | 288
hemoglobin level 10.3 g/dL | 0
hemoglobin level 8.5 g/dL | 264
upper GI bleeding concern | 288
lower GI bleeding concern | 288
pantoprazole drip started | 288
intravenous fluid resuscitation | 288
packed red blood cells transfused | 288
EGD revealed superficial punctate esophageal ulcers | 288
oozing blood | 288
clotted blood in gastric fundus | 288
hematochezia continued | 312
repeat EGD | 312
metoclopramide received | 312
punctate superficial oozing esophageal ulcers | 312
superficial linear gastric ulcerations | 312
biopsy not performed | 312
heparin infusion | 312
Hemospray applied | 312
cessation of bleeding | 312
hematochezia stopped | 312
Hb stabilized | 312
crusted vesicular lesions on upper lip | 312
crusted vesicular lesions on lateral aspect of tongue | 312
HSV suspected | 312
IV acyclovir started | 312
buccal ulceration swabbed | 312
HSV-1 PCR positive | 312
HSV-1 IgG 4.97 index | 312
HSV IgM not detected | 312
Helicobacter pylori stool antigen negative | 312
Helicobacter pylori serologies negative | 312
blood counts stabilized | 312
repeat EGD performed | 624
normal esophageal mucosa | 624
discharged | 624
