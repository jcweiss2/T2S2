58 years old | 0
male | 0
found on the floor of his apartment | -1
loose bowel movements | -24
denies change in stool color | -24
denies blood in diarrhea | -24
no abdominal pain | -24
no nausea | -24
no vomiting | -24
no recent antibiotics use | -24
no fever | -24
no cough | -24
no chest pain | -24
no dyspnea | -24
not hospitalized within the past year | -8760
never traveled outside the United States | -0
diagnosed with Crohn's disease | -33600
multiple bowel resections | -33600
not on steroids | 0
treated with Vedolizumab | -576
treated with infliximab | -576
stopped infliximab | -576
physical examination showed emaciated patient | 0
blood pressure 78/50 | 0
heart rate 98 | 0
respiratory rate 22 | 0
temperature 99° F | 0
lung exam showed crackles over the right lung | 0
abdominal exam were unremarkable | 0
cardiovascular exam were unremarkable | 0
elevated WBCs count | 0
chest X ray with multiple opacities in the right lung field | 0
IgE level was 205 | 0
HIV was negative | 0
admitted to intensive care unit | 0
septic shock caused by pneumonia | 0
started on Vancomycin | 0
started on Aztreonam | 0
started on Levofloxacin | 0
started on vasopressors | 0
clinical picture didn't improve | 24
sputum and blood cultures were negative | 24
CT of the chest | 72
opacification within the entirety of the right lung with air bronchograms | 72
bronchoscopy | 96
normal mucosa without lesions in the upper and lower airways | 96
bronchoalveolar lavage | 96
cultures were negative for bacteria | 96
cultures were negative for tuberculosis | 96
cultures were negative for fungi | 96
bronchial washing cytology showed acute inflammation | 96
filariform larvae | 96
serology was positive for Strongyloides antibodies | 96
started on ivermectin | 96
condition improved significantly | 120
discharged in good condition | 168