28 years old| 0
male | 0
farmer | 0
presented with ingestion of two fresh tablets of Celphos (AlP) | -4
vomiting | -4
pain in the abdomen | -4
agitated | -4
anxious | -4
irritable | -4
pulse rate not palpable | -4
blood pressure not recordable | -4
heart rate 110/min | -4
respiratory rate 28/min | -4
oxygen saturation 95% | -4
ECG shows sinus tachycardia | -4
T wave inversion in lead 3 | -4
managed with IV crystalloids | -4
IV magnesium sulphate 1 gm stat and 8 hourly | -4
IV calcium gluconate 8 hourly | -4
IV hydrocortisone 100 mg stat and 12 hourly | -4
IV dopamine | -4
noradrenaline | -4
immediate gastric lavage performed with potassium permanganate | -4
activated charcoal kept in the stomach | -4
activated charcoal repeated 8 hourly | -4
routine investigations normal at admission | 0
arterial blood gas analysis shows metabolic acidosis | 0
pH 7.2 | 0
HCO3 8 mmol/L | 0
PCO2 33 mmol/L | 0
metabolic acidosis correction performed | 0
intubated | 0
shifted to ICU | 0
BP 60-80 mmHg systolic at 6 hours | 6
PR 120/min at 6 hours | 6
RR 20/min at 6 hours | 6
input/output 3L/300 ml over next 24 hours | 24
developed monomorphic ventricular tachycardia on day 2 | 48
DC cardio-version of synchronised 150 J | 48
converted to NSR | 48
IV amiodarone 150 mg bolus | 48
IV amiodarone infusion continued till next 48 hours | 48
NSR maintained till discharge | 48
cardiac biomarkers raised on day 2 | 48
cardiac biomarkers normalised by day 14 | 336
BP 70/50 mmHg to 90/60 mmHg till day 4 | 96
blood urea 100 mg/dl on day 4 | 96
serum creatinine 4.5 mg/dl on day 4 | 96
urine output 400 ml/24 hours on day 4 | 96
AST/ALT 80/90 IU/L on day 4 | 96
ALP 200 U/L on day 4 | 96
S bilirubin 2.5 mg/dl on day 4 | 96
BP 100/70 mmHg on day 5 | 120
PR 110/min on day 5 | 120
RR 22/min on day 5 | 120
TLC 14000/mm3 with polymorphonuclear leucocytosis on day 5 | 120
urea 200 mg/dl on day 5 | 120
S. creatinine 7.5 mg/dl on day 5 | 120
urine output 400 ml/24 hours on day 5 | 120
ABG pH 7.1 on day 5 | 120
ABG HCO3 10 mmol/L on day 5 | 120
haemodialysis performed on day 5 | 120
haemodialysis performed on day 7 | 168
blood urea 70 mg/dl after day 7 haemodialysis | 168
creatinine 4.0 mg/dl after day 7 haemodialysis | 168
urine output 1200 ml/24 hours after day 7 haemodialysis | 168
extubated on day 6 | 144
shifted to SDU on day 8 | 192
vitals normal | 192
liver functions improving | 336
kidney functions improving | 336
liver and kidney functions near normal by day 14 | 336
discharged on day 14 | 336
