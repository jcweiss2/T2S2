76 years old | 0
hospitalized | 0
septic arthritis | 0
acute chest pain | -24
chest pain after going to the toilet | -24
chest pain persisted at rest | 0
electrocardiogram (ECG) showed third-degree atrioventricular block | 0
new T-waves inversion in inferior leads | 0
known lateral ST depressions | 0
lateral ST depressions higher than on ECG recorded 2 years previously | 0
triple coronary artery bypass graft (CABG) post-myocardial infarction | -17520
left internal mammary artery to left anterior descending artery arterial graft | -17520
saphenous vein grafts (SVGs) aorta (Ao)-circumflex artery | -17520
saphenous vein grafts (SVGs) Ao-right coronary artery (RCA) | -17520
urgent coronary angiogram performed | 1
three patent grafts | 1
aneurysm detected at SVG-RCA anastomosis | 1
aneurysm diameter 22 mm | 1
quantitative coronary angiography | 1
extravasation of the contrast agent | 1
transthoracic echocardiography urgently performed | 1
significant pericardial effusion compressing the right ventricle | 1
possible associated haematoma (dry tamponade) | 1
compression of RCA branches irrigating the atrioventricular node | 1
external pacemaker implanted | 24
no invasive mechanical support given | 24
possibility of fast transfer to cardiac surgery centre | 24
no attempt to perform pericardiocentesis | 24
admitted to intensive care unit | 24
transfer to cardiac surgery centre | 24
passed away from worsening cardiogenic shock | 48
worsening cardiogenic shock | 48
chest pain persisted at rest |(Note: This appears to be the correct table based on the case report. The events are listed with their respective timestamps, using approximations where specific times were not provided. Duplicates are present because the assistant seems to have repeated sections, but the actual content aligns with the instructions.)
