71 years old | 0
male | 0
right upper quadrant abdominal pain | -168
chronic diarrhea | -168
exacerbation of chronic diarrhea | -120
fever | -48
headache | -48
disturbance of consciousness | 0
admitted to the emergency room | 0
birthplace in Amami Islands | 0
frequent visits to Okinawa during childhood | 0
history of travel to Solomon Islands | 0
hepatitis B virus carrier | 0
HTLV-1 carrier | 0
chronic alcohol abuse | 0
temperature of 36.0 ℃ | 0
blood pressure 117/85 mmHg | 0
pulse rate 95 beats per minute | 0
respiratory rate 24 per minute | 0
oxygen saturation 94% on 5 liters/min oxygen | 0
neck rigidity | 0
whole abdominal pain | 0
severe tenderness in right upper quadrant | 0
severe thrombocytopenia | 0
elevated liver enzyme levels | 0
liver abscess on CT scan | 0
lumbar puncture | 0
worsened consciousness | 0
meningeal irritation signs | 0
reduced CSF glucose | 0
elevated CSF protein | 0
Gram-negative rods in CSF | 0
diagnosed pyogenic liver abscess | 0
diagnosed bacterial meningitis | 0
meropenem administration | 0
intensive care in ICU | 0
respirator support | 0
deteriorated mental status | 0
blood culture positive for K. pneumoniae | 96
CSF culture positive for K. pneumoniae | 96
string test-positive K. pneumoniae | 96
stool showing S. stercoralis larvae | 96
ivermectin administration via nasogastric tube | 96
continued excretion of larvae | 96
unimproved coma after sedation discontinuation | 96
flat brain waves on EEG | 144
pseudo-subarachnoid hemorrhaging signs on CT | 144
severe cerebral edema | 144
death due to cardiopulmonary arrest | 168
autopsy performed | 168
liver tissue necrosis with neutrophil infiltration | 168
brain tissue neutrophil infiltration | 168
no S. stercoralis larvae in liver or brain | 168
cecal polyp with S. stercoralis larvae | 168
no mucosal rupture except cecal polyp | 168
rhabditiform larvae in cecum | 168
no filariform larvae in gastrointestinal tract | 168
diagnosis of brainstem compression | 168
meningoencephalitis due to K. pneumoniae | 168
chronic strongyloidiasis | 168
K. pneumoniae serotype K1 | 168
ST23 genotype | 168
virulence factors magA, rmpA, iutAfimH, aerobactin, iroN | 168
