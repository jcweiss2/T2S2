72 years old | 0
male | 0
hypertension | 0
alcohol abuse | 0
acute change in mental status | -168
unsteady gait | -168
meningitis twelve years prior | -105120
acting oddly | -168
febrile | 0
tachycardic | 0
head imaging unremarkable | 0
chest imaging unremarkable | 0
left band shift | 0
no leukocytosis | 0
fever | 0
nuchal rigidity | 0
altered mental status | 0
lumbar puncture | 0
increased CSF total protein | 0
increased CSF WBC | 0
increased CSF neutrophils |) 0
decreased CSF glucose | 0
admitted to ICU | 0
septic shock | 0
intravenous ceftriaxone | 0
intravenous vancomycin | 0
intravenous dexamethasone | 0
Streptococcus pneumoniae speciation | 24
completed antibiotic therapy | 336
recurrent meningitis | 0
alcoholism | 0
no predisposing infection | 0
negative HIV 4th Generation test | 0
negative ANA screen | 0
elevated total protein | 0
low albumin | 0
mild anemia | 0
elevated serum creatinine | 0
unprovoked pneumococcal infection | 0
increased monoclonal gammopathy | 0
elevated IgG | 0
elevated β2-microglobulin | 0
no osseous lytic lesions | 0
normal serum calcium | 0
hypercellular bone marrow | 0
monoclonal IgG lambda restricted plasma cells | 0
multiple myeloma diagnosis | 0
transferred to acute rehab | 504
neurological deficits | 504
fevers | 504
leukocytosis | 504
transferred back to inpatient medical floor | 504
broad-spectrum antibiotics | 504
sepsis of unknown source | 504
Candida auris in blood cultures | 504
intravenous micafungin | 504
negative subsequent cultures | 840
delayed chemotherapy start | 840
resolved active infections | 840
induction chemotherapy with CyBorD regimen | 840
changed chemotherapy regimen to lenalidomide, bortezomib, and dexamethasone | 840
complete remission | 840
no recurrent infections | 840
