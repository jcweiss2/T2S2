68 years old | 0 | 0 
male | 0 | 0 
type 1 diabetic | 0 | 0 
hypertensive | 0 | 0 
on amlodipine | 0 | 0 
operated for treatment of right inguinal hernia | -7200 | -7200 
admitted to the emergency room | 0 | 0 
abdominal pain | -72 | 0 
ketoacidosis decompensation | -72 | 0 
uremic syndrome | -72 | 0 
conscious patient | 0 | 0 
hemodynamically stable | 0 | 0 
dyspneic | 0 | 0 
febrile at 39,6 °C | 0 | 0 
right lumbar tenderness | 0 | 0 
oliguric | 0 | 0 
diuresis at 300 ml/24h | 0 | 0 
altered renal function | 0 | 0 
creatinine at 92 mg/l | 0 | 0 
urea at 3,1 g/l | 0 | 0 
K+ at 6.9 mmol/l | 0 | 0 
Na+ at 123 mmol/l | 0 | 0 
blood sugar at 6.5 g/l | 0 | 0 
alkaline reserves at 8 mEq/l | 0 | 0 
infectious syndrome | 0 | 0 
CRP at 418 mg/l | 0 | 0 
white blood cells at 26000/ml | 0 | 0 
hemoglobin at 12,3 g/dl | 0 | 0 
leucocyturia 320,000 | 0 | 0 
hematuria at 120,000 | 0 | 0 
single anatomical right kidney | 0 | 0 
emphysematous pyelonephritis | 0 | 0 
renal abscess | 0 | 0 
pneumoperitoneum | 0 | 0 
admitted to intensive care | 0 | 0 
dialysis sessions | 0 | 72 
insulin therapy | 0 | 72 
antibiotic therapy | 0 | 48 
ceftriaxone | 0 | 48 
metronidazole | 0 | 48 
surgical drainage of abscesses | 48 | 48 
right double J stent | 48 | 0 
favorable evolution | 48 | 120 
decrease of the infectious syndrome | 48 | 120 
apyrexia | 48 | 48 
chronic renal failure | 120 | 0 
creatinine plateau of 20 mg/l | 120 | 0 
discharged | 240 | 240 
oral antibiotics | 240 | 0 
abdominopelvic CT | 672 | 672 
clear regression of the bubbles of air | 672 | 672 
double J catheter removed | 1008 | 1008