35 years old | 0
male | 0
admitted to the hospital | 0
left leg pain | -24
redness | -24
swelling | -24
visited the Department of Dermatology | -24
focused enhanced computed tomography | -24
cellulitis | -24
Cefdinir | -24
symptoms deteriorated | -12
re-visited the Department of Dermatology | -12
biochemistry analysis | -12
multiple organ dysfunction | -12
history of recurrent cellulitis | 0
obese since childhood | 0
employed in home demolition | 0
Glasgow Coma Scale score 15 | 0
blood pressure 174/65 mmHg | 0
heart rate 108 beats per minute | 0
respiratory rate 30 breaths per minute | 0
SpO2 98% | 0
body temperature 36.7℃ | 0
redness | 0
swelling | 0
tenderness | 0
venous gas analysis | 0
pH 7.352 | 0
PCO2 28.8 mmHg | 0
PO2 61.7 mmHg | 0
HCO3- 15.5 mmol/L | 0
lactate 6.2 mmol/L | 0
electrocardiogram | 0
sinus tachycardia | 0
chest roentgenogram | 0
cardiac enlargement | 0
biochemical analysis | 0
white blood cell count 6800/μL | 0
neutrophil 96% | 0
lymphocyte 2% | 0
monocyte 2% | 0
hemoglobin 14.0 g/dL | 0
platelet count 9.0×10^4/μL | 0
C-reactive protein 12.8 mg/dL | 0
aspartate aminotransferase 315 IU/L | 0
alanine aminotransferase 93 IU/L | 0
glucose 78 mg/dL | 0
blood urea nitrogen 26.0 mg/dL | 0
creatinine level 1.34 mg/dL | 0
creatinine phosphokinase 9670 IU/L | 0
activated partial thromboplastin time 38.7 s | 0
international normalized ratio of prothrombin time 1.83 | 0
fibrinogen 261 mg/dL | 0
fibrinogen degradation product 21.4 mg/dL | 0
sepsis | 0
multiple organ failure | 0
left leg infection | 0
Ringer's lactate | 0
linezolid | 0
meropenem | 0
tracheal intubation | 0
surgical exploration | 12
necrotic soft tissue infection | 12
left leg amputation not performed | 12
oligouria | 24
renal replacement therapy not performed | 24
died of multiple organ failure | 96
culture of surgical material | 96
Streptococcus dysgalactiae | 96
blood culturing not performed | 0