57 years old | 0
woman | 0
generalized anxiety disorder | -4320
choreiform movements | -168
presented to Emergency Department | 0
oral bleeding | -24
vaginal bleeding | -24
anxiety with worsening in the last 8 months | -5760
chorea diagnosed 46 days prior | -1104
choreiform movements worsened over the past 3 days | -72
levetiracetam 750 mg twice daily | -168
valproic acid 250 mg 3 times daily | -168
admitted 7 weeks prior for traumatic subacute right frontoparietal subdural hematoma | -1176
methicillin-susceptible Staphylococcus aureus bacteremia | -1176
Glasgow Coma Scale 15 | -1176
choreiform movements of arms, legs, and trunk | -1176
involuntary movements started 6 months prior | -4320
family history of abnormal movements | -4320
dystonia ruled out | -1176
denial of antipsychotic use | -1176
denial of antidepressant use | -1176
evaluation for hereditary hemochromatosis | -1176
evaluation for malignancy | -1176
evaluation for vasculitis | -1176
evaluation for Wilson’s disease | -1176
evaluation for atypical parkinsonism | -1176
evaluation for Pantothenate kinase-associated neurodegeneration | -1176
evaluation for Huntington’s disease | -1176
initiation of clonazepam 0.5 mg twice daily | -1176
initiation of levetiracetam 250 mg twice daily | -1176
increased levetiracetam to 750 mg twice daily | -1176
increased clonazepam to 0.5 mg 3 times daily | -1176
valproic acid 250 mg 3 times daily added on prior hospitalization day 22 | -1176
platelet count 139,000 μL prior to VPA initiation | -1176
platelet count 90,000 μL at VPA initiation | -1176
discharge with genetic testing outpatient | -1176
GCS 15 at discharge | -1176
platelet count 122,000 μL at discharge | -1176
clonazepam 0.5 mg twice daily at discharge | -1176
levetiracetam 750 mg twice daily at discharge | -1176
valproic acid 250 mg 3 times daily at discharge | -1176
blood pressure 131/91 mm Hg | 0
heart rate 120 beats/min | 0
respiratory rate 16 breaths/min | 0
temperature 36.5°C | 0
GCS 15 on admission | 0
atraumatic contusions | 0
ecchymosis throughout chest | 0
ecchymosis throughout abdomen | 0
ecchymosis throughout back | 0
ecchymosis throughout upper extremities | 0
ecchymosis throughout lower extremities | 0
ecchymosis in left periorbital area | 0
clonazepam discontinued post-discharge | -168
CT head showing left temporal frontal subdural hematoma | 0
acute subdural hematoma along interhemispheric falx | 0
mass effect on right lateral ventricle | 0
3 mm right-to-left midline shift | 0
large-amplitude choreiform movements | 0
admitted to intensive care unit | 0
white blood cells 14.6×10⁶/µL | 0
red blood cells 2.75×10⁶/µL | 0
platelets 4,000/μL | 0
hemoglobin 7.3 g/dL | 0
hematocrit 23.1% | 0
prothrombin time 15.7 seconds | 0
partial thromboplastin time 30.4 seconds | 0
fibrinogen 467 mg/dL | 0
valproic acid level 26.3 μg/mL | 0
valproic acid held on admission | 0
hematology data 15 days prior within normal limits | -360
decreased maximum amplitude on TEG 33.4 mm | 0
evaluation for disseminated intravascular coagulation | 0
evaluation for heparin-induced thrombocytopenia | 0
positive heparin-PF4-related antibody | 0
negative serotonin release assay | 0
no heparin therapy in prior admission | -1176
VPA level decreased to <10 μg/mL on hospital day 2 | 48
fibrinogen decreased to 367 mg/dL | 48
hemoglobin decreased to 5.3 g/dL | 48
CT head stable subdural hematomas | 48
mild improvement in midline shift | 48
hematology consultation on hospital day 1 | 24
methylprednisolone 60 mg intravenous 3 times daily | 24
acute decrease in platelet count on hospital day 4 | 96
intravenous immune globulin 1 g/kg ordered | 96
VPA discontinued | 0
clonazepam not re-initiated | 0
levetiracetam continued | 0
platelet counts improved over next 3 weeks | 504
altered mental status | 0
urinary tract infection | 0
Escherichia coli bacteremia | 0
sepsis | 0
discharged on hospital day 21 | 504
platelet count 108,000 at discharge | 504
GCS 14 at discharge | 504
