29 years old | 0
female | 0
admitted to the ICU | 0
high fever | -72
signs of damage to multiple organs | -72
caesarian section | -72
G1 P0 A1 | 0
pregnancy at 37 wk and 6 d | -216
hip position | -216
labor admission | -216
breeched position of the fetus | -72
spinal anesthesia | -72
healthy baby delivered | -72
fever | -24
peak body temperature of 38.4 °C | -24
chills | -48
shortness of breath | -48
intermittent tingling on both sides of the lower abdomen | -48
abdominal distension | -48
temperature of 40 °C | -48
heart rate of 115 beats/min | -48
blood pressure of 147/84 mmHg | -48
respiratory rate of 20 times/min | -48
oxygen saturation of 92% | -48
white blood cells 10.29 × 10^9/L | -72
white blood cells 14.83 × 10^9/L | -24
neutrophils 83.2% | -24
lymphocytes 9.9% | -24
procalcitonin of 5.19 μg/L | -48
Gram-negative bacteria detected in blood culture | -48
intestinal obstruction | -48
upper gastrointestinal bleeding | -48
pulmonary embolism | -48
CT-scan with contrast | -48
multiple small intestine and colorectal expansion | -48
abdominal and pelvic effusion | -48
peritonitis | -48
increased uterine volume | -48
intermixed high and low intrauterine density | -48
shadow of a partial filling defect in the bilateral lower pulmonary artery | -48
gastrointestinal decompression | -48
coffee-color liquid came out of the gastric tube | -48
post-vaginal dome puncture | -48
light-yellow ascites | -48
latent blood experiment positive | -48
gastrointestinal bleeding confirmed | -48
white blood count > 20.00 × 10^9/L | -24
wheeze | -96
SpO2 68% | -96
disseminated intravascular coagulation | -96
fibrinogen 4.03 g/L | -96
D-dimer determination 23.70 mg/L FEU | -96
fibrin degradation products 59.53 mg/mL | -96
antithrombin III 56.20% | -96
increased serum sodium ion concentration of 164 mmol/L | -96
C. kerstersii detected by mNGS | -48
C. kerstersii detected by blood culture | -48
clindamycin treatment | -48
levofloxacin treatment | -48
metronidazole treatment | -48
piperacillin-tazobartan treatment | -48
meropenem treatment | 0
low-molecular-weight heparin treatment | 0
rehydration | 0
body temperature returned to normal | 96
respiratory rate returned to normal | 96
heart rate returned to normal | 96
oxygenation of the lung returned to normal | 96
gastrointestinal bleeding stopped | 96
abdominal distension relieved | 96
gastrointestinal function recovered | 96
transferred back to the obstetrics department | 96
symptoms completely relieved | 168