54 years old | 0
male | 0
admitted to the Accident and Emergency Department | 0
ventral hernia | -720
ventral hernia increased in size | -672
ventral hernia became stony, hard, painful, and irreducible | -168
vomiting | -168
absolute constipation | -168
road traffic accident | -175200
dysarthria | -175200
socially inactive | -175200
dehydrated | 0
pulse rate of 104 beats/minute | 0
blood pressure within normal range | 0
huge ventral hernia (25x30 cm) | 0
tense and tender | 0
bulging more on right abdomen | 0
skin discoloration | 0
bowel sounds not audible | 0
rectal examination unremarkable | 0
leukocytosis | 0
chest x-ray no air under diaphragm | 0
abdominal x-ray dilated bowel loops with few air fluid levels | 0
diagnosis of strangulated ventral hernia | 0
resuscitation with isotonic fluids | 0
intravenous cefuroxime | 0
intravenous metronidazole | 0
shifted for operation within 2 hours from presentation | 0
laparotomy | 0
entire small bowel and part of large bowel protruding in hernial sac | 0
hemorrhagic fluid | 0
constriction at abdominal wall | 0
pressure over mesentery | 0
tight neck of sac (5x5 cm) | 0
hernial sac opened | 0
offensive fluid | 0
gangrenous bowel | 0
gangrenous mesentery | 0
gangrenous omentum | 0
hemorrhagic fluid shower upon opening sac | 0
gangrenous jejunum | 0
gangrenous ileum | 0
gangrenous cecum | 0
gangrenous ascending colon | 0
gangrenous proximal half of transverse colon | 0
constriction divided | 0
viability trial (100% oxygen, warm sponging) | 0
clear demarcation line established | 0
gut totally black | 0
gut foul smelling | 0
gut lost sheen and luster | 0
no peristalsis | 0
mesentery black | 0
mesenteric vessels gangrenous | 0
patient condition not good during anesthesia/surgery | 0
decision to resect gangrenous bowel | 0
decision to resect gangrenous omentum | 0
gangrenous sac excised | 0
60 cm proximal jejunum remaining | 0
anastomosis to transverse colon | 0
primary anastomosis | 0
direct hernia repair without mesh | 0
histopathology gangrenous bowel with clear margins | 0
postoperative course uneventful | 0
total parenteral nutrition (TPN) | 0
enteral feeding | 0
episodes of diarrhea | 0
enteral feed increased gradually | 0
discharged from hospital | 720
short bowel syndrome | 720
combination enteral and normal diet | 720
mixed consistency stool 4-5 times/day | 720
weight loss 30 kg | -2160
dietary issues managed with dietitian | 720
