34 years old | 0
female | 0
African | 0
admitted to the hospital | 0
fever | -168
new painful blisters | -168
rash | -168
HIV infection | -8760
Combivir | -8760
Kaletra | -8760
supportive care | -120
pain relieving medications | -120
vitamins | -120
micronutrients | -120
acetylsalicylic acid | -120
acetaminophen | -120
consulted a general practitioner | -120
cefuroxime | -96
azithromycin | -96
fluconazole | -96
rash began | -96
rash expanded | -72
painful blisters | -72
higher fevers | -72
malaise | -72
conscious | 0
oriented | 0
normotensive | 0
sinus tachycardia | 0
dry lips | 0
dry tongue | 0
dehydration | 0
conjunctival injection | 0
no abnormalities in chest examination | 0
no abnormalities in abdominal examination | 0
blisters | 0
TEN suspected | 0
dermatologist consulted | 0
burn surgeon consulted | 0
transferred to ICU | 0
central venous access secured | 0
fluid resuscitation initiated | 0
former antimicrobial therapy stopped | 0
CRP increased | 0
leucocytes not increased | 0
serum protein elevated | 0
LDH concentration elevated | 0
no pathological findings in chest X-ray | 0
cultures of blood, urine and wound unrevealing | 0
blisters disinfected | 0
blisters covered with Acticoat | 0
dressings changed every 3 days | 0
intermittent high fever | 0
Avalox started | 0
Ecalta started | 0
former anti-viral HIV therapy continued | 0
polymerase chain reaction testing for viruses | 72
dengue virus DNA detected | 72
antimicrobials stopped | 120
fever decreased | 120
wounds recovered | 120
discharged | 432
follow-up examination | 432
no secondary deficits | 432