79 years old | 0
female | 0
ventilator use | 0
transferred to ICU | 0
biliary sepsis | 0
treated with combined antibiotics | -168
supportive treatment | -168
severely ill | 0
jaundiced | 0
heart problems | 0
hypothyroidism | 0
diabetes mellitus | 0
high total bilirubin (10.94 mg/dL) | 0
high direct bilirubin (9.67 mg/dL) | 0
high CRP (269.48 mg/L) | 0
abdominal ultrasound | 0
MRI evaluation | 0
large cyst (14.7 × 6.2 cm) in left liver lobe | 0
gastric compression | 0
bile duct obstruction | 0
large stone in distal CBD | 0
piperacillin-tazobactam | 0
amikacin | 0
levothyroxine | 0
insulin therapy | 0
supportive treatments | 0
MRI review by senior radiologist | 0
large cyst possibly pancreatic pseudocyst | 0
decision for biliary drainage | 0
bedside PTBD in ICU | 0
transabdominal US guidance | 0
bile fluid aspiration | 0
guide wire insertion | 0
PTBD pigtail catheter insertion | 0
bile fluid from drain catheter | 0
catheter fixation | 0
cyst aspiration | 0
dark-brown cyst fluid | 0
infected cyst | 0
cyst fluid amylase (42 U/L) | 0
cyst fluid lipase (125 U/L) | 0
cyst fluid CEA (476.55 ng/mL) | 0
decreased bilirubin (3.38 mg/dL) | 144
decreased CRP (180.93 mg/L) | 144
breathing improvement | 144
ventilator mode change (CMV to CPAP) | 144
pigtail catheter dislodgement | 144
ERCP procedure | 144
cholangiogram showing large stone | 144
7-Fr double-pigtail stent placement | 144
EUS cyst evaluation | 144
difficult puncture location | 144
19-G FNA needle puncture | 144
guide wire insertion into cyst | 144
6-Fr cystotome use | 144
7-Fr double-pigtail stent insertion into cyst | 144
patient condition improvement | 144
spontaneous breathing | 144
discharge from ICU | 144
discharge from hospital | 168
repeat ERCP for CBD stone crushing | 720
SpyGlass Cholangioscopy DS System use | 720
pancreatic cyst size reduction | 720
pancreatic cyst stent maintained | 720
pancreatitis | 0
biliary obstruction | 0
acute pancreatitis | 0
chronic pancreatitis | 0
gallstone disease | 0
acute gallstone pancreatitis | 0
pancreatic fluid collection | 0
potential complications | 0
cyst fluid leakage | 0
multidisciplinary expert center | 0
