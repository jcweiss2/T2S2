46 years old | 0
male | 0
ulcerative colitis | 0
malaise | -72
fever | -72
loss of appetite | -72
admission to hospital | 0
blood pressure 124/46 mmHg | 0
heart rate 122 beats per min | 0
SpO2 98% | 0
respiratory rate 16/min | 0
body temperature 40.2°C | 0
alert | 0
chills | 0
nausea | 0
cardiac arrest | 0
chest compression | 0
tracheal intubation | 0
ventricular fibrillation | 0
defibrillation | 0
adrenaline administration | 0
resuscitation | 0
diagnosis of Brugada syndrome | 0
coved-type ST elevation in V1 and V2 | 0
hypercalcemia | 0
acetaminophen administration | 0
fever subsided | 0
improvement of coved-type ST elevation | 0
hypotension | 12
septic shock | 12
tazobactam-piperacillin administration | 12
vasopressors administration | 12
extubation | 48
fever reoccurrence | 120
liver abscess | 120
meropenem administration | 120
vancomycin administration | 120
puncture drainage | 120
infection control | 720
pilsicainide test | 720
implantable cardioverter defibrillator implantation | 720
discharge | 720
family history of sudden death | 0
high parathyroid hormone levels | 720
abnormal uptake in the anterior mediastinum | 720
tumor resection | 720
pathological diagnosis of ectopic parathyroid adenoma | 720
nonfunctional pituitary adenoma | 720
nonfunctional adrenal tumor | 720
multiple endocrine neoplasia type 1 | 720
electrocardiogram on October 4, 2021 | -365
electrocardiogram on June 28, 2021 | -365
electrocardiogram on March 24, 2021 | 0
electrocardiogram on September 25, 2017 | -1536