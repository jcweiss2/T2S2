75 years old | 0
    female | 0
    multiple left renal calculi | 0
    right upper ureteric calculus | 0
    abdominal X-ray | 0
    sonography | 0
    left PCNL | -48
    tract dilatation | -48
    severe bleeding | -48
    percutaneous nephrostomy drainage tube placed | -48
    clamped | -48
    transferred to our hospital | -24
    hemodynamically unstable condition | 0
    resuscitated | 0
    blood products transfused | 0
    emergency exploration deferred | 0
    acute kidney injury | 0
    serum urea 105 mg/dL | 0
    serum creatinine 5.77 mg/dL | 0
    noncontrast CT abdomen | 0
    PNDT traversing renal parenchyma | 0
    suspicion tip of PNDT in renal vein | 0
    hemodialysis | 0
    refractory hyperkalemia | 0
    electrocardiogram changes | 0
    bilateral urinary diversion planned | 0
    cystoscopy | 24
    right-sided double-J stent placed | 24
    left percutaneous nephrostomy placed | 24
    sepsis resolved | 24
    AKI resolved | 24
    CT renal angiography | 96
    dynamic renal scan | 168
    position of PNDT in renal vein confirmed | 96
    secondary thrombosis | 96
    no uptake in left kidney | 168
    left nephrectomy planned | 168
    laparoscopic left simple nephrectomy | 192
    thrombectomy | 192
    dense adhesions between mesocolic fat and Gerota's fascia | 192
    two renal arteries | 192
    tip of PNDT in renal vein | 192
    thrombus extending up to interaortocaval groove | 192
    renal arteries clipped | 192
    renal vein dissected in aortocaval groove | 192
    renal vein clipped | 192
    PNDT removed | 192
    no intraoperative complications | 192
    operative time 125 min | 192
    direct tract from renal cortex into renal vein | 192
    intra-abdominal drain removed | 240
    discharged | 288
    right ureteroscopic lithotripsy planned | 288
