80 years old | 0
female | 0
admitted to the intensive care unit | 0
dyspnea | -96
lethargy | -96
chest tightness | -96
denied cough | 0
denied hemoptysis | 0
denied fever | 0
denied gastrointestinal symptoms | 0
denied recent sick contacts | 0
denied traveling | 0
end-stage renal disease | 0
hypertension | 0
hemodialysis | 0
severe pulmonary hypertension | 0
chronic obstructive pulmonary disease | 0
former smoker | 0
15-pack year history of cigarette use | 0
no anti-coagulants | 0
no amiodarone | 0
no chemotherapeutic agents | 0
no recent nitrofurantoin use | 0
acute respiratory distress | 0
tachypnea | 0
hypoxemia | 0
oxygen saturation of 89% on room air | 0
improved to 95% on 2 liters of oxygen via nasal cannula | 0
afebrile | 0
temperature of 36.7°C | 0
blood pressure of 89/55 mmHg | 0
heart rate of 89 beats per minute | 0
lungs examination normal | 0
awake and alert | 0
normal cardiac examination | 0
normal abdomen examination | 0
no petechiae | 0
no bruising | 0
no gingival bleeding | 0
no oozing from intravenous access sites | 0
anemia | 0
hemoglobin level of 9.9 g/dL | 0
hemoglobin level of 13.3 g/dL at 1 month prior | -720
leukocytosis | 0
white blood cell count of 13.0×10³ cells/μL | 0
left shift | 0
neutrophil count of 10.8×10³ cells/μL | 0
serum lactate of 3.7 mmol/L | 0
arterial blood gas pH of 7.317 | 0
arterial blood gas pCO₂ of 57.7 mmHg | 0
arterial blood gas pO₂ of 40.2 mmHg |BAL performed in the left lower lobe | 0
BAL performed in the right lower lobe | 0
BAL cytology 4 1513 cells/mm³ WBCs | 0
segmented neutrophils 54% | 0
lymphocytes 44% | 0
red blood cells 111 250 million cells/mm³ | 0
antinuclear antibody negative | 0
cytoplasmic antineutrophilic cytoplasmic autoantibodies negative | 0
perinuclear antineutrophilic cytoplasmic autoantibodies negative | 0
rheumatoid factor negative | 0
echocardiogram showed severe pulmonary hypertension | 0
pulmonary artery systolic pressure of 78 mmHg | 0
PaO₂/FiO₂ ratio of 102 mmHg | 0
positive end expiratory pressure of 8 mmHg | 0
intravenous methylprednisolone 250 mg/day | 48
improvement in oxygenation | 72
PaO₂/FiO₂ ratio of 317 mmHg | 72
repeated fiberoptic bronchoscopy | 120
normal mucosa | 120
progressively clear returns on BAL | 120
decreased oxygen requirement | 120
septic shock | 0
died | 336
influenza A (H1N1) | 0
retrocardiac infiltrates | 0
left lower lobe infiltrates | 0
right upper lobe infiltrates | 0
right lower lobe nodule | 0
no pulmonary embolus | 0
airway erythema | 48
BAL bloody returns | 48
BAL negative for cultures | 48
blood cultures negative | 48
urine cultures negative | 48
vancomycin | 0
piperacillin-tazobactam | 0
azithromycin | 0
oseltamivir | 0
intubated | 0
mechanical ventilation | 0
pressors | 0
DAH diagnosis | 48
arterial blood gas pO₂ of 40.2 mmHg | 0
chest x-ray retrocardiac infiltrates | 0
nasopharyngeal swabs positive for influenza A | 0
clinical status deteriorated | 0
chest CT left lower lobe infiltrates | 0
chest CT right upper lobe infiltrates | 0
chest CT right lower lobe nodule | 0
chest CT no pulmonary embolus | 0
fiberoptic bronchoscopy day 2 | 48
BAL left lower lobe bloody returns | 48
BAL right lower lobe bloody returns | 48
BAL cytology 1513 cells/mm³ WBCs | 48
segmented neutrophils 54% | 48
lymphocytes 44% | 48
red blood cells 250 million cells/mm³ | 48
antinuclear antibody negative | 48
cytoplasmic antineutrophilic cytoplasmic autoantibodies negative | 48
perinuclear antineutrophilic cytoplasmic autoantibodies negative | 48
rheumatoid factor negative | 48
echocardiogram severe pulmonary hypertension | 48
pulmonary artery systolic pressure of 78 mmHg | 48
PaO₂/FiO₂ ratio of 102 mmHg | 48
positive end expiratory pressure of 8 mmHg | 48
repeated fiberoptic bronchoscopy day 5 | 120
BAL progressively clear returns | 120
