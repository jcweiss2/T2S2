male | 0
27 weeks of gestation | 0
small for gestational age | 0
signs of placental insufficiency | 0
primary cesarean delivery | 0
amniotic fluid clear | 0
newborn adaptation delayed | 0
respiratory support by CPAP mask | 0
transferred to neonatal intensive care unit | 0
administration of surfactant | 0
caffeine citrate | 0
empirical antibacterial therapy with piperacillin | 0
spironolactone | 0
hydrochlorothiazide | 0
sonography of central nervous system | 0
intracranial hemorrhages grade 1 | 0
intracranial hemorrhages grade 2 | 0
initial perianal smear negative | 0
colonization with multidrug-resistant Acinetobacter pittii | -336
open both-sided inguinal hernia repair | 0
awake caudal anesthesia | 0
blood pressure monitored noninvasively | 0
oxygen saturation monitored noninvasively | 0
heart rate monitored noninvasively | 0
sedated with propofol | 0
positioned in left lateral position | 0
spontaneous breathing maintained | 0
caudal anesthesia performed | 0
skin disinfected with Braunoderm | 0
surgical face masks worn | 0
sterile gloves worn | 0
caudal space identified with ultrasound | 0
22-gauge hollow needle with obturator | 0
1.15 mL/kg of 0.375% solution of ropivacaine instilled | 0
aspiration negative for blood and CSF | 0
epidural spread of local anesthetics confirmed | 0
sufficient analgesia confirmed | 0
surgery started | 0
surgery finished | 51
no further analgesics required | 51
neurology remained adequate | 51
fever up to 39°C | 12
elevated infect parameters in blood | 12
CRP 3 mg/dL | 12
IL-6 1477 pg/dL | 12
empiric broad antibacterial therapy initiated | 12
i.v. cefotaxime | 12
ampicillin | 12
gentamycin | 12
abdomen firm and painful | 12
abdominal sonography | 12
x-ray | 12
explorative laparotomy | 24
brain sonography | 48
signs of inflammatory process | 48
ventriculitis | 48
periventricular leukomalacia | 48
lumbar puncture | 48
increased cell counts | 48
protein increased | 48
lactate increased | 48
differential count | 48
polymorphonuclear leukocytes | 48
mononuclear leukocytes | 48
Gram stain assay | 48
Gram-instable rods | 48
microbiological culture | 48
antibacterial therapy switched | 48
meropenem | 48
vancomycin | 48
lumbar puncture repeated | 72
lactate still high | 72
cell counts decreased | 72
protein decreased | 72
blood cultures | 72
presence of Clostridium perfringens detected | 72
dexamethasone administered | 72
clinical condition deteriorated | 96
sonography exhibited cystic remodeling | 96
secondary brain edema grade 3 | 96
generalized epileptic seizures | 96
anticonvulsive therapy | 96
diazepam | 96
phenobarbital | 96
apnea | 120
severe disturbance of temperature homeostasis | 120
death | 168