25 years old | 0
male | 0
admitted to the hospital | 0
high-grade fever | -144
diffuse abdominal pain | -48
hematemesis | -48
anemia | 0
thrombocytopenia | 0
hyperbilirubinemia | 0
raised transaminases | 0
normal coagulation profile | 0
normal renal function | 0
hemoglobin 10 g/dl | 0
total leukocyte count 5300/cumm | 0
platelet count 15,000/cumm | 0
serum creatinine 1.0 mg/dl |
