seven years old | 0
male | 0
admitted to the hospital | 0
pre-B-ALL | -672
relapse of pre-B-ALL | -672
allogeneic HSCT | -672
hemoglobin 8.5 g/dl | 0
thrombocytes 13,000/μl | 0
WBC 940/μl | 0
neutrophils 50/μl | 0
CRP 6.83 mg/dl | 0
ferritin 182 μg/dl | 0
cachexia | 0
dry skin | 0
pallor | 0
multiple hematomas | 0
hepatosplenomegaly | 0
antibiotic prophylaxis with ceftriaxone | 0
antiviral prophylaxis with acyclovir | 0
antifungal prophylaxis with caspofungin | 0
pain in the left flank | 0
morphine treatment | 0
blinatumomab treatment started | 0
pain aggravated | 5
ultrasound scan | 5
somnolent and sleepy | 6
cerebral side effect of blinatumomab | 6
neurological condition worsened | 6
cerebral CT scan | 6
MRI scan | 6
multiple cerebral hemorrhages | 6
cardio-respiratory decompensation | 6
mechanical ventilation | 6
catecholamine therapy | 6
blinatumomab treatment stopped | 6
hemoglobin 6.7 g/dl | 6
thrombocytes 49,000/μl | 6
WBC 120/μl | 6
neutrophils 20/μl | 6
CRP 23.13 mg/dl | 6
ferritin 1439 μg/dl | 6
echocardiography | 6
multiple thrombi in the left and right ventricle | 6
thromboembolic events | 6
endocarditis | 6
septic embolisms | 6
antibiotic regimen intensified | 6
meropenem | 6
teicoplanin | 6
gentamicin | 6
CT scans of the thorax, abdomen, and pelvis | 12
multiple systemic thromboembolic lesions | 12
ischemia | 12
bleeding | 12
infarction | 12
bone marrow aspiration | 12
bone marrow aplasia | 12
lymphatic blasts | 12
cerebral pressure rising | 12
cerebral herniation | 24
died | 24
autopsy | 24
invasive mycosis of R. pusillus | 24
systemic fungal infection | 24
R. pusillus identified via PCR-based methods | 24