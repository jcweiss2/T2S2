60 years old | 0
female | 0
admitted to the emergency department | 0
migratory right lower quadrant pain | -24
diarrhea | -24
fevers | -24
rigors | -24
previous diverticulitis | -6720
hypertension | -6720
shocked | 0
blood pressure of 86/52 | 0
borderline tachycardiac at 95 bpm | 0
tender in the right lower quadrant | 0
guarding | 0
acute kidney injury (AKI) | 0
eGFR of 37 ml/min | 0
white cell count of 32.9 | 0
referred to the surgical team | 0
clinical diagnosis of acute appendicitis | 0
Alvarado score of nine | 0
urine microscopy showed >500 leucocytes | 0
non-contrast computer tomography (CT) | 0
malrotated right ectopic kidney | 0
perinephric stranding | 0
non-obstructing 6 mm calculus in renal pelvis | 0
treated with ampicillin | 0
reduced dose of gentamicin | 0
admitted to the intensive care unit (ICU) | 0
inotropic support | 0
urine and blood culture grew Escherichia coli | 24
repeat CT with contrast | 24
early renal abscess | 24
transferred to another hospital | 48
insertion of a ureteric stent | 72
improved post stent insertion | 96
discharged | 168
removal of stone and ureteric stent | 1008