20 years old | 0
African American female | 0
weight 75 kg | 0
height 1.75 meters | 0
body mass index 24.5 kg.m-2 | 0
admitted to the emergency room | 0
postictal state | 0
generalized tonic-clonic seizure | -1
new-onset headache | -1
blood pressures 170-140 and 120-90 mmHg | 0
prenatal care unremarkable | 0
medical history unremarkable | 0
hypertensive disorders negative | 0
seizure disorders negative | 0
platelet count 124,000 per cubic millimeter | 0
alkaline phosphatase 207 IU.L-1 | 0
alanine aminotransferase 60 IU.L-1 | 0
aspartate aminotransferase 50 IU.L-1 | 0
lactate dehydrogenase 353 IU.L-1 | 0
uric acid 7.4 mg.dL-1 | 0
Prothrombin Time (PT) 9.9 seconds | 0
fibrinogen 463 mg.dL-1 | 0
3+ urine protein | 0
International Normalized Ratio (INR) 0.9 | 0
Partial Thromboplastin Time (PTT) 29.2 seconds | 0
magnesium sulfate infusion started | 0
frequent neurological checks | 0
blood tests | 0
continuous fetal monitoring | 0
decision to delay head imaging | 0
blood pressures 160-140 and 100-80 mmHg | 1
hourly clinical examinations | 1
neurologically improving patient | 1
no seizure episodes | 1
denies headache | 1
denies visual disturbances | 1
betamethasone for fetal lung maturity | 1
platelet counts decreased to 97,000 per cubic millimeter | 3
HELLP syndrome possible | 3
repeat coagulation profile | 3
low PT | 3
elevated fibrinogen | 3
normal INR | 3
normal PTT | 3
decision to deliver the fetus | 3
urgent cesarean section | 3
Thromboelastography (TEG) performed | 3
TEG results normal | 3
Reaction (R) time 5.8 minutes | 3
Kinetics (K) time 1.8 minutes | 3
alpha angle 66.2 degrees | 3
Lysis index 30 (LY30) 0% | 3
Maximal Amplitude (MA) 66.2 mm | 3
spinal anesthesia performed | 4
hyperbaric 0.75% bupivacaine 14.25 mg | 4
intrathecal morphine 0.02 mg | 4
lumbar 3-4 intervertebral space | 4
20G needle introducer | 4
24G spinal needle | 4
adequate thoracic 4-sensory level block | 4
cesarean section proceeded uneventfully | 4
neonate’s appearance, pulse, grimace, activity, and respiration scores 7/7/7 | 4
neonate sent to neonatal intensive care unit | 4
patient hemodynamically stable | 4
blood pressures 140-130 mmHg to 90-60 mmHg | 4
no excessive bleeding during surgery | 4
blood loss estimated 700 mL | 4
patient recovered in recovery unit | 5
post-spinal anesthesia evaluation unremarkable | 5
frequent neurological checks | 5
platelet counts improving | 5
liver function tests improving | 5
patient discharged home | 120
no complications | 120