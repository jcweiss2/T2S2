baby boy | 0
born by emergency cesarean section | 0
severe preeclampsia in the mother | -72
gestational week 25 6/7 | 0
birthweight 665 g | 0
intubated in the delivery room | 0
transferred to the neonatal intensive care unit | 0
mechanical ventilation | 0
total parenteral nutrition | 24
minimal enteral nutrition with breast milk | 24
delayed meconium passage | 48
abdominal distension | 48
increased gastric residuals | 48
necrotizing enterocolitis | 48
gastric free drainage | 144
broad-spectrum antibiotic therapy | 144
perforated NEC | 144
operation | 144
short bowel syndrome | 144
thyroid screening tests | 336
serum levels of fT4 0.87 ng/dL | 336
TSH 0.061 mIU/L | 336
cortisol 5.75 µg/dL | 336
serum total bilirubin level 12.12 mg/dL | 336
direct reacting bilirubin 11.48 mg/dL | 336
enteral levothyroxine 5 µg/kg/day | 336
no response to treatment | 336
enteral dose of levothyroxine 10 µg/kg/day | 336
poor absorption of the drug | 336
rectal levothyroxine treatment | 432
fT4 levels increased | 441
bilirubin levels decreased | 441
died | 1872
severe bronchopulmonary dysplasia | 1872
surgical NEC | 1872
short bowel syndrome | 1872
sepsis | 1872