76 years old | 0
male | 0
admitted to the hospital | 0
bloody diarrhea | -96
diarrhea about 6 times per day | -96
intermittent abdominal pain | -96
vomiting | -96
dizziness | -96
generalized weakness | -96
watery foul-smelling diarrhea | -2160
generalized weakness | -2160
weight loss | -2160
celiac disease | -43680
gluten-free diet | -43680
non-compliant to gluten-free diet | -2904
afebrile | 0
tachycardic |#FFRejected
severely hypotensive | 0
cachectic | 0
severely dehydrated | 0
hyperactive bowel sounds | 0
diffuse abdominal tenderness | 0
microcytic hypochromic anemia | 0
metabolic acidosis | 0
hypoalbuminemia | 0
hypokalemia | 0
acute renal failure | 0
severe coagulopathy | 0
septic shock due to gastrointestinal infection | 0
hemolytic uremic syndrome | 0
gastrointestinal malignancy | 0
ischemic colitis | 0
blood culture | 0
urine culture | 0
stool culture | 0
CT abdomen and pelvis without contrast | 0
no acute intraabdominal process | 0
admitted to MICU | 0
intravenous fluids | 0
antibiotics | 0
vancomycin | 0
piperacillin-tazobactam | 0
sodium bicarbonate drip | 0
fresh frozen plasma | 0
electrolyte supplementation | 0
emergent hemodialysis | 0
hypotension | 0
anion-gap metabolic acidosis | 0
ARF | 0
improvement within 24 hours | 24
ferritin level 49.9 ng/mL | 24
low serum iron 24 ug/dL | 24
normal total iron-binding capacity 256 ug/dL | 24
low iron saturation 9.38% | 24
iron deficiency anemia | 24
thyrotropin normal | 24
vitamin B12 normal | 24
folate levels normal | 24
total bilirubin normal | 24
lactate dehydrogenase normal | 24
peripheral blood smear normal | 24
fecal leukocytes negative | 24
Clostridium difficile toxin PCR negative | 24
ova and parasites negative | 24
intravenous antibiotics discontinued | 48
persistent diarrhea | 48
colonoscopy | 48
EGD | 48
normal colonic mucosa | 48
normal rectal mucosa | 48
flattened mucosa | 48
mucosal nodularity in duodenum | 48
duodenal biopsies inflammation | 48
intraepithelial lymphocytosis | 48
subtotal villous blunting | 48
diagnosed with celiac crisis | 48
intravenous vitamin K | 48
parenteral nutrition | 48
methylprednisolone | 48
clinical improvement | 48
transferred to general medicine floor | 48
gluten-free diet initiated | 48
oral budesonide | 48
oral steroid discontinued | 240
discharged | 240
gluten-free diet | 240
improvement of malabsorptive symptoms | 240
adherence to gluten-free diet | 8760
asymptomatic at 12-month follow-up | 8760
