baby boy was born by emergency cesarean section | -1
severe preeclampsia in the mother | -1
birthweight of 665 g | -1
intubated in the delivery room | -1
transferred to the neonatal intensive care unit | -1
mechanical ventilation | 0
total parenteral nutrition (TPN) started | 0
minimal enteral nutrition with breast milk started | 0
delayed meconium passage | 1
abdominal distension with increased gastric residuals | 1
laboratory and radiological findings compatible with NEC | 1
minimal enteral feeding discontinued | 1
gastric free drainage initiated | 1
broad-spectrum antibiotic therapy initiated | 1
operated on due to perforated NEC | 6
long segment of intestine resected | 6
stoma formed | 6
TPN continued | 6
minimal enteral feeding started | 13
TPN support could not be discontinued | 13
thyroid screening tests revealed low fT4 and TSH levels | 14
cortisol level was 5.75 µg/dL | 14
serum total bilirubin level was 12.12 mg/dL | 14
direct reacting bilirubin (DB) was 11.48 mg/dL | 14
enteral levothyroxine 5 µg/kg/day started | 21
fT4 level decreased | 28
enteral levothyroxine dose increased to 10 µg/kg/day | 28
fT4 levels did not increase | 28
rectal levothyroxine treatment started | 35
fT4 levels increased | 44
bilirubin levels decreased | 44
baby died on postnatal 77th day | 77
cause of death was severe bronchopulmonary dysplasia, surgical NEC, short bowel syndrome, and sepsis | 77