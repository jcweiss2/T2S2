13 years old | -3600
female | -3600
diagnosed with CESD | -3600
hepatomegaly | -3600
headaches | -3600
feeling of pressure in the right epigastrium | -3600
increasing jaundice | -3600
abnormal bilirubin | -3600
abnormal lipid profile | -3600
abnormal α1-antitrypsin | -3600
hospitalized | 0
laparoscopic cholecystectomy | 0
symptomatic gallstones | 0
chronic and florid fibroplastic cholecystitis | 0
Child-Pugh A/B cirrhosis | 0
Lab-MELD 14 | 0
esophageal varices | 0
solitary fundal varix | 0
hepatosplenomegaly | 0
thrombocytopenia | 0
vitamin D deficiency | 0
calcium deficiency | 0
discharged | 24
readmitted | 120
subjective increase in abdominal circumference | 120
tiredness | 120
scleral jaundice | 120
nausea | 120
pruritus | 120
lack of appetite | 120
Child-Pugh C | 120
Lab-MELD score 18 | 120
hepatic encephalopathy | 120
rifaximin | 120
esophageal varices | 120
fundal varices | 120
elevated transaminases | 120
pancytopenia | 120
abnormal clotting tests | 120
discharged | 144
readmitted | 168
acute onset of epigastric pain | 168
febrile urinary tract infection | 168
E. coli sepsis | 168
parenteral antibiotics | 168
readmitted | 192
compensated cirrhosis | 192
splenomegaly | 192
repeat ligature of esophageal varices | 192
exclusion of relevant fundal varices | 192
vomited blood | 216
emergency endoscopy | 216
Histoacryl treatment | 216
esophageal stent | 216
clipping of an acute Forrest Ia bleed | 216
severe coagulopathy | 216
hemorrhagic shock | 216
diffuse nosebleed | 216
tamponade | 216
clotting factor replacement | 216
severe hypoalbuminemia | 216
dried blood test | 216
reduced acid lipase | 216
reduced beta-galactosidase | 216
apoptosis marker M30 | 216
overall cell death marker M65 | 216
multiorgan failure | 240
died | 240
increased troponin I | 240
increased myoglobin | 240