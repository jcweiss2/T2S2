52 years old | 0
male | 0
Malay | 0
financial consultant | 0
admitted to the hospital | 0
HCV infection | -672
liver cirrhosis | -672
portal hypertension | -672
grade 1 esophageal varices | -672
HIV infection | -672
baseline HCV RNA load was 374000 IU/mL | -672
CD4 count was 76 cell/uL | -672
CD8 was 588 cell/uL | -672
HIV viral load was 1210 copies/mL | -672
HAART regime | -672
Tenvir-EM | -672
efavirenz | -672
alanine aminotransferase was within normal range | -672
follow up | -168
relatively well | -168
severe epigastric pain | -72
breathlessness | -72
nausea | -72
vomiting | -72
no fever | -72
no cough | -72
no diarrhea | -72
no chest pain | -72
conscious | 0
Glasgow coma scale of 14/15 | 0
lethargic | 0
dehydrated | 0
blood pressure was 90/42 mmHg | 0
pulse rate was 133 beats per minute | 0
temperature was 36° Celsius | 0
tachypneic | 0
respiratory rate of 36 per minute | 0
oxygen saturation was 92% | 0
mildly icteric | 0
no flapping tremor | 0
minimal crepitations | 0
reduced vocal resonance | 0
bibasally | 0
soft abdomen | 0
moderate ascites | 0
pitting edema | 0
cardiovascular examination was insignificant | 0
severe metabolic acidosis | 0
arterial blood gas pH of 7.08 | 0
HCO3- of 12 mmol/L | 0
base excess of -16.9 mmol/L | 0
pCO2 of 32 mmHg | 0
lactate level was 12.4 mmol/L | 0
serum ammonia was 116 mmol/L | 0
liver enzyme | 0
ALT was 55mmol/L | 0
bilirubin 37 mmol/L | 0
infective parameters | 0
white blood cell count was 21 × 109 | 0
C-reactive protein was 4.0 mmol/L | 0
amylase was unremarkable | 0
chest radiograph showed minimal interstitial opacities | 0
electrocardiogram revealed normal sinus rhythm | 0
no ischemic changes | 0
intubated | 0
intravenous amoxicillin/clavulanic acid | 0
intravenous metronidazole | 0
continuous veno-venous hemofiltration | 0
antiretroviral therapy was discontinued | 0
peritoneal fluid analysis | 24
abdominal computed tomography scan | 24
repeated CD4 and CD8 cell counts | 24
blood cultures grew gram-negative rod Escherichia coli | 24
septicemic shock | 24
multiorgan dysfunction | 24
lactic acid level remained high | 48
deterioration in liver function | 48
deteriorated | 72
succumbed to his illness | 72