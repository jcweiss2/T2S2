50 years old | 0
male | 0
admitted to the hospital | 0
distortion of the oral commissure | -72
dizziness | -72
headache | -72
malaise | -72
vomiting | -72
shallow nasolabial sulcus on the left side | -72
weakness in closing the left eye | -72
no diplopia | 0
no dysdipsia | 0
no hemiplegia | 0
no limb numbness | 0
lucid | 0
alert | 0
acute upper respiratory tract infection | -72
peripheral facial neuritis | -72
tuberculosis diagnosed | -350400
tuberculosis cured | -350400
no history of immunodeficiency | 0
no history of major trauma | 0
no toxic exposure | 0
no smoking | 0
no alcoholism | 0
no drug abuse | 0
no hereditary disease | 0
family denied unpasteurized buttermilk consumption | 0
blood pressure 135/85 mmHg | 0
temperature 36.5°C | 0
pulse rate 85 bpm | 0
no signs of meningismus | 0
no other neurological irregularities | 0
white blood cell count 10.61×10^9/L | 0
fasting blood glucose 6.3 mmol/L | 0
glycosylated hemoglobin 6.1% | 0
normal serum creatinine | 0
normal cholesterol | 0
normal C-reactive protein | 0
normal creatine kinase | 0
normal procalcitonin | 0
normal blood coagulation parameters | 0
negative HIV antibodies | 0
negative Treponema pallidum antibodies | 0
emergency head CT no abnormalities | 0
chest CT fibrotic streaks in both lungs | 0
dexamethasone 10 mg/day IV | 0
headache | 72
dysdipsia | 72
malaise | 72
fever 39.2°C | 72
neck stiffness | 72
slowness of the pharyngeal reflex | 72
peripheral facial paralysis | 72
facial nerve affected | 72
glossopharyngeal nerve affected | 72
meninges affected | 72
head CT re-examination no abnormalities | 72
somnolence | 96
aphagia | 96
slurred speech | 96
brain MRI multiple abnormal foci in the brainstem | 96
CSF opening pressure 245 mmH2O | 96
CSF white blood cell count 8.35×10^8/L | 96
CSF potassium 2.5 mmol/L | 96
CSF chloride 144 mmol/L | 96
CSF glucose 3.0 mmol/L | 96
CSF microprotein 2.19 g/L | 96
no organisms on Gram stain | 96
no organisms on India ink stain | 96
no organisms on acid-fast stain | 96
transferred to ICU | 96
physical cooling with ice blanket | 96
ice cap | 96
ceftriaxone 2g IV every 12 hours | 96
ganciclovir 0.25g IV every 12 hours | 96
intracranial decompression with mannitol | 96
symptomatic treatment | 96
supportive treatment | 96
negative influenza A and B antigens | 120
negative anti-Toxoplasma antibodies | 120
L. monocytogenes isolated from blood culture | 120
identified by mass spectrometry | 120
no CSF culture abnormality | 120
CSF genome sequencing found L. monocytogenes | 120
respiratory failure | 144
mechanical ventilation | 144
ampicillin 1g IV every 8 hours | 144
amikacin 0.4g IV every 12 hours | 144
meropenem 2g IV every 8 hours | 144
transferred to standard ward | 1440
walk normally | 1440
eat normally | 1440
central respiratory insufficiency | 1440
intermittent mechanical ventilation | 1440
satisfied with treatment | 1440
satisfied with recovery | 1440
