54 years old | 0
male | 0
autism | 0
bipolar disorder | 0
intellectual disability | 0
urinary incontinence | 0
admitted to the hospital | 0
scrotal swelling | -24
fever | -24
temperature of 101.2F | 0
tachycardic | 0
heart rate of 111 beats/min | 0
respiratory rate was 16 breaths/min | 0
saturating at 100% on room air | 0
disheveled | 0
disoriented | 0
not following commands | 0
leukocytosis | 0
neutrophil predominance of 74% | 0
bandemia of 5% | 0
acute renal injury | 0
creatinine of 1.38 mg/dL | 0
lactatemia of 1.8 mmol/L | 0
pyuria | 0
WBC >50 cells/hpf | 0
leukocyte esterase concentration large | 0
RBC 10-25 cells/hpf | 0
started on empiric intravenous vancomycin | 0
started on empiric piperacillin/tazobactam | 0
ultrasound of the testicles | 0
diffuse scrotal wall thickening | 0
right testes measured 3.8 × 1.3 × 2.5 cm | 0
left testes measured 3.6 × 1.7 × 2.4 cm | 0
normal echogenicity | 0
normal echotexture | 0
no masses or areas of architectural distortion | 0
normal blood flow pattern | 0
no hydrocele | 0
no varicocele | 0
distended urinary bladder | 0
ultrasound of the kidneys | 0
moderate hydronephrosis of the right kidney | 0
CT abdomen and pelvis | 0
abscess at the base of the penis | 0
measuring 3.8 × 5.2 × 5.2 cm | 0
causing urinary bladder distention | 0
bilateral hydronephrosis | 0
septic shock | 24
transferred to the medical intensive care unit | 24
norepinephrine initiated | 24
interventional radiology guided aspiration of the perineal abscess | 48
placement of a suprapubic catheter | 48
purulent, sanguinous fluid aspirated | 48
abscessogram | 48
collapsed, amorphous cavity | 48
blood cultures remained negative | 72
cultures from the drainage positive for gram positive cocci | 72
Aerococcus urinae identified | 96
norepinephrine discontinued | 96
returned to the medicine floor | 96
repeat CT of the pelvis | 120
near-complete resolution of the peripenile abscess | 120
persistent cavity and output | 120
catheter remained in place | 120
repeat CT and fluoroscopic guided tube check | 168
removal of the drainage catheter | 168
failed a trial of voiding | 168
retention of 400 mL | 168
suspected urethral strictures | 168
discharged to his group home | 168
follow-up with his urologist | 168
completed treatment with oral amoxicillin/clavulanate | 336
two weeks total of antimicrobials | 336