62 years old | 0
female | 0
admitted to the emergency department | 0
alleged acute myocardial infarction | 0
fever | -144
abdominal pain | -144
abdominal computed tomography scan | -144
liver abscess | -144
hepatic venous thrombosis | -144
empirical antibiotics | -144
pus drained | -144
Klebsiella oxytoca isolated | -144
chest pain | -120
dyspnea | -120
electrocardiography | -120
ST elevation | -120
poor R progression | -120
elevated troponin I | -120
anxious patient | 0
acute respiratory distress | 0
blood pressure 91/62 mmHg | 0
temperature 37.7℃ | 0
respiratory rate 28 breaths per minute | 0
oxygen saturation 88% | 0
decreased breath sounds | 0
diffuse crackles | 0
regular rhythm | 0
no gallops or murmurs | 0
B-type natriuretic peptide level 1,512 pg/mL | 0
white blood cell count 18,600/mm3 | 0
C-reactive protein level 14.44 mg/dL | 0
troponin I normalized | 0
severely impaired LV function | 0
ejection fraction 30% | 0
akinesia in the mid- to distal portion of the LV chamber | 0
Takotsubo cardiomyopathy suspected | 0
coronary angiography | 0
normal epicardial coronary vessels | 0
systolic blood pressure dropped to 70 mmHg | 0
hypotension | 0
fluid resuscitation | 0
vasopressors | 0
dobutamine | 0
diuretic support | 0
hemodynamically stable | 120
improved symptoms | 120
improved chest radiographic findings | 120
persistent apical ballooning | 168
ejection fraction 18% | 168
medical treatment for heart failure | 168
beta-blocker | 168
nitrate | 168
diuretics | 168
angiotensin-converting enzyme inhibitor | 168
persistent LV dysfunction | 504
cardiac magnetic resonance imaging | 504
no signs of tissue hyperenhancement | 504
no scarred myocardial tissue | 504
ejection fraction 36% | 840
apical thrombus | 840
full-dose heparin | 840
oral anticoagulation therapy with warfarin | 840
no embolic event | 840
persistent akinesia of the LV apex | 2160
slightly improved contractility of the mid-ventricular wall segment | 2160
ejection fraction 40% | 2160
apical thrombus completely resolved | 2160