22 years old | 0
female | 0
admitted to the hospital | 0
persistent high fever | -120
systemic joint pain | -120
low saturation of pulse oximetry oxygen | -120
appearance of blastic cell | -120
low platelet count | -120
given acetaminophen | -120
given antibacterial agent | -120
complained of high fever | -120
complained of joint pain | -120
body temperature 37.8°C | 0
SpO2 99% | 0
no systemic superficial lymphadenopathy | 0
no skin eruption | 0
white blood cell count 6680/μL | 0
atypical lymphocytes 44% | 0
hemoglobin 15.2 g/dL | 0
hematocrit 43.5% | 0
platelet count 2.6 × 10^4/μL | 0
PT 16.9 sec | 0
PT-INR 1.59 | 0
APTT 71.8 sec | 0
Fibrinogen 160.4 mg/dL | 0
FDP 137.6 μg/mL | 0
total protein 5.1 g/dL | 0
albumin 2.8 g/dL | 0
AST 537 IU/L | 0
ALT 256 IU/L | 0
LDH 5574 IU/L | 0
total bilirubin 5.4 mg/dL | 0
direct bilirubin 4.7 mg/dL | 0
ALP 1174 IU/L | 0
triglyceride 362 mg/dL | 0
BUN 68.6 mg/dL | 0
Cre 2.67 mg/dL | 0
uric acid 13.3 mg/dL | 0
C-reactive protein 17.78 mg/dL | 0
serum ferritin 23,700 ng/mL | 0
soluble IL-2 receptor 35,300 U/mL | 0
bilateral pneumonia | 0
bilateral pleural effusion | 0
mild cardiomegaly | 0
intra-abdominal lymph node swelling | 0
hepatosplenomegaly | 0
bone marrow examination | 0
atypical lymphoid cells | 0
active histiocytes | 0
hemophagocytosis | 0
flow cytometric analysis | 0
CD8-positive T-cells | 0
methylprednisolone pulse therapy | 0
chemotherapy with CHOPE | 24
EBV titers examined | 0
EBV-DNA viral load examined | 0
Southern blotting analysis | 0
T-cell receptor beta gene rearrangement | 0
diagnosis of systemic EBV+T-cell LPD of childhood | 0
treated with CHASE | 288
treated with high-dose methotrexate and AraC | 576
allo-HSCT | 1032
myeloablative conditioning | 1032
HLA-mismatched sibling donor | 1032
bone marrow transplantation | 1032
graft-versus-host disease prophylaxis | 1032
enrollment | 1296
acute grade II GVHD | 1568
treated with local therapy | 1568
skin GVHD flared to grade III | 2184
treated with PSL | 2184
discharged | 3168
PSL and FK506 tapered and stopped | 5088
in complete remission | 8760
EBV-DNA viral load not detected | 8760
serological change in EBV titers | 8760