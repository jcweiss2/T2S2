50 years old | 0
male | 0
admitted to the hospital | 0
tick bite | -168
generalized myalgias | -168
lethargy | -168
dizziness | -168
mitral valve prolapse | 0
chronic anxiety | 0
hyperlipidemia | 0
peak temperature of 101.5 °F | -24
systolic blood pressure of 80 mm Hg | -24
WBC count of 23.6 10E3/μL | -24
hemoglobin of 21.3 g/dL | -24
hematocrit of 63.4% | -24
erythrocyte sedimentation rate (ESR) of 1 mm/h | -24
venous doppler with compressible veins | -24
computed tomography of the chest with contrast | -24
transthoracic echocardiogram with ejection fraction of 56.4% | -24
electrocardiogram (EKG) with normal sinus rhythm | -24
Lyme titer negative | -24
intravenous (IV) aztreonam | -24
vancomycin | -24
levofloxacin | -24
pulseless electrical activity (PEA) arrest | -2
intubation | -2
return of spontaneous circulation | -2
extensive dusky mottling of all distal extremities | 0
cool to touch | 0
full and firm extremities | 0
lower extremity pulses appreciated with Doppler ultrasound | 0
capillary refill time more than 3 s | 0
right-sided leg lesion concerning for necrosis/vasculopathy | 0
IV vancomycin | 0
tazobactam-piperacillin | 0
doxycycline | 0
hypotensive requiring norepinephrine and vasopressin drips | 0
hemoglobin of 22.4 g/dL | 0
hematocrit of 65.1% | 0
WBC count of 34.5 10E3/μL | 0
platelets of 167 10E3/μL | 0
lactic acid of 7.5 mEq/L | 0
creatinine of 2.49 mg/dL | 0
evidence of liver injury due to shock | 0
aspartate aminotransferase (AST) of 433 IU/L | 0
alanine aminotransferase (ALT) of 477 IU/L | 0
alkaline phosphatase of 26 IU/L | 0
total bilirubin of 0.4 mg/dL | 0
direct bilirubin of 0.0 mg/dL | 0
serum albumin of <1.5 g/dL | 0
multiple albumin infusions | 0
serum calcium of 5.1 mg/dL | 0
intravenous calcium supplementation | 0
fibrinogen of 118 mg/dL | 0
ddimer of 16.17 μg/ml | 0
fibrin split products of >40 μg/ml | 0
disseminated intravascular coagulation | 0
worsening diffuse edema of extremities | 24
ankle-brachial index could not be done | 24
arterial doppler of bilateral lower extremities | 24
four-compartment right lower extremity fasciotomy | 48
right lateral thigh fasciotomy | 48
right forearm fasciotomy | 48
application of vacuum-assisted closures (VAC) | 48
below-knee amputation of the right lower extremity | 168
multiple wound VAC changes | 168
eventual closure of wounds | 720
creatinine of 1.2 mg/dL | -24
creatinine of 2.5 mg/dL | 0
creatinine of 6.61 mg/dL | 24
renal replacement therapy | 24
continuous renal replacement therapy | 24
intermittent hemodialysis | 168
furosemide drip | 168
creatinine of 1.03 mg/dL | 168
infectious workup negative | 0
complements, C3 of 31.4 mg/dL | 0
complements, C4 of 5.5 mg/dL | 0
C3 and C4 levels normalized | 24
serum immunoglobulin G (IgG) of 148 mg/dL | 0
serum immunoglobulin A (IgA) of 32 mg/dL | 0
serum immunoglobulin M (IgM) of 19 mg/dL | 0
serum protein electrophoresis | 24
immunofluorescence | 24
monoclonal gammopathy of unknown significance (MGUS) | 24
anti-nuclear antibody (ANA) titer of 1:640 | 0
workup for connective tissue disorders negative | 0
hemoglobin of 8.5 g/dL | 720
hematocrit of 26.7% | 720
fungemia with Candida albicans | 720
IV micafungin | 720
discharged to an acute rehab | 720
idiopathic systemic capillary leak syndrome (SCLS) | 0