24 years old | 0 | 0 
primigravida | 0 | 0 
37 weeks of gestation | 0 | 0 
admitted to the hospital | 0 | 0 
high grade fever | -72 | 0 
decreased urine output | -72 | 0 
yellowish discolouration | -72 | 0 
altered sensorium | -72 | 0 
disoriented | 0 | 0 
febrile | 0 | 0 
icteric | 0 | 0 
sub-conjunctival haemorrhages | 0 | 0 
fine basal crepitations | 0 | 0 
receiving intravenous artesunate | -72 | 0 
receiving ceftriaxone | -72 | 0 
receiving doxycycline | -72 | 0 
anaemia | -72 | 0 
jaundice | -72 | 0 
deranged liver function | -72 | 0 
coagulopathy | -72 | 0 
thrombocytopenia | -72 | 0 
increased total leucocyte count | -72 | 0 
elevated blood urea nitrogen | -72 | 0 
elevated serum creatinine | -72 | 0 
singleton pregnancy | 0 | 0 
adequate liquor | 0 | 0 
umbilical artery systolic-diastolic ratio of 2:1 | 0 | 0 
mild hepato-splenomegaly | 0 | 0 
non-reassuring fetal heart rate | 0 | 0 
aspiration prophylaxis | 0 | 0 
high-risk consent | 0 | 0 
rapid sequence intubation | 0 | 0 
cricoid pressure | 0 | 0 
thiopental | 0 | 0 
succinylcholine | 0 | 0 
right internal jugular vein cannulation | 0 | 0 
left radial artery cannulation | 0 | 0 
anaesthesia maintained with isoflurane | 0 | 2 
N2O-O2 mixture | 0 | 2 
atracurium | 0 | 2 
delivery of a 2.25 kg baby | 2 | 2 
fentanyl | 2 | 2 
oxytocin infusion | 2 | 24 
hypotension | 2 | 24 
blood loss | 2 | 24 
packed red blood cells transfusion | 2 | 24 
fresh frozen plasma transfusion | 2 | 24 
platelets transfusion | 2 | 24 
noradrenaline infusion | 2 | 24 
mild acidosis | 2 | 2 
normal electrolytes | 2 | 2 
normal serum glucose | 2 | 2 
intensive care unit | 2 | 144 
post-operative analgesia | 2 | 144 
ultrasound guided bilateral transverse abdominis plane block | 2 | 144 
pulmonary haemorrhage | 48 | 48 
coagulopathy | 48 | 48 
blood products transfusion | 48 | 48 
bed side fibre-optic bronchoscopy | 48 | 48 
erythematous mucosa | 48 | 48 
blood clots | 48 | 48 
active oozing | 48 | 48 
diffuse bleeding | 48 | 48 
broncho alveolar lavage | 48 | 48 
Factor VIIa administration | 48 | 48 
bleeding cessation | 48 | 60 
reduction of inspired oxygen fraction | 48 | 60 
bilateral non-homogeneous opacities | 48 | 48 
clear chest radiograph | 60 | 60 
acute kidney injury | 48 | 144 
severe hyperbilirubinemia | 48 | 144 
haemolytic uremic syndrome | 48 | 144 
high serum lactate dehydrogenase | 48 | 48 
schistocytes in peripheral blood | 48 | 48 
nephrology opinion | 48 | 48 
plasmapheresis | 72 | 120 
dialysis | 72 | 120 
altered mental status | 0 | 144 
diffuse cerebral oedema | 72 | 72 
cerebroprotective measures | 72 | 144 
head elevation | 72 | 144 
not rotating neck | 72 | 144 
maintain serum sodium | 72 | 144 
keeping blood partial pressure of carbondioxide | 72 | 144 
stress ulcer prevention | 2 | 144 
deep vein thrombosis prophylaxis | 2 | 144 
glycemic control | 2 | 144 
reducing fever | 96 | 144 
improving consciousness | 96 | 144 
inotropic support tapered | 96 | 144 
improving urine output | 96 | 144 
improving liver function test | 96 | 144 
improving coagulation parameters | 96 | 144 
improving Pao2/Fio2 ratio | 96 | 144 
extubation | 144 | 144 
discharged from the hospital | 168 | 168