78 years old | 0
male | 0
Caucasian | 0
admitted to the hospital | 0
esophageal rupture | -672
sudden onset respiratory distress | -1
chest pain | -1
back pain | -1
hypotensive | -1
tachycardic | -1
evaluated in the emergency department | 0
COPD | -672
atrial fibrillation | -672
Clostridium difficile infection | -672
empyema with mediastinitis | -672
esophageal repair | -672
gastrostomy tube insertion | -672
born in the U.S | -77760
no history of recent travel | 0
blood pressure 100/60 mmHg | 0
heart rate 80/min | 0
respirations 16/min | 0
temperature 99°F | 0
decreased bilateral air entry upon lung auscultation | 0
dullness to percussion of the right lung | 0
admitted to the intensive care unit | 0
diagnosis of acute respiratory distress secondary to acute diastolic decompensation | 0
started on 50% oxygen via mask | 0
ordered to have nothing by mouth | 0
placed on enoxaparin | 0
amiodarone | 0
digoxin | 0
respiratory failure | 1
intubated | 1
mild leukocytosis of 13.8 K/uL | 1
85% neutrophils | 1
hemoglobin 9.1 g/dL | 1
hematocrit 27.6% | 1
platelet 468.0 K/uL | 1
serum chemistries were within normal limits | 1
urine cultures | 1
sputum cultures | 1
three sets of blood cultures | 1
treated empirically for septic shock with intravenous vancomycin | 1
cefepime | 1
clindamycin | 1
computed tomography demonstrated persistent esophageal leakage of contrast | 2
bronchopulmonary fistula | 2
A. israelii positive blood culture | 2
esophageal stent placement | -24
A. israelii infection | -24
discharged | 168