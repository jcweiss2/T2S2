37 years old | 0
male | 0
admitted to the hospital | 0
pain | 0
open postoperative wound | 0
enterocutaneous fistulas | 0
high-degree obesity | -672
bariatric surgery | -672
distal gastrectomy | -672
Roux-en-Y gastric bypass | -672
Braun anastomosis | -672
Shalimov plug | -672
adhesive small bowel obstruction | -72
emergency surgery | -72
relaparotomy | -72
adhesiolysis | -72
nasointestinal intubation | -72
emergency surgery | -55
relaparotomy | -55
adhesiolysis | -55
nasointestinal intubation | -55
gastroenteroanastomosic leakage | -48
peritonitis | -48
surgical wound dehiscence | -48
total parenteral nutrition | -48
fistuloclysis | -48
fever | -24
bowel content in wound | -24
surgical wound dehiscence | -24
fistula output increased | -24
emergency relaparotomy | -17
bypass gastroenterostomy | -17
septic shock | -17
multiple enteroatmospheric fistulas | -17
abdominal wall phlegmon | -17
emergency relaparotomy | -4
collateral enteroenteric anasthomosis | -4
weight loss | -120
abdominal wall wound | 0
wound edges with granulation tissue | 0
wound bottom with small bowel loops | 0
enterocutaneous fistula | 0
Kehr’s T-tube | 0
gastroenteric anastomosis leakage | 0
enteral feeding tube | 0
small bowel lumens with enteric contents | 0
bile | 0
recess in anterior abdominal wall | 0
drainage tube | 0
skin inflammation | 0
maceration | 0
hyperemia | 0
fistulas output | 0
anemia | 0
hypoproteinemia | 0
hypoalbuminemia | 0
hypokalemia | 0
hyperlactataemia | 0
elevated fibrinogen | 0
pulmonary embolism | 0
free fluid in pleural cavity | 0
atelectasis | 0
abdominal wall defect | 0
thrombosis of femoral vein | 0
hepatomegaly | 0
liver steatosis | 0
free liquid in abdomen | 0
fistulography | 0
contrast catheterization | 0
afferent small bowel loops | 0
efferent small bowel loops | 0
gastroenteric leakage | 0
enteroenteroanastomosis | 0
intensive care management | 0
electrolyte imbalance correction | 0
sepsis control | 0
nutritional support | 0
therapy of thromboembolic complications | 0
wound treatment | 0
active aspiration | 0
skin protection | 0
gastric contents aspiration | 0
nasogastric tube | 0
reconstructive surgery | 2160
laparotomy | 2160
distal gastrectomy | 2160
resection of small bowel | 2160
Roux-gastrojejunostomy | 2160
transversostomy | 2160
midline laparotomy | 2160
revision of abdomen | 2160
adhesions separation | 2160
entero-enteric anastomoses | 2160
enterocutaneous fistulas | 2160
gastric fistula | 2160
transverse colon fistula | 2160
stomach mobilization | 2160
gastroenterostomy | 2160
bowel resection | 2160
Roux-en-Y gastric bypass | 2160
colostomy | 2160
postoperative therapy | 2160
total parenteral nutrition | 2160
infusion | 2160
secretion suppression | 2160
thromboembolic prevention | 2160
wound dressing | 2160
uneventful recovery | 2160
wound healing | 2175
sutures removal | 2175
discharge | 2181
laparotomy | 8760
adhesiolysis | 8760
colostomy closure | 8760
transversodescendostomy | 8760
post-surgery period | 8760
discharge | 8769