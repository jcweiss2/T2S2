56 years old | 0
man | 0
multiply recurrent ventral hernia | 0
open recurrent umbilical hernia repair with Atrium C-QUR mesh | -720
seroma formation | -720
open wound | -720
wound vacuum therapy | -720
multiple washouts | -720
mesh excision | -720
repeat ventral hernia repair with Alloderm mesh | -720
medial component separation | -720
recurrence | -672
significant pain | -672
discomfort associated with large ventral hernia defect | -672
preoperative body mass index of 31 | 0
significant lateral retraction of bilateral rectus abdominis muscles | 0
tobacco chewer | -720
hypertension | 0
multiply operated abdomen | 0
combined endoscopic bilateral component separation | 0
open recurrent giant ventral incisional hernia repair with Strattice mesh | 0
extensive open lysis of adhesions | 0
100 cm2 dermatolipectomy | 0
peak airway pressures in high 20s | 0
progressive oliguric | 24
elevated creatinine level of 3.1 | 24
potassium level of 7.1 | 24
transfer to intensive care unit | 24
intraabdominal pressures elevated to high 30s | 24
diagnosis of abdominal compartment syndrome | 24
intubation | 24
paralysis | 24
nasogastric tube decompression | 24
voided 1600 mL of urine | 26
creatinine normalized to 0.8 mg/dL | 36
potassium within normal limits | 36
bladder pressures declined to normal | 36
peak airway pressure improved to mid-20s | 36
intubated and paralyzed through postoperative day 2 | 24
paralytic medication discontinued | 72
continuous positive airway pressure trials | 96
extubated | 120
trickle-tube feeds | 96
ambulatory with abdominal binder | 120
clear liquid diet | 144
regular diet | 168
transferred to floor | 144
discharged | 192
home oxygen requirement | 192
stable urine output | 192
stable electrolytes | 192
stable creatinine level | 192
stable oxygen saturations | 192
