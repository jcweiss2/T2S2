36 years old | 0
female | 0
admitted to the hospital | 0
abdominal pain | 0
diarrhea | 0
mucus blood | 0
pus | 0
recurrent tenesmus attacks | 0
ulcerative colitis | -8760
mesalazine | -8760
prednisone | -8760
anuria | -216
vomiting | -216
diarrhea | -216
fecal microbiota transplantation | -216
dyspnea | 0
cold clammy limbs | 0
increased pulse rate | 0
abdominal cavity pressure of 25 mmHg | 0
grade IV abdominal hypertension | 0
dark colored urine | 0
bloody fluid | 0
total colonic wall thickening | 0
erosions in luminal surface of colon | 0
hyperemia | 0
friability | 0
bleeding | 0
ulcerations | 0
white blood count of 40.77 × 10^9/L | 0
red blood count of 2.41 × 10^12/L | 0
hemoglobin of 60 G/L | 0
sequential organ failure assessment scores of 10 | 0
suspicious thin perforations at rectosigmoid colon | 0
massive ascites | 0
septic shock | 0
colonic perforation | 0
acute renal failure | 0
disseminated intravascular coagulation | 0
severe anemia | 0
urgent total proctocolectomy | 24
ileostomy | 24
massive ascites | 24
total colonic necrosis | 24
edema | 24
dilatation of small intestine | 24
mucosal inflammation | 24
necrosis | 24
hemorrhage | 24
antibacterial therapy | 24
anticoagulant therapy | 24
nutritional support treatment | 24
thrombosis in the trunk of portal vein | 168
thrombosis in the intrahepatic branches | 168
thrombosis in the superior mesenteric vein | 168
thrombosis in the splenic vein | 168
discharged from the hospital | 720