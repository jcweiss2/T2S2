male | 0
infant | 0
birth weight 3562 grams | 0
gestation 39 4/7 weeks | 0
appropriate for gestational age | 0
vaginal delivery | 0
spontaneous rupture of membrane | -11
meconium stained amniotic fluid | 0
perinatal asphyxia | 0
Apgar scores 2, 6, 9 | 0
oral and endotracheal suction | 0
positive pressure ventilation | 0
orally intubated | 0
mechanical ventilation | 0
admission diagnosis severe respiratory distress | 0
meconium aspiration syndrome | 0
perinatal depression | 0
suspected neonatal sepsis | 0
intubation | 0
ventilator support | 0
surfactant meconium lavage | 0
surfactant replacement therapy | 0
antibiotics for neonatal sepsis prophylaxis | 0
ampicillin | 0
gentamicin | 0
umbilical venous catheter placement | 0
umbilical arterial catheter placement | 0
initial UVC position confirmed | 0
UVC tip at T9 | 0
initial blood workup for sepsis negative | 0
respiratory status improving | 0
hypoxia resolving | 0
respiratory acidosis resolving | 0
weaned to minimal settings | 0
preparation for extubation | 0
liver enlargement noted | 144
abdominal X-ray | 144
mildly elevated liver enzymes | 144
febrile | 144
hemodynamically stable | 144
presumptive diagnosis of disseminated neonatal HSV infection | 144
Acyclovir started | 144
HSV polymerase chain reaction pending | 144
blood culture and blood cell parameters repeated | 144
antibiotics coverage continued | 144
extubation failed | 168
upper airway edema | 168
worsening respiratory status | 168
abdominal girth increased | 168
liver enzyme increased | 168
UVC tip at T10 | 168
UVC migrated into liver | 168
abdominal distension | 168
ascites | 168
obstructive uropathy | 168
progressive worsening of respiratory status | 168
abdominal girth increased | 192
liver size increased | 192
X-ray of chest and abdomen | 192
small lung volume | 192
compressed by gasless abdomen | 192
huge liver | 192
marked abdominal distension | 192
ascites | 192
liver enzymes markedly increased | 192
AST 929 U/L | 192
ALT 380 U/L | 192
total/D bilirubin 4.1/1.5 g/dL | 192
lactate dehydrogenase 1861 IU/L | 192
abdominal ultrasound | 192
computed tomography | 192
ascites confirmed | 192
huge liver with echogenic mass | 192
mild left hydroureter/hydronephrosis | 192
obstructive uropathy | 192
intrahepatic biliary duct dilatation | 192
TPN extravasation via UVC suspected | 192
UVC infusion stopped | 192
UVC removed | 192
peripheral intravenous access obtained | 192
dextrose with electrolytes started | 192
pediatric surgeon consulted | 192
exploratory laparotomy | 192
clot removal | 192
ascites drainage | 192
Penrose drain placement | 192
paracentesis confirmed TPN extravasation | 192
peritoneal fluid analysis | 192
protein 1213 mg/dL | 192
triglyceride 591 mg/dL | 192
glucose 539 mg/dL | 192
HSV polymerase chain reaction negative | 240
IV Acyclovir discontinued | 240
repeat blood culture negative | 240
IV ampicillin and gentamicin discontinued | 264
clinical status improved | 240
surgically draining ascites | 240
removal of peritoneal blood clots | 240
exploratory laparotomy | 240
Penrose drain placed | 240
removed 5 days later | 336
elevated liver enzymes dropped | 240
hematuria resolved | 336
enteric nutrition started | 288
full enteric feedings | 336
extubated to room air | 456
nipple feeding started | 600
breast and bottle feeding | 600
Similac Advance | 600
liver laceration resolved | 672
liver mass resolved | 672
obstructive uropathy resolved | 672
ascites resolved | 672
abdominal ultrasound normal | 648
small residual liver mass | 648
discharge home | 672