68 years old | 0
male | 0
admitted to the hospital | 0
superior digestive tract hemorrhage | 0
type 2 diabetes | 0
high blood pressure | 0
cholecystectomy | 0
dental extraction | 0
first episode of bleeding | -1
rushed to the Emergency Room | 0
diagnostic endoscopy | 0
endoscopic hemostasis treatment using clips | 0
bleeding temporarily stopped | 0
lost consciousness | 0
orotracheal intubation | 0
admitted to Intensive Care Unit | 0
altered mental status (Glasgow Coma Scale – 12) | 0
ventilator support | 0
hemodynamic state stable | 0
blood pressure 100/60 mmHg | 0
hemoglobin 6.3 g/dL | 0
hematocrit 22% | 0
blood urea 94 mg/dL | 0
blood creatinine 0.7 mg/dL | 0
lactic acid 4.5 mmol/l | 0
glycemia 350 mg/dL | 0
activated partial thromboplastin time 38 seconds | 0
international normalized ratio 0.8 | 0
transaminases 9.9 U/L | 0
direct bilirubin 0.13 mg/dL | 0
total bilirubin 0.3 mg/dL | 0
serum total protein 5 g/dL | 0
serum albumin 28 g/L | 0
transfused with whole blood | 0
transfused with fresh frozen plasma | 0
continuous saline infusion | 0
colloid infusion | 0
hemostatic agents administered | 0
prokinetic agents administered | 0
proton pump inhibitor (Pantoprazole) continuous infusion | 0
osmotic diuretic therapy | 0
pulmonary congestion | 0
possible cerebral edema | 0
weaned from ventilator | 48
four more episodes of bleeding | 24
endoscopic hemostasis attempted | 24
chest CT angiography performed | 72
prolonged prothrombin time | 72
transfusion with fresh frozen plasma | 72
transfusion with cryoprecipitate | 72
clinical investigations to rule out hemophilia | 72
blood sample sent to external laboratory | 72
low plasma value of FVIII (12%) established | 96
diagnosis of hemophilia | 96
infusion of FVIII (3000 IU every 12 hours for three days) | 96
transfusion of FVIII concentrate increased plasma value to 50% | 96
5th hemostasis endoscopic attempt | 96
clinical status significantly improved | 96
peripheral blood smear analysis | 96
hypochromic microcytic red blood cells | 96
hospital acquired infection | 96
broad-spectrum antibiotic therapy | 96
transferred to Department of Gastroenterology | 168
discharged | 168
