46 years old | 0
male | 0
deceased donor kidney transplantation | -19200
basiliximab | -19200
extended-release tacrolimus (Tac, 2.5 mg/day) | -19200
mycophenolic acid (MPA, 720 mg bid) | -19200
prednisone (5 mg/day) | -19200
creatinine level of 1.13 mg/dL | -19200
productive cough | -96
diarrhea | -96
MPA reduced to 1,080 mg/day | -96
amoxicillin/clavulanic acid therapy | -96
non-resolution of symptoms | -72
MPA reduced to 720 mg/day | -72
Tac reduced to 2 mg/day | -72
azithromycin therapy | -72
SARS-CoV-2 RNA positive | -48
admitted to hospital | -48
body temperature of 38.8°C | -48
persistent cough | -48
diarrhea | -48
chest X-ray left basal opacity | -48
chest X-ray right infra-hilar reticulonodular interstitial pattern | -48
leukocytopenia | -48
thrombocytopenia | -48
hypokalemia | -48
elevated C-reactive protein | -48
elevated lactate dehydrogenase | -48
MPA withdrawn | -48
Tac reduced to 1.5 mg/day | -48
Tac withdrawn | -48
hydroxychloroquine therapy | -48
respiratory status deterioration | -48
renal function deterioration | -48
transferred to ICU | -48
dyspnea | 0
peripheral blood oxygenation 93% under 15 L/min O2 | 0
tachycardia | 0
hypotension | 0
diarrheic stool passage | 0
elevated acute phase reactants | 0
hyperleukocytosis | 0
thrombocytopenia | 0
raised D-dimers | 0
hypokalemia | 0
hyponatremia | 0
sepsis biomarkers negative | 0
no hydronephrosis | 0
normal Doppler graft parameters | 0
hematuria (3+) | 0
proteinuria (2+) | 0
leukocyturia | 0
chest CT suggestive of COVID-19 pneumonia | 0
chest CT bacterial pneumonia features | 0
intubation | 2
high-flow nasal cannula oxygen therapy | 0
respiratory rate 40/min | 0
O2 saturation 89% | 0
PaO2/FiO2 117 | 0
noninvasive mechanical ventilation | 96
oxygen therapy | 96
remission of respiratory insufficiency | 96
stage 3 acute kidney injury | 0
creatinine peak 2.65 mg/dL | 312
creatinine returned to baseline | 456
oliguria | 0
polyuria | 48
normal urine output | 96
severe hyponatremia | 0
inadequate response to hypertonic saline | 0
prednisone replaced with methylprednisolone 16 mg/day | 0
methylprednisolone i.v. pulse therapy (50 mg/day) | 48
methylprednisolone i.v. pulse therapy (100 mg/day) | 72
Tac reintroduced 1.5 mg/day | 528
Tac increased to 2.5 mg/day | 576
discharged home | 672
hydroxychloroquine therapy | 0
lopinavir/ritonavir therapy | 0
meropenem therapy | 0
linezolid therapy | 0
trimethoprim/sulfamethoxazole therapy | 0
caspofungin therapy | 0
negative bacterial cultures | 0
negative blood cultures | 0
negative urine cultures | 0
neutrophilia | 0
broad-spectrum antibacterial therapy | 0
antifungal prophylaxis | 0
resolution of neutrophilia | 0
radiological improvement | 0
dehydration | 0
fluid loss from diarrhea | 0
hesitance in fluid administration | 0
elevated D-dimers | 0
elevated lactate dehydrogenase | 0
elevated ferritin | 0
low platelet counts | 0
prophylactic anticoagulation with enoxaparin | 0
absent dysmorphic erythrocytes | 0
absent red blood cell casts | 0
absent nephrotic range proteinuria | 0
rapid kidney function resolution | 0
moderate tubular dysfunction | 0
polyuria | 0
pre?renal cause of decreased urine output | 0
no renal replacement therapy | 0
tubular dysfunction from drug toxicity | 0
tubular dysfunction from viral infiltration | 0
kidney function recovery | 0
SARS-CoV-2 PCR negative | 528
LPVr introduction | 0
Tac plasma level 2.1 ng/mL | 576
Tac plasma level 4.1 ng/mL | 576
hypertension | 0
impaired glucose tolerance | 0
lymphopenia | 0
cytokine storm | 0
low?dose pulse methylprednisolone | 0
negative procalcitonin | 0
negative lactate | 0
clinical risk factors | 0
laboratory risk factors | 0
favorable ICU evolution | 0
good renal function control | 0
anti?rejection drug management | 0
drug interactions | 0
graft rejection avoided | 0
glucocorticoid use debate | 0
cytokine storm treatment | 0
creatinine rising trend | 0
mechanical ventilation | 0
elevated C?reactive protein | 0
Tac reintroduction | 0
Tac plasma levels monitored | 0
Tac safely increased | 0
empirical antibiotherapy | 0
prophylactic antifungal therapy | 0
superimposed infection suspicion | 0
AKI development | 0
prerenal etiology | 0
renal etiology | 0
dehydration contributor | 0
hypercoagulative status | 0
renal thrombosis absence | 0
tubular dysfunction | 0
drug toxicity | 0
viral infiltration | 0
kidney biopsy consideration | 0
Tac plasma levels consideration | 0
unknown long?term kidney consequences | 0
written informed consent | 0
compliance with ethics policy | 0
World Medical Association Declaration of Helsinki | 0
no conflicts of interest | 0
no funding sources | 0
case report drafting | 0
critical revision | 0
supervision | 0
approval of final manuscript | 0
supplementary data | 0
