74 years old | 0
male | 0
hypertension | 0
insulin-dependent diabetes mellitus type 2 | 0
diabetic retinopathy | 0
weight loss | -672
iron deficiency anemia | -672
tumor in the colon ascendens | -672
liver metastases | -672
right hemicolectomy | -672
low-grade pT3cN0 adenocarcinoma | -672
absence of metastases in 24 excised lymph nodes | -672
lymphovascular growth | -672
no vascular or perineural growth | -672
activated BRAF mutation | -672
loss of expression of MLH1 and PMS2 | -672
mismatch repair-deficient (MMR-D)/microsatellite-instable (MSI) tumor | -672
initiated therapy with pembrolizumab | 0
symptoms of a cold | 168
leukocytosis | 168
increase in C-reactive protein | 168
dry coughing | 528
no fever | 528
increase in AST and ALT | 528
ICI-induced hepatitis grade 2 | 528
initiated prednisolone therapy | 528
second dose of pembrolizumab not given | 528
dyspnea | 696
elevation of troponin T | 696
septal hypokinesia | 696
somnolence | 720
difficulty walking | 720
dysarthria | 720
hoarseness | 720
pain in neck and right leg | 720
difficulty raising right leg | 720
increased dose of prednisolone | 720
computed tomography did not show signs of stroke | 720
increased creatine kinase and myoglobin levels | 720
ICI-induced myositis suspected | 720
antibodies against acetylcholine receptor and titin present | 720
albumin present in cerebrospinal fluid | 720
myasthenia gravis (MG) | 720
unable to sit up | 816
severe dysarthria and dysphagia | 816
absent reflexes | 816
intubated | 816
given methylprednisolone | 816
given intravenous immunoglobulins | 816
given infliximab | 888
felt better | 888
better muscle strength in hands | 888
carbon dioxide retention | 936
noninvasive ventilation | 936
sinus bradycardia | 936
died | 936
autopsy showed significant stenosis of right coronary artery | 936
no fibrosis or signs of recent myocardial infarction | 936
tongue softened | 936
no surgical complication after hemicolectomy | 936
metastasis in right liver lobe | 936
inflammatory infiltration of lymphocytes in intercostal musculature, diaphragm, cervical musculature, and tongue | 936
fibrosis in one area of heart | 936
inflammatory infiltrate in small area of heart | 936
hepatocellular cancer (HCC) in liver | 936
fibrosis stage 2-3 in porta field | 936
cause of death determined as respiratory insufficiency due to polymyositis | 936