33 years old | 0
male | 0
alcohol use disorder | 0
seizures | 0
presented to the emergency room | 0
hypothermic | 0
tachypneic | 0
Bi-level Positive Airway Pressure ventilation | 0
computed tomography of the abdomen and pelvis | 0
cirrhotic liver | 0
extremely large volume ascites | 0
bilateral pleural effusions | 0
admitted to the step down unit | 0
anion gap metabolic acidosis | 0
sepsis | 0
urinary tract infection | 0
cirrhosis | 0
hypoxemic respiratory failure | 0
thoracentesis | 0
paracentesis | 0
melena | -144
gastroenterology consulted | -144
interventional radiology consulted | -144
TIPS procedure | -216
MELD score calculated | -216
MELD score 19 | -216
platelet transfusion | -216
TIPS procedure performed | -216
ultrasound-guided access through the right internal jugular vein | -216
angiography | -216
hepatic venography | -216
TIPS puncture needle rotated and advanced to the portal vein | -216
guidewire inserted | -216
angiographic catheter advanced into the portal vein | -216
balloon catheter dilation | -216
stent deployed | -216
portal pressure measured for gradient reduction | -216
venography repeated | -216
variceal bleeding stopped | -216
somnolent | 0
systolic blood pressure in the 80s | 0
rapid response called | 0
hemoglobin decreased | 0
white blood cell count elevated | 0
red blood cells transfused | 0
CT abdomen performed | 0
shunt patent | 0
decreased enhancement of the liver within posterior segments | 0
dense material within the lesser sac | 0
dense material along the lateral border of the liver | 0
intraperitoneal hemorrhage | 0
upgraded to the intensive care unit | 0
5% albumin administered | 0
cryoprecipitate transfused | 0
fresh frozen plasma transfused | 0
multiple transfusions | 0
coagulopathy | 0
prolonged INR/PT | 0
prolonged aPTT | 0
hematology consulted | 0
intravenous vitamin K administered | 0
cryoprecipitate transfused for fibrinogen | 0
platelet count maintained above 50,000 | 0
cyanocobalamin administered | 0
ferrous sulfate supplementation | 0
folic acid supplementation | 0
prothrombin complex concentrate recommended | 0
another angiogram performed | 384
no active extravasation | 384
post-TIPS venogram performed | 384
patent TIPS shunt | 384
hemoglobin stabilized | 384
hematocrit stabilized | 384
discharged | 384
referred for transfer to a liver transplant center | 384
denied transfer | 384
follow up as an outpatient | 384
hemoperitoneum | 0
inadvertent puncture of the liver capsule | 0
intraperitoneal hemorrhage occurred | 0
bleeding diathesis | 0
