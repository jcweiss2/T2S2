19 years old | 0
    male | 0
    presented to the emergency department (ED) | 0
    motor vehicle accident | 0
    conscious upon admission | 0
    no abnormal symptoms in airways | 0
    normal lung examination | 0
    blood pressure 130/85 mmHg | 0
    pulse rate 130 beats per minute | 0
    no free fluid detected in FAST scan | 0
    BMI 36.3 | 0
    morbid obesity | 0
    no tenderness to palpation on spinal column | 0
    no symptoms of laceration in chest and abdomen | 0
    no abdominal guarding and tenderness | 0
    normal perineal examination | 0
    normal pelvic examination | 0
    normal distal pulses | 0
    deformity in distal third of left forearm | 0
    left lower extremity crash injury | 0
    left leg nearly amputated below knee | 0
    severe muscle and skin damage | 0
    nerves and vessels cut | 0
    history of suicide attempt | 0
    history of psychological disorders | 0
    treated with valproate | 0
    nasogastric tube (NGT) insertion | 0
    foley catheter insertion | 0
    normal chest x-ray | 0
    normal pelvic radiograph | 0
    normal brain CT scan | 0
    planned limb amputation | 0
    below knee amputation performed | 0
    aggressive soft-tissue debridement performed | 0
    serial examinations performed | 0
    hydration performed to prevent kidney damage | 0
    NGT pulled out | -24
    tachypnea | 0
    sinus tachycardia with heart rate 150 beats per minute | 0
    upper abdominal pain | 0
    NGT reinsertion | 0
    pain alleviation | 0
    situation improvement | 0
    tendency to eating | 0
    previous lack of appetite | 0
    transferred to operating room | 24
    suspicion of gastrointestinal bleeding | 24
    suspicion of ischemia | 24
    suspicion of necrosis | 24
    coffee ground secretions in drained fluid | 24
    midline laparotomy performed | 24
    gastric dilation detected | 24
    gastric discoloration detected | 24
    gastric decompression performed | 24
    external compression of stomach | 24
    discoloration disappearance | 24
    suspicious areas necessitated | 24
    lack of improvement | 24
    transferred to operating room for second laparotomy | 48
    total gastrectomy performed | 48
    Roux-en-Y esophagojejunostomy performed | 48
    transferred to ICU | 48
    condition improved during following three days | 48
    surgical debridement performed three times | 72
    infection of amputation stump not controlled | 72
    above-knee amputation due to severe infection | 96
    tachypnea on 5th post-operative day | 120
    re-elevated heart rate | 120
    anuria | 120
    leukocytosis | 120
    elevated creatinine levels | 120
    metabolic acidosis | 120
    blood culture performed | 120
    urine culture performed | 120
    bilateral patchy pulmonary infiltrations | 120
    infectious disease consultation performed | 120
    imipenem administered | 120
    ciprofloxacin administered | 120
    vancomycin administered | 120
    severe sepsis treated | 120
    creatinine level adjusted | 120
    hemodialysis performed | 120
    creatinine elevation | 120
    anuria | 120
    lack of response to crystalloid administration | 120
    high suspicion of anastomosis leakage | 144
    contrast study performed | 144
    gastrografin used | 144
    contrast not detected in intestinal lumen | 144
    failure to rule out anastomosis leakage | 144
    transferred to operating room again | 144
    anastomoses found normal | 144
    no leakage detected | 144
    died three days later | 168
    multi-organ failure | 168