63 years old | 0
female | 0
relapsed AML | -672
diabetes mellitus | -672
induction chemotherapy | 0
cytarabine | 0
clofarabine | 0
allogeneic stem cell transplantation | 0
loose stools | 144
diffuse abdominal pain | 144
Clostridium difficile infection | 144
oral metronidazole | 144
abdominal pain persisted | 168
abdominal pain localized to right lower quadrant | 168
neutropenia | 168
afebrile | 168
abdominal and pelvic CT scan | 168
segmental hypoenhancing area in mid appendix | 168
minimal surrounding fat stranding | 168
concern for appendicitis | 168
broad-spectrum intravenous antibiotics | 168
meropenem | 168
right lower quadrant abdominal pain continued | 192
localized peritoneal signs | 192
repeat CT scan | 192
stable inflammation of appendix | 192
adjacent loop of small bowel with thickened wall | 192
no extraluminal air | 192
no drainable fluid collections | 192
appendectomy | 216
laparoscopic approach | 216
necrotic appendix | 216
necrotic terminal ileum | 216
ileocecectomy | 216
primary stapled anastomosis | 216
intensive care unit | 216
extubated | 240
fever | 288
tachypnea | 384
hypoxia | 384
re-intubated | 384
CT scan of chest | 384
peripheral cavitary lesions | 384
bronchoalveolar lavage | 384
pathological diagnosis of zygomycosis | 432
Hematoxylin and eosin (H&E)-stained sections | 432
ischemic changes | 432
hemorrhage | 432
thrombosed vessels | 432
broad irregular aseptate hyphae | 432
Gomori methenamine silver (GMS)-stained sections | 432
wide ribbon-like aseptate hyphae | 432
antifungal therapy | 432
amphotericin B | 432
fungal overgrowth in surgical wound | 480
culture of bronchoalveolar lavage | 480
Absidia spp. | 480
disseminated angioinvasive zygomycosis | 480
severe hypotension | 528
vasopressors | 528
deteriorating clinical condition | 528
transition to comfort care | 528
expired | 576