54 years old | 0
    man | 0
    sent to the emergency department by his family doctor | 0
    evaluation of a new cardiac murmur | 0
    gastroesophageal reflux disease | 0
    degenerative disc disease | 0
    lived in a home with his wife | 0
    rarely consumed alcohol | 0
    denied smoking | 0
    denied using other substances | 0
    subacute onset of subjective fevers | -336
    subacute onset of chills | -336
    arthritis of his right knee | -336
    arthritis of his left wrist | -336
    erythema | -336
    pain | -336
    swelling | -336
    visited a walk-in clinic | -336
    prescribed naproxen | -336
    temperature was 37.1°C | 0
    pulse was 80 beats per minute | 0
    blood pressure was 109/62 mm Hg | 0
    respiratory rate was 24 breaths per minute | 0
    oxygen saturation was 97% on room air | 0
    grade III to VI early diastolic murmur | 0
    faint crackles to the lung bases | 0
    mild swelling | 0
    pain to his right knee | 0
    pain to his left wrist | 0
    no erythema | 0
    no rash on his skin | 0
    no rash on mucosal surfaces | 0
    point-of-care ultrasonography of the lungs and heart | 0
    diffuse bilateral B-lines | 0
    pulmonary edema | 0
    aortic regurgitation | 0
    neutrophil-dominant leukocytosis of 22 cells × 10⁹/L | 0
    hemoglobin of 126 g/L | 0
    platelets of 164 × 10⁹/L | 0
    creatinine of 137 μmol/L | 0
    increased from a baseline of 90 μmol/L | 0
    C-reactive protein was 209 mg/L | 0
    liver enzymes within normal limits | 0
    chest radiography showed pulmonary edema | 0
    electrocardiography showed complete heart block | 0
    ventricular escape rate | 0
    transthoracic echocardiography showed bicuspid aortic valve | 0
    severe aortic insufficiency | 0
    aortic root abscess | 0
    moderate mitral insufficiency | 0
    transesophageal echocardiography confirmed aortic root abscess | 0
    fistula from the right ventricle to the aortic root | 0
    blood cultures drawn before empiric administration of intravenous ceftriaxone | 0
    blood cultures drawn before empiric administration of vancomycin | 0
    Neisseria gonorrhoeae identified | 0
    diagnosed gonococcal endocarditis | 0
    testing showed susceptibility to azithromycin | 0
    testing showed susceptibility to ceftriaxone | 0
    stopped vancomycin | 0
    prescribed oral azithromycin | 0
    continued ceftriaxone | 0
    did not obtain oral samples for gonococcal testing | 0
    did not obtain genital samples for gonococcal testing | 0
    did not obtain rectal samples for gonococcal testing | 0
    HIV tests negative | 0
    syphilis tests negative | 0
    hepatitis B tests negative | 0
    hepatitis C tests negative | 0
    admitted to the cardiac intensive care unit | 0
    care led by intensivists | 0
    guidance from infectious disease services | 0
    guidance from nephrology services | 0
    guidance from cardiovascular surgery services | 0
    underwent modified Bentall procedure | 0
    surgical aortic valve replacement | 0
    insertion of a bioprosthetic valve | 0
    concomitant aortic root repair | 0
    intraoperative findings showed fistula between the aortic root and the right ventricle | 0
    extensive destruction of the left ventricular outflow tract | 0
    required venous–arterial extracorporeal membrane oxygenation | 0
    inotropic support for 2 days after surgery | 48
    remained in complete heart block | 0
    requiring temporary transvenous pacing | 0
    aortic valve tissue gram stain negative for bacteria | 0
    aortic valve tissue culture negative for bacteria | 0
    16S rRNA gene sequencing confirmed Neisseria gonorrhoeae | 0
    valvular pathology showed active purulent process | 0
    neutrophilic infiltration | 0
    reported contact only with his wife | 0
    did not recall genitourinary symptoms | 0
    did not recall pharyngeal symptoms | 0
    did not recall rectal symptoms | 0
    informed local public health services | 0
    postoperative course complicated by acute tubular necrosis | 0
    required continuous renal replacement therapy | 0
    underwent implantation of a dual-chamber permanent pacemaker | 336
    continued administration of ceftriaxone for 28 days after valve replacement | 672
    transitioned from continuous renal replacement therapy to intermediate hemodialysis | 0
    discharged home | 0
    kidney function improved | 2016
    stopped hemodialysis | 2016
    remained well at nephrology follow-up | 8016
    two months after cardiovascular surgery | 1344
    eleven months after initial presentation | 8016
    