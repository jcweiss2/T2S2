67 years old | 0
African American | 0
female | 0
obesity | -672
chronic active smoker | -672
chronic obstructive pulmonary disease | -672
obstructive sleep apnea | -672
severe pulmonary hypertension | -672
atrial fibrillation | -672
type 2 diabetes | -672
hypertension | -672
dyslipidemia | -672
hypercapnic hypoxic respiratory failure | -672
mechanical ventilation | -672
discharged to rehabilitation facility | -672
admitted to the hospital | 0
generalized weakness | 0
light-headedness | 0
shortness of breath | 0
dry cough | 0
denies subjective fevers | 0
denies chills | 0
denies headache | 0
denies photophobia | 0
denies sputum production | 0
denies nausea | 0
denies vomiting | 0
denies diarrhea | 0
denies dysuria | 0
denies vaginal discharge | 0
denies recent travel | 0
denies exposure to pets | 0
simvastatin | -672
metformin | -672
glipizide | -672
valsartan | -672
labetalol | -672
diltiazem | -672
warfarin | -672
fluticasone/salmeterol | -672
albuterol | -672
hypotension | 0
tachypnea | 0
O2 saturation | 0
pulse | 0
temperature | 0
conjunctival pallor | 0
dry mucous membranes | 0
arrhythmic heart sounds | 0
tricuspid murmur | 0
bilateral crackles | 0
wheezing | 0
nontender abdomen | 0
ascites | 0
edema | 0
decreased peripheral pulses | 0
no skin ulcers | 0
no meningeal signs | 0
no focal deficits | 0
cefepime | 0
vancomycin | 0
leukocyte count | 0
neutrophils | 0
no bandemia | 0
platelets | 0
acute kidney injury | 0
creatinine | 0
hyperglycemia | 0
lactate | 0
International normalized ratio | 0
HIV test | 0
urinalysis | 0
chest computed tomography | 0
abdominal computed tomography | 0
right pleural effusion | 0
right-sided atelectasis | 0
cardiomegaly | 0
moderate ascites | 0
enlarged caliber hepatic veins | 0
transesophageal echocardiogram | 0
ejection fraction | 0
severe tricuspid regurgitation | 0
mild mitral regurgitation | 0
no endocarditis | 0
cytology | 0
peritoneal fluid | 0
pleural fluid | 0
blood cultures | 0
urine cultures | 0
no vasopressors | 24
Gram-negative bacilli | 24
vancomycin discontinued | 24
Sphingobacterium multivorum | 96
resistant to ceftazidime | 96
resistant to trimethoprim/sulfamethoxazole | 96
intermediate susceptibility to meropenem | 96
intermediate susceptibility to piperacillin/tazobactam | 96
ciprofloxacin | 96
negative urine culture | 96
negative peritoneal fluid culture | 96
negative pleural fluid culture | 96
discharged | 240
follow-up | 336
follow-up | 672
clinically stable | 336
clinically stable | 672