22 years old | 0
male | 0
admitted to hospital | 0
fevers | -24
headache | -24
generalized myalgia | -24
non-productive cough | -72
denies photophobia | 0
denies neck stiffness | 0
denies urinary symptoms | 0
denies bowel symptoms | 0
recently well before presentation | -24
Q fever | -672
febrile | 0
tachycardic | 0
no increased work of breathing | 0
chest clear on auscultation | 0
abdomen soft and non-tender | 0
progressive onset of severe epigastric pain | 24
vomiting | 24
septic shock | 24
transferred to intensive care unit | 24
noradrenaline infusion | 24
intravenous piperacillin-tazobactam | 24
ischaemic hepatitis | 24
acute kidney injury | 24
disseminated intravascular coagulopathy | 24
screening for hepatitis B | 24
screening for hepatitis C | 24
screening for HIV | 24
lumbar puncture not performed | 0
abdominal ultrasound | 24
contrast enhanced CT abdomen/pelvis | 24
blood culture revealed N. meningitidis | 72
intravenous benzylpenicillin | 72
clinically improved | 240
discharged from hospital | 240
represented to hospital | 264
mild intermittent left upper quadrant abdominal pain | 264
systemically well | 264
left upper quadrant tender on palpation | 264
abdominal ultrasound | 264
splenic necrosis | 264
CT abdomen/pelvis | 264
extensive splenic necrosis | 264
abscess formation | 264
CT angiogram | 264
percutaneous drainage of splenic abscess | 264
conscious sedation | 264
percutaneous catheter inserted | 264
thick altered blood drained | 264
no growth from collection | 264
recovered well from procedure | 264
discharged | 294
post-splenectomy vaccines | 294
antibiotics prophylaxis | 294