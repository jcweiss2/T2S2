70 years old | 0
female | 0
admitted to the hospital | 0
painless jaundice | -4320
weight loss | -4320
poor appetite | -4320
computed tomography of the chest, abdomen and pelvis | -4320
magnetic resonance cholangiopancreatography | -4320
endoscopic ultrasound | -4320
endoscopic retrograde cholangiopancreatography | -4320
positive emission topography scan | -4320
diagnostic laparoscopy | -4320
open appendectomy for appendicitis | -30240
admitted to the intensive care unit | 0
nasojejunal feeding tube | 0
enteral nutrition commenced | 6
vasopressor support not required | 6
feed rate increased | 24
transferred to the surgical ward | 24
high nasogastric output | 24
osmotic laxative prescribed | 24
oral intake introduced | 48
nausea | 120
vomiting | 120
central abdominal pain | 120
mild tachycardia | 120
central abdominal tenderness | 120
computed tomography scan | 120
large volume of fluid in distal thoracic esophagus and stomach | 120
nasojejunal feeding tube located in efferent small bowel loop | 120
small bowel obstruction | 120
faecalisation | 120
adhesions | 120
laparotomy | 144
small bowel distension | 144
serosal tears | 144
full thickness tear | 144
faecal and feed contamination of the peritoneum | 144
decompression of small bowel | 144
extensive washout | 144
enterotomy repair | 144
nasojejunal feeding tube replaced with standard large bore nasogastric tube | 144
central venous catheter placed | 144
total parenteral nutrition commenced | 144
inotropic support | 144
acute kidney injury | 144
antifungal treatment added to antibiotic regimen | 144
wound dehiscence | 240
intra-abdominal collection | 240
percutaneously inserted drains | 240
oral intake resumed | 360
nourishing fluids continued | 360
wound dehiscence required dressing changes | 360
negative-pressure wound therapy | 360
discharged | 888
follow-up in outpatient clinic | 1008
full diet resumed | 1008