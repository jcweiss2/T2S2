17 years old | 0
    male | 0
    Caucasian | 0
    throat pain | -168
    odynophagia | -168
    acute promyelocytic leukemia (M3) | 0
    daunorubicin | 0
    vesanoid | 0
    extensive necrotic lesion in M. palatoglossus | 0
    necrotic lesion in soft palate | 0
    necrotic lesion in uvula | 0
    necrotic lesion in right tonsil | 0
    unpleasant odor | 0
    biopsy | 0
    culture | 0
    chronic diffuse inflammation | 0
    necrotic areas | 0
    numerous bacteria | 0
    Enterococcus spp | 0
    Staphylococcus aureus | 0
    Candida SP | 0
    noma-like lesion | 0
    ceftazidime | 0
    amicacin | 0
    vancomycin | 0
    fluconazole | 0
    penicillin G | 0
    pneumonia | 24
    sepsis | 24
    intensive care unit | 24
    total recovery | 1080
    extensive loss of soft palate tissue | 1080
