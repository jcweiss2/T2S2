68 years old | 0
female | 0
resident of a long-term nursing facility | 0
dementia | 0
presented to the ED | 0
new onset vomiting | -72
new onset diarrhea | -72
memory loss | 0
denied nausea | 0
denied abdominal pain | 0
denied bleeding |"0
denied fevers | 0
bilateral leg swelling | 0
vague leg discomfort | 0
increased diuretic dose | -72
increased lower extremity edema | -72
denied focal leg pain | 0
denied redness | 0
denied trauma | 0
denied rash | 0
denied shortness of breath | 0
denied chest pain | 0
nonalcoholic fatty liver disease | 0
cirrhosis | 0
chronic kidney disease stage III | 0
insulin-dependent type 2 diabetes | 0
never smoked cigarettes | 0
no history of alcohol abuse | 0
no history of substance abuse | 0
afebrile | 0
heart rate 55 | 0
BP 96/43 mm Hg | 0
respiratory rate 16 breaths/min | 0
oxygen saturation 96% on room air | 0
BMI 36 kg/m² | 0
alert and conversant | 0
oriented to self and place only | 0
dry mucous membranes | 0
anicteric sclera | 0
regular heart rate | 0
no S3 | 0
normal JVP | 0
clear lungs | 0
benign abdomen | 0
negative stool hemoccult | 0
pitting lower extremity edema to knees | 0
no focal tenderness | 0
no erythema | 0
no common findings of cirrhosis | 0
hemoglobin 8.7 g/dL | 0
WBC 12,400/μL | 0
91% segmental neutrophils | 0
no bands | 0
platelets 77,000/μL | 0
sodium 138 mM | 0
potassium 4.4 mM | 0
bicarbonate 15 mM | 0
BUN 72 mg/dL | 0
creatinine 4.16 mg/dL | 0
total bilirubin 1.9 mg/dL | 0
aspartate aminotransferase 63 u/L | 0
alanine aminotransferase 34 u/L | 0
INR 2.1 | 0
ammonia 94 umol/L | 0
venous lactate 1.6 mmol/L | 0
ECG sinus bradycardia | 0
chest radiograph multiple nodular densities | 0
hypotensive (BP 78/34 mm Hg) | 0
received fluid resuscitation | 0
empiric broad-spectrum antibacterials | 0
admitted to the hospital | 0
received IV fluids | 0
normal lactic acid level | 0
negative blood cultures | 0
negative urine cultures | 0
unable to produce sputum | 0
nasal swab negative for MRSA | 0
vancomycin stopped after 48 hours | 48
liver enzymes elevated | 0
ultrasound consistent with cirrhosis | 0
echocardiogram normal systolic and diastolic function | 0
progressive oliguric renal failure | 0
dialysis initiated | 0
developed hypoxic respiratory failure | 72
admitted to ICU | 72
intubated | 72
follow-up chest X-ray worsening | 120
mechanical ventilation | 72
pressors | 72
vancomycin resumed | 72
piperacillin/tazobactam continued | 72
CVVHD initiated | 72
respiratory function stabilized | 168
PEEP 5 cm H2O | 168
FiO2 40% | 168
unable to wean from ventilator | 168
waxing and waning encephalopathy | 168
hypotensive | 168
pressor-dependent | 168
stress-dose steroids | 168
thrombocytopenia | 168
anemia | 168
coagulopathy | 168
transitioned to comfort care | 432
died | 432
hepatic cirrhosis | 432
massive abdominal ascites | 432
esophageal varices | 432
intratubular oxylate crystals | 432
nodular glomerulosclerosis | 432
arterial and arteriolar nephrosclerosis | 432
aortocoronary atherosclerosis | 432
mild cardiomegaly | 432
myocyte hypertrophy | 432
acute and chronic pancreatitis | 432
lung consolidation | 432
septated hyphae with acute angle branching | 432
invasive pulmonary aspergillosis | 432
organizing pulmonary thromboemboli | 432
