62 years old | 0
male | 0
admitted to the hospital | 0
central chest pain | 0
ECG performed | 0
no ST elevation | 0
well perfused | 0
normotensive | 0
sinus rhythm | 0
70 b.p.m. | 0
normal heart sounds | 0
no added sounds or murmurs | 0
clear chest | 0
no arm claudication | 0
good pulses in both upper limbs | 0
normal full blood count | 0
raised fibrinogen | 0
raised troponin T | 0
raised brain natriuretic peptide | 0
coronary angiogram performed | 0
significant left main coronary artery disease | 0
three-vessel disease | 0
patent right brachio-cephalic artery | 0
left ventricular ejection fraction 30% | 0
hypokinesia in inferior and anterior segments | 0
surgical revascularization | 0
LIMA to LAD | 0
saphenous venous graft to intermediate | 0
saphenous venous graft to posterior descending artery | 0
unstable during anaesthetic induction | 0
ST-elevation | 0
urgent initiation of surgery | 0
mixed cardiogenic and distributive shock | 48
intra-aortic balloon pump | 48
high doses of inotropes | 48
weaned after 7 days | 55
septic | 55
inotropic support restarted | 55
empiric antibiotic coverage initiated | 55
meropenem | 55
profound hypokinesia in mid-distal LAD territory | 55
deteriorating echocardiographic picture | 55
transferred to catheterization laboratory | 55
chronic total occlusion of left subclavian artery | 55
peak systolic gradient 60 mmHg | 55
percutaneous coronary intervention | 55
sirolimus-eluting stent in LMS-LAD | 55
paclitaxel-eluting balloon inflation in proximal circumflex artery | 55
comprehensive invasive functional assessment | 55
pressure wire | 55
fractional flow reserve | 55
absolute flow | 55
occlusion of LIMA | 55
coils deployment | 55
Micro Vascular Plug device | 55
complete occlusion of LIMA | 55
improved significantly | 72
weaned from inotropic support | 72
weaned from ventilator | 72
discharged to ward | 720
discharged home | 720
intense rehabilitation | 720
EF 40% | 2160
hypokinesia of inferior wall | 2160
normalization of anterior wall contractility | 2160
prediabetes | -100000
heavy smoker | -100000
acne | -672 
minocycline | -672 
increased WBC count | 0
eosinophilia | 0
systemic involvement | 0
diffuse erythematous or maculopapular eruption | 0
pruritis | 0
DRESS syndrome | 0
fever persisted | 0
rash persisted | 0
discharged | 24