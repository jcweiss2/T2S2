64 years old | 0
male | 0
Japanese | 0
multiple myeloma | -18240
admitted to the hospital | 0
septic shock | 0
febrile episode | 0
lumargia | -6720
L1-2 compression fracture | -6720
blood pressure 82/60 mmHg | 0
heart rate 78/min | 0
body temperature 39.1℃ | 0
respiration rate 20/min | 0
SpO2 95% | 0
no clear focus of infection | 0
no muscular pain | 0
massive myolysis | 0
elevated creatinine kinase | 0
CK 3582 U/L | 0
skeletal muscle | 0
multiple myeloma stage IIIA | -18240
IgG λ type | -18240
melphalan treatment | -18240
prednisolone treatment | -18240
VAD treatment | -18240
vincristine treatment | -18240
doxorubicin treatment | -18240
dexamethasone treatment | -18240
BD treatment | -18240
bortezomib treatment | -18240
thalidomide treatment | -18240
lenalidomide treatment | -4320
IgG increased | -4320
Morganella morganii bacteremia | 0
rehydration | 0
central venous catheterization | 0
catecholamine infusion | 0
dopamine 3 mg/kg/h | 0
meropenem treatment | 0
cervical to pelvis CT | 0
no clear findings | 0
hypotension | 48
oliguria | 48
renal impairment | 48
hemodialysis | 48
endotoxin absorption | 48
respiratory failure | 48
mechanical ventilation | 48
multi-organ failure | 72
death | 72
elevated CK level | 72
CK 19790 U/L | 72
M. morganii sensitive to broad spectrum beta-lactams | 0
M. morganii resistant to cefotiam, minomycin, and ciprofloxacin | 0
outpatient clinic visit | -144
routine follow-up examination | -144
intravenous immunoglobulin | -144