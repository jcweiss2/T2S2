68 years old | 0
male | 0
admitted to the hospital | 0
dyspnea | 0
femoral neck fracture | 0
tonsil cancer | -120 months
radiation therapy | -120 months
recurrent aspiration | -120 months
refused nasogastric tube | -120 months
refused percutaneous endoscopic gastrostomy | -120 months
malnutrition | -120 months
transferred to hospital | 0
aspiration pneumonia | 0
nothing per oral | 0
vegetable soup with solid materials | 5
respiratory failure | 5
shock | 5
intubated | 5
transferred to ICU | 5
bronchoscopy | 5
extracted vegetables | 5
recovered from pneumonia | 10
difficulty liberating from ventilator | 10
recommended tracheostomy | 10
family refused tracheostomy | 10
percutaneous dilatational tracheostomy | 60
discharged to nursing hospital | 72
home ventilator | 72
fever | 2160
dyspnea | 2160
visited ER | 2160
transferred to another hospital | 2160
chest CT | 2160
pneumonia | 2160
no evidence of TEF | 2160
visited ER again | 2268
secretion from tracheostomy tube | 2268
suspiciously similar to enteral feeding materials | 2268
chest CT | 2268
revealed TEF | 2268
continuous leakage of ventilator circuit | 2268
changed T-tube to endotracheal tube | 2268
inflated balloon to maximum | 2268
bronchoscopy | 2268
oval-shaped TEF | 2268
2 cm in diameter | 2268
located on left side of proximal trachea | 2268
NG tube visible through TEF | 2268
consulted radiologist | 2268
consulted gastroenterologist | 2268
consulted pulmonary interventionist | 2268
consulted chest surgeon | 2268
esophageal stent insertion impossible | 2268
endosponge and endoluminal vacuum therapy not agreed | 2268
no stent available for large trachea | 2268
recommended primary closure operation | 2268
improving malnutrition via PEG insertion | 2268
liberation of home ventilator | 2268
family refused PEG procedure | 2268
gave up on primary treatment of TEF | 2304
discharged to nursing hospital | 2304
withdrew from further life-sustaining treatment | 2304
admitted to ICU | 2592
planned esophagogastroscopy and PEG | 2592
routine scope could not enter esophagus | 2592
esophagus inlet stenosis | 2592
complication caused by radiation therapy | 2592
PEG procedure impossible | 2592
thinner scope investigated esophagus | 2592
balloon of endotracheal tube in esophagus | 2592
discussed jejunostomy | 2592
pneumonia | 2592
septic shock | 2592
died | 2616