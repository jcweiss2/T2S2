Here is the table of events and timestamps:

male | 0
infant | 0
born | 0
25-year-old | 0
primigravida | 0
pregnancy was uncomplicated | 0
well before delivery | 0
spontaneous onset of labor | 0
hospital attendance | 0
fetal distress | -2
cardiotocography | -2
ventouse-assisted delivery | -2
male infant | -2
born with a birth weight of 3940 grams | -2
required immediate resuscitation | -2
mask ventilation | -2
intubated at 8 minutes of age | -8
ongoing poor respiratory effort | -8
transferred to the neonatal intensive care unit (NICU) | -8
synchronized intermittent positive pressure ventilation (SIPPV) | -8
minimal pressures | -8
no additional oxygen requirement | -8
empirical antibiotics | -8
gentamicin | -8
benzyl penicillin | -8
presumed early-onset sepsis | -8
respiratory support | -8
weaned | -8
extubated at 13.5 hours of age | -13.5
initial full blood counts | -18
neutropenia | -18
significant left shift | -18
inflammatory markers | -18
C-reactive protein (CRP) | -18
60 mg/L | -18
procalcitonin | -18
68.55 µg/L | -18
lumbar puncture | -23
normal cell count | -23
negative for a range of pathogens | -23
meningococcus | -23
placental surface eSwab | -23
light pure growth of an organism | -23
Gram-negative diplococci | -23
Matrix-Assisted Laser Desorption/Ionization-Time Of Flight (MALDI-TOF) mass spectrometry | -23
Neisseria meningitidis | -23
molecular testing | -23
in-house real-time polymerase chain reaction (PCR) assay | -23
N. meningitidis ctrA and porA genes | -23
real-time PCR assay | -23
common genogroups (serotypes) | -23
B, C, W, and Y | -23
placental isolate | -23
confirmed the detection of a meningococcus genogroup (Serogroup) W clonal complex 11 (CC11) organism | -23
blood cultures | -29
negative | -29
pre–antibiotic treatment | -29
heel-prick blood in EDTA | -34.5
presence of N. meningitidis genogroup W DNA | -34.5
real-time PCR assays | -34.5
no antibiotics were given to the mother | 0
maternal bloods | 0
elevated leucocyte count | 0
21.1×10^9/L | 0
neutrophil count | 0
18.1×10^9/L | 0
mother remained completely well | 0
baby remained well | 0
discharged home from the NICU | 8
day 8 of life | 8
contact tracing | 8
14 staff members | 8
2 parents | 8
3 grandparents | 8
chemoprophylaxis | 8
ciprofloxacin | 8
vaccination | 8
quadrivalent conjugate meningococcal vaccine | 8
counseling | 8
probable ascending infection | 0
materno-fetal transmission | 0
early-onset neonatal sepsis | 0
invasive meningococcal disease (IMD) | 0
neonatal IMD | 0
early-onset sepsis (EOS) | 0
within the first 7 days of life | 0
blood cultures were negative | 0
presence of meningococcal DNA | 0
fetal bloodstream >5 hours postdelivery | 0
funisitis | 0
chorioamnionitis | 0
fetal and maternal inflammatory process | 0
Neisseria species | 0
commensals of the female genital tract | 0
nontypeable strains of N. meningitidis | 0
vaginal specimens | 0
N. meningitidis W CC11 | 0
clusters of urethritis | 0
Australia | 0
IMD rates due to N. meningitidis W | 0
significant case fatality rates | 0
public health concern | 0
heightened vigilance | 0
appropriate treatment and control measures | 0