78 years old | 0
male | 0
admitted to the hospital | 0
red, tender and hot swelling lump on his left breast | -744
pus discharge | -744
treated in the primary care | -744
Flucloxacillin 500 mg TDS | -744
sinus discharging pus | -720
residual abscess | -720
bilateral simple gynecomastia | -2628
Hypertension | 0
Atrial Fibrillation | 0
Diabetes | 0
Hyperlipidaemia | 0
Allopurinol | 0
Amlodipine | 0
Warfarin | 0
large bilateral gynecomastia | 0
abscess/inflammatory mass | 0
ultrasound scan | 0
large abscess in the left retroareolar region | 0
aspiration | 0
mammogram | 24
well-marginated, round 60 mm mass | 24
overlying skin thickening | 24
simple gynecomastia | 24
irregular vascularised hypoechoic mass | 48
enlarged and morphologically abnormal lymph nodes | 48
core biopsy | 72
grade 2 Invasive ductal carcinoma | 72
oestrogen receptor positive | 72
MDT meeting | 72
primary bridging hormone treatment | 72
Tamoxifen 20 mg tablets | 72
staging investigations | 96
no distant metastasis | 96
downstage the tumour | 96
hormone treatment | 120
no real response with Tamoxifen | 216
listed for mastectomy and axillary clearance | 216
mastectomy | 240
axillary clearance | 240
chest wall involvement | 240
final surgical histology | 240
no cellular response to Tamoxifen | 240
tumour size increased | 240
muscle involvement | 240
metastases in lymph nodes | 240
tumour emboli | 240
post-operative MDT | 264
GnRH analogue plus an aromatase inhibitor | 264
adjuvant endocrine treatment | 264
post-mastectomy radiotherapy | 264
chemotherapy | 264
Fluorouracil, Epirubicin, Cyclophosphamide and Docetaxel | 288
six-cycle regime | 288
neutropenic sepsis | 408
omit the final cycle | 408
Radiotherapy and dual anti-hormone treatment | 432
discharged | 480