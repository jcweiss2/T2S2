79 years old | 0
female | 0
hypertension | 0
severe aortic stenosis | 0
chronic heart failure | 0
admitted to the hospital | 0
TAVR | 0
temporary TVP wires placement | 0
transferred to the ICU | 0
extubated | 0
stable condition | 0
TTE performed | 24
decision to remove the pacer wires | 24
removal of pacer wires | 24
became diaphoretic | 24.5
hypotensive | 24.5
resuscitated with intravenous fluid boluses | 24.5
started on a norepinephrine drip | 24.5
BP increased | 25
stat TTE performed | 25
moderate pericardial effusion | 25
excessive respiratory variation of the mitral inflow velocities | 25
mild RV collapse | 25
cardiac tamponade physiology | 25
emergency pericardiocentesis | 25
180 ml of sanguineous fluid drained | 25
pericardial drain left in place | 25
RV rupture | 25
stable | 72
draining minimal amount of fluid | 72
repeat TTE | 72
no new pericardial effusion | 72
decision to remove the pericardial drain | 72
removal of pericardial drain | 72
developed similar acute symptoms | 72.3
hemodynamically unstable | 72.3
emergent TTE | 72.3
reaccumulation of pericardial fluid | 72.3
pericardiocentesis | 72.3
200 ml of frank blood drained | 72.3
coronary angiogram | 72.5
aortic root aortogram | 72.5
transesophageal echocardiography | 72.5
good valve function | 72.5
transferred back to the ICU | 72.5
plan to continue conservative management | 72.5
pericardial catheter clamped | 144
TTE performed | 146
no accumulation of pericardial fluid | 146
drain removed | 146
vital signs monitored | 146
transferred from the ICU to step-down | 170