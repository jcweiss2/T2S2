16 years old | 0
male | 0
admitted to the hospital | 0
sore throat | -24
fatigue | -24
myalgias | -24
fever | -24
left forearm soreness | -24
temperature of 39.1°C | 0
heart rate of 143 beats per min | 0
normal respiratory rate | 0
normal pulse oximetry | 0
normal blood pressure | 0
dry mucus membranes | 0
mild cervical lymphadenopathy | 0
mild erythema of the posterior pharyngeal wall | 0
elevated creatinine level | 0
vancomycin | 0
ceftriaxone | 0
forearm soreness evolved into a swollen, tender, and erythematous area | 48
hypotension | 48
tachycardia | 48
unresponsive to a fluid challenge | 48
transferred to the pediatric Intensive Care Unit | 48
ionotropic support | 48
intra-arterial access | 48
transaminitis | 48
increased bilirubin | 48
C-reactive protein | 48
leukocytosis | 48
coagulation profile consistent with DIC | 48
medical toxicology department consulted | 48
diagnosis of loxoscelism | 48
vesicular areas over a darkening, necrotic-appearing base | 72
skin swab from the lesion submitted for ELISA | 72
ELISA positive for Loxosceles venom | 72
dyspneic | 120
mild pulmonary edema | 120
echocardiogram showed acceptable function with an ejection fraction of 55% | 120
hemoglobin dropped precipitously | 144
LDH increased | 144
bilirubin increased | 144
plasma free hemoglobin increased | 144
intravascular hemolysis | 144
packed red blood cells transfused | 144
methylprednisolone initiated | 144
tachycardia with diffuse T-wave changes on electrocardiogram | 144
myocarditis | 144
B-type natriuretic peptide elevated | 144
troponin-I elevated | 144
creatine kinase-muscle/brain levels elevated | 144
cardiac magnetic resonance imaging demonstrated myocarditis | 144
intravenous immunoglobulins initiated | 144
bumetanide administered | 144
hemoglobin reached a nadir of 5.9 gm/dL | 168
further transfusions | 168
plasmapheresis performed | 192
hematological laboratory results normalized | 192
discharged home | 480
follow-up outpatient echocardiogram was normal | 1440