63 years old | 0 | 0 
female | 0 | 0 
admitted to the hospital | 0 | 0 
general body malaise | -48 | 0 
diarrhea | -48 | 0 
vomiting | -48 | 0 
influenza-like symptoms | -48 | 0 
confusion | 0 | 0 
splenectomy | -77496 | -77496 
idiopathic thrombocytopenic purpura | -77496 | -77496 
menometrorhagia | -77496 | -77496 
vaccinated with PPV23 | -672 | -672 
fever | 0 | 48 
hypotension | 0 | 48 
bradycardia | 0 | 48 
tachypnea | 0 | 48 
decreased oxygen saturation | 0 | 48 
cyanosis | 0 | 48 
severe sepsis | 0 | 48 
volume therapy | 0 | 48 
broad-spectrum antimicrobial therapy | 0 | 48 
hydrocortisone | 0 | 48 
white blood cell count | 0 | 0 
neutrophils | 0 | 0 
hemoglobin | 0 | 0 
thrombocytes | 0 | 0 
C-reactive protein | 0 | 0 
P-lactate | 0 | 0 
aB-P-O2 | 0 | 0 
aB-P-CO2 | 0 | 0 
aB-pH | 0 | 0 
Streptococcus pneumococcal urinary antigen test | 0 | 0 
disseminated intravascular coagulation | 48 | 48 
microthrombi | 48 | 48 
blood cultures showed growth of S. pneumoniae | 48 | 48 
antimicrobial treatment changed to penicillin G | 48 | 48 
suspicion of endocarditis | 72 | 72 
trans-thoracic echocardiography | 72 | 72 
modest hypokinesia of the apical part of the left ventricle | 72 | 72 
ejection fraction of 45% | 72 | 72 
necrosis of the fingertips and toes | 72 | 216 
renal insufficiency | 72 | 216 
hemodialysis | 72 | 216 
antibiotic therapy altered to ceftriaxone | 96 | 96 
leucocytes decreased | 96 | 96 
CRP decreased | 96 | 96 
fever dissolved | 96 | 96 
tracheal secret for culture | 96 | 96 
culture was negative | 96 | 96 
transferred from the ICU to the medical department | 216 | 216 
antibiotics stopped | 216 | 216 
serological analysis of the pneumococcal isolate | 216 | 216 
serotype 12F | 216 | 216 
discharged | 528 | 528 
oral dicloxacillin | 528 | 538 
necrotic fingers and toes amputated | 774 | 774 
readmitted with severe sepsis | 1296 | 1296 
sepsis regimen and ceftriaxone therapy | 1296 | 1296 
transesophageal echocardiography | 1296 | 1296 
endocarditis with several moving elements on the aortic valve | 1296 | 1296 
blood cultures showed growth of S. pneumoniae | 1296 | 1296 
antimicrobial treatment altered to penicillin G | 1296 | 1296 
treated conservatively with penicillin G | 1296 | 1476 
recovered | 1476 | 1476 
antipneumococcal-12F-antibodies measured | -432 | 876 
antibody response to serotype 12F | -432 | 876 
antibody levels to 12F | -432 | 876 
serological tests of the pneumococcal capsule polysaccharides | -432 | 876 
vaccination coverage for the individual patient | 0 | 0 
vaccination is no guarantee against infection | 0 | 0 
need for titer cut-offs for the remaining pneumococcal serotypes | 0 | 0 
laboratory answers to the clinicians should be more detailed | 0 | 0 
patients at increased risk of IPD | 0 | 0 
compromised immune function | 0 | 0