57 years old | 0
    female | 0
    family history of mitral valve prolapse | 0
    presented to the hospital | 0
    altered mental status | 0
    fatigue | -168
    generalized weakness | -168
    episodes of nonbloody vomiting | -168
    diarrhea | -168
    denied chest pressure | 0
    denied chest pain | 0
    denied fever | 0
    denied history of intravenous drug use | 0
    heart rate of 135 beats per minute | 0
    thin | 0
    dry | 0
    lethargic | 0
    Janeway lesions over palms | 0
    Janeway lesions over soles | 0
    Osler nodes | 0
    splinter hemorrhages | 0
    regular heart rhythm | 0
    no murmurs | 0
    white blood cell count of 17,000/mm³ | 0
    hemoglobin of 11.7 g/dL | 0
    platelets 89,000/mm³ | 0
    point of care troponin of 0.28 ng/mL | 0
    sinus tachycardia | 0
    nonspecific ST-wave changes | 0
    blood cultures drawn | 0
    intravenous fluids | 0
    empiric intravenous antibiotics (ceftriaxone and vancomycin) | 0
    follow-up troponin returned at 0.85 | 0
    heparin drip initiated | 0
    chest pain free | 0
    persistent sinus tachycardia | 0
    no ST-segment changes | 0
    subacute infarcts in cerebral hemispheres | 0
    infarctions in kidney | 0
    infarctions in spleen | 0
    heparin drip stopped | 0
    transthoracic echocardiogram (TTE) ordered | 0
    cardiology consulted | 0
    blood cultures positive for methicillin-sensitive Staphylococcus aureus | 0
    TTE showed ejection fraction (EF) of 55% | 0
    no vegetations | 0
    experienced chest pain | 72
    repeat EKG showing diffuse ST-segment elevation | 72
    PR depression consistent with pericarditis | 72
    treated with nonsteroidal anti-inflammatory drugs | 72
    symptomatic relief | 72
    repeat TTE showed EF of 35% to 40% | 72
    severe diffuse hypokinesis of apical wall | 72
    possible vegetation on mitral valve | 72
    transesophageal echocardiogram (TEE) scheduled on day 4 | 96
    TEE confirmed EF of 30% to 35% | 96
    severe hypokinesis | 96
    medium-sized, 1.3 cm (L) × 1.0 cm (W), mobile vegetation on mitral valve | 96
    moderate to severe mitral valve regurgitation | 96
    cardiothoracic surgery consulted | 96
    developed shortness of breath | 96
    decompensated into cardiogenic shock | 96
    placed on vasopressor support | 96
    troponin trended up to 49.50 ng/mL | 96
    emergent cardiac catheterization | 96
    no signs of atherosclerotic coronary artery disease | 96
    100% occlusion of proximal LAD artery | 96
    transferred to cardiac intensive care unit | 96
    underwent mitral valve replacement | 144
    coronary artery bypass grafting (CABG) | 144
    gross specimen showed vegetations involving mitral valve leaflets | 144
    discharged to rehabilitation center | 336
    intravenous antibiotics (cefazolin) | 336
    metoprolol tartrate | 336
    furosemide | 336
    potassium chloride | 336
    repeat TTE on postoperative day 1 showed EF of 10% | 24
    EF improved to 20% on postoperative day 5 | 120
    witnessed seizure | 504
    went into pulseless electrical activity (PEA) | 504
    CPR performed | 504
    return of spontaneous circulation | 504
    potassium of 8 | 504
    elevated troponins | 504
    lactic acid | 504
    CT scan of brain showed evolution of ischemic infarctions | 504
    no acute components | 504
    no hemorrhagic components | 504
    TTE postcardiac arrest showed EF of 20% | 504
    cardiac arrest likely secondary to seizure causing hyperkalemia | 504
    PEA arrest | 504
    no structural changes in TTE | 504
    no dynamic changes in TTE | 504
    terminally extubated | 504
    