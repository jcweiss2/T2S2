22 years old | 0
male | 0
admitted to the hospital | 0
septic shock | 0
aspiration pneumonia | 0
central venous line insertion | 0
somnolent | -5
intubation | -5
arterial catheter insertion | -5
emergency room admission | -5
intensive care unit entry | 5
sepsis | 14
septic shock deterioration | 14
SvO2 measurement | 14.25
SvO2 100% | 14.25
pO2 198 mmHg | 14.25
SvO2 control measurement | 14.5
pO2 200 mmHg | 14.5
arterial blood gas analysis | 14.583
SaO2 98% | 14.583
pO2 90–111 mmHg | 14.583
chest X-ray | 14.833
central venous catheter tip on left heart | 14.833
echocardiography | 15.25
no aortic catheter positioning | 15.25
vena cava superior not seen | 15.25
ECG venous pressure-like curve | 16
C-wave before R-wave | 16
computed tomography | 16.5
catheter in upper left pulmonary vein | 16.5
partial anomalous pulmonary venous return diagnosis | 16.5
conservative treatment | 0
hospital discharge | 336
1-year follow-up | 8784
no significant past medical history | 0
normal venous pO2 (30–40 mmHg) | 0
normal arterial pO2 (75–100 mmHg) | 0
normal venous pCO2 (40–50 mmHg) | 0
normal arterial pCO2 (35–45 mmHg) | 0
catheter tip next to aortic arch | 0
jugular vein insertion confirmation | 0
mean venous pressure 16 mmHg | 0
atypical venous pressure curve | 0
PAPVR prevalence (0.4–0.7%) | 0
asymptomatic PAPVR | 0
conservative management | 0
pulmonary hypertension risk | 0
right heart failure risk | 0
no rerouting needed | 0
no atrial septal defect | 0
no persistent left superior vena cava | 0
no persistent foramen ovale | 0
no other cardiac anomalies | 0
no symptoms post-discharge | 336
no stenosis post-treatment | 336
normal follow-up examination | 336
normal blood gas values post-discharge | 336
