male | 0 | 0 
10 years old | 0 | 0 
admitted to the hospital | 0 | 0 
born | -8760 | -8760 
birth weight 2100 g | -8760 | -8760 
birth length 48 cm | -8760 | -8760 
prominent forehead | -8760 | 0 
relative macrocephaly | -8760 | 0 
limb asymmetry | -8760 | 0 
5th finger clinodactyly | -8760 | 0 
2/3 toe syndactyly | -8760 | 0 
hypomethylation of the 11p15 region | -510 | -510 
genetic examination | -510 | -510 
diagnosis of SRS | -510 | -510 
delayed motor development | -384 | 0 
walked independently | -336 | -336 
hepatic dysfunction | -408 | -408 
increased concentration of alanine aminotransferase | -408 | -408 
increased concentration of aspartate aminotransferase | -408 | -408 
increased creatine kinase level | -408 | -408 
diagnosis of Duchenne muscular dystrophy | -408 | -408 
genetic test | -408 | -408 
mutation of the maternal DMD gene | -408 | -408 
corticosteroids treatment | -192 | 0 
prednisone treatment | -192 | -96 
deflazacort treatment | -96 | 0 
G-CSF treatment | -144 | 0 
sepsis | -144 | -144 
hypoglycaemia | -144 | -144 
neurological symptoms | -144 | -144 
low glucose level | -144 | -144 
urological care | -144 | 0 
hypospadias | -144 | 0 
cardiological diagnostics | -12 | -12 
episodes of sinus tachycardia | -12 | -12 
heart murmur | -12 | -12 
propranolol treatment | -12 | 0 
growth hormone deficiency | -12 | -12 
rhGH treatment | 0 | 18 
growth hormone therapy | 0 | 18 
impaired glucose tolerance | 12 | 12 
insulin resistance | 12 | 12 
discontinuation of rhGH therapy | 18 | 18 
weight gain | 12 | 18 
obesity | 12 | 18 
progressive muscle weakness | 18 | 18 
shortening of 6MT | 18 | 18 
weakened gait | 18 | 18 
discontinuation of rhGH therapy | 18 | 18 
bone density test | 12 | 12 
low bone mineral density | 12 | 12 
scoliosis | 0 | 0 
regular assessment of bone mineral density | 0 | 0 
dual-energy X-ray absorptiometry | 12 | 12 
behavioural therapy | 12 | 18 
physical rehabilitation | 12 | 18 
withdrawal from therapy | 18 | 18