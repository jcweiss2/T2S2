44 years old| 0
    man| 0
    presented to the emergency department| 0
    progressive right lower-extremity pain| -8
    untreated atrial fibrillation| 0
    ulcerative colitis| 0
    ongoing treatment with mesalamine| 0
    agitated| 0
    unable to get comfortable on the stretcher| 0
    severe right lower-extremity pain| 0
    diaphoretic| 0
    tachycardic| 0
    hypertensive| 0
    afebrile| 0
    edematous right lower extremity| 0
    pulseless right lower extremity| 0
    insensate right lower extremity| 0
    no crepitus| 0
    deep vein thrombosis| 0
    workup for pulmonary embolism| 0
    computed tomography (CT) pulmonary angiogram ordered| 0
    right lower-extremity crepitus| 24
    CT extended to include abdomen, pelvis, and lower extremities| 24
    general surgery consulted| 24
    intramuscular air in the proximal right thigh| 24
    intrafascial air in the proximal right thigh| 24
    air tracking up into the pelvis and abdomen| 24
    colonic wall thickening| 24
    contained perforation| 24
    decision to urgently take patient to operating room| 24
    episodes of cardiac arrest| 24
    successfully resuscitated| 24
    stabilized for surgery| 24
    exploratory laparotomy| 24
    fasciotomy| 24
    possible amputation| 24
    disarticulation| 24
    exploratory laparotomy performed| 24
    pneumatosis| 24
    contained colonic perforation| 24
    induration around descending colon| 24
    omental stranding around descending colon| 24
    subtotal colectomy performed| 24
    retroperitoneum hemorrhagic| 24
    retroperitoneum friable| 24
    scrotum evaluated| 24
    perineum evaluated| 24
    right lower extremity blisters| 24
    blisters extending to groin| 24
    incision made over proximal right thigh| 24
    hissing of gas released| 24
    gas bubbles in tissues| 24
    foul-smelling odor| 24
    necrotic muscle| 24
    no active bleeding in extremity| 24
    hip disarticulated| 24
    extremity placed in pathology tray| 24
    cultures of devitalized tissues sent to microbiology| 24
    necrotic muscle debulked| 24
    transferred to intensive care unit| 24
    multiple vasopressors| 24
    multiorgan failure| 24
    succumbed| 24
    Clostridium septicum in tissue cultures| 24
    low-grade mucinous carcinoma| 24
    metastatic deposits in omentum| 24
    gas gangrene| 24
    necrotizing soft-tissue infection| 24
    gastrointestinal malignancy| 24