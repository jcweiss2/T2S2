48 years old | 0
male | 0
admitted to the hospital | 0
asthenia | -216
fever | -216
night sweats | -216
weight loss | -216
cough | -120
dyspnea on exertion | -120
pancytopenia | -168
severe neutropenia | -168
low hemoglobin | -168
low leukocyte count | -168
low lymphocyte count | -168
low monocyte count | -168
low platelet count | -168
bacterial pneumonia | -168
hospitalized in semi-intensive care unit | 0
all blood cultures negative | 0
serum galactomannan test negative | 0
bone marrow aspirate | 0
lymphoid cells with morphology resembling hairy cells | 0
immunophenotyping by flow cytometry | 0
expression of CD19 | 0
expression of CD20bright | 0
expression of CD11c | 0
expression of CD25 | 0
expression of CD103 | 0
expression of CD123 | 0
monoclonality demonstrated by light chain restriction | 0
classic HCL | 0
deterioration of general condition | 168
worsening of dyspnea | 168
persistent fever | 168
septic shock of pulmonary origin | 168
ARDS | 168
acute renal injury | 168
hemodialysis | 168
orotracheal intubation | 168
broad-spectrum antibiotics | 168
meropenem | 168
liposomal amphotericin B | 168
vancomycin | 168
subcutaneous Filgrastim | 168
IFN-α | 168
BRAF V600E mutation negative | 168
progressive weaning of vasoactive drugs | 216
extubation | 216
increasing neutrophil count | 216
packed red blood cell units | 216
recovery of clinical status | 216
resolution of acute renal failure | 216
cladribine | 336
complete recovery of blood counts | 504
satisfactory general condition | 504
good quality of life | 504
bone marrow biopsy | 2160
complete response | 2160