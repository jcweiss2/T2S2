27 years old | 0
male | 0
fell from 4 m height | -75
impaling injury | -75
U shaped metallic bar penetrated the left side of the pelvis | -75
bystanders lifted the patient | -75
EMS arrived | -75
patient was hemodynamically stable | -75
severe pain | -75
evaluation and stabilization of the deformed right lower extremity | -75
transported to the tertiary hospital | -75
airway patent | 0
bilateral good air entry | 0
blood pressure 110/70 | 0
pulse rate 98 | 0
respiratory rate 12 | 0
temperature 36.9 °C | 0
oxygen saturation 99% | 0
Glasgow coma scale 15 | 0
initial evaluation and management | 0
Focused Assessment Sonography for trauma (FAST) | 0
inconclusive FAST | 0
deformity of the right thigh | 0
distal pulses intact | 0
rectal examination negative for blood | 0
rectal examination negative for masses | 0
rectal examination negative for foreign body | 0
prophylactic antibiotic | 0
tetanus toxoid | 0
pelvic and abdominal X-ray assessment | 0
fracture of the right femur | 0
protruded metal bar cut | 0
computerized tomography (CT) scan | 0
metallic bar entered from the left side of the pelvis | 0
no exit site appreciated | 0
bar passed through the left iliac bone | 0
comminuted fracture in the supra-acetabular region | 0
overlying hematoma | 0
surgical emphysema in the soft tissue | 0
bar passed through the junction between the descending and the sigmoid colon | 0
extravasation of the rectally administered contrast | 0
large amount of free air in the upper part of the abdomen | 0
bar traversed the soft tissue behind the rectus muscle | 0
soft tissue contusions | 0
small metal density fragment | 0
exploratory laparotomy | 0
removal of the metallic bar | 0
repair of the sigmoid colon | 0
thorough irrigation | 0
abdomen closed | 0
intramedullary nailing for the fractured femur | 0
fever | 96
tachycardia | 96
tachypnea | 96
desaturation | 96
low white blood cells (WBC) count | 96
intubated | 96
admitted to the Intensive care unit (ICU) | 96
broad spectrum antibiotic | 96
chest and abdominal CT scan | 96
blood culture | 96
methicillin sensitive staphylococcus aureus bacteremia | 96
extubated | 120
transferred back to the ward | 144
abdominal wound infection | 240
pus collection | 240
drained and sent to bacteriology testing | 240
culture result positive for Escherichia Coli | 240
antibiotic changed | 240
wound managed and closed | 288
discharged home | 336