74 years old | 0
    woman | 0
    type 2 diabetes mellitus | 0
    presented to the emergency department | 0
    fever | -120
    jaundice | -120
    right upper quadrant abdominal pain | -120
    traveled to America from Ecuador | -120
    unintentional weight loss | -6720
    abdominal pain (diffuse) | -120
    vomiting (no blood or bile) | -120
    denied chest pain | 0
    denied dyspnea | 0
    denied melena | 0
    denied hematochezia | 0
    denied dysuria | 0
    denied hematuria | 0
    no history of cigarette, alcohol, or substance abuse | 0
    no family history of cancer | 0
    elevated serum alkaline phosphatase (800 IU/L) | 0
    elevated serum creatinine (3.83 mg/dL) | 0
    elevated INR (1.4) | 0
    elevated serum lactate dehydrogenase (471 U/L) | 0
    leukocytosis (17,300 cells/µL) | 0
    predominant monocytosis | 0
    marked thrombocytopenia (10,000/µL) | 0
    macrocytic anemia | 0
    hemoglobin 9 g/dL | 0
    mean corpuscular volume 102.4 fL | 0
    no blasts identified | 0
    diagnosis of sepsis | 0
    admitted to ICU | 0
    treated with broad-spectrum antibiotics | 0
    ultrasound imaging showed cholelithiasis | 0
    thickened gallbladder wall | 0
    positive sonographic Murphy sign | 0
    dilated common bile duct (17 mm) | 0
    ERCP showed purulence and stone in common bile duct | 0
    stone removed | 0
    no sphincterotomy (due to thrombocytopenia) | 0
    plastic stent placed in common bile duct | 0
    progressive leukocytosis | 0
    continued fevers | 0
    laparoscopic cholecystectomy | 0
    Jackson-Pratt drain insertion | 0
    gallbladder appeared gangrenous intraoperatively | 0
    received 1.8 liters crystalloid fluid | 0
    received two units of platelets | 0
    received one unit of irradiated PRBCs | 0
    continued fever | 0
    progressive leukocytosis (80,000 cells/µL) | 0
    clinical appearance of sepsis | 0
    active treatment discontinued | 0
    made comfortable | 0
    histopathology showed myeloblasts, promyelocytes, myelocytes | 0
    granulocytic sarcoma diagnosis | 0
    immunohistochemistry positive for lysozyme, CD68, CD33, HLA-DR | 0
    subsets positive for CD117, myeloperoxidase, CD56 | 0
    negative for CD34 | 0
    acute myelomonocytic leukemia (AML M5) diagnosis | 0