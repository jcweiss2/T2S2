74 years old | 0
male | 0
hypertension | 0
insulin-dependent diabetes mellitus type 2 | 0
diabetic retinopathy | 0
referred to surgery department | 0
8-kg weight loss | 0
iron deficiency anemia | 0
computed tomography | 0
magnetic resonance imaging |9 0
tumor in colon ascendens | 0
3 liver metastases | 0
right hemicolectomy | 0
low-grade pT3cN0 adenocarcinoma | 0
absence of metastases in 24 excised lymph nodes | 0
lymphovascular growth | 0
no vascular growth | 0
no perineural growth | 0
activated BRAF mutation in exon 15 | 0
V600E | 0
loss of expression of MLH1 | 0
loss of expression of PMS2 | 0
mismatch repair-deficient tumor | 0
microsatellite-instable tumor | 0
initiated therapy with pembrolizumab | 0
Keytruda | 0
first infusion of pembrolizumab | 168
symptoms of a cold | 168
leukocytosis | 168
white blood cell count 13.49 ×10^9/L | 168
slight increase in C-reactive protein | 168
dry coughing | 528
no fever | 528
increase in AST | 528
increase in ALT | 528
ICI-induced hepatitis grade 2 | 528
initiated prednisolone therapy | 528
decrease in C-reactive protein | 528
decrease in AST | 528
increased white blood cells | 528
increased neutrophils | 528
not given second dose of pembrolizumab | 528
acutely hospitalized due to dyspnea | 696
elevation of troponin T | 696
echocardiography showed septal hypokinesia | 696
no dynamic change in troponin T | 696
developed somnolence | 696
difficulty walking | 696
dysarthria | 720
hoarseness | 720
pain in neck | 720
pain in right leg | 720
difficulty raising right leg | 720
increased prednisolone dose | 720
computed tomography showed no stroke | 720
increased creatine kinase | 720
increased myoglobin levels | 720
ICI-induced myositis suspected | 720
gradual decrease in creatinine levels | 720
antibodies against acetylcholine receptor | 720
antibodies against titin | 720
albumin in cerebrospinal fluid | 720
unable to sit up | 816
pain in neck | 816
pain in shoulders | 816
severe dysarthria | 816
dysphagia | 816
unable to attain saturation without oxygen | 816
absent reflexes in biceps | 816
absent reflexes in brachioradialis | 816
absent reflexes in triceps | 816
absent reflexes in patellar tendons | 816
absent reflexes in Achilles tendons | 816
transferred to intensive care unit | 816
intubated | 840
suspected immunological involvement of intercostal musculature | 840
methylprednisolone therapy | 840
intravenous immunoglobulins | 840
infliximab therapy | 888
better muscle strength in hands | 912
carbon dioxide retention | 936
noninvasive ventilation | 936
sinus bradycardia | 936
death | 936
significant stenosis of right coronary artery | 936
no fibrosis | 936
no signs of recent myocardial infarction | 936
softened tongue | 936
no surgical complication after hemicolectomy | 936
liver metastases | 936
hepatocellular cancer | 936
fibrosis stage 2-3 in porta field | 936
respiratory insufficiency due to polymyositis | 936
pronounced inflammatory infiltration | 936
fibrosis in heart | 936
inflammatory infiltrate in heart | 936
no colorectal metastases in liver | 936
HCC positive for hepatocytes | 936
negative for glypican | 936
negative for CDX2 | 936
negative for CK20 | 936
negative for CK7 | 936
