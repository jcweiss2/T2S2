62 years old | 0
male | 0
progressive debilitating fatigue | 0
diffuse skin lesions | 0
generalized lymphadenopathy | 0
anemia | 0
peripheral blood blasts (25%) | 0
extensive axillary lymphadenopathy | 0
mediastinal lymphadenopathy | 0
inguinal lymphadenopathy | 0
splenomegaly | 0
flow cytometry monocytic precursors (CD56, CD123) | 0
bone marrow biopsy 37% blasts | 0
blasts expressed CD7 | 0
blasts expressed CD33 | 0
blasts expressed CD38 | 0
blasts expressed CD56 | 0
blasts expressed CD71 | 0
blasts expressed CD117 | 0
blasts expressed CD123 | 0
blasts expressed HLA-DR | 0
blasts negative for CD3 | 0
blasts negative for CD4 | 0
blasts negative for CD10 | 0
blasts negative for CD19 | 0
blasts negative for CD34 | 0
blasts negative for MPO | 0
blasts negative for TdT | 0
skin biopsy consistent with BPDCN | 0
inguinal node aspiration consistent with BPDCN | 0
started on tagraxofusp | 0
tagraxofusp for 8 cycles over 6 months | 0
recurrent scalp lesion | 168
recurrent BPDCN on biopsy | 168
Hyper-CVAD given | 168
hospitalized for neutropenic fever | 168
hospitalized for progressive hypoxia | 168
broad-spectrum antibiotics | 168
steroid course for drug-induced pneumonitis | 168
CSF analysis 76% blasts | 168
intrathecal methotrexate started | 168
CD34+ allogenic stem cell transplant | 216
fludarabine conditioning | 216
melphalan conditioning | 216
engraftment syndrome | 216
Staphylococcal epidermidis bacteremia | 216
Clostridium difficile infection | 216
angioedema | 216
generalized exanthematous pustulosis | 216
bone marrow recurrence (47.5% blasts) | 216
CSF positive for disease | 216
admitted for recurrent disease | 216
vyxeos given | 216
intrathecal methotrexate continued | 216
bone marrow complete response to vyxeos | 672
neutropenic fever | 672
pseudomonas infection | 672
sepsis | 672
succumbed to overwhelming infection | 672
passed away | 672
