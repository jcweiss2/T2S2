40 years old | 0
male | 0
Colombian | 0
living in Switzerland | 0
railway manufacturer | 0
admitted to the emergency department | 0
1-week history of persistent frontal headache | -168
progressive worsening of symptoms | -168
taking over-the-counter painkillers | -168
paracetamol | -168
NSAID | -168
chronic lower back pain | -6720
lumbar disc herniation | -6720
NSAID for chronic lower back pain | -6720
1-month trip to Colombia | -4320
vaccinated for yellow fever | -4320
no known exposure to cattle | -4320
no known exposure to rodents | -4320
no known exposure to tick bites | -4320
no known contact with tuberculosis-infected people | -4320
neurological examination | 0
laboratory work-up | 0
NSAIDs suspended | 0
opioid analgesics administered | 0
quick pain relief | 0
discharged | 24
diagnosis of tension-type headache | 24
paracetamol prescribed | 24
ibuprofen prescribed | 24
tramadol prescribed | 24
reappearance of headache | 24
fever sensation | 24
episode of diarrhoea | 24
physical examination | 24
temperature of 38.1°C | 24
lumbar puncture | 24
cerebrospinal fluid analysis | 24
neutrophilic meningitis | 24
elevated protein levels | 24
hypoglycorrhachia | 24
empirical treatment of dexamethasone | 24
empirical treatment of ceftriaxone | 24
CSF bacterial culture | 24
multiplex PCR assay | 24
contrast-enhanced computed brain tomography | 24
ibuprofen and other prescribed analgesics replaced by morphine | 48
rapid pain relief | 48
discharged | 72
diagnosis of aseptic meningitis | 72
recurrent headaches | 96
fever | 96
neck pain | 96
photophobia | 96
phonophobia | 96
loss of appetite | 96
fatigue | 96
hospitalised | 96
second lumbar puncture | 96
lymphocytic predominance | 96
persistence of high protein levels | 96
slightly lower blood glucose | 96
empirical treatment with intravenous acyclovir | 96
empirical treatment with amoxicillin | 96
empirical treatment with ceftriaxone | 96
thorough diagnostic workup | 96
eubacterial PCR | 96
panfungal PCR | 96
tuberculosis enzyme-linked immunospot assay | 96
CSF direct examination for acid-fast bacilli | 96
CSF PCR for Mycobacterium tuberculosis complex | 96
fourth-generation HIV test | 96
Syphilis screening | 96
tick-borne encephalitis serology | 96
Borrelia burgdorferi serology | 96
PCR in the CSF for B. burgdorferi | 96
lymphocytic choriomeningitis serology | 96
West Nile virus serology | 96
Toscana virus serology | 96
mumps IgG serology | 96
discontinuation of anti-infective therapies | 120
discontinuation of ibuprofen | 120
temporal relationship between ibuprofen use and symptom worsening | 120
symptoms resolution after ibuprofen discontinuation | 144
fever waning | 144
complete resolution of symptoms | 168
follow-up | 720
no headache recurrence | 720
no neurological sequela | 720