36 weeks gestation | 0
female | 0
caucasian | 0
newborn | 0
spontaneous vaginal delivery | 0
thick meconium | 0
tracheal suctioning | 0
positive pressure ventilation | 0
nasal continuous positive airway pressure | 0
marked pallor | 0
normocytic normochromic anemia | 0
10.6 g/dL hemoglobin | 0
31.9% hematocrit | 0
C-reactive protein normal | 0
kidney function tests normal | 0
serum electrolyte levels normal | 0
no signs of hemolysis | 0
no fetomaternal hemorrhage | 0
chorioamnionitis | 0
intravenous antibiotics | 0
blood transfusion | 0
stable | 2
no respiratory distress | 2
spontaneous breathing | 2
oral feeding started | 48
breast feeding | 48
formula feeding | 48
irritable | 72
lethargic | 72
severe dehydration | 72
25% body weight loss | 72
hyperchloremic metabolic acidosis | 72
hypernatremic dehydration | 72
loose watery bloodless stools | 72
mucus in stools | 72
nil per os | 72
volume expansion with normal saline | 72
fluid and sodium bicarbonate replacement therapy | 72
total parenteral nutrition | 72
central venous line | 72
weight loss | 96
hyponatremia | 96
metabolic acidosis | 96
urinary catheterization | 96
profuse diarrhea | 96
high sodium requirements | 96
stool output 120 ml/kg/day | 96
stool reducing substance negative | 96
fecal pH 8 | 96
Na+ concentration in stools 83 mmol/L | 96
fecal ion gap <50 | 96
secretory diarrhea | 96
octreotide | 456
no improvement | 456
cholestasis | 456
catheter-related sepsis | 456
exhaustive etiological investigation | 456
blood cultures normal | 456
stool cultures normal | 456
urine cultures normal | 456
metabolic screen normal | 456
immunoreactive trypsinogen levels normal | 456
renal testing normal | 456
hepatic testing normal | 456
endocrinological testing normal | 456
serum cow milk IgE levels normal | 456
immunodeficiency testing normal | 456
autoimmune enteropathy testing normal | 456
cerebral ultrasound normal | 456
abdominal ultrasound normal | 456
cardiac ultrasound normal | 456
renal ultrasound normal | 456
endoscopy | 288
duodenal biopsy | 288
unspecific inflammatory enteropathy | 288
duodenal biopsy | 744
microvillus atrophy | 744
PAS staining normal | 744
EM examination normal | 744
DNA sequencing | 744
compound heterozygous mutations of MYO5B gene | 744
MVID diagnosis | 744
genetic counseling | 744
discharged home | 744
TPN | 744
liver function deterioration | 1200
septic shock | 2160
catheter-related infection | 2160
death | 2160