35 years old | 0
male | 0
admitted to the hospital | 0
polydipsia | -168
generalized weakness | -168
light headedness | -168
visual disturbances | -168
diabetic ketoacidosis | 0
rhabdomyolysis | 0
blood glucose of 600 mg/dL | 0
arterial blood pH of 7.26 | 0
beta-hydroxybutyrate level of greater than 46.8 mg/dL | 0
anion gap of 27 mmol/L | 0
hemoglobin A1c of 11% | 0
mild leukocytosis at 12,250 cells/mcl | 0
treated with intravenous fluids | 0
treated with insulin infusion | 0
transferred to the medical floor | 48
subcutaneous insulin | 48
fever of 101.6 °F | 48
mental status severely altered | 48
unable to follow multistep commands | 48
unable to tell time on a standard clock | 48
unaware of where he was | 48
unaware of hospitalization | 48
unaware of the current President of the United States | 48
auditory hallucinations | 48
visual hallucinations | 48
generalized muscle soreness | 48
neck stiffness | 48
impaired finger to nose testing | 48
dysconjugate gaze | 48
no nuchal rigidity | 48
Kernig’s sign negative | 48
Brudzinski’s sign negative | 48
chest radiograph showed no acute cardiopulmonary pathology | 48
computed tomography imaging of the head was negative | 48
magnetic resonance imaging of the brain with and without contrast was negative | 48
lumbar puncture | 48
cerebrospinal fluid analysis showed elevated protein | 48
cerebrospinal fluid analysis showed normal glucose | 48
cerebrospinal fluid analysis showed 14 red blood cells | 48
cerebrospinal fluid analysis showed 10 white blood cells | 48
Gram stain of CSF showed no organisms | 48
Herpes virus PCR in CSF was negative | 48
Enterovirus PCR in CSF was negative | 48
blood cultures sent | 48
urine cultures sent | 48
urine analysis revealed large blood | 48
urine analysis revealed 2 red blood cells per high power field | 48
myoglobinuria | 48
initial creatine kinase was measured at 19,154 U/L | 48
empirically started on vancomycin | 48
empirically started on cefepime | 48
mental status gradually improved | 96
hallucinations resolved | 96
creatine kinase rose to 118,400 U/L | 96
weakness improved | 96
muscle tenderness was mild | 96
vastus lateralis muscle biopsy | 96
muscle biopsy showed only rare hypotrophic fibers | 96
muscle biopsy showed no evidence of rhabdomyolysis | 96
muscle biopsy showed no evidence of myopathy | 96
muscle viral myositis and paraneoplastic panel sent | 96
vancomycin stopped | 96
cefepime stopped | 96
continued to improve | 96
creatine kinase started to gradually decrease | 96
muscle tenderness resolved | 96
discharged home | 264
no neurological deficits | 264
CSF results returned positive for IgM antibodies to West Nile Virus | 264
CSF results returned positive for IgG antibodies to West Nile Virus | 264
muscle viral and paraneoplastic panel returned negative | 264