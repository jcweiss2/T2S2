male | 0
preterm | 0
extremely low birth weight | 0
26 weeks of gestation | 0
chronic hypertension | -672
premature prolonged rupture of membranes | -288
latency antibiotics | -288
intravenous ampicillin | -288
oral amoxicillin | -288
azithromycin | -288
chorioamnionitis | -120
ampicillin | -120
trichomonas infection | -672
treated | -672
group B streptococcal culture | -672
negative | -672
spontaneous vaginal delivery | 0
950 g | 0
positive pressure ventilation | 0
intubation | 0
APGAR scores | 0
6 | 0
3 | 0
4 | 0
admitted to the neonatal intensive care unit | 0
arterial cord blood gas pH | 0
6.96 | 0
pCO2 | 0
76 mm Hg | 0
base excess | 0
-15.9 mmol/L | 0
venous cord blood gas pH | 0
7.17 | 0
pCO2 | 0
42 mm Hg | 0
base excess | 0
-12.7 mmol/L | 0
mixed metabolic and respiratory acidosis | 0
high ventilator support | 0
respiratory acidosis | 0
improved | 0
ventilator adjustments | 0
surfactant administration | 0
persistent metabolic acidosis | 0
leukopenia | 0
thrombocytopenia | 0
elevated C-reactive protein | 0
21.1 mg/L | 0
blood culture | 0
ampicillin | 0
gentamicin | 0
hypotensive | 4.5
rapidly deteriorated | 4.5
fluid resuscitation | 4.5
pressors | 4.5
dopamine | 4.5
dobutamine | 4.5
repeat blood culture | 4.5
tracheal aspirate | 4.5
died | 5.5
parents declined autopsy | 5.5
blood cultures | 12
positive | 12
gram-positive cocci | 12
S. gallolyticus | 12
MALDI-TOF | 12
tracheal aspirate culture | 12
negative | 12
placental pathology | 12
acute chorioamnionitis | 12
fetal membranes | 12