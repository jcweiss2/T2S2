70 years old | 0
man | 0
transferred to the hospital | 0
rapid onset consciousness disorder | 0
fever | 0
nausea | 0
vomiting | 0
atopic dermatitis | 0
colon cancer | 0
mitral valve stenosis | 0
ischemic cardiomyopathy | 0
resection of the sigmoid colon | -26208
sigmoid cancer | -26208
adjuvant chemotherapy | -26208
mitral valve replacement | -17520
bioprosthetic valve | -17520
coronary artery bypass | -17520
local recurrence in the pelvis | -4320
totally implantable central venous access device inserted | -4320
chemotherapy started | -4320
impaired consciousness | 0
Glasgow Coma Scale E3V4M5 | 0
blood pressure 90/70 mmHg | 0
heart rate 120 beats/min | 0
respiratory rate 24 breaths/min | 0
oxygen saturation 96% | 0
body temperature 38.4℃ | 0
no rash | 0
no redness at the site of the totally implantable central venous access device | 0
high inflammation state | 0
white blood cells 21,300/mm3 | 0
C-reactive protein 44.8 mg/dL | 0
procalcitonin 85.7 ng/mL | 0
renal dysfunction | 0
creatinine 2.73 mg/dL | 0
blood urea nitrogen 56.7 mg/dL | 0
liver dysfunction | 0
total bilirubin 3.3 mg/dL | 0
Aspartate transaminase 284 IU/L | 0
Alanine transaminase 133 IU/L | 0
disseminated intravascular coagulopathy | 0
DIC | 0
platelet 1.7×104/mm3 | 0
D-dimer 240 μg/mL | 0
prothrombin time 43% | 0
high lactate levels 11.2 mmol/L | 0
plain CT of the chest | 0
plain CT of the abdominal areas | 0
local recurrence at the pelvis showed no change | 0
Gram-positive cluster-forming cocci in urine | 0
antimicrobial therapy initiated | 0
meropenem | 0
linezolid | 0
intravenous fluids | 0
norepinephrine | 0
hypotension | 0
mechanical ventilator support | 0
admitted to the ICU | 0
totally implantable central venous access device removed | 48
no abscess found at the surgical site | 48
prosthetic valve endocarditis suspected | 48
transthoracic echocardiograms | 72
MRSA detected in blood cultures | 72
MRSA detected in urine culture | 72
prolonged state of shock | 72
multiple organ failure | 72
renal failure | 72
hepatic failure | 72
hematologic failure | 72
central nervous system failure | 72
antimicrobial therapy changed to linezolid and clindamycin | 72
intravenous immune globulin administered | 72
transesophageal echocardiogram performed | 72
vegetation at the prosthetic mitral valve | 72
diagnosed with PVE caused by MRSA | 72
antimicrobial therapy changed from linezolid to daptomycin | 96
persistent fever | 144
elevation of CRP | 144
whole-body enhanced CT performed | 144
multiple cerebral emboli | 144
cerebral abscesses | 144
bilateral renal infarctions | 144
renal abscesses | 144
spleen infarction | 144
antimicrobial therapy changed from daptomycin to linezolid | 144
recovered from persistent shock | 192
weaned off mechanical ventilation | 192
TEE performed | 264
enlargement of the vegetation | 264
abscess around the prosthetic valve | 264
surgery for PVE required | 264
transferred to the hospital for mitral valve re-replacement | 264
mitral valve re-replacement with bioprosthetic valve performed | 312
intraoperative valve culture positive for MRSA | 312
antimicrobial therapy continued with linezolid | 312
cerebral infarction | 672
TEE revealed vegetation on the mitral valve | 672
recurrent PVE diagnosed | 672
antimicrobial therapy changed to vancomycin and rifampicin | 672
blood cultures negative after surgery | 672
intravenous antimicrobial therapy continued for four weeks | 672
antimicrobial therapy changed to oral sulfamethoxazole/trimethoprim and rifampicin | 672
bedridden | 672
transferred to a long-term-care sanatorium | 672
antibiotic susceptibility pattern of MRSA | 672
resistance to gentamycin | 672
sensitivity to clindamycin | 672
sensitivity to minocycline | 672
sensitivity to levofloxacin | 672
sensitivity to sulfamethoxazole/trimethoprim | 672
sensitivity to vancomycin | 672
sensitivity to teicoplanin | 672
sensitivity to linezolid | 672
sensitivity to daptomycin | 672
MLST conducted | 672
ST8 | 672
agr l | 672
SCCmec type IVl | 672
CoaIII | 672
PVL-negative | 672
ACME-negative | 672
tst-1 positive | 672
sec positive | 672
sel positive | 672
other virulence genes negative | 672
concluded CA-MRSA/J strain caused PVE | 672
