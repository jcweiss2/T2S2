23 years old | 0
female | 0
abdominal pain | -8
nausea | -8
vomiting | -8
major depression | -7560
bulimia nervosa | -7560
frequent vomiting after binge eating | -7560
suicide attempts | -7560
ate a large quantity of food | -10
abdominal distension | -10
tenderness | -10
no rebound tenderness | -10
abdominal computed tomography (CT) | -10
gastric distension | -10
normal blood test results | -10
joint general surgery consultation | -10
declined hospitalization | -10
warned of possible complications | -10
self-discharge | -10
returned home | -3
re-visited emergency room | 0
persistent abdominal pain | 0
mental confusion | 0
unconscious | 0
severe abdominal distension | 0
abdominal rigidity | 0
pale legs | 0
no auscultation sounds | 0
no dorsalis pedis pulse | 0
shock suspected | 0
low blood pressure | 0
high heart rate | 0
high aspiration rate | 0
high temperature | 0
metabolic acidosis | 0
electrolyte imbalance | 0
severe hypoglycemia | 0
acute renal failure | 0
sodium bicarbonate treatment | 0
abdominal X-ray | 0
gastrointestinal tract filled with food | 0
no bowel gas | 0
abdominal CT | 0
stomach dilation | 0
esophagus dilation | 0
duodenum dilation | 0
endotracheal intubation | 1
Foley catheter insertion | 1
no urine output | 1
emergency hemodialysis | 1
central venous catheter insertion | 1
radial artery conduit placement | 1
nasogastric tube insertion | 1
blockage near esophagus | 1
impossible to insert nasogastric tube | 1
surgical decompression | 6
gastrotomy | 6
food and body fluid drainage | 6
gastric bleeding | 6
low blood pressure | 6
acidosis worsened | 6
electrolyte imbalance exacerbated | 6
hemoglobin decreased | 6
sodium bicarbonate administration | 6
insulin administration | 6
calcium chloride administration | 6
epinephrine administration | 6
continued bleeding | 6
erythrocyte transfusion | 6
fresh frozen plasma transfusion | 6
abdomen closure | 7
cardiopulmonary resuscitation (CPR) | 7
pulseless electrical activity | 7
additional epinephrine administration | 7
vasopressin administration | 7
transfer to intensive care unit (ICU) | 7
no urine output | 7
continued transfusion | 7
disseminated intravascular coagulation (DIC) | 7
low hemoglobin | 7
high prothrombin time | 7
high activated partial thromboplastin time | 7
low platelet count | 7
death | 10