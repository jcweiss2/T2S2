33 years old | 0
    female | 0
    chronic hypersensitivity pneumonitis | 0
    progressively increasing dyspnea | 0
    treated with high-dose glucocorticoids | -72 (assuming treatment started weeks before admission)
    treated with azathioprine | -72
    enlisted for lung transplantation | -72
    lung transplantation | 0
    explantation of donor lungs | -10 (surgery took 10 hours, so explantation started 10 hours before admission)
    secretions in main bronchi | -10
    bacterial culture sent | -10
    clamshell incision | -10
    sequential lung transplant | -10
    induction immunosuppression with basiliximab | -10
    induction immunosuppression with methylprednisolone | -10
    surgery completed in 10 hours | -10
    shifted to ICU | 0
    continued immunosuppression with methylprednisolone | 0
    continued immunosuppression with tacrolimus | 0
    histopathological examination showing chronic hypersensitivity pneumonitis | 0
    required FiO2 0.4 for 24 hours | 0
    chest radiograph showing bilateral diffuse alveolar opacities | 0
    echocardiography showing normal ejection fraction | 0
    primary graft dysfunction considered | 0
    antibody-mediated rejection considered | 0
    hospital-acquired infection considered | 0
    direct crossmatch negative | 0
    started on colistin IV | 0
    started on colistin nebulized | 0
    started on vancomycin | 0
    extubated on second postoperative day | 48
    preemptive NIV administered | 48
    MDR Klebsiella pneumoniae cultured from bronchial swabs | 0
    MDR Klebsiella pneumoniae in blood culture | 0
    MDR Klebsiella pneumoniae in BAL fluid | 0
    persistent fever | 0
    respiratory failure not improving | 0
    tigecycline added | 24 (assuming started after initial 24 hours)
    vancomycin stopped | 24
    tacrolimus withheld | 24
    basiliximab withheld | 24
    immunosuppression maintained with prednisolone | 24
    blood culture grew MDR Klebsiella pneumoniae after 7 days | 168
    developed bilateral empyema | 168
    fosfomycin added | 168
    intrapleural irrigation with colistin | 168
    partial clearing of lung opacities | 168
    weaned off NIV | 168
    oxygen via high-flow nasal cannula | 168
    oxygen via nasal prongs | 168
    acute onset hypotension on 12th postoperative day | 288
    fresh blood in chest drains | 288
    surgical re-exploration | 288
    right ventricle puncture by sternal wire | 288
    repair of cardiac injury | 288
    continued deterioration postoperatively | 288
    increasing alveolar opacities | 288
    subcutaneous air collection | 288
    succumbed to septic shock | 336 (14 days after surgery)
    hospital-acquired pneumonia | 336
    lung biopsy showed no graft rejection | 288
    donor colonization with MDR Klebsiella pneumoniae | -10
    donor had traumatic brain injury | -672 (assuming donor injury occurred weeks before)
    donor mechanically ventilated | -672
    donor FiO2 0.21 | -672
    donor chest radiograph unremarkable | -672
    donor bronchoscopy unremarkable | -672
    donor fit for lung donation | -672
    recipient postoperative complications | 0
    recipient developed empyema | 168
    recipient developed septic shock | 336
    recipient's lung fibrosis | 0
    recipient's chronic hypersensitivity pneumonitis | 0
    recipient's immunosuppression complications | 0
    recipient's infection with MDR Klebsiella pneumoniae | 0
    recipient's surgical complication (cardiac injury) | 288
    recipient's death due to septic shock | 336
    