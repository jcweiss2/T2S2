39 years old | 0
businessman | 0
presented to ICU | 0
acute onset severe abdominal pain | -24
vomiting | -24
binge drinking | -24
chronic alcoholic | -87600
irregularly treated hypertension | -17520
normal baseline creatinine values | 0
no history of chest pain suggesting myocardial infarction | 0
no history of chest trauma | 0
conscious | 0
restless | 0
distended abdomen | 0
tender abdomen | 0
shock | 0
high total leukocyte count | 0
high serum creatinine | 0
high lipase | 0
septic shock | 0
multiple episodes of septic shock | 0
acute kidney injury | 0
raised intra-abdominal pressure | 0
treated with broad-spectrum antibiotics | 0
treated with anti-fungals | 0
treated with vasopressor | 0
treated with inotropes | 0
mechanical ventilation | 0
tracheostomy | 0
enteral nutrition | 0
renal replacement therapy | 0
multiple percutaneous drainages | 0
timely necrosectomy | 0
drain necrotic abdominal content | 0
calcification of mitral leaflet | 2016
calcification of myocardium | 2016
grade I diastolic dysfunction of left ventricle | 2016
ring calcification around left ventricle | 2016
non-specific ST-T changes | 2016
normal cardiac enzyme markers | 2016
normal serum calcium levels | 0
normal serum phosphorus levels | 0
initiation of cardiac calcification | 1008
multi-drug-resistant complicated intra-abdominal infection | 2016
septic shock leading to death | 2016
succumbed to illness | 2016
