51 years old | 0
male | 0
admitted to the hospital | 0
history of asthma | 0
found unconscious at home | -2
swallowed agricultural pesticide | -2
intubated | 2
loss of consciousness | 2
Glasgow Coma Scale (GCS) score of 8 | 2
blood pressure 65/40 mmHg | 2
metabolic acidosis | 2
treated with normal saline | 2
treated with norepinephrine infusion | 2
treated with bicarbonate | 2
treated with hydrocortisone | 2
treated with N-acetylcysteine (NAC) | 2
ingestion of hexaflumuron 10% | -2
Glasgow Coma Scale (GCS) score of 5 | 4
blood pressure 78/36 mmHg | 4
pulse rate 80 beats/min | 4
axillary temperature 37.2°C | 4
respiratory rate 22 cycles/min | 4
intubated and mechanically ventilated | 4
cherry-colored skin | 4
bedside blood glucose level 204 mg/dL | 4
fluid therapy | 4
cardiac monitoring | 4
norepinephrine infusion | 4
hydrocortisone administration | 4
NAC administration | 4
paraclinical evaluations | 4
urine immunoassay positive for tricyclic antidepressant | 4
electrocardiogram | 4
magnesium sulfate administration | 4
echocardiographic finding | 4
transferred to intensive care unit | 7
blood pressure 80/50 mmHg | 7
re-administered normal saline | 7
venous blood gas (VBG) values | 7
bicarbonate administration | 7
norepinephrine infusion discontinued | 30
magnesium sulfate discontinued | 30
serum creatinine level 2.6 mg/dl | 30
low urinary volume | 30
furosemide administration | 30
fluid therapy continued | 30
bicarbonate administration continued | 30
improved on the third day | 52
bicarbonate infusion discontinued | 52
not ready for withdrawal of ventilator support | 52
clinical evidence of pulmonary edema | 52
treated with morphine | 52
treated with furosemide | 52
echocardiogram indicators normal | 52
evidence of pneumonia | 52
antibiotic treatment started | 52
pulmonary x-ray showed broncho-vascular markings | 52
pulmonary x-ray showed para-cardiac opacity | 52
patchy opacity in both lungs | 52
uniform opacity in the inferior and right inferior zones of right lung | 52
blood and urine cultures performed | 52
urine culture positive for Ecoli | 52
no germ grew in blood culture | 52
developed fever | 52
underwent treatment | 52
did not respond appropriately | 52
bradycardia | 72
hypotension | 72
cardiac arrest | 72
cardiopulmonary resuscitation | 72
death | 72