48 years old | 0
male | 0
admitted to the hospital | 0
headache | 0
subarachnoid hemorrhage | 0
untreated hypertension | -672
no smoking history | 0
no family history of thrombotic disease | 0
surgical titanium clipping for left intracranial aneurysms | 0
transferred from the intensive care unit to the general ward | 72
receiving rehabilitation | 72
high grade fever | 120
chills | 120
nausea | 120
ceftriaxone | 120
vancomycin | 120
hypotensive | 144
tachycardia | 144
temperature 37.4 | 144
blood pressure 62/52 | 144
heart rate 110/min | 144
respiratory rate 26 breaths/min | 144
oxygen saturation 68% | 144
cold limbs | 144
cyanosis | 144
tachypnea | 144
leukocytosis | 144
elevated liver enzymes | 144
elevated serum creatinine | 144
C-reactive protein 29.33 | 144
protein C level normal | 144
pyuria | 144
bacteriuria | 144
acute focal bacterial nephritis | 144
septic shock | 144
intravenous fluid resuscitation | 144
antimicrobials | 144
vasopressors | 144
methylprednisolone | 144
anticoagulant therapy | 144
continuous hemodiafiltration | 144
Enterobacter aerogenes | 168
high-grade fever | 168
DIC | 168
platelet transfusion | 168
extensive purpura | 192
purpura fulminans | 192
skin biopsy | 192
necrosis | 192
bullae | 192
thrombosis | 192
limb amputation | 216
hypotension improved | 216
low platelet levels improved | 216
persistent fever | 216
chills | 216
all devices changed | 216
blood cultures | 216
persistent bacteremia | 216
transfusion dependent | 216
anemia | 216
low platelet levels | 216
platelets transfused | 216
red blood cells transfused | 216
condition worsened | 432
died | 456
autopsy | 456
multiple abscesses | 456
thrombosis | 456
lung | 456
intestinal tract | 456
kidney | 456