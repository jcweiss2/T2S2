51 years old | 0
    male | 0
    admitted to the hospital | 0
    emphysema on the skin | 0
    right thigh local tenderness | 0
    back local tenderness | 0
    septic shock | 0
    blood pressure 100/50mmHg | 0
    mean arterial pressure 68mmHg | 0
    heart rate 110bpm | 0
    body temperature 39.0°C | 0
    fluid resuscitation with 2500ml Ringer's lactate | -3
    tobacco abuse | 0
    nickel allergy | 0
    sciatica of the right leg | -2160
    cortisone injections | -2160
    oral non-steroidal anti-inflammatory drugs | -2160
    emergency surgery | 0
    right hemipelvectomy | 0
    double-transverse transversostoma | 0
    debridement into healthy tissue | 0
    soft tissue necrosis | 0
    muscle necrosis | 0
    phlegmonous inflammation of subcutaneous and muscular tissue | 0
    empirical antibiotic fourfold therapy | 0
    Meropenem | 0
    Linezolid | 0
    Penicillin G | 0
    Clindamycin | 0
    postoperative CT scan showing acicular foreign body in upper rectum | 24
    rectoscopy | 24
    toothpick removal | 24
    no clinical improvement | 24
    second control CT showing peritonitis and free intraabdominal air | 48
    immediate laparotomy | 48
    sigmoid colon perforation | 48
    peritonitis | 48
    sigmoid colon resection | 48
    proctosigmoidectomy (Hartmann's procedure) | 48
    three further wound revisions | 72
    rotation flap surgery | 72
    ESBL-Escherichia coli identified | 72
    antibiotic therapy deescalated to Meropenem monotherapy | 120
    Levofloxacin 500mg orally twice a day | 360
    Levofloxacin discontinued | 432
    mobilized with forearm crutches | 432
    transferred to rehabilitation | 1008
    