40 years old | 0
male | 0
admitted to the hospital | 0
motorcycle collision | -1
hypotensive | 0
alert | 0
left needle thoracostomy | 0
decreased breath sounds | 0
intubated | 0
massive transfusion protocol activated | 0
left chest deformity | 0
left chest tube placed | 0
>2000 cc blood | 0
left thoracotomy | 1
multiple comminuted rib fractures | 1
multiple large pulmonary lacerations | 1
left diaphragm injury | 1
bilateral hemothoraces | 1
fragment of bone abutting the pericardium | 1
clamshell thoracotomy | 1
pericardium incised | 1
heart intact | 1
tractotomy | 1
pulmonary hemorrhage controlled | 1
left chest packed | 1
exploratory laparotomy | 1
superficial splenic lacerations | 1
left humerus fracture | 1
left scapula fracture | 1
hypotensive | 2
systolic blood pressures in the low 80s mmHg | 2
hypoxic | 2
massive transfusion | 2
38 packed red blood cells | 2
36 plasma | 2
4 units of platelets | 2
hospital's blood supply exhausted | 2
prognosis poor | 2
vasopressors started | 2
resuscitation continued | 2
failed to respond to additional fluid resuscitation | 4
hemorrhage controlled | 4
empiric hydrocortisone 100 mg | 4
hydrocortisone every 8 h | 4
stabilized | 6
systolic blood pressures into the 150s mmHg | 6
vasopressors weaned | 6
fluids decreased | 6
history of hypopituitarism | -10000
levothyroxine | -10000
hydrocortisone | -10000
returned to the operating room | 48
washout | 48
rib fixation | 48
closure of left chest | 48
extubated | 144
left bronchopulmonary fistula | 150
pulmonary embolism | 150
heparin-induced thrombocytopenia | 150
discharged | 1104
follow-up | 8760
recovered | 8760
returned to work | 8760
no respiratory difficulty | 8760