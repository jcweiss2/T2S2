16 years old | 0 | 0 | Factual
primigravida | 0 | 0 | Factual
admitted to the emergency room | 0 | 0 | Factual
pregnancy diagnosis of 37.6 weeks of gestation | -672 | 0 | Factual
viable intrauterine pregnancy | -672 | 0 | Factual
fetal heart rate of 143 beats per minute | -672 | 0 | Factual
fetus situated longitudinally with cephalic presentation | -672 | 0 | Factual
back to the left | -672 | 0 | Factual
cervix 6 cm dilated | -672 | 0 | Factual
70% effaced | -672 | 0 | Factual
station +1 | -672 | 0 | Factual
intact membranes | -672 | 0 | Factual
mild edema of the extremities | -672 | 0 | Factual
normal osteotendinous reflexes | -672 | 0 | Factual
obstetrical ultrasound | -672 | 0 | Factual
pregnancy of 37+0 weeks of gestation | -672 | 0 | Factual
posterior body placenta maturation grade III | -672 | 0 | Factual
amniotic fluid index of 8.7 cm | -672 | 0 | Factual
biophysical profile of 8/8 | -672 | 0 | Factual
Hadlock of 34.2% | -672 | 0 | Factual
weight of 3033 grams | -672 | 0 | Factual
labor monitoring | 0 | 5 | Factual
spontaneous rupture of the membranes | 0 | 0 | Factual
effective labor | 0 | 5 | Factual
4 contractions every 10 minutes | 0 | 5 | Factual
contractions lasted 40 to 45 seconds | 0 | 5 | Factual
no need for uterotonic agents | 0 | 5 | Factual
live newborn delivered | 5 | 5 | Factual
Apgar scores of 7 and 9 | 5 | 5 | Factual
gestational age of 40 weeks | 5 | 5 | Factual
height 48 cm | 5 | 5 | Factual
weight of 2650 grams | 5 | 5 | Factual
placenta came out with normal characteristics | 5 | 5 | Factual
grade III uterine inversion | 5 | 5 | Factual
manual reinversion maneuvers performed | 5 | 5 | Factual
total blood loss of 1200 mL | 5 | 5 | Factual
uterine atony | 5 | 5 | Factual
oxytocin used | 5 | 5 | Factual
carbetocin used | 5 | 5 | Factual
misoprostol used | 5 | 5 | Factual
persistent uterine inversion | 5 | 5 | Factual
exploratory laparotomy | 5 | 5 | Factual
reinversion successful | 5 | 5 | Factual
persistent uterine atony | 5 | 5 | Factual
persistent postpartum hemorrhage | 5 | 5 | Factual
Hayman hemostatic suture placed | 5 | 5 | Factual
no response to Hayman suture | 5 | 5 | Factual
bilateral ligation of the anterior trunk of the hypogastric artery | 5 | 5 | Factual
immediate recovery of uterine tone | 5 | 5 | Factual
cessation of postpartum hemorrhage | 5 | 5 | Factual
uterus regained tone in approximately 5 minutes | 5 | 10 | Factual
postligation bleeding of 50 mL | 10 | 10 | Factual
transfusion of 2 bags of packed red blood cells | 10 | 10 | Factual
gasometry showed a hemoglobin level of 7 g | 10 | 10 | Factual
transfer to recovery room | 10 | 10 | Factual
transfer to medical intensive care unit | 10 | 10 | Factual
normal diet | 24 | 24 | Factual
ambulation | 24 | 24 | Factual
spontaneous uresis | 24 | 24 | Factual
normal peristalsis | 24 | 24 | Factual
breastfeeding | 24 | 24 | Factual
discharge on the second day | 48 | 48 | Factual
no postoperative complications | 48 | 48 | Factual