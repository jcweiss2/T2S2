25 years old | 0
    male | 0
    admitted to the hospital | 0
    collapse during marathon | -12
    severe hypotension | -12
    unrecordable blood pressure | -12
    intravenous fluids initiated | -12
    confused | 0
    Glasgow Coma Score of 10 | 0
    temperature of 105.4°F | 0
    sweaty | 0
    tachycardic (heart rate 160 bpm) | 0
    systolic blood pressure 90 mm Hg | 0
    elevated creatinine phosphokinase (CPK) 515 U/l | 0
    creatinine 228 μmol/l | 0
    elevated white blood cells 12.3 × 10^9/l | 0
    elevated neutrophils 8.0 × 10^9/l | 0
    elevated haemoglobin 17.8 g/dl | 0
    platelets 254 × 10^9/l | 0
    urea 5.90 mmol/l | 0
    potassium 4.66 mmol/l | 0
    random glucose 4.08 mmol/l | 0
    INR 1.12 | 0
    CPK 515 U/l | 0
    ALP 110 U/l | 0
    ALT 34 U/l | 0
    GGT 29 U/l | 0
    bilirubin 7.4 μmol/l | 0
    lactate 1.8 mmol/l | 0
    drugs of abuse screen negative | 0
    urine myoglobin test negative | 0
    resuscitated with fluids | 0
    low blood pressure requiring ephedrine for 6 hours | 0
    CT scan of brain normal | 0
    started on co-amoxiclav | 0
    elevated CPK 178,850 U/l on day one | 24
    elevated ALT 143 U/l on day one | 24
    transferred to general ward | 24
    ALT peaked at 2,912 U/l on day two | 48
    liver screen normal | 48
    negative viral screen | 48
    negative autoimmune screen | 48
    mildly raised ferritin 621 ng/ml | 48
    ultrasound of liver normal | 48
    discontinued antibiotics | 48
    started intravenous NAC 100 mg/kg 16-hourly | 48
    discharged home | 72
    follow-up with improving CPK and ALT | 72
