83 years old | 0
male | 0
admitted to the hospital | 0
leg ecchymosis | 0
anuric | 0
rhabdomyolysis-induced AKI | 0
sepsis | 0
acute prostatitis | 0
syncope | -12
fell to the ground | -12
lying on the floor | -12
increased urea | 0
increased creatinine | 0
increased myoglobin | 0
increased CPK | 0
increased LDH | 0
increased CRP | 0
increased PCT | 0
increased total bilirubin | 0
increased direct bilirubin | 0
increased AST | 0
increased ALT | 0
increased PSA | 0
increased white blood cell count | 0
volume expansion | 0
diuretic treatment | 0
antibiotic treatment | 0
furosemide | 0
femoral central venous catheter | 0
HFR-Supra | 0
endogenous reinfusion | 0
hydrophobic resin | 0
adsorbent cartridge | 0
low flux polyphenylene membrane | 0
high-dose furosemide | 0
intravenous fluids | 0
24-h urine output 300 mL | 96
24-h urine output 2,400 mL | 192
furosemide tapered | 192
antibiotic therapy | 0
piperacillin/tazobactam | 0
meropenem | 0
E. coli resistant to piperacillin/tazobactam | 0
myoglobin reduction | 120
CPK reduction | 120
LDH reduction | 120
CRP reduction | 120
PCT reduction | 120
HFR-Supra sessions | 120
blood flow 250 mL/min | 0
endogenous ultrafiltrate flow 14 L | 0
low molecular weight heparin | 0
enoxaparin | 0
femoral hemodialysis catheter removed | 144
right jugular central venous catheter | 144
on-line hemodiafiltration | 144
high-flux hemodialysis | 144
Phylter HF 17G dialyzer | 144
dialysis no longer required | 504
discharge | 504
urea 96 mg/dL | 504
creatinine 3.06 mg/dL | 504
CRP 3.2 mg/dL | 504
total bilirubin 0.81 mg/dL | 504
ASL 27 IU/L | 504
ALT 25 IU/L | 504
PSA 61 ng/mL | 504
white blood cells count 6,300 cells/µL | 504
urea 89 mg/dL | 1296
creatinine 2.41 mg/dL | 1296
GFR 24 mL/min | 1296