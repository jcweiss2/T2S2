51 years old | 0
female | 0
admitted to the hospital | 0
general convulsions | 0
diazepam | 0
partial vigilance | 0
vital signs and physical examination were normal | 0
hypertension | -672
ramipril | -672
diabetes mellitus | -672
fast and long-acting insulin | -672
personality disorder | -672
flufenazide | -672
alcohol abuse | -672
laboratory exams | 0
tests for alcohol and drugs were negative | 0
pyometra | 0
extraneous body inside the uterine cavity | 0
focal epileptic activity | 0
levetiracetam | 0
valproate | 0
propofol | 0
phenytoin | 0
intubation | 0
admission to the intensive care unit | 0
endoscopic removal of the extraneous body | 24
antibiotic treatment with clindamycin and gentamicin | 24
septic shock | 120
hypotension | 120
norepinephrine | 120
epinephrine | 120
sustained ventricular tachycardia | 132
amiodarone | 132
DC-shock | 132
diffuse ST-segment elevation | 137
shark-fin sign | 137
echocardiogram | 137
severe reduction of left ventricular function | 137
akinesia of the apex and periapical segments | 137
apical ballooning | 137
coronary angiography | 144
mild stenosis of the mid-left anterior descending artery | 144
Tako-Tsubo syndrome | 144
mild troponin elevation | 144
substitution of phenytoin with levetiracetam | 144
stop of vasopressors | 144
single antiplatelet therapy with aspirin | 144
beta-blockers | 144
ramipril | 144
extubation | 216
discharge from ICU | 216
progressive resolution of the ST-segment elevation | 240
recovery of the left-ventricular function | 240
discharge | 600
asymptomatic | 4320
no further cardiovascular event | 4320