36 years old | 0
male | 0
admitted to the hospital | 0
hypotension | 0
altered mental status | 0
ingestion of unknown quantity of medication | -1
ingestion of metformin | -1
ingestion of trazodone | -1
empty pill bottle found | 0
volume resuscitation initiated | 0
lactic acidosis | 0
hyperkalemia | 0
normal transaminase | 0
normal troponin | 0
normal creatine kinase | 0
undetectable serum acetaminophen | 0
undetectable serum salicylate | 0
normal blood glucose | 0
hypoglycemia | 1
dextrose administered | 1
octreotide administered | 1
acute dialysis catheter placed | 1
hemodialysis initiated | 3.5
norepinephrine drip started | 4
worsening hypotension | 4
worsening mental status | 4
worsening lactic acidosis | 4
intubated | 5
vasoplegia | 5
high doses of norepinephrine | 5
high doses of vasopressin | 5
high doses of epinephrine | 5
high doses of phenylephrine | 5
echocardiography | 5
normal left ventricular function | 5
normal right ventricular function | 5
bicarbonate pushes | 5
bicarbonate drip | 5
hydroxocobalamin administered | 5
methylene blue administered | 6
transient improvement in blood pressure | 6
CRRT attempted | 7
CRRT discontinued | 7
VA ECMO support initiated | 19
cannulation | 19
peripheral cannulation | 19
VA ECMO support | 19
CRRT reinitiated | 20
shock resolved | 48
decannulation | 48
vasopressors discontinued | 48
lactic acid normalized | 96
mental status improved | 96
extubated | 96
discharged | 480
metformin level 678 μg/mL | 0
trazodone level 2.1 μg/mL | 0
mCPP found in urine | 0
mCPP not found in serum | 0
metformin level 309 μg/mL | 5.5
metformin level 255 μg/mL | 10.5
metformin level 219 μg/mL | 11.5
urine metformin level 2224 μg/mL | 12
trazodone level 2.4 μg/mL | 5.5
trazodone level 1.1 μg/mL | 10.5
trazodone level 0.8 μg/mL | 11.5
urine trazodone level 3.6 μg/mL | 12