34 years old | 0
male | 0
Marfan syndrome | -8760
admitted to the hospital | 0
dyspnea | -72
tachycardia | 0
fever | 0
infective endocarditis | 0
heart rate 118 beats/min | 0
blood pressure 92/45 mmHg | 0
peripheral oxygen saturation 85% | 0
body temperature of 38.6°C | 0
COVID-19 infection | -72
positive real-time polymerase chain reaction test for COVID-19 | 0
moved to a negative-pressure room in the ICU | 0
high-resolution computed tomography of the chest | 0
bilateral ground glass opacities | 0
interlobular septal thickening | 0
dependent consolidation | 0
transthoracic echocardiography | 0
mechanical bileaflet prosthetic valve | 0
suspected vegetations on the leaflets | 0
dehiscence of the aortic root | 0
para-aortic abscess | 0
moderate aortic regurgitation | 0
no pericardial effusion | 0
CT aortogram | 0
contrast leakage in the mediastinum | 0
anemia | 0
leukocytosis | 0
thrombocytopenia | 0
high procalcitonin | 0
high interleukin-6 | 0
meropenem | 0
vancomycin | 0
remdesivir infusion | 0
urgent cardiac surgery | 0
EuroSCORE II 10.82% | 0
negative-pressure operating room | 0
cardiopulmonary bypass | 0
CytoSorb hemoadsorber | 0
myocardial protection | 0
moderate hypothermia | 0
antegrade Custodiol crystalloid cardioplegia | 0
alpha-stat blood gas management | 0
redo sternotomy | 0
thorough cleaning of the pus | 0
extraction of the previous valve graft | 0
creation of a neo-annulus | 0
redo Bentall procedure | 0
porcine root | 0
intraoperative epinephrine | 0
intraoperative norepinephrine | 0
red blood cells transfusion | 0
fresh frozen plasma transfusion | 0
platelet apheresis transfusion | 0
postoperative ventilation | 48
weaned from the ventilator | 48
inotropes | 48
inflammatory markers improvement | 48
hemodynamic parameters improvement | 48
discharged | 120 
Note: The time stamp is an approximation based on the text and may not be exact. The events that happened before admission to the hospital are assigned a negative time stamp, and the events that happened after admission are assigned a positive time stamp. The time stamp 0 is assigned to the events that happened at the time of admission or have no specific time mentioned.