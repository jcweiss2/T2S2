49 years old | 0
female | 0
hepatocellular carcinoma | 0
end-stage hepatitis B liver cirrhosis | 0
MELD score 14 | 0
Child-Pugh class B | 0
hypertension | 0
medications for hypertension | 0
blood type A | 0
Rh+ | 0
ABO compatible donor | 0
donor son | 0
anesthesia induced | 0
fentanyl | 0
thiopental sodium | 0
vecuronium | 0
oxygen | 0
air | 0
desflurane | 0
neuromuscular block | 0
atracurium | 0
hemodynamic monitoring | 0
surgery proceeded | 0
piggyback technique | 0
preservation of caval flow | 0
reperfusion of graft liver | 0
right posterior sectionectomy | 0
improved right hepatic venous flow | 0
graft blood flow did not improve | 0
intractable bleeding | 0
hypovolemia | 0
cardiac arrest | 0
chest compression | 0
epinephrine | 0
volume resuscitation | 0
fluid management system | 0
cardiopulmonary resuscitation | 0
spontaneous circulation | 0
normal sinus rhythm | 0
arterial blood gas analysis | 0
coagulation profiles | 0
serum potassium level elevated | 0
serum calcium level decreased | 0
hematocrit level decreased | 0
oozing continued | 0
surgical hemostasis | 0
stop surgery | 0
intensive medical treatment | 0
planned second operation | 0
gauze packing | 0
transferred to surgical intensive care unit | 0
operation time 1,270 minutes | 0
crystalloid infused | 0
5% albumin infused | 0
colloid infused | 0
leukocyte depleted red blood cell infused | 0
leukocyte depleted platelet concentrate infused | 0
cell saver blood infused | 0
fresh frozen plasma infused | 0
cryoprecipitate infused | 0
urine output | 0
estimated blood loss | 0
metabolic acidosis | 24
azotemia | 24
severe hypoxemia | 24
fraction of inspired oxygen 1.0 | 24
mechanical ventilation | 24
positive end-expiratory pressure | 24
pulmonary congestion | 24
echocardiography | 24
cardiac physiology normal | 24
cardiac function normal | 24
cardiac structure normal | 24
anuria | 31
continuous renal replacement therapy | 31
brain tomography | 31
no abnormal finding | 31
VV ECMO initiated | 48
cardiologist evaluation | 48
no cardiac support needed | 48
central cannula removed | 48
Swan-Ganz catheter removed | 48
drainage cannula placed | 48
return cannula placed | 48
CAPIOX emergent bypass system | 48
circuit primed | 48
CAPIOX EBS oxygenator kit | 48
CRRT continued | 48
VV ECMO circulation | 48
sweep gas flow | 48
heparin not used | 48
antithrombin injected | 48
activated clotting time measured | 48
ECMO treatment | 48
patient's condition improved | 72
SpO2 95% | 72
FiO2 0.3-0.4 | 72
FiO2 1.0 | 72
second LT | 72
deceased donor LT | 72
warm ischemic time | 72
cold ischemic time | 72
perioperative ABGA profiles | 72
coagulation profiles | 72
preoperative chest radiograph | 72
pulmonary congestion | 72
bilateral pleural effusions | 72
MELD score 30 | 72
ECMO support | 72
CRRT support | 72
discontinued CRRT | 72
restarted CRRT | 72
anesthesia management | 72
femoral arterial blood pressure | 72
pulmonary arterial pressure | 72
cardiac output monitoring | 72
core temperature monitored | 72
fluid heated | 72
peripheral vascular access removed | 72
warm blanket | 72
humidifier | 72
patient's limbs covered | 72
room temperature maintained | 72
anesthetic management | 72
SpO2 stable | 72
FiO2 0.5 | 72
tidal volume | 72
respiratory rate | 72
PEEP | 72
body temperature maintained | 72
compartment syndrome | 72
abdominal closure | 72
total administered volume | 72
crystalloid | 72
colloid | 72
5% dextrose water | 72
cell saver autotransfusion | 72
leukocyte-depleted red blood cell | 72
fresh frozen plasma | 72
plateletpheresis | 72
cryoprecipitate | 72
hematocrit level maintained | 72
no severe oozing | 72
no acute massive bleeding | 72
no hypotensive episode | 72
urine not excreted | 72
sedation maintained | 72
midazolam | 72
fentanyl | 72
CRRT restarted | 72
ECMO continued | 72
body temperature maintained | 72
forced-air warmer | 72
heated humidifier | 72
pre-warmed fluid | 72
Glasgow coma scale | 72
pupil size | 72
light reflex | 72
limb movement | 72
orientation | 72
pupil dilatation | 72
light reflex normal | 72
neurologic abnormalities | 72
ECMO weaning | 104
bypass flow reduced | 104
oxygen flow reduced | 104
FiO2 increased | 104
ABGA performed | 104
ECMO removed | 106
PaO2/FiO2 ratio improved | 106
PaCO2 level similar | 106
ventilatory demand decreased | 106
PaO2/FiO2 stabilized | 106
SpO2 over 90% | 106
FiO2 0.6 | 106
laparotomy wound closure | 132
liver congestion | 133
hepatic drainage failed | 133
surgical decompression | 133
stenosis at intrahepatic IVC | 138
stenting | 138
graft failure | 138
long-term use of high dose vasopressor | 138
leg necrosis | 138
sepsis | 138
fentanyl stopped | 138
cisatracurium stopped | 138
eye opening | 138
low grade motor responses | 138
no further improvement | 138
expired | 168
multi-organ failure | 168
graft failure | 168
uncontrolled sepsis | 168