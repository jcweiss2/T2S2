80 years old | 0 | 0 
male | 0 | 0 
admitted to the hospital | 0 | 0 
urinary tract infection | -120 | 0 
fever | -120 | 0 
dysuria | -120 | 0 
clean catch urine specimen | -120 | -120 
urine analysis | -120 | -120 
leukocyte esterase | -120 | -120 
bacteria | -120 | -120 
Escherichia coli | -120 | -120 
cephalexin | -120 | -48 
rash | -48 | 0 
sloughing of the skin | -24 | 0 
discontinued cephalexin | 0 | 0 
transferred to BICU | 0 | 0 
chronic obstructive pulmonary disease | 0 | 0 
type 2 diabetes mellitus | 0 | 0 
coronary artery disease | 0 | 0 
hypertension | 0 | 0 
hypothyroidism | 0 | 0 
depression | 0 | 0 
end-stage renal disease | 0 | 0 
hemodialysis | 0 | 0 
myocardial infarctions | 0 | 0 
ischemic cardiomyopathy | 0 | 0 
atrial fibrillation | 0 | 0 
hydrocodone/acetaminophen | 0 | 0 
levothyroxine | 0 | 0 
escitalopram | 0 | 0 
carvedilol | 0 | 0 
guaifenesin | 0 | 0 
docusate | 0 | 0 
calcitriol | 0 | 0 
albuterol | 0 | 0 
amiodarone | 0 | 0 
pulmonary infiltrates | 24 | 24 
respiratory failure | 24 | 24 
intubated | 24 | 24 
difficulty swallowing | 24 | 24 
endotracheal tube | 24 | 24 
toxic epidermal necrolysis syndrome | 0 | 0 
body surface area skin detachment | 0 | 0 
cutaneous erythema | 0 | 0 
blister formation | 0 | 0 
hemorrhagic eruptions | 0 | 0 
stomatitis | 0 | 0 
conjunctivitis | 0 | 0 
full-thickness necrosis | 0 | 0 
blood pressure | 0 | 0 
respiratory rate | 0 | 0 
temperature | 0 | 0 
white blood cell count | 0 | 0 
neutrophils | 0 | 0 
platelet count | 0 | 0 
serum creatinine | 0 | 0 
venous serum lactate | 0 | 0 
oxygen saturation | 0 | 0 
pain | 0 | 0 
peripheral blood cultures | 24 | 24 
skin surveillance cultures | 24 | 24 
urine culture | 24 | 24 
chest radiograph | 24 | 24 
right pleural effusion | 24 | 24 
right lower and left basilar opacities | 24 | 24 
norepinephrine | 24 | 120 
vasopressin | 24 | 120 
albumin | 24 | 120 
lactated Ringer’s | 24 | 120 
tetanus–diphtheria toxoids vaccine | 24 | 24 
gentamicin | 24 | 72 
fluconazole | 24 | 120 
WBC | 48 | 48 
SCr | 48 | 48 
venous serum lactate | 48 | 48 
random serum gentamicin level | 48 | 48 
supportive continuous renal replacement therapy | 48 | 120 
fluconazole | 48 | 120 
Gram’s stain | 48 | 48 
tracheal aspirate | 48 | 48 
Pseudomonas aeruginosa | 48 | 48 
gentamicin | 96 | 96 
amiodarone | 96 | 96 
wide complex tachycardia | 96 | 96 
physical examination | 120 | 120 
sloughing of skin | 120 | 120 
culture and sensitivity results | 120 | 120 
Pseudomonas aeruginosa | 120 | 120 
gentamicin | 120 | 120 
expired | 144 | 144 
cardiac arrest | 144 | 144 
multisystem organ failure | 144 | 144 
autopsy | 144 | 144 
necrotizing bronchopneumonia | 144 | 144 
SCORTEN | 144 | 144 
predicted mortality | 144 | 144