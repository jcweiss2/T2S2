29 years old | 0
female | 0
gravida I para I | 0
admitted to the hospital | 0
right hip and flank pain | -504
right flank bruising | -504
pain started | -672
uncomplicated spontaneous vaginal delivery | -168
severe right flank pain | -168
Crohn’s disease | -4320
Methadone | -672
Azathioprine | -672
acute flares | -730
severe abdominal pain | -730
vomiting | -730
bloody diarrhea | -730
Infliximab infusions | -730
stopped Infliximab infusions | -168
mild acute flares | -168
oral prednisone | -168
copper intrauterine device | -672
no history of sexually transmitted diseases | -672
fever | 0
pulse 177 bpm | 0
blood pressure 106/62 mmHg | 0
white blood cell count 50 000 cells/mm3 | 0
elevated platelet count 717 mcL | 0
hemoglobin 6.0 g/dL | 0
lactic acid level 5.2 mmol/L | 0
elevated alkaline phosphatase 207 unit/L | 0
no acute abnormalities on chest X-ray | 0
large complex air-fluid collection | 0
diagnosed with severe sepsis | 0
retroperitoneal abscess | 0
taken to the operating room | 0
incision, drainage, and debridement | 0
ileal perforation | 0
ileal resection | 0
transferred to the intensive care unit | 0
intubated | 0
OR cultures grew Escherichia coli | 0
OR cultures grew Beta Hemolytic Group C Streptococcus | 0
IV Meropenem | 0
IV Vancomycin | 0
IV Clindamycin | 0
additional debridement | 24
irrigation of the necrotizing soft-tissue infection | 24
wound vacuum-assisted closure device | 24
transferred to the medical floor | 96
worsening sepsis | 168
tachycardia | 168
tachypnea | 168
fever | 168
leukocytosis 62 000 cells/mm3 | 168
acute respiratory failure | 168
exploratory laparotomy | 216
intraperitoneal abscess | 216
transverse colon staple line leak | 216
purulence | 216
drainage of the abscess | 216
repair of the leak | 216
omentum patch | 216
Enterococcus faecalis | 216
Candida albicans | 216
Vancomycin | 216
Micafungin | 216
transferred to the medical floor | 264
continued to improve | 264
discharged to long-term acute care | 336
IV antibiotic therapy | 336
aggressive wound management | 336
left the long-term care facility | 840