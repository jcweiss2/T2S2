45 years old | 0
female | 0
presented to first ED | -168
7-day history of fevers | -168
headache | -168
arthralgias | -168
nausea | -168
fatigue | -168
neck pain | -168
tachycardic at first ED | -168
afebrile at first ED | -168
no rash at first ED | -168
normal labs | -168
unremarkable CT | -168
diagnosed with viral illness | -168
discharged from first ED | -168
presented to second ED | 0 (since it's part of the admission process)
worsening confusion | 0
combativeness | 0
dyspnea | 0
ataxia | 0
