19 years old | 0
male | 0
admitted to the hospital | 0
fever | -144
headache | -144
nausea | -144
vomiting | -144
leukocytosis | 0
neutrophils | 0
thrombocytopenia | 0
elevated aspartate transaminase | 0
elevated alanine transaminase | 0
elevated C-reactive protein | 0
anti-HIV test negative | 0
sepsis | 0
admitted to the intensive care unit | 0
sepsis protocol performed | 0
blood sample collected | 0
broad-spectrum antibiotic therapy started | 0
ceftriaxone administered | 0
metronidazole administered | 0
oxacillin administered | 0
mechanical ventilation | 0
brain CT scan performed | 0
heterogeneous collection with air foci | 0
partial sagittal sinus thrombosis | 0
paranasal sinus CT scan performed | 0
right frontal, maxillary and ethmoidal sinus disease | 0
soft tissue drainage performed | 12
neurosurgical drainage performed | 168
gram-positive cocci identified | 24
anticoagulation initiated | 24
enoxaparin administered | 24
S. constellatus identified | 24
antimicrobial therapy changed | 24
vancomycin administered | 24
metronidazole continued | 24
sensory improvement | 672
discharged | 720
follow-up | 4320
no sequelae | 4320