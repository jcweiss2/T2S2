29 years old|0
male|0
admitted to the hospital|0
unresponsive|-120
out-of-hospital cardiac arrest|0
initiated cardiac pulmonary resuscitation|0
ventricular fibrillation|0
defibrillator-delivered electrical shocks (200 J and 300 J)|0
intubated|0
sinus tachycardia (120 bpm)|0
no chest pain|0
no palpitations|0
no syncope|0
no sudden cardiac death prior to admission|0
blood pressure 122/70 mmHg|0
temperature 38.5 °C|0
pulse 102 bpm|0
respiratory rate 22 bpm|0
small amount of moist rales in the lungs|0
normal general physical examinations|0
no history of previous disease|0
family history of Brugada syndrome|0
no family history of sudden cardiac death|0
post-arrest ECG typical type 1 Brugada pattern|0
coved-type ST-segment elevations > 2 mm in V1 to V2|0
negative T-wave in two right precordial leads|0
elevated white blood cell count (21.9 × 109/L)|0
elevated neutrophil count (92.7%)|0
low hemoglobin level (71 g/L)|0
elevated creatine kinase (4600 IU/L)|0
elevated CK-MB (75 IU/L)|0
elevated urea (36 mmol/mL)|0
elevated creatinine (1079 µmol/mL)|0
elevated serum alanine transaminase (296 IU/L)|0
elevated aspartate aminotransferase (426 IU/L)|0
elevated total bilirubin (40.9 µmol/L)|0
elevated direct bilirubin (12.8 µmol/L)|0
elevated procalcitonin (22 ng/mL)|0
elevated D-dimer (7141 ng/mL)|0
elevated fibrinogen degradation products (93 µg/mL)|0
prolonged activated partial thromboplastin time (91.4 s)|0
elevated brain natriuretic peptides (5623 ng/L)|0
normal electrolytes|0
echocardiography no structural disease|0
chest radiography pulmonary infection|0
head CT no infarction or hemorrhage|0
diagnosis of Brugada syndrome|0
diagnosis of NYHF IV|0
diagnosis of multiple organ dysfunction syndrome|0
diagnosis of sepsis|0
diagnosis of hypoxic ischemic encephalopathy|0
induced-hypothermia protocol|0
sedation|0
analgesia|0
continuous renal replacement therapy|0
Linezolid injection 600 mg twice a day for 7 days|0
Sulperazon injection 3 g twice a day|0
Mycamine injection 50 mg twice a day|0
correcting water-electrolyte balance|0
correcting acid-base balance|0
nutritional support|0
protecting hepatorenal function|0
tracheotomy performed|480
no further episodes of VT/VF|480
various ECG changes in the same lead during treatment|0
refused ICD for secondary prevention of SCD|480
brother received Reveal LINQ ICM for primary prevention of SCD|480
recommended genetic testing|480
no arrhythmia episodes after discharge|864
good physical condition 3 years later|26208
subsequent ECGs normal sinus rhythm|864
brother's remote monitoring no ventricular arrhythmia|864
brother's ECG sinus rhythm during follow-up|864
fever for more than 9 days|0
pulmonary infection|0
sepsis|0
education and lifestyle measures for prevention of arrhythmia events|0
informed about precipitating factors|0
fever treated immediately with antipyretics|0
multidisciplinary team cooperation|0
