40 years old | 0  
    male | 0  
    Graves’ disease | -175200  
    paroxysmal atrial flutter | -175200  
    admitted to the hospital | 0  
    resuscitation | 0  
    cardiac arrest | 0  
    ventricular fibrillation | 0  
    no risk factors for ischemic heart disease | 0  
    electrocardiogram showed atrial fibrillation | 0  
    ventricular extra systoles | 0  
    q-waves in anterior leads | 0  
    in hospital heart monitoring showed paroxysmal complete heart block | 0  
    elevated troponin-T | 0  
    elevated creatine kinase myocardial band | 0  
    elevated total CK | 0  
    chest X-ray showed cardiomegaly | 0  
    transthoracic echocardiography disclosed dilatation of left ventricle | 0  
    left ventricular ejection fraction 25-30% | 0  
    hypofunction of right ventricle | 0  
    inferoseptal akinesia | 0  
    coronary angiography showed normal coronary arteries | 0  
    cardiac magnetic resonance imaging confirmed inferoseptal akinesia | 0  
    late gadolinium enhancement in subendocardial pattern | 0  
    implantation of Cardiac-Resynchronization-Therapy-Defibrillator device | 0  
    anticoagulants | 0  
    antiarrhythmics | 0  
    statin | 0  
    heart failure therapy | 0  
    muscle weakness for 2 years | -17520  
    elevated total CK tracing back to 2014 | -17520  
    muscle strength testing confirmed proximal weakness | 0  
    no signs of rheumatic/neurologic disease | 0  
    followed by cardiologists and neurologists | 0  
    progressive muscular weakness | 0  
    repetitive supraventricular arrhythmias | 0  
    repetitive ventricular arrhythmias | 0  
    elevated cardiac enzymes | 0  
    elevated muscle enzymes | 0  
    serological tests for myositis-specific autoantibodies negative | 0  
    anti-HMGCR negative | 0  
    ANA negative | 0  
    genetics for neuromuscular diseases negative | 0  
    whole-body PET-CT normal | 0  
    pulmonary function tests normal | 0  
    muscle biopsy showed fiber variability | 0  
    muscle biopsy showed cell necrosis compatible with immune-mediated necrotizing myopathy | 0  
    initiation of prednisolone 75 mg/day | 0  
    improved physical performance | 0  
    addition of methotrexate 15-25 mg/week | 0  
    prednisolone tapered | 0  
    continued clinical improvement | 0  
    stable LVEF of 35% | 0  
    experienced worsening of muscle weakness | 0  
    experienced dyspnea | 0  
    rising total CK | 0  
    X-ray revealed pulmonary congestion | 0  
    condition improved transitorily on diuretics | 0  
    increased MTX to 25 mg/week | 0  
    brought to intensive care in cardiogenic shock | 0  
    decompensated severe biventricular failure | 0  
    stabilized by inotropic support | 0  
    stabilized by diuretics | 0  
    stabilized by amiodarone | 0  
    upregulation of CRT pace | 0  
    glucocorticoids | 0  
    TTE depicted biventricular hypofunction/dilatation | 0  
    LVEF 10-15% | 0  
    cardiac PET-CT showed nonviable perfusion defect | 0  
    myocardial biopsy revealed mild to moderate hypertrophy | 0  
    replacement fibrosis | 0  
    alcian-positive matrix indicating presence of glycosaminoglycans | 0  
    endothelial proliferation | 0  
    few inflammatory cells | 0  
    recent loss of myocytes | 0  
    addition of cyclosporine 200 mg/day | 0  
    addition of mycophenolate mofetil 2 g/day | 0  
    prednisolone 15 mg/day | 0  
    stable peripheral muscle function | 0  
    no convincing cardiac effect | 0  
    testing for AMA | 0  
    AMA present in high titers | 0  
    diagnosis of cardiomyopathy related to AMA-associated inflammatory myositis | 0  
    initiation of rituximab therapy | 0  
    no cardiac improvement | 0  
    severe chronic renal impairment | 0  
    liver failure | 0  
    not a candidate for heart transplantation | 0  
    death in cardiogenic and septic shock | 0  
    death | 0  
    
