46 years old | 0
male | 0
benign prostatic hyperplasia | -672
end-stage renal disease | -672
hemodialysis | -672
peritonitis | 0
septic shock | 0
pneumoperitoneum | 0
diagnostic laparoscopy | 0
gross bilious contamination | 0
perforation of the anterior duodenal bulb | 0
modified Graham patch | 0
endoscopic leak test | 0
open approach | 0
midline laparotomy | 0
Graham patch reconstruction | 0
repeat endoscopic leak test | 0
abdomen irrigation | 0
drains placement | 0
abdomen closure | 0
intra-abdominal abscess | 168
percutaneous drainage | 168
Helicobacter pylori | 0
triple therapy | 0
discharged | 216
hematochezia | 744
symptomatic anemia | 744
transfusion | 744
computed tomography angiography | 744
inferior vena cava thrombus | 744
intraluminal air formation | 744
duodenal-caval fistula | 744
upper endoscopy | 744
clots | 744
bleeding | 744
exploratory laparotomy | 768
Kocher maneuver | 768
duodenal-caval fistula identification | 768
Pringle maneuver | 768
right renal artery ligation | 768
right renal vein ligation | 768
right ureter ligation | 768
transesophageal echocardiography | 768
intraoperative ultrasound | 768
thrombectomy | 768
venorrhaphy | 768
duodenal perforation repair | 768
nasogastric tube placement | 768
abdomen temporary closure | 768
AbThera wound vacuum device | 768
intensive care unit | 768
re-exploration | 792
open cholecystectomy | 792
right nephrectomy | 792
abdomen temporary closure | 792
AbThera device | 792
intensive care unit | 792
abdomen opening | 816
duodenal repair inspection | 816
omentum patch placement | 816
pyloric exclusion | 816
gastrostomy | 816
gastrojejunostomy | 816
enterolysis | 816
nasojejunal tube placement | 816
distal feeding tube placement | 816
drains placement | 816
abdomen closure | 816
hemorrhagic shock | 1008
intraluminal bleeding | 1008
anomalous duodenal artery | 1008
angioembolization | 1008
subhepatic fluid collection | 1092
percutaneous drainage | 1092
bleeding | 1216
angioembolization | 1216
discharged | 1680