37 years old | 0
    female | 0
    vaginal delivery | -96
    twins | -96
    lateral episiotomy | -96
    HIV serology | -96
    hepatitis serology | -96
    vaginal swabs | -96
    urine culture | -96
    discharged | -72
    abdominal pain | 0
    septic shock | 0
    axillary temperature 36°C | 0
    blood pressure 80/30 mmHg | 0
    tachycardia 130/min | 0
    marbling | 0
    cold limbs | 0
    free intra-abdominal fluid | 0
    fluid resuscitation | 0
    catecholamine use | 0
    noradrenaline 0.5-2 μg/kg/min | 0
    tachypnea 30 cycles/min | 0
    unspecific bowel infection | 0
    imipenem 1g | 0
    amikacin 20 mg/kg | 0
    teicoplanin 400 mg | 0
    hemoglobin 9.2 g/dL | 0
    leukocytes 1540×10³/μL | 0
    platelet count 104000/μL | 0
    C-reactive protein 340 mg/dL | 0
    creatinine 1.92 mg/dL | 0
    albumin 1.2 g/dL | 0
    cytolysis | 0
    ALT 120 UI/L | 0
    AST 146 UI/L | 0
    cholestasis | 0
    metabolic acidosis pH 7.12 | 0
    arterial lactate 8.9 mmol/L | 0
    SOFA score 9 | 0
    exploratory laparotomy | 0
    purulent fluid | 0
    venous congestion | 0
    bladder inspection | 0
    uterus inspection | 0
    adnexa inspection | 0
    bowel inspection | 0
    normal appendix | 0
    peritoneal lavage | 0
    pelvic drain | 0
    mesenteric ischemia suspicion | 0
    heparin 50 mg | 0
    CT scan abdomen | 0
    intraperitoneal free fluid | 0
    paralytic ileus | 0
    fluid culture | 0
    blood culture | 0
    Group A streptococci | 0
    intensive care transfer | 0
    multiorgan failure | 0
    disseminated intravascular coagulation | 0
    death | 12
    