26 years old | 0
G1P1 | 0
routine prenatal care | -672
serologies were all negative or nonreactive | -672
spontaneous labor | -8
spontaneous rupture of membranes | -8
delivery | 0
male | 0
appropriate for gestational age | 0
2.92 kg | 0
no resuscitation was required | 0
Apgar's scores were normal | 0
admitted for normal newborn cares | 0
respiratory distress | 5
grunting | 5
lethargic | 5
hypoglycemic | 5
blood glucose: 26 mg/dL | 5
oxygen was initiated via nasal cannula | 5
concern for bacterial sepsis | 5
IV access was obtained | 5
empiric administration of ampicillin and gentamicin | 5
chest X-ray revealed bibasilar infiltrates | 5
complete blood count revealed severe leukopenia | 5
white blood cell count: 2.3 × 10e9/L | 5
NICU referral was made | 5
transport team intubated the infant | 5
fluid resuscitation was started | 5
progressive respiratory failure | 5
poor perfusion | 5
lactic metabolic acidosis | 12
leukopenia with severe neutropenia | 12
absolute neutrophil count: 500 × 10e9/L | 12
thrombocytopenia | 12
platelet count 111 × 10e9/L | 12
no coagulopathy | 12
no evidence of other end organ dysfunction | 12
chest radiograph revealed continued infiltrates | 12
blood culture grew gram-negative rods | 12
evaluation for other infectious foci | 12
lumbar puncture | 12
urinary catheterization | 12
tracheal aspiration | 12
cerebrospinal fluid analysis showed normal white blood cell count | 12
elevated red blood cell count | 12
normal protein and glucose concentrations | 12
negative Gram's stain | 12
urinalysis was unremarkable | 12
tracheal aspirate showed few gram-negative rods | 12
fewer than 25 polymorphonuclear cells | 12
persistent pulmonary hypertension | 12
progressive septic shock | 12
continued hypotension | 12
poor perfusion | 12
infectious diseases consultation was obtained | 12
antibiotics were broadened to include meropenem | 12
fluid resuscitation | 12
multiple vasoactive medications | 12
inhaled nitric oxide | 12
improve oxygenation | 12
persistent fetal circulation | 12
blood and tracheal cultures revealed P. multocida | 12
organism was susceptible to all agents tested | 12
ampicillin | 12
ceftriaxone | 12
levofloxacin | 12
penicillin | 12
trimethoprim-sulfa | 12
azithromycin | 12
cerebral spinal fluid and urine cultures were both negative | 12
subsequent blood cultures were negative | 12
multiple pets in the parents' home | 12
two cats | 12
one dog | 12
family members denied any history of bites or scratches | 12
maternal vaginal culture was obtained | 12
maternal vaginal culture was positive for P. multocida | 12
mother did not endorse any vaginal symptoms | 12
molecular diagnostic studies were performed | 12
positive cultures from the patient's blood and tracheal aspirate | 12
maternal vaginal specimen | 12
initial identification as P. multocida | 12
matrix-assisted laser desorption ionization–time of flight (MALDI-TOF) mass spectrometry | 12
16S rRNA gene sequencing | 12
polymerase chain reaction (PCR) | 12
Applied Biosystems 3130 Genetic Analyzer | 12
GenBank database | 12
basic local alignment search tool (BLAST) algorithm | 12
P. multocida, subspecies septica | 12
100% match | 12
National Center for Biotechnology Information (NCBI) nucleotide BLAST function | 12
three separate sequences of the three bacterial isolates were a 100% match | 12
neonatal EOS with pneumonia | 12
vertical transmission from the mother | 12
maternal vaginal colonization | 12
related to pet exposure in her home | 12
no specimens from those animals were obtained | 12
Infectious Diseases Service recommended treatment of the mother | 12
amoxicillin-clavulanic acid | 12
10-day course | 12
mother sought infectious diseases consultation | 12
subsequent pregnancies | 12
vaginal colonization testing | 12
infant made steady clinical progress | 120
ventilator and cardiovascular support were weaned | 120
hemodynamically stable | 120
without need for respiratory support | 120
neutropenia quickly resolved | 120
thrombocytopenia initially worsened | 120
nadir of 36 × 10e9/L | 120
one transfusion | 120
eventual normalization | 120
C-reactive protein levels peaked | 60
174 mg/L | 60
normalization | 168
antibiotic therapy was narrowed | 168
ceftazidime | 168
gentamicin | 168
synergy | 168
completed a 14-day course of antibiotics | 168
single agent ceftazidime | 168
infant was discharged to home | 408
with his parents | 408
infancy was without noted morbidities | 408