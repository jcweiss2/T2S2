63 years old | 0
female | 0
168 cm height | 0
53 kg weight | 0
papillary thyroid carcinoma | -9720
resection | -9720
radiotherapy | -9720
stenosis of the esophagus | -8760
repeated aspiration | -8760
respiratory insufficiency | -8760
pneumonia | -8760
purulent pleurisy | -8760
pleurectomy | -8760
restrictive ventilation pattern | -8760
recurrent nerve palsy | -8760
percutaneous endoscopic gastrostomy | -8760
tracheostoma | -8760
home ventilation | -8760
decreased mobility | -8760
secondary depression | -8760
fixed mandible | -8760
limited mouth opening | -8760
stented left axis vertebralis | -4380
stenosis of the internal axis carotis | -4380
arterial hypertension | -4380
secondary lactase deficiency | -4380
esophageal stenosis dilation | -120
fistula between the esophagus and tracheal membrane | -120
decreasing general condition | 0
admitted to the University of Erlangen | 0
examined by chiefs and consultants | 0
deemed too unstable for open surgery | 0
inability to open the mouth | 0
recurrent nerve palsy | 0
minimal invasive orthograde approach impossible | 0
referred to the surgical intensive care unit | 15
pneumonia by 4-multiresistente gramnegative Pseudomonas aeruginosa | 15
veno-venous extracorporeal membrane oxygenation | 15
partial thromboplastin time of 60 seconds | 15
preseptic status | 15
ventilated through a tracheostoma | 15
thoracic computed tomography | 16
big fistula of the tracheal membrane | 16
tracheal cannula ended shortly beneath the lower limit of the mediastinal fistula | 16
decision to try endobronchial stenting | 17
plan to close the fistula with a pedicled omentum majus replacement | 17
surgical plastic needed an abutment and a secured continuous airway replacement | 17
procedure performed | 17
vv-ECMO began to be partly ineffective | 17
high volume input of physiological saline | 17
oral approach only allowed a small flexible bronchoscope | 17
approach for the upper part of the trachea had to be performed through the percutaneous tracheostoma | 17
retrograde stenting performed in four steps | 17
Step I | 17
Step II | 18
Step III | 19
Step IV | 20
successful retrograde stenting | 20
lungs not aerated | 20
spontaneous breathing work increased | 20
vv-ECMO support reduced | 20
lungs became re-aerated | 20
patient woke up | 20
patient could communicate with her family | 20
infections continued to be severe | 20
spontaneous work of breathing never exceeded a tidal ventilation of 170 mL per breath | 20
reduction of intravenous saline injection limited | 20
vv-ECMO support reduced | 20
patient died | 360
cause of death: pulmonary infection | 360