10 years old | 0
male | 0
diagnosed with high-risk early T-cell precursor acute lymphoblastic leukemia | 0
treated according to LAL SEHOP-PETHEMA 2013 protocol | 0
developed an early CNS relapse | -336
treated according to the InteReALL HR 2010 with bortezomib protocol | -336
neutropenic for four weeks | -672
receiving prophylaxis with cefepime | -672
receiving prophylaxis with cotrimoxazole | -672
receiving prophylaxis with fluconazole | -672
treated with acyclovir for herpes simplex virus type 1 skin infection | -672
developed an intense holocranial headache | 0
cranial computed tomography scan showed a hypodense lesion in the right temporal lobe | 0
lumbar puncture was performed | 0
cefepime was replaced by meropenem and vancomycin | 0
developed septic shock signs | 24
transferred to the pediatric intensive care unit | 24
inotropic and vasoactive support | 24
antimicrobial spectrum was broadened with gentamycin and caspofungin | 24
blood analysis showed a progressive increase of C reactive protein and procalcitonin | 24
hematological analysis showed pancytopenia due to chemotherapy | 24
microbiological blood tests ruled out bacteremia and fungemia | 24
all herpes viruses were negative | 24
urine and stool cultures were also negative | 24
biochemical analysis of the cerebrospinal fluid was strictly normal | 24
B. cereus was detected in microbiologic study | 24
electroencephalogram showed a diffuse slowing of brain activity | 72
cranial magnetic resonance was performed | 96
showed two hyperintense lesions in T2 and FLAIR sequences | 96
parietal lesion presented ring-enhancing after gadolinium administration | 96
small hemorrhagic foci dispersed throughout the parenchyma were observed | 96
diagnosis of B. cereus abscess | 96
treated with meropenem, vancomycin, and gentamycin | 96
evolved favorably with no headache or findings on neurological examination | 336
control magnetic resonance showed a decrease in the size of the lesion | 336
vancomycin and acyclovir were suspended | 504
meropenem was maintained over six weeks | 504