43 years old | 0
male | 0
admitted to hospital | 0
cough | -168
high fever | -168
anosmia | -168
nasopharyngeal PCR swab | 0
SARS-CoV-2 positive | 0
gout | 0
hypertension | 0
chronic kidney disease | 0
unprovoked lower limb venous thromboembolism | -1728
lupus anticoagulant positive | -1728
B2-glycoprotein IgG negative | -1728
anti-cardiolipin IgM negative | -1728
homocysteine normal | -1728
anti-thrombin III normal | -1728
protein C levels normal | -1728
intubation | 24
respiratory failure | 24
dual vasopressors | 24
norepinephrine | 24
vasopressin | 24
continuous renal replacement therapy | 24
COVID-19 acute respiratory distress syndrome | 24
prone-positioning | 24
paralysis | 24
cytokine release syndrome | 48
interleukin-6 level | 48
D-dimer | 48
ferritin | 48
Lactate dehydrogenase | 48
Aspartate transaminase | 48
H-score | 48
tocilizumab | 48
hydrocortisone | 48
heparin infusion | 48
lower gastrointestinal bleeding | 408
high-volume diarrhoea | 408
rectal tube insertion | 408
CT mesenteric angiogram | 408
embolisation | 408
bleeding | 432
repeated CTMA | 432
second embolisation | 432
colonoscopy | 480
endostasis | 480
right-sided hemicolectomy | 480
segmental resection of the terminal ileum | 480
extensive ulceration of the terminal ileum | 480
colitis of the caecum and ascending colon | 480
HIV screening negative | 480
Clostridium difficile testing negative | 480
tissue bacterial culture | 480
fungal cultures | 480
acid-fast smears negative | 480
molecular testing for tuberculosis negative | 480
serology for cytomegalovirus IgM negative | 480
blood PCR for cytomegalovirus negative | 480
histological analysis for viral inclusions negative | 480
stool PCR for SARS-CoV-2 negative | 480
swab taken per stoma negative for SARS-CoV-2 PCR | 480
discharged | 720