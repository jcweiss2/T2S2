69 years old | 0
male | 0
intractable esophageal dysmotility | -672
gastroesophageal reflux | -672
aspiration | -672
dysphagia | -672
distorted gastroesophageal anatomy | -672
distended intrathoracic post-Collis gastroplasty gastric segment | -672
failed fundoplication | -672
endoscopic esophageal dilations | -672
temporary relief of dysphagia | -672
Ivor Lewis esophagectomy | 0
upper midline abdominal incision | 0
right posterolateral thoracotomy | 0
anastomotic leak | 48
mediastinitis | 48
sepsis | 48
return to operating theatre | 48
intensive care unit | 48
complicated recovery | 48
discharged from hospital | 1290
swelling over the right costal margin | 2628
erythema over the right costal margin | 2628
pain over the right costal margin | 2628
costal osteomyelitis | 2628
noncontrast CT | 2628
clindamycin | 2628
no change in symptoms | 3108
surgical intervention | 3150
magnetic resonance imaging (MRI) | 3150
enhancing collection overlying the sixth rib | 3150
phlegmonous changes | 3150
oblique sinus tract | 3150
rib fracture | 3150
elective surgical debridement | 3164
tissue samples | 3164
growth of C. albicans | 3164
discharged with treatment plan | 3170
oral clindamycin | 3170
surgical wound remained tender | 3190
swollen | 3190
warm | 3190
oral fluconazole | 3190
readmitted | 3200
intravenous fluconazole | 3200
clindamycin | 3200
skin breakdown | 3200
cellulitis | 3200
further debridement | 3210
resection of right anterior fifth and sixth ribs | 3210
good recovery | 3280
6-month course of oral fluconazole | 3280