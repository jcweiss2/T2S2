23 years old | 0
    acute lymphoblastic leukemia | 0
    normal karyotype pre-B | 0
    no molecular risk factors | 0
    second complete remission | 0
    FLAM protocol chemotherapy | 0
    fludarabine phosphate | 0
    cytarabine | 0
    mitoxantrone hydrochloride | 0
    first consolidation treatment | 0
    PALG ALL6 protocol | 0
    cyclophosphamide | 0
    cytarabine | 0
    pegaspargase | 0
    fever (39°C) | 48
    abdominal pain | 48
    diarrhea | 48
    piperacillin/tazobactam | 48
    fluconazole | 48
    nifuroxazide | 48
    temperature returned to normal | 72
    symptoms receded | 96
    condition improved | 96
    fever (38°C) | 192
    abdominal pain | 192
    diarrhea | 192
    decrease in blood count parameters | 192
    granulocytopenia | 192
    WBC 0.1–0.0 G/l | 192
    excluded bacteria in peripheral blood | 192
    excluded neutropenic enterocolitis | 192
    excluded pseudomembranous enteritis | 192
    no Clostridium difficile in feces | 192
    medical therapy modified | 192
    meropenem | 192
    metronidazole | 192
    itraconazole | 192
    granulocyte-colony stimulating factors | 192
    filgrastim | 192
    temperature returned to normal | 336
    abdominal pain subsided | 336
    nifuroxazide continued | 336
    G-CSF continued | 336
    agranulocytosis | 336
    four asymptomatic days | 432
    delayed second cycle of chemotherapy introduced | 432
    fever (39°C) | 468
    abdominal pain | 468
    diarrhea | 468
    Candida albicans in feces culture | 468
    metronidazole supplemented | 468
    ketoconazole | 468
    piperacillin/tazobactam | 468
    vancomycin | 468
    granulocyte-colony stimulating factors | 468
    agranulocytosis | 468
    Enterobacter cloacae detected | 468
    improvement of general condition | 468
    reduction of abdominal pain | 468
    fever | 552
    vomiting | 552
    acute pain in right epigastrium | 552
    acalculous gallbladder | 552
    overdistention | 552
    wall thickening (14 mm) | 552
    pericholecystic fluid | 552
    acalculous cholecystitis | 552
    medical therapy continued | 552
    broad spectrum antibiotic regimen | 552
    G-CSF | 552
    intravenous fluids | 552
    fasting | 552
    condition deteriorated | 576
    renal failure | 576
    liver failure | 576
    qualified for life-saving surgery | 576
    laparoscopic cholecystectomy | 576
    platelet concentrate transfused | 576
    platelet count increased to 43 G/l | 576
    lymphocyte infiltration of gallbladder mucous membrane | 576
    hyperemia | 576
    no neutrophil infiltrations | 576
    no leukemia cells (TdT–, CD34–) | 576
    no bacteria | 576
    no fungal cells | 576
    bile culture showed no micro-organisms | 576
    moved to intensive care ward | 576
    broad spectrum antibiotic regimen | 576
    G-CSF | 576
    erythrocyte concentrate transfusions | 576
    PC transfusions | 576
    fever (38°C) | 624
    lower values of peripheral blood pressure | 624
    chest X-ray demonstrated atelectatic-inflammatory changes | 624
    parenchymatous-interstitial changes | 624
    intensive respiratory rehabilitation | 624
    imipenem/cilastatin sodium | 624
    vancomycin | 624
    metronidazole | 624
    teicoplanin | 624
    ketoconazole | 624
    supplemented with ciprofloxacin hydrochloride | 624
    co-trimoxazole | 624
    patient's condition improved | 624
    no abdominal symptoms related to cholecystectomy | 672
    no abdominal pain | 672
    no diarrhea | 672
    permitted to eat | 744
    light diet well tolerated | 744
    marked improvement in peripheral blood | 816
    G-CSF discontinued | 864
    antibiotic therapy discontinued | 912
    transferred to Department of Hematology | 912
    discharged from hospital | 960
    good general condition | 960

    23 years old | 0
    acute lymphoblastic leukemia | 0
    normal karyotype pre-B | 0
    no molecular risk factors | 0
    second complete remission | 0
    FLAM protocol chemotherapy | 0
    fludarabine phosphate | 0
    cytarabine | 0
    mitoxantrone hydrochloride | 0
    first consolidation treatment | 0
    PALG ALL6 protocol | 0
    cyclophosphamide | 0
    cytarabine | 0
    pegaspargase | 0
    fever (39°C) | 48
    abdominal pain | 48
    diarrhea | 48
    piperacillin/tazobactam | 48
    fluconazole | 48
    nifuroxazide | 48
    temperature returned to normal | 72
    symptoms receded | 96
    condition improved | 96
    fever (38°C) | 192
    abdominal pain | 192
    diarrhea | 192
    decrease in blood count parameters | 192
    granulocytopenia | 192
    WBC 0.1–0.0 G/l | 192
    excluded bacteria in peripheral blood | 192
    excluded neutropenic enterocolitis | 192
    excluded pseudomembranous enteritis | 192
    no Clostridium difficile in feces | 192
    medical therapy modified | 192
    meropenem | 192
    metronidazole | 192
    itraconazole | 192
    granulocyte-colony stimulating factors | 192
    filgrastim | 192
    temperature returned to normal | 336
    abdominal pain subsided | 336
    nifuroxazide continued | 336
    G-CSF continued | 336
    agranulocytosis | 336
    four asymptomatic days | 432
    delayed second cycle of chemotherapy introduced | 432
    fever (39°C) | 468
    abdominal pain | 468
    diarrhea | 468
    Candida albicans in feces culture | 468
    metronidazole supplemented | 468
    ketoconazole | 468
    piperacillin/tazobactam | 468
    vancomycin | 468
    granulocyte-colony stimulating factors | 468
    agranulocytosis | 468
    Enterobacter cloacae detected | 468
    improvement of general condition | 468
    reduction of abdominal pain | 468
    fever | 552
    vomiting | 552
    acute pain in right epigastrium | 552
    acalculous gallbladder | 552
    overdistention | 552
    wall thickening (14 mm) | 552
    pericholecystic fluid | 552
    acalculous cholecystitis | 552
    medical therapy continued | 552
    broad spectrum antibiotic regimen | 552
    G-CSF | 552
    intravenous fluids | 552
    fasting | 552
    condition deteriorated | 576
    renal failure | 576
    liver failure | 576
    qualified for life-saving surgery | 576
    laparoscopic cholecystectomy | 576
    platelet concentrate transfused | 576
    platelet count increased to 43 G/l | 576
    lymphocyte infiltration of gallbladder mucous membrane | 576
    hyperemia | 576
    no neutrophil infiltrations | 576
    no leukemia cells (TdT–, CD34–) | 576
    no bacteria | 576
    no fungal cells | 576
    bile culture showed no micro-organisms | 576
    moved to intensive care ward | 576
    broad spectrum antibiotic regimen | 576
    G-CSF | 576
    erythrocyte concentrate transfusions | 576
    PC transfusions | 576
    fever (38°C) | 624
    lower values of peripheral blood pressure | 624
    chest X-ray demonstrated atelectatic-inflammatory changes | 624
    parenchymatous-interstitial changes | 624
    intensive respiratory rehabilitation | 624
    imipenem/cilastatin sodium | 624
    vancomycin | 624
    metronidazole | 624
    teicoplanin | 624
    ketoconazole | 624
    supplemented with ciprofloxacin hydrochloride | 624
    co-trimoxazole | 624
    patient's condition improved | 624
    no abdominal symptoms related to cholecystectomy | 672
    no abdominal pain | 672
    no diarrhea | 672
    permitted to eat | 744
    light diet well tolerated | 744
    marked improvement in peripheral blood | 816
    G-CSF discontinued | 864
    antibiotic therapy discontinued | 912
    transferred to Department of Hematology | 912
    discharged from hospital | 960
    good general condition | 960