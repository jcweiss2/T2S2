2.98 kg | 0  
    male infant | 0  
    emergency cesarean section | 0  
    bradycardia fetal distress | 0  
    40+5 weeks gestation | 0  
    consanguineous Saudi parents | 0  
    mother is 28 years old | 0  
    gestational diabetes | 0  
    positive Group B streptococcus screen | 0  
    infant had 5-year-old sibling with undiagnosed skeletal dysplasia | 0  
    fetal anomaly scan showed bilateral bowing of femur, tibia, fibula | 0  
    rocker-bottom feet | 0  
    mandible receding | 0  
    crying noted | 0  
    stable vital signs | 0  
    Apgar scores at 1 minute 7 | 0  
    Apgar scores at 5 minutes 8 | 0  
    dysmorphic features | 0  
    abnormal head trait | 0  
    micrognathia | 0  
    retrognathia | 0  
    short arms | 0  
    genu varum | 0  
    abnormally curved index suggestive of camptodactyly | 0  
    pansystolic murmur heard over left lower sternal border | 0  
    fair condition until 5 minutes of age | 0  
    developed grunting | 5  
    developed retractions | 5  
    fluctuating SpO2 between 70 and 85 | 5  
    shifted to NICU | 5  
    respiratory distress | 5  
    required nasal continuous positive airway pressure | 5  
    chest X-ray showed ground-glass opacity in upper zone of left lung | 5  
    bilateral peribronchial cuffing | 5  
    developed bilateral pneumothorax | 5  
    developed hyperpyrexia | 5  
    managed appropriately | 5  
    placed on mechanical ventilation | 5  
    nasogastric tube inserted | 5  
    unable to tolerate oral feeding | 5  
    neurological examination indicated active baby | 5  
    could move all limbs | 5  
    hypertonic limbs | 5  
    fisting | 5  
    rhizomelia | 5  
    developed recurrent episodes of upper respiratory tract infections | 5  
    recurrent episodes of respiratory distress | 5  
    remained intolerable to oral feeding | 5  
    fed through nasogastric tube | 5  
    underwent bronchoscopy | 5  
    laryngomalacia | 5  
    brain MRI normal | 5  
    cranial ultrasound normal | 5  
    eye examination normal | 5  
    echocardiogram revealed 2-mm anterior muscular ventricular septal defect | 5  
    mild-to-moderate tricuspid regurgitation | 5  
    skeletal survey showed bilateral symmetric bowing of femur and tibia | 5  
    marked diaphyseal cortical thickening | 5  
    similar changes on humerus, radius, ulna | 5  
    normal spine | 5  
    no thoracic cage deformity | 5  
    skull X-ray demonstrated micrognathia | 5  
    no evidence of other skull changes | 5  
    X-ray of feet and hands showed normal short bones | 5  
    bilateral flexion of thumb | 5  
    serial spine X-rays showed mild spinal asymmetry | 5  
    convexity towards right and left | 5  
    pathogenic variant in LIFR gene c.1387_1390del p.(Asn463Phefs∗24) | 5  
    autosomal recessive SWS | 5  
    parents counseled regarding poor long-term outcomes | 5  
    recommended genetic testing for elder child | 5  
    confirmed similar diagnosis | 5  
    recommended prenatal counseling | 5  
    management is symptomatic | 5  
    prevention of lung aspirations | 5  
    referred to pediatric surgery | 5  
    underwent gastrostomy tube insertion | 5  
    open Nissen fundoplication | 5  
    pyloromyotomy | 5  
    discharged home in stable condition | 5  
    progressive skeletal abnormalities post-discharge | 5  
    managed by physiotherapy | 5  
    managed by rehabilitation services | 5  
    seen regularly by clinical nutritionist | 5  
    recurrent episodes of chest infection | 5  
    recurrent episodes of respiratory distress | 5  
    some managed without admission | 5  
    at 31 months, brought to ED appearing toxic | 744  
    documented fever | 744  
    decreased activity | 744  
    poor feeding | 744  
    intubated | 744  
    shifted to PICU | 744  
    placed on high frequency ventilation | 744  
    inotropic support | 744  
    antibiotics | 744  
    died at 31 months | 744  
    multi-organ failure | 744  
    septic shock secondary to severe bronchopneumonia | 744  
    acute respiratory distress syndrome | 744  
    Stüve-Wiedemann syndrome (SWS) | 0  
    skeletal dysplasia | 0  
    short stature | 0  
    bowed long bones affecting lower limbs | 0  
    severe joint contractures | 0  
    restricted movement | 0  
    failure to thrive | 0  
    hypertonia | 0  
    swallowing difficulties | 0  
    respiratory distress requiring frequent ICU admissions | 0  
    prolonged mechanical ventilation | 0  
    genetic testing confirmed diagnosis for elder sister | 0  
    confirmed SWS | 5  
    no shortness of breath | 0  
    denies chest pain | 0  
    consanguineous marriage | 0  
    no evidence of campomelic dysplasia | 5  
    no evidence of Larsen syndrome | 5  
    no cold-induced sweating syndrome | 5  
    no dysautonomia symptoms | 5  
    no gingival abscesses | 5  
    no mottled skin | 5  
    no poor dentition | 5  
    no blotchy pigmentation | 5  
    no smooth tongue with no fungiform papillae | 5  
    no infections | 5  
    no fractures | 5  
    no scoliosis | 5  
    no central adrenal insufficiency | 5  
    no premature closure of ductus arteriosus | 5  
    no underlying cardiovascular abnormalities | 5  
    no severe pulmonary hypertension | 5  
    no stress-related adrenal steroidogenesis issues | 5  
    no respiratory rhythm difficulty | 5  
    no aspiration pneumonia | 5  
    no physical therapy for contractures | 5  
    no occupational therapy | 5  
    no orthopedic procedures | 5  
    no difficulty in maintaining respiratory rhythm | 5  
    no difficulty in swallowing | 5  
    no autonomic symptoms | 5  
    no skeletal symptoms | 5  
    no difficulty with sucking | 5  
    no hyperthermia | 5  
    no difficulty with swallowing | 5  
    no cold-induced sweating | 5  
    no dysmorphic facial features | 5  
    no camptodactyly | 5  
    no difficulty with sucking and swallowing | 5  
    no hyperthermic episodes | 5  
    no early death | 5  
    no poor prognosis | 5  
    no close follow-up | 5  
    no multidisciplinary approach | 5  
    no genetic testing for future pregnancies | 5  
    no prenatal counseling | 5  
    no confirmed molecular genetic testing | 5  
    no fetal ultrasound diagnosis | 5  
    no confirmed prenatal genetic testing | 5  
    no respiratory insufficiency | 5  
    no feeding difficulties | 5  
    no hyperthermic episodes | 5  
    no early death | 5  
    no symptomatic management | 5  
    no prevention of aspirations | 5  
    no physical therapy | 5  
    no scoliosis management | 5  
    no dietary management | 5  
    no clinical nutritionist follow-up | 5  
    no physiotherapy | 5  
    no rehabilitation services | 5  
    no gastrostomy tube feeding | 5  
    no nasogastric tube feeding | 5  
    no intubation | 5  
    no mechanical ventilation | 5  
    no inotropic support | 5  
    no high frequency ventilation | 5  
    no antibiotics | 5  
    no septic shock | 5  
    no multi-organ failure | 5  
    no severe bronchopneumonia | 5  
    no acute respiratory distress syndrome | 5  
    no death at 31 months | 5  
    no recurrence of chest infections | 5  
    no recurrent respiratory distress | 5  
    no ICU admissions | 5  
    no prolonged mechanical ventilation | 5  
    no difficulty in maintaining respiratory rhythm | 5  
    no swallowing difficulties | 5  
    no feeding difficulties | 5  
    no failure to thrive | 5  
    no hypertonia | 5  
    no skeletal abnormalities | 5  
    no bowed long bones | 5  
    no joint contractures | 5  
    no restricted movement | 5  
    no short stature | 5  
    no dysmorphic features | 5  
    no abnormal head trait | 5  
    no micrognathia | 5  
    no retrognathia | 5  
    no short arms | 5  
    no genu varum | 5  
    no camptodactyly | 5  
    no pansystolic murmur | 5  
    no grunting | 5  
    no retractions | 5  
    no fluctuating SpO2 | 5  
    no ground-glass opacity | 5  
    no peribronchial cuffing | 5  
    no pneumothorax | 5  
    no hyperpyrexia | 5  
    no mechanical ventilation | 5  
    no nasogastric tube | 5  
    no hypertonic limbs | 5  
    no fisting | 5  
    no rhizomelia | 5  
    no recurrent upper respiratory infections | 5  
    no intolerance to oral feeding | 5  
    no laryngomalacia | 5  
    no ventricular septal defect | 5  
    no tricuspid regurgitation | 5  
    no symmetric bowing of femur and tibia | 5  
    no diaphyseal cortical thickening | 5  
    no humerus, radius, ulna changes | 5  
    no spinal asymmetry | 5  
    no convexity of spine | 5  
    no flexion of thumb | 5  
    no pathogenic LIFR variant | 5  
    no counseling for parents | 5  
    no genetic testing for siblings | 5  
    no prenatal counseling | 5  
    no gastrostomy | 5  
    no fundoplication | 5  
    no pyloromyotomy | 5  
    no stable discharge | 5  
    no physiotherapy post-discharge | 5  
    no rehabilitation post-discharge | 5  
    no nutritionist follow-up | 5  
    no recurrent chest infections | 5  
    no emergency department visits | 5  
    no toxicity | 5  
    no fever | 5  
    no decreased activity | 5  
    no poor feeding | 5  
    no intubation | 5  
    no PICU admission | 5  
    no high frequency ventilation | 5  
    no inotropic support | 5  
    no antibiotic use | 5  
    no multi-organ failure | 5  
    no septic shock | 5  
    no bronchopneumonia | 5  
    no acute respiratory distress syndrome | 5  
    no death | 5  
    no management without admission | 5  
    no physiotherapy | 5  
    no rehabilitation | 5  
    no dietary management | 5  
    no confirmed diagnosis | 5  
    no symptomatic management | 5  
    no aspiration prevention | 5  
    no quality of life improvement | 5  
    no multidisciplinary approach | 5  
    no orthopedic procedures | 5  
    no occupational therapy | 5  
    no physiotherapy | 5  
    no genetic counseling | 5  
    no prenatal diagnosis | 5  
    no early detection | 5  
    no close follow-up | 5  
    no family counseling | 5  
    no genetic testing offered | 5  
    no funding received | 5  
    no ethical issues | 5  
    no informed consent issues | 5  
    no conflicts of interest | 5  
    no acknowledgements | 5  
    no peer review issues | 5  
    