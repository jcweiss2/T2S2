72 years old | 0
female | 0
admitted to the hospital (ventral hernia repair) | 0
bulging mass on low abdomen | -120
severe abdominal pain | -120
septic shock | -120
exploratory laparotomy | -120
extensive intestinal adhesions | -120
severe intraperitoneal contamination | -120
removal of mesh | -120
blunt dissection | -120
placement of three open drain systems | -120
postoperative EAF | -120
systemic infection | -120
two EAFs developed | -120
well-controlled hypertension | 0
well-controlled diabetes | 0
no intestinal obstruction | 0
no abnormalities on complete blood cell count | 0
no abnormalities on cardiac markers | 0
no abnormalities on coagulation profile | 0
fasting with full caloric parenteral nutrition | 0
electrolyte repletion | 0
antacids | 0
octreotide | 0
frequent surgical wound dressing | 0
protection of surrounding tissue from enteric effluent | 0
EAF output > 1000 mL/d | 0
severe contamination by enteric effluent | 0
vacuum-assisted closure (VAC) dressings | 0
unable to initiate enteral nutrition | 0
rubber drains inserted into intestinal lumens | 0
fistula output < 500 mL/d | 0
fistula output returned to > 1000 mL/d with EN attempt | 0
insufficient rubber drain diameter | 0
attempted endoscopic stent insertion | 0
expulsion of stents | 0
implanted two vascular grafts | 792
anastomoses between intestinal openings and vascular grafts | 792
no fistula output post-operation | 792
elemental EN initiated on 5th POD | 792
leakage after EN initiation | 792
output < 300 mL/d | 792
patient comfortable clinically and emotionally | 792
discharged on 16th POD after graft implantation | 864
VAC dressing management | 864
EAF resection two months after discharge | 2928
involved distal jejunum | 2928
involved sigmoid colon | 2928
