39 years old | 0
female | 0
palpable mass on right breast | -168
Hodgkin lymphoma | -6336
chemotherapy | -6336
mantle field radiation | -6336
inflammatory colitis | -6336
mesalazine | -336
breast cancer | 0
invasive ductal carcinoma | 0
triple-negative phenotype | 0
MIB1 85% | 0
staging CT scan | 0
neoadjuvant chemotherapy | 0
paclitaxel | 0
carboplatin | 0
port-à-cath insertion | 48
subcutaneous cellulitis | 96
colliquative necrosis | 96
fever | 96
elevated white blood cell count | 96
neutrophilia | 96
elevated C-reactive protein | 96
broad-spectrum i.v. antibiotic therapy | 96
piperacillin/tazobactam | 96
daptomycin | 96
PORT rimotion | 96
necrosectomy | 96
defervescence | 120
improvement in subcutaneous cellulitis | 120
improvement in blood works | 120
febrile seizure | 144
WBC rise | 144
worsening of skin lesion | 144
second necrosectomy | 144
peripheral blood cultures | 144
skin plug | 144
i.v. catheter tip positivity for Klebsiella pneumoniae | 144
antibiotic therapy modification | 144
meropenem | 144
levofloxacin | 144
chest/abdomen CT scan | 144
mediastinitis | 144
bilateral pleural effusion | 144
left pulmonary atelectasis | 144
thoracoscopy | 144
pleural and mediastinal drainage | 144
sepsis | 144
broad-spectrum antibiotic and antifungal therapy | 144
hemodynamic support | 144
non-invasive ventilation | 144
intensive inflammatory infiltrate | 144
neutrophils | 144
PG diagnosis | 144
systemic methylprednisolone | 144
topical cyclosporine | 144
seriate chest X-ray | 168
progressive resolution of mediastinitis | 168
progressive resolution of pleural effusion | 168
wound improvement | 168
scar | 168
progressive normalization of blood count | 168
progressive normalization of flogosis index | 168
breast ultrasound | 240
no change in the dimension of the lump | 240
multidisciplinary meeting | 240
right mastectomy | 240
axillary dissection | 240
breast surgical wound healing | 240
fibroelastosis | 240
chronic inflammation | 240
isolated neoplastic cells | 240
negative axillary nodes | 240
restaging brain/chest/abdomen CT | 240
negative for distant metastasis | 240
BRCA and p53 mutation tests | 240
negative | 240
autologous skin graft | 432
no further complications | 432
PICC implant | 432
chemotherapy with carboplatin and paclitaxel | 432
dose reduction | 432
good tolerance | 720
follow-up | 720