80 years old | 0
female | 0
Caucasian | 0
admitted to the hospital | 0
arterial hypertension | -8760
dyslipidemia | -8760
type 2 diabetes mellitus | -8760
ischemic cardiomyopathy | -8760
preserved ejection fraction | -8760
chronic hepatitis B virus infection | -8760
progressive fatigue | -216
malaise | -216
anorexia | -216
cough with blood-streaked sputum | -840
peripheral edema | -840
denied fever | -840
denied weight loss | -840
denied arthralgia | -840
denied skin rash | -840
multifocal pneumonia | -48
acute kidney injury | -48
iron deficiency anemia | -48
serum creatinine 5.69 mg/dL | -48
hemoglobin 7.6 g/dL | -48
IV fluid administration | -48
amoxicillin-clavulanate | -48
azithromycin | -48
piperacillin-tazobactam | -24
elevated erythrocyte sedimentation rate | -24
negative ANCA | -24
negative anti-GBM antibodies | -24
negative antistreptolysin O antibodies | -24
normal C3 and C4 levels | -24
microscopic hematuria | -24
subnephrotic proteinuria | -24
bilateral nodular infiltrates | -24
hemoptysis | -24
bronchoscopy | -24
bronchoalveolar lavage | -24
alveolar macrophages | -24
polymorphonuclear cells | -24
hemosiderin-laden macrophages not identified | -24
renal replacement therapy | 0
pale | 0
afebrile | 0
blood pressure 130/70 mm Hg | 0
pulse rate 87 beats/min | 0
tachypneic | 0
oxygen saturation 94% | 0
fine crackles | 0
peripheral edema | 0
no rash | 0
MPO-ANCA 121.1 U/mL | 48
PR3-ANCA 312.6 U/mL | 48
anti-GBM antibody 202 U | 48
rheumatoid factor 26 IU/mL | 48
normal C3 and C4 levels | 48
negative antinuclear antibody | 48
negative cryoglobulins | 48
negative anti-dsDNA | 48
IV high-dose methylprednisolone | 48
oral prednisolone | 48
pulses of IV cyclophosphamide | 48
plasma exchange | 48
entecavir 0.5 mg weekly | 48
renal biopsy | 144
cellular crescents | 144
focal fibrinoid necrosis | 144
mildly interstitial fibrosis | 144
moderate inflammatory infiltrate | 144
no vasculitis | 144
linear deposition of immunoglobulin G | 144
along the GBM | 144
progressive improvement | 168
resolution of hypoxemia | 168
no recurrence of cough | 168
no recurrence of blood-streaked sputum | 168
renal function did not improve | 168
chest CT scan | 240
resolution of pulmonary infiltrates | 240
discharged | 816
oral glucocorticoid therapy gradually reduced | 816
HBV viral load undetectable | 4320
abdominal ultrasound | 4320
normal liver morphology | 4320
liver stiffness value compatible with F0-F1 | 4320
dialysis-dependent | 8760
no relapse of DAH | 8760
ANCA and anti-GBM antibody titers remain negative | 8760