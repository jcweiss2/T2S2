25 years old | 0
    male | 0
    admitted to the hospital | 0
    high-grade fever | -144
    diffuse abdominal pain | -48
    hematemesis | -48
    anemia | 0
    thrombocytopenia | 0
    hyperbilirubinemia | 0
    raised transaminases | 0
    normal coagulation profile | 0
    normal renal function | 0
    hemoglobin 10 g/dl | 0
    total leukocyte count 5300/cumm | 0
    platelet count 15,000/cumm | 0
    serum creatinine 1.0 mg/dl |
### 8 Ways to Get More Sleep

If you want to live a long and healthy life, you need to make sure you get enough sleep. The problem is that most people don't get nearly enough. According to a recent poll, 1 in 3 Americans aren't getting the recommended 7 to 9 hours of sleep each night. That's not good for your physical or mental health. Here's how to fix that. 1. Stop using electronics before bed. The blue light from your devices messes with your circadian rhythms and makes it harder to fall asleep. So put down the phone or tablet at least an hour before bedtime. 2. Go to bed and wake up at the same time each day. If you can establish a regular sleep schedule, your body will start to adapt and make it easier to fall asleep each night. 3. Avoid caffeine and other stimulants before bed. They can stay in your system for hours, so avoid them in the afternoon. 4. Make sure your bedroom is dark, quiet, and cool. These conditions are optimal for sleeping. 5. Exercise regularly. Physical activity helps you sleep better, but don't do it too close to bedtime. 6. Wind down before bed. Read a book or take a bath to relax. 7. Don't eat a heavy meal before bed. Your body needs time to digest, so eat at least a few hours before bedtime. 8. See a doctor if you have persistent sleep problems. Insomnia can be a sign of other health issues. The bottom line is that sleep is essential for good health. If you're not getting enough, take steps to improve your sleep habits today. Your body and mind will thank you.