70 years old | 0
male | 0
admitted to the hospital | 0
complaint of persistent cough | -72
cough lasted for three months | -72
taking statin | -8760
taking anti-hypertensive drugs | -8760
stable vital signs | 0
no significant physical examination findings | 0
chest computed tomographic (CT) scan | 0
positron emission tomography (PET) | 0
malignant lung mass in the left lower lobe (LLL) | 0
multiple mediastinal lymph nodes | 0
bone metastases | 0
cancer at stage IV | 0
bronchoscopy | 0
irregular mucosal changes | 0
protruding mass at the orifice of the LLL | 0
invasive mucinous lung adenocarcinoma | 0
positive for thyroid transcription factor 1 (TTF-1) | 0
routine mutation profiling | 0
epidermal growth factor receptor mutations | 0
anaplastic lymphoma kinase (ALK) or ROS proto-oncogene 1 (ROS1) fusions | 0
PD-L1 tumor proportion score (TPS) 100% | 0
initiated first-line pembrolizumab monotherapy | 0
pembrolizumab 200 mg intravenously administered every three weeks | 0
first response evaluation | 24
slight increase in the size of primary tumor mass | 24
slight increase in the mediastinal lymph nodes | 24
continued with an additional two cycles of treatment | 48
cough difficult to control | 48
use of antitussives | 48
use of inhaled bronchodilators | 48
use of systemic corticosteroids | 48
follow-up chest CT and PET scans | 96
marked enlargement of both the primary lung tumor | 96
marked enlargement of the mediastinal lymph nodes | 96
newly developed bone metastases | 96
carcinoembryonic antigen level elevated | 96
discontinued frontline treatment | 96
switched to cytotoxic chemotherapy | 96
pemetrexed and carboplatin | 96
next-generation sequencing (NGS) | 96
KRAS (p.G12V) mutation | 96
TP53 (p.E286K) mutation | 96
STK11 (p.Y36fs*) mutation | 96
developed pneumonia | 120
elevated serum C-reactive protein | 120
elevated procalcitonin levels | 120
chest CT scan showed definite bronchial obstruction | 120
intensive care with broad-spectrum antibiotics | 120
mechanical ventilation | 120
pneumonia quickly progressed to sepsis | 144
patient succumbed | 144