60 years old | 0 | 0 
male | 0 | 0 
admitted to the hospital | 0 | 0 
fever | -48 | 0 
abdominal pain | -48 | 0 
edema of the scrotum | -48 | 0 
edema of the penis | -48 | 0 
edema of the perineum | -48 | 0 
edema of the right gluteal region | -48 | 0 
hypertension | 0 | 0 
osteoporosis | 0 | 0 
hemorrhoids | 0 | 0 
blood pressure 103/62 mmHg | 0 | 0 
heart rate 135/min | 0 | 0 
oxygen saturation 88% | 0 | 0 
white blood cell count 13.11/μL | 0 | 0 
C-reactive protein level 61.4 mg/dL | 0 | 0 
serum creatinine 4.3 mg/dL | 0 | 0 
blood urea 157 mg/dL | 0 | 0 
blood sugar 142 mg/dL | 0 | 0 
procalcitonin 8.53 ng/mL | 0 | 0 
CT of the abdomen and the pelvis | 0 | 0 
inflammatory infiltration of the subcutaneous tissues of the hypogastrium and the penis | 0 | 0 
liquefaction and presence of gas in the subcutaneous tissues of the scrotum, the perineum, and the right gluteal region | 0 | 0 
RT-PCR test for SARS-CoV-2 | 0 | 0 
negative RT-PCR test for SARS-CoV-2 | 0 | 0 
diagnosed with FG | 0 | 0 
qualified to undergo surgery | 0 | 0 
antibiotic therapy using meropenem | 0 | 432 
antibiotic therapy using metronidazole | 0 | 432 
antibiotic therapy using linezolid | 0 | 432 
resection of the necrotic tissues | 24 | 24 
bilateral orchiectomy | 24 | 24 
excision of the penile and scrotal skin | 24 | 24 
transferred to the ICU | 24 | 24 
mechanical ventilation | 24 | 552 
broad-spectrum antibiotics | 24 | 552 
supportive and nutritional therapies | 24 | 552 
colostomy | 48 | 48 
wound debridement | 48 | 552 
negative pressure wound therapy | 48 | 552 
sedation discontinued | 120 | 120 
recovered consciousness | 120 | 120 
extubated | 120 | 120 
able to breathe on his own with oxygen on low flow | 120 | 552 
hemodynamically stable | 120 | 552 
diuresis stimulated using a small dose of furosemide | 120 | 552 
inflammatory markers decreased significantly | 168 | 168 
culture of the pus material showed Escherichia coli and Pseudomonas aeruginosa | 168 | 168 
antibiotic therapy modified to include cephazolin | 168 | 576 
NPWT discontinued | 168 | 168 
transferred to the Department of Plastic Surgery | 240 | 240 
free-skin grafts applied to the debrided areas | 240 | 240 
discharged | 1104 | 1104 
received continous nursing care | 1104 | 1104 
free-skin graft care | 1104 | 1104 
regular dressing changes | 1104 | 1104 
testosterone supplementation | 1104 | 1104 
physiotherapy | 1104 | 1104 
follow-up in the urological and surgical clinic | 1104 | 1104 
colostomy reversal | 1104 | 1104 
wound closure | 1104 | 1104 
application of the free-skin graft to the right gluteal area | 1104 | 1104