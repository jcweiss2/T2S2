58 years old | 0
male | 0
admitted to the hospital | 0
fever | -168
fatigue | -168
cough | -168
shortness of breath | -168
oxygen saturation 70% | 0
intubated | 0
bilateral diffuse pulmonary infiltrates | 0
interstitial thickening | 0
bilateral basal consolidation | 0
COVID-19 positive | 0
pancytopenia | 0
WBC 2.6 × 10^3/μL | 0
ANC 1.8 × 10^3/μL | 0
Hgb 12.1 g/dL | 0
platelet count 85 × 10^3/μL | 0
acute kidney injury | 0
serum creatinine level 120 μmol/L | 0
transaminitis | 0
ALT 170.2 U/L | 0
AST 330 U/L | 0
LDH 857 U/L | 0
hydroxychloroquine 400 mg | 0
azithromycin 500 mg | 0
IL-6 1,843 pg/mL | 0
D-dimer 73.37 mg/L | 0
ferritin 2,166.0 μg/L | 0
tocilizumab 400 mg | 0
methylprednisone 40 mg | 0
IVIG 0.4 g/kg | 0
severe sepsis | 0
vasopressors | 0
broad-spectrum antibiotics | 0
antifungals | 0
SLED | 0
G-CSF | 0
persistent pancytopenia | 384
WBC 0.5 × 10^3/μL | 384
ANC 0.3 × 10^3/μL | 384
Hgb 8.4 g/dL | 384
platelet count 74 × 10^3/μL | 384
peripheral blood smear pancytopenia | 384
red cell agglutination | 384
atypical lymphoid cells | 384
hairy cells | 384
bone marrow examination | 384
BM aspirate hypocellular | 384
trilineage hematopoiesis decreased | 384
infiltrated with atypical lymphoid cells | 384
hairy cells | 384
BM core biopsy mildly hypercellular | 384
interstitial infiltration | 384
focal areas of diffuse extensive infiltration | 384
decreased erythropoiesis | 384
decreased granulopoiesis | 384
increased megakaryocytes | 384
hairy cells positive for CD20 | 384
hairy cells positive for DBA.44 | 384
hairy cells positive for PAX5 | 384
hairy cells positive for annexin A1 | 384
hairy cells positive for cyclin D1 | 384
hairy cells positive for CD25 | 384
V600E-mutant BRAF protein positive | 384
flow cytometry on BM aspirate | 384
monotypic B cells | 384
CD45 positive | 384
CD19 positive | 384
CD20 positive | 384
CD10 positive | 384
CD79b positive | 384
CD11c positive | 384
CD103 positive | 384
CD25 positive | 384
CD200 positive | 384
cBCL2 positive | 384
IgM positive | 384
lambda light chain restriction | 384
CD23 negative | 384
CD5 negative | 384
CD123 negative | 384
CD43 negative | 384
IgD negative | 384
FISH analysis normal | 384
cytogenetic analysis normal | 384
BRAF gene mutation analysis positive | 384
multidisciplinary team meeting | 384
decision to wait for full COVID-19 recovery | 384
discharged | 720