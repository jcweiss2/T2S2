47 years old | 0
male | 0
HCV-related cirrhosis | -672
hepatocarcinoma | -672
admitted to the hospital | -216
spontaneous bacterial peritonitis | -216
partial portal vein thrombosis | -216
liver transplantation | -72
antimicrobial prophylaxis | -72
tacrolimus | 0
mycofenolate mofetil | 0
prednisone | 0
discharged | 336
fever | 336
malaise | 336
moderate hepatic dysfunction | 336
readmitted | 336
magnetic resonance cholangiography | 336
biliary leak | 336
bilioma | 336
ascites | 336
vancomycin | 336
piperacillin/tazobactam | 336
fluconazole | 336
bilioma drained percutaneously | 336
bile sample sent to laboratory | 336
septic shock | 432
admitted to ICU | 432
mechanical ventilation | 432
inotropic support therapy | 432
new blood cultures | 432
tracheal aspirate | 432
linezolid | 432
meropenem | 432
tacrolimus withdrawal | 432
fluconazole stopped | 432
anidulafungin | 432
bilateral pneumonia | 432
surgical drainage of hepato-biliary ducts | 432
C. norvegensis isolated | 432
Enterococcus faecalis isolated | 432
identification and susceptibility assay | 432
MICs of fluconazole and voriconazole | 432
ESBL producing Klebsiella pneumoniae | 576
clinical conditions improved | 720
resolution of fever | 720
hemodynamic stability | 720
weaning from MV | 720
blood cultures negative | 720
bile cultures negative for C. norvegensis | 1008
trans-esophageal echocardiography | 1008
fundus oculi examination | 1008
linezolid stopped | 1008
meropenem continued | 1008
anidulafungin continued | 1008
bile tract repaired | 1008
tacrolimus re-started | 1008
discharged | 2160
asymptomatic during follow-up | 8760