46 years old | 0
female | 0
tracheotomy | -2160
pneumonia | -2160
intracerebral bleeding | -2160
hospitalized | -2160
transferred to rehabilitation center | -1440
massive hemorrhage | -1440
tracheal suction | -1440
cyanosis | -1440
respiratory failure | -1440
shocks | -1440
cuff air maximally expanded | -1440
bleeding did not stop | -1440
tube removed | -1440
suction consistently carried out | -1440
cuffed endotracheal intubation tried | -1440
attempt failure due to visual obstruction | -1440
cuffed endotracheal tube inserted | -1440
cuff expanded | -1440
tube moved up | -1440
bleeding stopped | -1440
transferred to intensive care center | -1440
blood test carried out | -1440
hemoglobin decreased from 10.9 g/dl to 8.9 g/dl | -1440
cervical CT carried out | -1440
no special abnormality identified | -1440
bronchoscopy did not show endotracheal area due to blood clot | -1440
complete examination not done due to risk of re-bleeding | -1440
conservative treatment continued | -1440
transfemoral angiography | -1320
innominate artery small luminal outpouching to trachea | -1320
diagnosis of TIAF | -1320
transferred to thoracic surgery unit | -1320
operation for TIAF | -1320
tracheoplasty with bypass graft | -1320
rupture area 1×0.5 cm observed | -1320
innominate artery rebuilt | -1320
artificial blood vessel connected right subclavian artery and right aorta | -1320
tracheoplasty done using fifth costal cartilage | -1320
tracheostenosis | -720
inflammation | -720
bronchoscopy carried out due to wheezing and tachypnea | -720
endotracheal balloon dilatation conducted | -720
no improvement in symptoms | -720
replacement of Montgomery T-tube | -720
rehabilitation continued | -720
transferred to rehabilitation center | -720
patient survives without further complications | -720
surgery carried out | -720
eleven months since surgery | -720
