45 years old | 0
    male | 0
    presented to the emergency department | 0
    upper abdominal pain | -72
    nausea | -72
    vomiting | -72
    tender to palpation | 0
    no muscle guarding | 0
    high-grade infection | 0
    no pneumoperitoneum | 0
    widespread thickening of the gastric wall | 0
    no signs of perforation | 0
    admitted | 0
    diffuse erythema | 0
    edema of the gastric wall | 0
    acute severe gastritis | 0
    gastric ischemia considered | 0
    malignancy considered | 0
    H2-blocker | 0
    cefuroxime | 0
    metronidazole | 0
    deteriorated into septic shock | 24
    multiple organ failure | 24
    high serum lactate | 24
    diagnostic laparoscopy | 24
    widespread irreversible gastric ischemia | 24
    laparotomy | 24
    total gastrectomy | 24
    no primary anastomosis | 24
    admitted to intensive care unit | 24
    hemodynamic support | 24
    continuous veno-venous hemofiltration | 24
    unstable condition | 24
    anastomoses conducted | 72
    Roux-Y esophagojejunostomy | 72
    suspicion of streptococcal toxic shock syndrome | 72
    multi-organ involvement | 72
    cultures confirmed | 72
    pathological examination confirmed | 72
    phlegmonous gastritis | 72
    group A Streptococcus | 72
    recovered | 336
    discharged | 336
    
    
    <|end_header_id|>