22 years old | 0
male | 0
admitted to intensive care unit | 0
high-grade fever | -72
hypoxic respiratory failure | 0
ventilatory support | 0
elevated white blood cell count | 0
elevated procalcitonin (PCT) | 0
elevated troponin | 0
myocarditis | 0
pneumonia |6 0
sepsis | 0
fever | -72
sore throat | -72
generalized weakness | -72
myalgia | -72
abdominal pain | -72
outpatient treatment | -72
no relief | -72
admitted to the floors | -72
tachycardia (heart rate: 118/min) | 0
febrile spikes (Tmax: 102.7°F) | 0
unremarkable systemic examination | 0
normal oral cavity examination | 0
no petechiae | 0
no muscle tenderness | 0
past history of rheumatic fever | -87600
penicillin prophylaxis | -87600
stopped penicillin prophylaxis | -76680
no history of heart ailments | 0
no recurrence of joint pains | 0
leukocytosis (20.3 × 10³) | 0
blood cultures sampled | 0
intravenous antibiotics started | 0
became tachypneic | 24
became tachycardic | 24
chest pain | 24
electrocardiogram showed global ST depression | 24
elevated troponin I | 24
intubated due to respiratory distress | 24
2D echo showed new onset global hypokinesia | 24
normal 2D echo at admission | 0
continued febrile spikes | 0
antimicrobials upgraded (suspecting pneumonia, sepsis, myocarditis) | 24
negative blood cultures | 24
negative throat swab for H1N1 | 24
negative diphtheria | 24
persistence of febrile spikes | 24
typical rise in evening fever | 24
upper abdominal pain | 24
tachycardia | 24
repeat 2D echo normalized | 168
troponin I decreased | 168
maintained hemodynamics | 0
contrast-enhanced CT chest and abdomen showed bilateral basal consolidation | 168
elevated baseline PCT level | 0
ruled out infective causes (Leptospira, dengue, malaria, HIV, HCV, HbsAg, scrub typhus, Brucella) | 168
negative ANA | 168
negative ANA profile | 168
negative rheumatoid arthritis | 168
negative C-ANCA | 168
negative P-ANCA | 168
negative antistreptolysin O titers | 168
transesophageal echocardiography negative for infective endocarditis | 168
antibiotics upgraded to colistin | 168
Acinetobacter isolated from bronchoalveolar lavage cultures | 168
continued febrile spikes | 168
episodes of pulmonary edema | 168
elevated serial PCT levels | 168
failed extubation | 168
reintubated | 168
repeat CT chest consistent with prior findings | 168
negative septic PCR panel | 168
inconclusive bone marrow biopsy | 168
inconclusive bone marrow cultures | 168
elevated C-reactive protein | 168
elevated serum ferritin (>1200) | 168
initiated steroids | 168
initiated NSAIDs | 168
febrile spikes subsided | 168
PCT levels decreased after steroids | 168
extubated | 312
steroids tapered | 480
discharged | 480
Still's disease | 480
negative rheumatoid factor | 168
negative ANA (confirmatory) | 168
elevated IL-1, IL-6, IL-18, TNF, macrophage colony-stimulating factors | 480
NSAIDs treatment | 480
steroids treatment | 480
antirheumatic agents | 480
biologic agents (IL-1 inhibitors, IL-6 inhibitors, TNF inhibitors) | 480
plasma exchange | 480
intravenous immunoglobulins | 480
no shortness of breath | 0
denies chest pain (initial) | 0
