67 years old | 0
    male | 0
    presented to the emergency department | 0
    worsening dyspnea | -96
    irritating cough | -96
    expectoration of brownish sputum | -96
    general weakness | -96
    metabolic syndrome | 0
    diabetes | 0
    hyperlipidemia | 0
    intermittently uses PPI | 0
    subfebrile | 0
    complained of nausea | 0
    no vomiting | 0
    negated diarrhea | 0
    negated chest pain | 0
    no loss of taste | 0
    no loss of smell | 0
    blood saturation 92% O2 without oxygen | 0
    borderline blood pressure 115/60 mm Hg | 0
    mild tachycardia around 100 rpm | 0
    rapid test positive for COVID-19 | 0
    PCR test confirmed COVID-19 | 0
    chest X-ray showed bilateral pneumonia | 0
    elevation of CRP 168.9 mg/L | 0
    leukocytes 4.0 10^9/L | 0
    PCT 7.13 μg/L | 0
    Hb 143 g/L | 0
    thr 272 10^9/L | 0
    INR 0.93 | 0
    decompensated diabetes mellitus (glycemia 18.9 mmol/L) | 0
    normal renal function | 0
    normal liver function | 0
    acutely admitted to COVID-19 ward | 0
    barrier regime treatment | 0
    antibiotic therapy started | 0
    corticoids added | 0
    bronchodilators added | 0
    LMWH added | 0
    diabetic medication adjusted | 0
    shortness of breath | 0
    irritating cough | 0
    desaturation up to 76% O2 | 0
    transfer to intensive care unit | 0
    deep venous thrombosis excluded | 0
    pulmonary embolism excluded | 0
    HFNO therapy introduced | 0
    corticoids continued | 0
    antibiotics continued | 0
    LMWH dose increased | 0
    progression on day 6 | 144
    severe hypoxemia | 144
    transfer to anesthesiology and resuscitation department | 144
    intubation | 144
    tracheostomy | 144
    escalation of ATB | 144
    nutrition via nasogastric tube | 144
    circulatory support with vasopressors | 144
    condition improved | 144
    catecholamines withdrawn | 144
    febrile episodes subsided | 144
    inflammatory markers decreased | 144
    sedatives discontinued | 144
    regained consciousness | 144
    low muscle strength | 144
    noninfectious from day 21 | 504
    transfer to rehabilitation care planned | 504
    sudden rapid deterioration on day 23 | 552
    circulatory instability | 552
    tachypnea | 552
    fibrillation | 552
    massive enterorrhagia | 552
    hemoglobin drop to 81 g/L | 552
    septic shock | 552
    intubation | 552
    circulatory resuscitation | 552
    catecholamines up to 40 mL/h | 552
    multiple blood substitutes | 552
    hemostatic therapy started | 552
    LMWH discontinued | 552
    abdominal ultrasound performed | 552
    undilated small-bowel loops | 552
    meteoric colon | 552
    borderline width 6–7 cm | 552
    no obvious wall thickening | 552
    no free fluid in abdominal cavity | 552
    gastrofibroscopy performed | 552
    colonoscopy performed | 552
    normal mucosa from esophagus to D2 part of duodenum | 552
    no signs of bleeding | 552
    colonoscopy to hepatic flexure | 552
    clarity of colon wall aggravated | 552
    presence of intestinal contents with coagula | 552
    no source of bleeding | 552
    no mural lesion | 552
    CT angiography of abdomen | 552
    liquid content in cecum | 552
    suspected coagulum in sigmoid colon and ampulla recti | 552
    cecum distended to 80 mm | 552
    sigmoideum distended to 60 mm | 552
    no wall thickening | 552
    no clear source of bleeding | 552
    acute abdominal revision | 552
    midline laparotomy | 552
    free of effusion | 552
    distended colon | 552
    cecum with hemorrhagic filling | 552
    small bowel free of blood | 552
    desufflation of cecum over appendix stump | 552
    hemorrhagic filling verified | 552
    revision of small intestine | 552
    enterotomy in terminal ileum | 552
    filled with enteral contents only | 552
    no signs of bleeding | 552
    right-sided hemicolectomy | 552
    ileotransversoanastomosis | 552
    histological examination revealed ischemic enteritis | 552
    ischemic colitis | 552
    mucosal ulcerations | 552
    no evidence of infectious inflammation | 552
    no IBD inflammation | 552
    no Dieulafoy lesion | 552
    no dysplasia | 552
    no malignancy | 552
    postoperative stabilization | 552
    weaning without complications | 552
    adjustment of intestinal passage | 552
    enteral nutrition via nasogastric probe | 552
    hospitalized until day 42 | 1008
    transfer to post-acute intensive care unit | 1008
    readmitted for recurrent GIT bleeding | 1008
    colonoscopy showed small ulceration | 1008
    managed conservatively | 1008
    hemodynamic therapy | 1008
    transferred back to post-acute care | 1008
    no further signs of bleeding | 1008