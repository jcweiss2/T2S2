34 years old | 0
man | 0
primary refractory acute myeloblastic leukemia | -8760
multiple relapses | -8760
allogeneic bone marrow transplant from cord blood | -648
delayed engraftment | -648
prolonged severe neutropenia | -648
vancomycin-resistant Enterococcus bacteremia | -648
Streptococcus viridans bacteremia | -648
Streptococcus mitis bacteremia | -648
treated with tedizolid | -648
treated with cefepime | -648
treated with Flagyl | -648
treated with daptomycin | -648
acute abdominal pain | 0
filgrastim | 0
prophylaxis with acyclovir | 0
prophylaxis with Bactrim | 0
prophylaxis with caspofungin | 0
fever to 38.2°C | 0
tachycardia to 155 | 0
hypotension to 99/81 | 0
tachypnea to 36 | 0
ill appearing | 0
distended abdomen | 0
localized peritonitis | 0
white cell count 0.2 x 109 /L | 0
absolute neutrophil count (ANC) of zero | 0
anemia with hemoglobin 7 g/L | 0
thrombocytopenia with platelet count 10 x 109 /L | 0
lactic acid 3.1 mmol/L | 0
CT scan showing segmental ischemia of the small bowel | 0
exploratory laparotomy | 0
ischemic bowel segment identified | 0
small bowel resection | 0
primary anastomosis | 0
norepinephrine | 0
vasopressin | 0
admitted to intensive care unit | 0
pressors weaned | 24
extubated | 24
transferred to floor | 48
diet advanced | 72
passed flatus | 72
new fevers | 96
increased abdominal pain | 96
lactic acidosis | 96
respiratory decompensation | 96
neutropenic | 96
white cell count 0.1x 109 /L | 96
ANC 0 | 96
lactic acid 3.7 mmol/L | 96
amphotericin B (AmBisome) started | 96
repeat CT scan showing necrotic small bowel | 96
invasive fungal forms in omental specimen | 96
invasive fungal forms in small intestinal resection specimen | 96
angioinvasion | 96
hemorrhage | 96
transmural ischemic necrosis | 96
mucormycosis diagnosis | 96
amphotericin B added | 96
discussion with family and oncology team | 96
decision for comfort measures | 96
patient died | 120
white cell count 0.2 x 109 /L |
