69 years old | 0
male | 0
hypertension | 0
CKD stage 5 | 0
hemodialysis | 0
consumed 6 bilimbi fruits | -48
uncontrollable hiccups | -45
malaise | -45
abdominal discomfort | -45
two episodes of macroscopic hematuria | -45
nausea | -24
vomiting | -24
hiccups persisted | -24
abdominal discomfort persisted | -24
significant asthenia | 0
decreased level of consciousness | 0
dysarthria | 0
myoclonus of the upper limbs | 0
generalized tonic-clonic seizures | 0
subsequent seizures | 0
transferred to a referral emergency service | 0
refractory seizures | 0
mechanical ventilation | 0
orotracheal intubation | 0
sedation | 0
Richmond Agitation Sedation Scale score -3 | 0
hemodynamically stable | 0
blood pressure 110/60 mm Hg | 0
heart rate 68 bpm | 0
diffuse ecchymoses | 0
hemoglobin 13.1 g/dL | 0
hematocrit 39.3% | 0
white blood cells 13,600/mL | 0
band form count 3% | 0
platelets 179,000/mL | 0
urea 86.8 mg/dL | 0
serum creatinine 7.11 mg/dL | 0
serum sodium 139 mEq/L | 0
serum potassium 3.93 mEq/L | 0
computed tomography head hypoattenuation | 0
lumbar puncture transparent cerebrospinal fluid | 0
red blood cells 22 | 0
normal glucose | 0
normal white blood cells | 0
normal proteins | 0
negative bacterial test | 0
negative China ink test | 0
negative fungi analysis | 0
negative acid-fast staining | 0
transferred to intensive care unit | 0
phenytoin | 0
midazolam | 0
SLEDD initiated | 0
SLEDD discontinued due to hypotension | 0
indwelling urinary catheter | 0
macroscopic hematuria | 0
hemodynamic worsening | 72
norepinephrine | 72
hemoglobin 12.5 g/dL | 72
hematocrit 38.8% | 72
white blood cells 16,700/mL | 72
band form count 8% | 72
platelets 180,000/mL | 72
CRP 320 mg/dL | 72
antibiotic therapy piperacillin-tazobactam | 72
septic shock | 72
ventilator-associated tracheobronchitis | 72
seizures persisted | 96
attempts to reduce sedatives | 96
further tests ordered | 96
SLEDD discontinued | 96
diagnostic hypothesis CNS vasculitis | 96
immunosuppression methylprednisolone | 96
negative rheumatic disease search | 96
EEG epileptogenic activity | 120
thiopental added | 120
family confirmed bilimbi consumption | 120
EEG confirmed epileptogenic activity | 192
decreased paroxysmal activity | 192
thiopental continued | 192
midazolam continued | 192
valproic acid continued | 192
intensify hemodialysis | 192
EEG improvement | 240
thiopental decreased | 240
midazolam decreased | 240
valproic acid increased | 240
increased norepinephrine | 288
fever 38.5°C | 288
white blood cells 21,500/mL | 288
band form count 9% | 288
CRP 107 mg/dL | 288
lactate 3.9 mmol/L | 288
diagnostic hypothesis septic shock | 288
antibiotics meropenem | 288
vancomycin | 288
gentamicin | 288
samples collected | 288
multidrug-resistant Klebsiella pneumoniae | 288
tigecycline started | 288
conscious | 336
responsive | 336
no sedatives | 336
decreasing norepinephrine | 336
persistent myoclonus lower limbs | 336
no new seizures | 336
SLEDD maintained | 336
worsening clinical status | 552
increased vasoactive drugs | 552
continued hemodialysis | 552
fever | 552
leukocytosis | 552
increased CRP | 552
death | 648
circulatory failure | 648
