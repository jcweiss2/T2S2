78 years old | 0
male | 0
West Virginia resident | 0
admitted to the hospital | 0
generalized weakness | -264
fever | -264
chills | -264
gout | 0
hypertension | 0
hypothyroidism | 0
chronic kidney disease stage 3 | 0
automobile mechanic | 0
outdoor gardener | 0
tick bite | -720
decreased appetite | -264
fever and chills | -264
inability to ambulate | -240
severe weakness | -240
febrile | 0
tachycardic | 0
tachypneic | 0
irregular rhythm | 0
palpable liver | 0
leukopenia | 0
thrombocytopenia | 0
acute kidney injury | 0
transaminitis | 0
viral hepatitis panel negative | 0
neutrophils with toxic changes | 0
computed tomographic scan | 0
bilateral perinephric stranding | 0
IV ceftriaxone | 0
oral doxycycline | 24
ferritin elevated | 0
inflammatory markers high | 0
bone marrow biopsy | 72
dexamethasone | 72
serum cytomegalovirus PCR negative | 72
Epstein-Barr virus quantitative positive | 72
blood culture positive | 72
gram-positive cocci | 72
IV ampicillin-sulbactam | 72
bone marrow biopsy results | 96
neutrophils with intracellular organisms | 96
hemophagocytosis | 96
peripheral smear | 96
intracellular organisms | 96
serum PCR positive for A phagocytophilum | 96
oral doxycycline | 0
oral amoxicillin-clavulanate | 0
discharged | 504
follow-up visit | 1008
symptoms improved | 1008
Facklamia ignava | 264
anaplasmosis | 0
hemophagocytic lymphohistiocytosis | 0