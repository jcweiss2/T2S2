septuagenarian man | 0
male | 0
admitted to the hospital | 0
medication-controlled hypertension | -72
malaise | -72
gait unsteadiness | -72
left arm weakness | -72
fever | -72
vomiting | -72
headache | -72
lethargic | 0
reactive pupils | 0
full extraocular movements | 0
intact corneal reflexes |0
CT brain unremarkable | 0
blood cultures unremarkable | 0
no prior ophthalmic records |0
loss of oculocephalic movements |24
small pupils |24
intact corneal reflexes |24
no ophthalmology consult |24
severe lethargy |48
left hemiplegia |48
right gaze preference |48
poor gag reflex |48
intubation |48
ICU admission |48
CT brain showing infarction |48
CSF neutrophilic pleocytosis |48
CSF cultures negative |48
blood cultures negative |48
empiric treatment |48
EEG with epileptiform discharges |48
Dilantin administration |48
MRI brain |48
CSF India ink negative |48
CSF fungal culture negative |48
serological studies |120
EEE IgM positive in serum |120
CSF IgM negative |120
other serology negatives |120
progressive decline in consciousness |48
loss of brainstem reflexes |72
left pneumothorax |72
gastrointestinal hemorrhage |72
bilateral pulmonary edema |72
recurrent fevers |48
septic shock |72
consultants' differential diagnosis |48
MRI findings consistent with meningoencephalitis |48
expired |168
