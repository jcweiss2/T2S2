58 years old | 0
female | 0
productive cough | -120
fatigue | -120
fever | -120
diarrhea | -120
diffuse rhonchi | 0
blood pressure 156/95 mm Hg | 0
heart rate 130 beats/min | 0
oxygen saturation 82% | 0
respiratory rate 24 breaths/min | 0
temperature 38.7°C | 0
lower lobe–predominant bilateral infiltrates | 0
intubated | 0
hypoxic respiratory failure | 0
acute respiratory distress syndrome | 0
sinus tachycardia | 0
1-mm upsloping ST-segment elevations | 0
mild diffuse PR interval depressions | 0
diffuse ST-T wave changes | 0
initial troponin I level negative | 0
leukopenia | 0
absolute lymphocyte count of 1.04 K/mm3 | 0
SARS-CoV-2 RNA detected | 0
diabetes mellitus type 2 | -6720
hypertension | -6720
dyslipidemia | -6720
denies travel | 0
father ill with similar symptoms | -120
ST-segment elevation myocardial infarction | 0
stress cardiomyopathy | 0
myopericarditis | 0
akinetic middle to distal anterior segments | 0
moderately hypokinetic middle and distal inferolateral segments | 0
hyperdynamic basal segments | 0
apical ballooning | 0
left ventricular ejection fraction 20% | 0
distal third or apical right ventricular free wall akinetic | 0
hyperdynamic RV basal wall motion | 0
RV function mildly reduced | 0
admitted to intensive care unit | 0
medical therapy for acute coronary syndrome | 0
dual antiplatelet therapy | 0
anticoagulation with continuous intravenous heparin | 0
hydroxychloroquine therapy | 0
azithromycin | 0
cardiogenic shock | 24
central venous oxygen saturation 42% | 24
dobutamine | 24
cardiogenic shock improved | 72
central venous oxygen saturation 65% | 72
de-escalating need for dobutamine | 72
repeat echocardiogram | 144
improvement in overall wall motion | 144
LV ejection fraction 55% | 144
stress cardiomyopathy | 144
ECG no evidence of Q-wave myocardial infarction | 144
acute respiratory distress syndrome | 168
venovenous extracorporeal membrane oxygenation | 168
ECG remains free of evidence of active ischemia or infarction | 168
urgent coronary evaluation not warranted | 168
precautions to limit unnecessary testing | 168
future coronary evaluation recommended | 168