68 years old | 0
female | 0
admitted to the emergency room | 0
altered level of consciousness | 0
blood pressure 80/60 mm Hg | 0
pulse rate 112 beats/min | 0
respiratory rate 24 breaths/min | 0
body temperature 34.9°C | 0
chronic kidney disease | -8760
type 2 diabetes mellitus | -8760
treated with insulin | -8760
admitted for acute pyelonephritis | -1096
admitted for acute pyelonephritis | -728
admitted for acute pyelonephritis | -84
resided in a nursing hospital | -84
non-smoker | 0
no previous history of pulmonary disease | 0
elevated white blood cell count | 0
low hemoglobin | 0
normal platelets | 0
elevated blood urea nitrogen level | 0
elevated serum creatinine level | 0
fluid resuscitation | 0
catecholaminergic therapy | 0
septic shock | 0
metabolic acidosis | 0
lactate 5.9 mmol/L | 0
blood pH 6.965 | 0
bicarbonate 5.5 mmol/L | 0
urine microscopy showed many WBCs | 0
urine dipstick test positive for nitrite | 0
transferred to a medical intensive care unit | 0
received continuous renal replacement therapy | 0
received antibiotics | 0
dyspnea | 408
chest X-ray examination showed atelectasis | 408
urine cultures showed Escherichia coli | 408
chest computed tomography scan | 408
partial atelectasis in the right upper lobe | 408
prominent wall thickening and enhancement in the proximal portion of the RUL bronchus | 408
bronchoscopy | 456
inflammation of the RUL bronchus | 456
necrosis | 456
acid fast bacilli stain negative | 456
Mycobacterium tuberculosis DNA detection negative | 456
culture for MTB negative | 456
bronchoscopic biopsy showed fungal infection | 456
fungal infection with necrosis | 456
yeast-like fungus with positive periodic acid-Schiff stain | 456
Candida albicans grew from the endobronchial aspirate | 456
treated with fluconazole | 456
electrolyte imbalance | 504
uremia worsened | 504
considered dialysis treatment | 504
rejected dialysis treatment | 504
signed a do-not-resuscitate order | 504
died | 672
endobronchial fungal infection diagnosed | 456
Candida albicans infection diagnosed | 456
atelectasis of the RUL diagnosed | 408
obstruction of the main bronchus diagnosed | 408
immune deficiency suspected | 0
poorly controlled diabetes | -84
decreased immune function | 0
repeated pyelonephritis | -1096
repeated pyelonephritis | -728
repeated pyelonephritis | -84
fungal infection suspected | 408
Candida species suspected | 408
Aspergillus infection suspected | 408
invasive procedures considered | 456
non-culture diagnostic tests considered | 456
antigen detection assays considered | 456
antibody detection assays considered | 456
β-D-glucan detection assays considered | 456
PCR considered | 456
interventional bronchoscopy considered | 456
endobronchial ultrasound-guided transbronchial needle aspiration considered | 456
bronchoscopy performed | 456
culture performed | 456
tissue obtained | 456
diagnosis made | 456
treatment started | 456
patient deteriorated | 504
patient died | 672