67 years old | 0
male | 0
admitted to the hospital | 0
fever | -336
cough | -336
shortness of breath | -336
renal transplant | -70080
end-stage renal disease | -70080
diabetic nephropathy | -70080
hypertension | -70080
diabetes mellitus | -70080
antihypertensive therapy | -70080
insulin use | -70080
immunosuppressive therapy | -70080
creatinine value 138 μmol/L | -1464
normal chest CT scan | -1464
mycophenolate mofetil | 0
tacrolimus | 0
prednisone | 0
dyspnea | 0
body temperature 38.0°C | 0
respiratory rate 28 breaths/minute | 0
oxygen saturation 98% on 3 L via nasal cannula | 0
blood pressure 134/71 mmHg | 0
heart rate 101 beats/minute |===
pulmonary moist rale | 0
pitting edema in lower extremities | 0
white blood cell count 8.2×10^9 cells/L | 0
hemoglobin level 114 g/L | 0
platelet count 187×10^9 cells/L | 0
potassium ion 6.59 mmol/L | 0
creatinine 193 μmol/L | 0
C reactive protein 199 g/L | 0
HIV negative | 0
pleural effusion | 0
bilateral airspace opacities | 0
severe pneumonia | 0
methylprednisolone | 0
imipenem/cilastatin | 0
trimethoprim-sulfamethoxazole | 0
continuous venovenous hemodialysis | 0
mechanical ventilation | 24
transferred to ICU | 72
respiratory failure | 72
heart failure | 72
chest CT scan showing discrete scattered patchy consolidation | 72
sputum culture | 72
blood culture | 72
Candida albicans growth in sputum | 72
negative blood cultures from Day 1 to Day 8 | 0
teicoplanin | 72
caspofungin | 72
sepsis | 240
multiple organ failure | 240
T. asahii growth in blood cultures | 216
T. asahii growth in sputum | 216
death | 240
amphotericin B MIC 0.5 mg/L | 240
itraconazole MIC 0.125 mg/L | 240
fluconazole MIC 1 mg/L | 240
voriconazole MIC 0.06 mg/L | 240
5-fluorocytosine MIC 4 mg/L | 240
