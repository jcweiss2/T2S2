pancreatic adenocarcinoma with metastasis to the liver | 0
diastolic heart failure | 0
atrial fibrillation | 0
coronary artery disease | 0
severe hyponatremia | 0
pneumonia | 0
broad-spectrum antibiotics | 0
jugular vein distention | 0
lower extremity pitting edema | 0
mildly reduced systolic function | 0
septal flattening | 0
left atrial enlargement | 0
suspected MV vegetation | 0
severe mitral regurgitation | 0
tricuspid regurgitation | 0
elevated RV systolic pressure | 0
type 2 and type 3 pulmonary arterial hypertension | 0
ill-defined thickening in the TV leaflets | 0
leukocytosis | 0
recent urethral instrumentation | 0
blood cultures | 0
infectious disease specialist consultation | 0
TEE | 24
normal left ventricular size and function | 24
ejection fraction of 60%-65% | 24
normal RV size and function | 24
hypermobile interatrial septum | 24
no left atrial or left atrial appendage thrombus | 24
vegetations on the atrial aspect of MV leaflets | 24
severe mitral regurgitation | 24
systolic flow reversal in the pulmonary vein | 24
vegetation on the TV leaflet | 24
tricuspid regurgitation | 24
RVSP 47 mm Hg | 24
negative blood cultures | 48
negative polymerase chain reaction testing | 48
unremarkable workup for antiphospholipid syndrome | 48
discontinuation of broad-spectrum antibiotics | 48
start of enoxaparin | 72
computed tomography imaging of the head | 72
death | 168