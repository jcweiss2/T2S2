63 years old | 0
female | 0
smoker | 0
chronic obstructive pulmonary disease | 0
admitted to the emergency department | 0
dyspnea | 0
dysphasia | 0
vaccinated with 3rd dose of BNT162b2mRNA | -360
reverse transcription SARS-CoV-2 PCR positive | -336
percutaneous transluminal angioplasty | -192
left anterior tibial posterior occlusion | -192
conscious | 0
not cooperative | 0
lower extremity pulses not obtained | 0
arterial blood pressure 120/60 mm Hg | 0
heart rate 120/min | 0
respiratory rate 24/min | 0
body temperature 36.5℃ | 0
O2 saturation 90% | 0
12-lead ECG showed sinus tachycardia | 0
diffuse atherosclerosis | 0
many thrombotic events | 0
brain MRI revealed multiple embolic infarcts | 0
carotid Doppler ultrasonography showed stenosis of bilateral internal carotid arteries | 0
chest CTA revealed embolism in right lower lobe | 0
segmental pulmonary artery branches embolism | 0
minimal consolidation area in left lung lower lobe |A0
echocardiography showed pericardial effusion | 0
left ventricular ejection fraction 60% | 0
upper extremity Doppler ultrasonography showed acute thrombosis of ulnar vein | 0
lower extremity CTA showed undefined crural artery circulation | 0
subacute deep vein thrombosis in bilateral main femoral vein | 0
admitted to intensive care unit | 0
non-invasive mechanical ventilation applied | 0
pleural fluid drained | 0
enoxaparin sodium administered | 0
iloprost administered | 0
asetilsalisilik asit administered | 0
anticoagulant therapy continued | 0
D-Dimer high | 0
platelets normal | 0
hereditary coagulation disorders not tested | 0
PF4 antibodies not tested | 0
vasculitis markers negative | 0
antinuclear antibody negative | 0
anti-double stranded DNA negative | 0
perinuclear anti-neutrophil cytoplasmic antibodies negative | 0
echocardiography normal | 0
prolonged ECG normal | 0
acute arterial thrombosis in both lower extremities | 0
necrosis in both lower extremities | 0
lower extremities amputated below the knee | 0
transferred to service | 24
discharged home | 24
readmitted to another hospital | 72
died | 312
