33 years old | 0
male | 0
diabetic | 0
admitted to the hospital | 0
left thigh pain | -5
denied any history of recent trauma | 0
former smoker | 0
quit smoking | -336
no personal or family history of hypercoagulable disorders | 0
no illicit substance use | 0
no respiratory symptoms | 0
diffusely swollen left thigh | 0
cyanotic left thigh | 0
tender left thigh | 0
tense left thigh | 0
left leg cool to touch | 0
intact motor function | 0
intact sensory function | 0
palpable femoral pulse | 0
popliteal and posterior tibial artery signals present | 0
computed tomography angiography | 0
bilateral multifocal ground-glass opacities | 0
consolidation in the lower lobes of the lungs | 0
COVID-19 infection | 0
acute occlusion of the left mid-superficial femoral artery | 0
significant swelling in the left thigh musculature | 0
therapeutic anticoagulation with unfractionated heparin | 0
angiography of the lower extremity | 0
fasciotomy of the left thigh | 0
elevated pressures in the anterior and posterior compartments | 0
decompressive fasciotomy | 0
muscles of the left thigh compartment appeared healthy | 0
venous duplex ultrasound examination negative | 0
arterial flow demonstrated to be normal | 0
viral myositis suspected | 0
full-dose anticoagulation | 0
empirical treatment of COVID-19 infection with hydroxychloroquine and azithromycin | 0
polymerase chain reaction test results positive | 24
workup for hypercoagulable disorders negative | 24
creatine kinase levels normal | 0
improved after the initial operation | 24
left thigh improved | 24
left calf soft and nonedematous | 24
no respiratory symptoms during hospitalization | 0
acute-onset severe left calf pain | 216
elevated compartment pressures | 216
palpable distal pulses | 216
no concern for arterial thrombosis | 216
emergent four-compartment fasciotomy | 216
muscle in each compartment significantly edematous | 216
diabetic ketoacidosis | 216
acute kidney injury | 216
thrombocytopenia | 216
extensive bilateral subsegmental pulmonary embolism | 216
bilateral lower extremity iliofemoral and inferior vena cava thrombosis | 216
diffuse arterial thrombosis | 216
cold extremities bilaterally | 216
intact motor and sensory function | 216
pain in the right calf | 264
elevated compartment pressures | 264
right lower extremity four-compartment fasciotomy | 264
muscle edematous and dusky | 264
right thigh compartment syndrome | 312
three-compartment fasciotomy | 312
therapeutic anticoagulation | 0
prophylactic broad-spectrum antibiotics | 0
convalescent antibody plasma therapy | 384
left below-knee amputation | 624
right above-knee amputation | 624
discharged to a rehabilitation facility | 624