Here is the table of events and timestamps:

18 years old | 0
male | 0
admitted to the hospital | 0
fever | -72
rash | -72
urinary tract infection | -120
empirically started on cephalexin | -120
urine analysis was positive for large leukocyte esterase and bacteria | -120
culture grew Escherichia coli | -120
prescribed cephalexin 500 mg three times daily | -120
started to develop an extensive erythematous rash | -96
rash developed into sloughing of the skin | -96
discontinued cephalexin | -96
transferred to a local burn intensive care unit | -96
chronic obstuctive pulmonary disease | -672
type 2 diabetes | -672
coronary artery disease | -672
hypertension | -672
hypothyroidism | -672
depression | -672
end-stage renal disease | -672
hemodialysis | -672
hydrocodone/acetaminophen | -672
levothyroxine | -672
escitalopram | -672
carvedilol | -672
guaifenesin | -672
docusate | -672
calcitriol | -672
albuterol | -672
amiodarone | -672
difficulty swallowing | 0
intubated | 0
toxic epidermal necrolysis syndrome | 0
blood pressure 81/45 mm Hg | 0
respiratory rate 12 breaths/min | 0
temperature 36.8 °C | 0
white blood cell count 1.5 × 10^3/mm^3 | 0
platelet count 77,000/µL | 0
serum creatinine 2.12 mg/dL | 0
venous serum lactate 3.1 mmol/L | 0
oxygen saturation 99% on 6 L O2 | 0
pain 9/10 | 0
urine culture from a newly placed indwelling Foley catheter | 0
chest radiograph revealed right pleural effusion with right lower and left basilar opacities | 0
intubated | 0
norepinephrine and vasopressin drips for pressure support | 0
albumin 25% continuous infusion | 0
Lactated Ringer’s 300 mL/h | 0
tetanus–diphtheria toxoids vaccine intramuscularly | 0
gentamicin 120 mg IV | 0
fluconazole 100 mg IV | 0
WBC 5.4 × 10^3/mm^3 | 48
SCr 1.98 mg/dL | 48
venous serum lactate 1.8 mmol/L | 48
random serum gentamicin level 2.4 mg/dL | 48
gentamicin 120 mg IV | 72
supportive continuous renal replacement therapy | 72
fluconazole 200 mg IV every 24 h | 72
Gram’s stain of the tracheal aspirate | 72
heavy growth of pleomorphic Gram-negative rods and diphtheroid-like Gram-positive rods | 72
wide complex tachycardia | 96
amiodarone restarted | 96
gentamicin held | 96
sloughing of skin over his back, chest, upper extremities, abdomen, bilateral thighs, and buttocks | 120
culture and sensitivity results of the tracheal aspirate | 120
Pseudomonas aeruginosa | 120
sensitive to all anti-pseudomonal beta-lactams as well as gentamicin, tobramycin, amikacin, and colistin | 120
another 120 mg dose of gentamicin | 120
random gentamicin level returned under 2 mg/dL | 120
expired | 144