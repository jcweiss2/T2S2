36 years old | 0
Hispanic | 0
gravida 3 para 0 | 0
17 weeks' gestation | 0
lower abdominal pain | -48
intestinal gas | -24
pain persistent | 0
pain severe | 0
pain exacerbated by movement | 0
loss of appetite | 0
denied nausea | 0
denied emesis | 0
tachycardic (120 beats per minute) | 0
involuntary guarding in suprapubic region | 0
sterile speculum examination | 0
normal closed cervix | 0
spontaneous rupture of yellow purulent fluid | 0
posterior vaginal fornix | 0
posterior vaginal wall defect | 0
significant relief upon rupture | 0
white blood cell count elevated (18.7) | 0
neutrophilic shift (94%) | 0
transvaginal ultrasound | 0
5 cm × 2 cm complex collection | 0
posterior cul-de-sac | 0
multiloculated abscess | 0
appendicitis not top differential diagnosis | 0
pelvic magnetic resonance imaging | 0
right ovarian torsion | 0
abscess formation due to appendicitis | 0
antibiotic treatment with ceftriaxone | 0
antibiotic treatment with metronidazole | 0
general surgery consultation | 0
met criteria for sepsis | 24
decompensated with worsening hypotension | 24
decompensated with worsening pain | 24
multidisciplinary meeting | 24
vancomycin added | 24
diagnostic laparoscopy | 24
examination under anesthesia | 24
1 × 1 cm defect in posterior fornix | 24
expression of purulent yellow fluid | 24
appendix adherent to uterus | 24
abscess | 24
appendectomy | 24
right fallopian tube difficult to visualize | 24
ovary difficult to visualize | 24
acute inflammatory process | 24
adhesions in right lower quadrant | 24
no additional abnormalities | 24
right lower quadrant Penrose drain | 24
fetal status reassuring | 24
postoperative piperacillin–tazobactam | 24
Penrose drain removal | 120
regular diet | 120
fetal status remained reassuring | 120
discharged on postoperative day 5 | 120
oral cefpodoxime | 120
recovering appropriately at follow-up | 120
pelvic abscess | 0
acute nonperforated appendicitis | 0
peritoneovaginal fistula | 0
second trimester pregnancy | 0
endometriosis | 0
decidualization on pathology | 0
uncomplicated normal spontaneous vaginal delivery | 4016
healthy infant | 4016
no malformations | 4016
no neurological sequelae | 4016
no behavioral sequelae | 4016
