68 years old | 0
male | 0
admitted to the ICU | 0
septic shock | 0
hospital acquired pneumonia | 0
multiple organ dysfunction syndrome |@ 0
deteriorated kidney function | 0
eGFR 9.8 ml/min/1.73 m² | 0
blood urea 221 mg/dl | 0
blood creatinine 5.6 mg/dl | 0
regular hemodialysis | 0
tracheostomy tube placement | 0
massive bleeding around tube stoma | 0
oxygen saturation 62% | 0
disseminated intravascular coagulation (DIC) | 0
elevated d-dimer 3500 mcg/L | 0
thrombocytopenia 76,000/μL | 0
prolonged prothrombin time 20.8 s | 0
flexible bronchoscopy | 0
blood clots at larynx and proximal trachea | 0
forceps extraction | 0
blood clot at distal trachea | 0
cryoextraction | 0
bleeding after clot removal | 0
argon plasma coagulation (APC) | 0
FiO2 set to 40% | 0
APC at carina, anterior, and right lateral wall of distal trachea | 0
oxygen saturation 98% | 0
reevaluation bronchoscopy two days later | 48
no new blood clots | 48
discharged two months later | 1464
