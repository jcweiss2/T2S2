64 years old | 0
woman | 0
referred to hepatobiliary surgery department | 0
previously admitted to ICU in local hospital | -unknown
severe sepsis | -unknown
liver abscess | -unknown
conservative treatment with IV antibiotics | -unknown
investigations attributed liver abscess to foreign body migration | -unknown
transferred to our hospital for surgical exploration | 0
past medical history not remarkable for comorbidities | 0
past medical history not remarkable for surgical procedures | 0
past medical history not remarkable for psychiatric disorders | 0
well controlled hypertension | 0
vital signs stable | 0
mild pain in right upper quadrant | 0
mild pain in flank | 0
denied foreign body ingestion | 0
denied recent trauma | 0
abdominal clinical examination no abnormalities | 0
normal white blood cells count | 0
C-reactive protein 48 mg/dL | 0
haemoglobin 9.2 g/dL | 0
hematocrit 24% | 0
aspartate aminotransferase AST 45.4 IU/L |#%0
alanine aminotransferase ALT 49.5 IU/L | 0
computed tomography scan CT-scan demonstrated hypodense area in right lobe of liver | -unknown
hypodense area measured about 3 x 4 cm | -unknown
linear hyperdense feature adjacent to hypodense area | -unknown
abdominal ultrasonography US exhibited elongated hyperechoic structure in segment V of liver | -unknown
scheduled for selective laparotomy | 0
subcostal incision with midline extension | 0
intraoperative finding of scar on out surface of segment V | 0
loose adhesions between first part of duodenum and inferior surface of liver | 0
toothpick's migration from D1 to liver suggested | 0
intraoperative ultrasound scan utilized to locate and mark foreign body | 0
5 cm incision in liver capsule | 0
finger fracture technique of hepatic parenchyma used | 0
toothpick found measuring 5.5 cm-long | 0
embedded in tough fibroid tissue within hepatic parenchyma | 0
depth of about 4 cm from liver capsule | 0
abdomen closed | 0
no drains used | 0
spent two days on ward | 0
discharged uneventfully | 48
denied ingesting foreign body | 0
adhesions between duodenum and liver suggested toothpick migration | 0
clinical manifestations contingent on time, site, depth of perforation | 0
liver abscess induced by foreign body symptoms: pain | -unknown
liver abscess induced by foreign body symptoms: fever | -unknown
toothpick found accidentally in porta hepatic during laparoscopic cholecystectomy | -unknown
foreign body asymptomatic until abscess developed | -unknown
suspicion raised for cryptogenic liver abscess | 0
suspicion raised for episode of foreign body ingestion | 0
suspicion raised for recurrent general unspecific symptoms | 0
CT scan pivotal in discovering foreign bodies inside liver | -unknown
ultrasonography may reveal radio-lucent foreign bodies | -unknown
CT scan necessitated to confirm diagnosis | -unknown
CT scan sufficient to detect foreign body, abscess, make surgical decision | -unknown
clinical presentation similar to acute abdominal conditions | 0
diagnosis strategy required to determine cause of abscess | 0
successive methods of treatment | 0
written informed consent obtained | 0
case report exempt from ethical approval | 0
no sponsors for this case report | 0
no conflicts of interest | 0
aspartate aminotransferase AST 45.4 IU/L | 0
no sponsors for this case report |0
investigations attributed liver abscess to foreign body migration |
