48 years old | 0
man | 0
known diabetic | 0
presented with increasingly painful swelling in the back below the left shoulder | 0
low-grade fever | -1080
occasional cough | -1080
vaccinated with COVID-19 vaccine on left deltoid | -240
onset of swelling | -240
developed painful swelling on left arm | -240
swelling spread to shoulder | -240
swelling spread to scapular region | -240
decreased limb movements | -240
acute onset of fever | -168
acute onset of cough | -168
mucoid expectoration | -168
progressive deterioration of health | -168
received anti-tubercular drugs | -168
febrile (38.8°C) | 0
left arm swollen | 0
left arm tender | 0
reduced range of movement | 0
unable to raise arm above shoulder | 0
ultrasound confirmed abscess | 0
chest radiographs showed disseminated pulmonary pathology | 0
bilateral lung abscesses | 0
pleural effusions | 0
pus culture yielded Burkholderia pseudomallei | 0
treated with intravenous meropenem | 0
resolution of abscess | 552
decrease in respiratory symptoms | 552
discharged | 552
advised oral trimethoprim-sulfamethoxazole | 552
