73 years old | 0
female | 0
Ecuadorian indigenous ancestry | 0
admitted to the hospital | 0
intense and diffuse colicky abdominal pain | -48
abdominal distension | -48
inability to eliminate flatus | -48
hypothyroidism | -8760
conventional cholecystectomy | -7200
no prior history of colitis | 0
no prior history of gastrointestinal disease | 0
signs of peritonism | 0
increased polymerase chain reaction | 0
no leukocytosis | 0
no neutrophilia | 0
no acidosis | 0
mild hypokalemia | 0
obstructive abdomen | 0
non-surgical medical treatment | 0
analgesia | 0
bowel rest | 0
hydration | 0
clinical improvement | 24
gastrointestinal disturbances recurred | 96
pain | 96
distension | 96
inability to eliminate flatus | 96
colonoscopy | 168
numerous mucosal patches | 168
erosions | 168
edema | 168
lymphoplasmacytic infiltration | 168
eosinophiles | 168
congestion | 168
hemorrhage | 168
parasitic bodies | 168
phagocyted red blood cells | 168
E. histolytica trophozoites | 168
serum antibodies against E. histolytica | 168
negative | 168
metronidazole | 168
unfavorable evolution | 192
abdominal distension | 192
pain | 192
feeding intolerance | 192
persistent mild hypokalemia | 192
normal renal function | 192
normal liver function | 192
down trending leukocytes | 192
pneumoperitoneum | 336
colonic perforation | 336
exploratory laparotomy | 336
fecal peritonitis | 336
pneumoperitoneum | 336
phlegmonous descending colon | 336
massive colon dilation | 336
transmural perforations | 336
total colectomy | 336
ileostomy | 336
rectal stump closure | 336
hypotension | 336
sepsis | 336
fluids | 336
vasoactive drugs | 336
meropenem | 336
metronidazole | 336
tinidazole | 336
superficial surgical site infection | 432
carbapenem-resistant Klebsiella pneumoniae | 432
extended spectrum beta-lactamase producing Escherichia coli | 432
colistin | 432
wound opened | 432
serial dressing changes | 432
discharged | 720
mucosal ulceration | 720
edema | 720
congestion | 720
lymphoplasmacytic infiltration | 720
eosinophils | 720
macrophages | 720
necrotic areas | 720
granulation tissue | 720
E. histolytica trophozoites | 720
late closure of ileostomy | 720