history of methicillin-resistant Staphylococcus aureus (MRSA) impetigo at the forearm | -8760
history of right tibia fracture treated with intramedullary fixation (IMN) | -8760
interlocking screws removed due to skin irritation and pain | -840
redness and swelling at the surgical site | -672
diagnosed with stitch abscess | -672
cultures from the surgical site were positive for MRSA | -672
prescribed an oral antibiotic treatment | -672
discharged home | -672
returned to the ER with a fever and right groin pain | -504
discharged home with the diagnosis of viral infection | -504
returned to the ER with a systemic fever | -448
myalgia | -448
difficult and painful ambulation | -448
right forearm cellulitis | -448
right sudden onset uveitis | -448
systemic rash | -448
right hip lymphadenopathy | -448
increased CRP level | -448
elevated WBC count | -448
hepatic enzymes, lactic dehydrogenase (LDH), creatine phosphokinase (CPK) levels were also elevated | -448
radiograph of both hips in anterior-posterior view was unremarkable | -448
advised to start the treatment with intravenous (IV) antibiotics | -448
medical condition continued to deteriorate | -336
positron emission tomography-computed tomography (PET-CT) scan was conducted | -336
revealed OIM abscess with systemic manifestations | -336
blood cultures were positive for MRSA bacteria | -336
showed signs of hemodynamic deterioration | -336
admitted to the intensive care unit (ICU) | -336
underwent ultrasound-guided drainage | -336
underwent a full-body CT scan | -192
result showed further enlargement of the abscesses diameter | -192
persistent fever | -192
CRP level of 36 mg/dL | -192
WBC count of 20,000 | -192
consulting the orthopaedic team | -96
surgical intervention was considered | -96
special surgical plan was developed | -96
combined approach of Smith-Peterson and modified Stoppa was chosen | -96
surgery | 0
general condition was improving | 24
less frequent fever spikes were noticed | 24
decrease in CRP and WBC levels | 24
additional antibiotic treatment support for 6 weeks | 24
almost complete recovery | 1440
able to ambulate normally without any pain or functional limitations | 1440
returned to his daily activities | 1440