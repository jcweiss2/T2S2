73 years old | 0
male | 0
admitted to the hospital | 0
signs of infection at the surgical site on his left hip | 0
avascular necrosis | -7200
staged bilateral THA | -7200
empty sella syndrome | -7200
neurosurgical bleeding | -7200
penicillin allergy | -7200
adrenal insufficiency | -7200
drug addiction | -7200
aseptic loosening of his left hip | -4320
one-stage revision | -4320
purulent wound drainage | -360
elevation of markers of infection | -360
deep THA infection | -360
joint aspiration | -360
Escherichia coli | -360
ampicillin resistance | -360
open debridement and irrigation with prosthetic retention | -360
antibiotic therapy | -360
DAIR | -360
intravenous ciprofloxacin | -360
Staphylococcus epidermidis | -360
vancomycin | -168
rifampicin | -168
prosthetic dislocation | 720
two-stage revision | 720
placement of a cement spacer with antibiotics | 720
empirical IV meropenem | 720
trimethoprim/sulfamethoxazole | 720
S. epidermidis | 720
teicoplanin | 720
ciprofloxacin | 720
fever | 840
persistent wound drainage | 840
new surgical debridement | 840
spacer kept in place | 840
deep vein thrombosis | 840
intestinal ischemia | 840
resection of the transverse and small colon | 840
ICU | 840
Candida parapsilosis | 840
antifungals | 840
fluconazole | 840
discharged from the hospital | 840
reactivation of his chronic wound infection | 2520
fever | 2520
fistulous lesions | 2520
purulent spontaneous drainage | 2520
revision of the cement spacer | 2520
methicillin-sensitive S. aureus | 2520
E. coli | 2520
Acinetobacter baumannii | 2520
re-implantation arthroplasty procedure | 2736
femoral tumor stem | 2736
uncemented porous tantalum cup | 2736
3D printing | 2736
dislocation | 3060
reactivation of his chronic infection | 3060
DAIR | 3060
wide resection of necrotic tissue | 3060
retention of all components | 3060
S. maltophilia | 3060
levofloxacin | 3060
prosthesis dislocation | 3276
suppressive antibiotic therapy | 3276
no signs of reactivation of the chronic infection | 3600
discontinuing the suppressive antibiotic therapy | 3600