33 years old | 0
female | 0
Gravida 3 | 0
Para 2 | 0
unplanned pregnancy | -2800
Zoladex implant for endometriosis | -2800
polyhydramnios | -2800
antenatal ultrasounds normal | -2800
non-consanguineous marriage | 0
family history free of congenital malformation | 0
previous two pregnancies normal | 0
one normal boy | 0
one normal girl | 0
admitted to the hospital | 0
dysmorphic | 0
weight 2.370 kg | 0
length 47 cm | 0
microcephaly | 0
head circumference 29 cm | 0
severely deformed nose | 0
one stenotic nostril | 0
cul-de-sac detected | 0
hypotelorism | 0
cleft palate | 0
microphthalmia | 0
micrognathia | 0
respiratory distress | 0
admitted to NICU | 0
septic workup | 0
endotracheal intubation | 4
severe respiratory distress | 4
complete blood count normal | 4
blood electrolytes normal | 4
blood gases normal | 4
chest X-Ray normal | 4
echocardiogram abnormal | 4
atrial septal defect | 4
patent ductus arteriosus | 4
renal ultrasound normal | 4
brain ultrasound abnormal | 4
mild lateral ventricle dilatation | 4
absence of septum pellucidum | 4
three-dimensional computed tomography scan | 4
single midline mono-ventricle | 4
dorsal cyst of holoprosencephaly | 4
fused cerebral hemisphere and thalami | 4
no midline septum pellucidum | 4
no corpus callosum | 4
no flax cerebri | 4
mono-nostril | 4
hypotelorism | 4
lobar holoprosencephaly | 4
skeletal survey normal | 4
karyotype normal | 4
feeding started | 72
orogastric tube | 72
gram-negative sepsis | 336
Pseudomonas aeruginosa | 336
Disseminated Intravascular Coagulation | 336
death | 336
autopsy not mentioned | 336 
note: the time is estimated based on the text, and the unit is hour.