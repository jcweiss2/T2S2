34 years old | 0
male | 0
admitted to the hospital | 0
penile discharge | -504
blurred vision in the left eye | -504
left knee pain | -504
Neisseria gonorrhea isolated from penile discharge | -504
corneal ulcer OS | -504
best corrected visual acuity (BCVA) of counting fingers (CF) at 1 foot OS | -504
corneal scrapings of the ulcer negative for bacteria or fungi | -504
slit lamp examination unremarkable OD | -504
best corrected visual acuity (BCVA) of 20/20 OD | -504
dilated fundus examination revealed normal optic discs, macula, retinal vessels, and periphery in both eyes | -504
intensive topical treatment with moxifloxacin and natamycin | -504
healing of the corneal ulcer | -168
rapid progressive diminution of vision OD | -168
referred to the uveitis service | -168
BCVA of 20/400 OD | -168
BCVA of 20/60 OS | -168
slit lamp examination OD revealed inferior keratic precipitates | -168
intense anterior chamber inflammation with a 1-mm hypopyon | -168
dispersed pigment on the anterior lens capsule | -168
posterior subcapsular cataract | -168
4+ vitreous haze with no fundus view | -168
B scan revealed significant vitreous opacities with a flat retina | -168
healed corneal ulcer with large central scarring and no epithelial defect OS | -168
fundus examination OS was unremarkable | -168
serum testing was negative for syphilis | -168
serum testing was negative for angiotensin converting enzyme | -168
serum testing was negative for lysozyme | -168
serum testing was negative for tuberculosis (T spot) | -168
serum testing was negative for human immunodeficiency virus | -168
diagnosis of infective endophthalmitis | -168
scheduled for urgent vitreous biopsy and pars plana vitrectomy (PPV) OD | -168
intraoperative fundus examination revealed dense vitreous opacification | 0
peripheral retinitis | 0
vasculitis | 0
localized inferotemporal rhegmatogenous retinal detachment | 0
retinal tear | 0
endolaser applied to the retinal tear | 0
air-fluid exchange | 0
left aphakic | 0
vitreous cavity filled with perfluoropropane (C3F8) | 0
intravitreal vancomycin (1mg) and ceftazidime (2.25 mg) | 0
topical ofloxacin and prednisolone acetate | 0
oral levofloxacin and doxycycline | 0
repeat intravitreal vancomycin (1 mg), ceftazidime (2.25 mg) combined with dexamethasone (0.4 mg) | 48
vitreous tap and culture were positive for Staphylococcus capitis | 48
vitreous tap and culture were negative for toxoplasmosis | 48
vitreous tap and culture were negative for lymphoma | 48
vitreous tap and culture were negative for cytomegalovirus | 48
vitreous tap and culture were negative for herpes simplex virus | 48
vitreous tap and culture were negative for varicella zoster virus | 48
vitreous tap and culture were negative for fungal agents | 48
blood cultures were negative | 48
tranthoracic echocardiography was negative for vegetations | 48
anterior chamber reaction and vitreous haze continued to improve | 168
BCVA was CF OD (without aphakic correction) | 168
vitreous cavity showed minimal vitreous haze | 168
flat retina with no retinitis | 168
50% gas fill | 168
placement of a sulcus intraocular lens | 672
BCVA had improved to 20/80 OD | 672
retina remained flat with no vitreous cavity inflammation | 672