40 years old| 0
South Asian male| 0
emergency department presentation| 0
sudden altered consciousness| -120
high fever| -120
progressive shortness of breath| -120
febrile (39.6°C)| 0
heart rate 140 beats/minute| 0
oxygen saturation 72%| 0
thin and cachectic appearance| 0
weight 62 kg| 0
poor nutritional status| 0
numerous mouth ulcers| 0
scrotal swelling with redness and tenderness| 0
Candida mucositis diagnosis| 0
COVID-19 rtPCR test| 0
chest CT| 0
HIV screening| 0
HIV negative| 0
USG scrotal edema| 0
elevated inflammatory markers| 0
brain CT right basal ganglia infarct| 0
chest CT CO-RADS 5| 0
TLC 25×10^9/L| 0
hemoglobin 5.34 mmol/L| 0
platelets 128×10^9/L| 0
CRP 1750 mg/L| 0
procalcitonin 11 mcg/L| 0
INR 1.6| 0
HbA1c 11.3%| 0
serum creatinine 170 µmol/L| 0
serum potassium 6.2 mmol/L| 0
serum lactate 8 mmol/L| 0
blood sugar 24 mmol/L| 0
severe metabolic acidosis| 0
sepsis diagnosis| 0
multiple organ dysfunction| 0
brain infarction| 0
severe viral pneumonia| 0
respiratory failure| 0
uncontrolled DM| 0
oral candidiasis| 0
acute kidney injury| 0
hyperkalemia| 0
hyperlactatemia| 0
ICU admission| 0
GCS 13/15| 0
HFNC therapy| 0
anticoagulation with enoxaparin| 0
remdesivir therapy initiation| 0
broad-spectrum antibiotics (tigecycline, levofloxacin)| 0
anidulafungin therapy initiation| 0
insulin therapy| 0
electrolyte replenishment| 0
COVID-19 rtPCR positive| 24
left leg swelling| 24
iliofemoral DVT| 24
enoxaparin dose increased| 24
consciousness regained| 24
hemodynamic improvement| 24
ventilatory improvement| 24
fever subsided| 24
hyperglycemia controlled| 24
TLC 14×10^9/L| 24
oxygenation improvement| 24
weaned to nasal cannula| 24
CRP high| 24
procalcitonin high| 24
anti-cytokine therapy not initiated| 24
supine and self-prone positioning| 24
clinical deterioration| 168
GCS 5/15| 168
oxygen requirement increased| 168
hypotension requiring norepinephrine| 168
TLC 23×10^9/L| 168
refractory hypoglycemia| 168
dextrose 50% infusion| 168
remdesivir discontinued| 240
chest X-ray worsening bilateral infiltrates| 240
sputum culture Klebsiella pneumoniae| 240
sputum culture Candida albicans| 240
HAP diagnosis| 240
invasive mechanical ventilation| 240
antibiotics changed to meropenem, linezolid| 240
anidulafungin continued| 240
fever subsided| 240
TLC 15×10^9/L| 240
euglycemia achieved| 240
vasopressors weaned| 240
oxygen requirement decreased| 240
extubated| 288
HFNC continued| 288
ICU extended stay| 288
oxygenation deteriorated| 336
reintubation| 336
oxygen requirement 70%| 336
suspected PE| 336
CT angiogram no PE| 336
HRCT chest cavitary lesions| 336
pleural effusion| 336
necrotizing pneumonia| 336
lung abscess| 336
pleural drainage| 336
BAL Candida albicans| 336
meropenem continued| 336
linezolid continued| 336
anidulafungin continued| 336
clinical improvement| 432
extubated| 432
meropenem dose adjusted| 432
linezolid oral therapy| 432
voriconazole initiation| 432
weaned off HFNC| 528
oxygen support discontinued| 720
ICU stay until room air| 720
nutritional support| 720
anticoagulation titration| 720
DM control| 720
regular ward transfer| 888
chest X-ray improvement| 888
discharge| 1416
