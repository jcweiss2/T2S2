54 years old| 0
    woman | 0
    Roux-en-Y procedure | -105840
    exploratory laparotomy | -2160
    small bowel obstruction | -2160
    altered mental status | -72
    confusion | -72
    hallucinations | -72
    chest pain | -72
    blood pressure 119/78 mmHg | 0
    pulse 85 beats per minute | 0
    temperature 97.8 F° | 0
    respiratory rate 18/minute | 0
    SpO2 84% | 0
    Glasgow Coma Scale 13/15 | 0
    alert | 0
    awake | 0
    not oriented to person | 0
    not oriented to place | 0
    not oriented to time | 0
    lung exam bilateral coarse crackles | 0
    expiratory wheezes | 0
    cardiovascular exam regular rate and rhythm | 0
    normal S1 | 0
    normal S2 | 0
    no murmurs | 0
    no gallops | 0
    electrocardiogram normal sinus rhythm | 0
    no ST changes | 0
    no T wave changes | 0
    abdomen exam present bowel sounds | 0
    mild diffuse tenderness to palpation | 0
    3 cm abdominal wound | 0
    healing well | 0
    no surrounding erythema | 0
    no exudate | 0
    white blood cell count 11.8×10³/mm³ | 0
    total bilirubin 3.2 mg/dL | 0
    AST 131 U/L | 0
    ALT 178 U/L | 0
    ALK phosphate 339 IU/L |1
    urinalysis negative for infections | 0
    urine drug screen positive for opiates | 0
    urine drug screen positive for benzodiazepines | 0
    arterial blood gas pH 7.37 | 0
    PCO2 40.7 | 0
    PO2 56 | 0
    HCO3 23.3 | 0
    chest X-ray multi-lobar pneumonia | 0
    brain MRI right fronto-parietal infarct | 0
    brain MRI left cerebellar infarct | 0
    BiPAP placement | 0
    blood cultures drawn | 0
    IV antibiotics started | 0
    Vancomycin | 0
    Cefepime | 0
    Metronidazole | 0
    transfer to critical care unit | 0
    severe acute hypoxic respiratory failure | 24
    intubation | 24
    trans-esophageal echocardiogram | 24
    multi-lobar infarct diagnosis | 24
    Eustachian valve vegetations | 24
    diffuse hypokinesia | 24
    left ventricle ejection fraction 30% | 24
    patent foramen ovale | 24
    blood cultures Staphylococcus capitis | 24
    bronchoalveolar lavage culture Methicillin Resistant Staphylococcus Aureus | 24
    extubation | 168
    mental status improved | 168
    residual left facial droop | 168
    residual left upper extremity weakness | 168
    repeat transthoracic echocardiogram ejection fraction 45-50% | 168
    normal Eustachian valve | 168
    repeat blood cultures negative | 96
    discharge to skilled nursing facility | 168
    IV Vancomycin continued | 168
    Cefepime continued | 168
    antibiotics duration 6 weeks | 168
    repeat transthoracic echocardiogram prominent Eustachian valve | 672
    no vegetation | 672
    ejection fraction 55% | 672
    multi-lobar pneumonia | 0
    acute ischemic edema right posterior frontal parietal distribution | 0
    acute ischemic edema left cerebellar hemisphere | 0
    <|eot_id|>
    