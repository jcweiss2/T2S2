22 years old | 0
Japanese woman | 0
referred to the hospital | 0
persistent high fever | 0
systemic joint pain | 0
low saturation of pulse oximetry oxygen | 0
appearance of blastic cell | 0
low platelet count | 0
high fever (38.9°C) | -120
pain of several joints | -120
acetaminophen | -120
antibacterial agent | -120
healthy until the onset of disease | -120
nonconsanguineous parents | -120
no family history of similar disorders | -120
body temperature 37.8°C | 0
acetaminophen response | 0
SpO2 99% under O2 inhalation of 3 L/min | 0
no systemic superficial lymphadenopathy | 0
no skin eruption | 0
white blood cell count 6680/μL | 0
atypical lymphocytes 44% | 0
hemoglobin 15.2 g/dL | 0
hematocrit 43.5% | 0
platelet count 2.6 × 104/μL | 0
PT 16.9 sec | 0
PT-INR 1.59 | 0
APTT 71.8 sec | 0
Fibrinogen 160.4 mg/dL | 0
FDP 137.6 μg/mL | 0
total protein 5.1 g/dL | 0
albumin 2.8 g/dL | 0
AST 537 IU/L | 0
ALT 256 IU/L | 0
LDH 5574 IU/L | 0
total bilirubin 5.4 mg/dL | 0
direct bilirubin 4.7 mg/dL | 0
ALP 1174 IU/L | 0
TG 362 mg/dL | 0
BUN 68.6 mg/dL | 0
Cre 2.67 mg/dL | 0
UA 13.3 mg/dL | 0
CRP 17.78 mg/dL | 0
serum ferritin 23,700 ng/mL | 0
sIL-2R 35,300 U/mL | 0
CT scan bilateral pneumonia | 0
bilateral pleural effusion | 0
mild cardiomegaly | 0
intra-abdominal lymph node swelling | 0
hepatosplenomegaly | 0
bone marrow examination medium to large-sized atypical lymphoid cells | 0
active histiocytes with prominent hemophagocytosis | 0
flow cytometric analysis CD8-positive T-cells | 0
clonal T-cell lymphoproliferative disease | 0
EBV-associated disease | 0
hemophagocytosis | 0
multiorgan damages | 0
coagulopathy | 0
methylprednisolone pulse therapy | 0
CHOPE chemotherapy | 24
antibiotics for GPC and GNR | 0
blood culture | 0
transient abatement of fever | 0
another cycle of CHASE chemotherapy | 288
high fever flare-up | 288
pneumonia exacerbation | 288
PaO2 55 mmHg | 288
O2 inhalation 10 L/min | 288
moved to ICU | 288
CPAP | 288
BiPAP | 288
transient effects of CHASE | 288
third cycle of chemotherapy with high-dose MTX and AraC | 576
mPSL pulse | 576
reappearance of high fever | 576
exacerbation of pneumonia | 576
bone marrow suppression | 576
rhG-CSF use | 576
allo-HSCT required | 576
older brother as allo-BMT donor | 576
HLA-DRB1 allele mismatch | 576
MAC started | 864
ALT 64 IU/L | 864
LDH 355 IU/L | 864
sustained low-grade fever | 864
remaining lung infiltrative shadows | 864
conditioning regimen ETP 15 mg/kg | 864
CY 60 mg/kg | 864
TBI 12 Gy | 864
allo-BMT | 1104
BM cells 3.25 × 108/kg | 1104
GVHD prophylaxis FK506 | 1104
short-term MTX | 1104
engraftment at day 18 | 1296
Y-chromosome 99.3% | 1296
acute grade II GVHD of the skin | 672
controlled with local treatment | 672
no VOD | 672
no TMA | 672
no severe infections | 672
grade III GVHD flare-up | 1776
PSL commenced 1 mg/kg | 1776
skin GVHD cleared | 1776
AST 19 IU/L | 2400
ALT 34 IU/L | 2400
LDH 273 IU/L | 2400
ferritin 2078.3 ng/mL | 2400
sIL-2R 331 U/mL | 2400
EBV-DNA viral load <2.0 × 101 copies/106 cells | 2400
Southern blotting no clonality | 2400
CT scan no lymph node swelling | 2400
no hepatosplenomegaly | 2400
discharged from the hospital | 3456
PSL tapered | 8640
FK506 tapered | 12240
undetectable FK506 trough levels | 8640
complete remission | 3456
normal laboratory data | 26280
no EBV-DNA viral load | 26280
EBV titers VCA IgG ×640 | 26280
VCA IgM <×10 | 26280
VCA IgA ×10 | 26280
EA-DR IgG ×80 | 26280
EA-DR IgA <×10 | 26280
EBNA ×80 | 26280
successful allo-BMT | 1104
complete remission for 3 years | 26280
no EBV-DNA detection | 26280
