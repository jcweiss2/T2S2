62 years old | 0
male | 0
admitted to the hospital | 0
fever | -48
hypotension | -48
high-grade fever | -72
arthralgia | -72
generalized malaise | -72
shock identified | -72
systolic blood pressure 72 mmHg | -72
heart rate 110 beats per minute | -72
pain in lateral aspect of right elbow | -72
transferred to our hospital | -72
tachypneic | 0
blood pressure 102/66 mmHg | 0
heart rate 114 beats per minute | 0
respiratory rate 28 breaths per minute | 0
febrile 38.5°C | 0
required oxygen | 0
oxygen saturation 94% on 3 L/min cannula | 0
chest examination no abnormalities | 0
abdominal examination no abnormalities | 0
lateral aspect of right elbow erythematous | 0
lateral aspect of right elbow visibly swollen | 0
tenderness on palpation | 0
entered state of shock | 0
disseminated intravascular coagulation (DIC) | 0
multiple organ failure (MOF) | 0
intensive care required | 0
blood cultures obtained | 0
Streptococcus pyogenes in blood cultures | 0
right arm evaluated with CT | 0
examined by surgeon | 0
fasciotomy performed | 0
debridement performed | 0
necrotizing fasciitis | 0
streptococcal toxic shock syndrome (STSS) diagnosed | 0
initial contrast-enhanced abdominal CT no IPA | 0
intubation required | 0
emergency surgery for right arm | 0
hemodynamic instability | 0
vasopressors | 0
antibiotics | 0
fluid management | 0
ventilation support | 0
became afebrile | 360
high-grade fever | 816
hypotension | 816
tachycardia | 816
leukocytosis | 816
evidence of MOF | 816
vasopressors to maintain hemodynamic stability | 816
abdominal CT demonstrated left IPA | 816
no pathological findings in right arm | 816
no pathological findings in chest | 816
no pathological findings in abdomen | 816
other sources of infection ruled out | 816
Klebsiella pneumoniae in blood cultures | 816
critically ill | 816
drainage of primary IPA not performed | 816
intravenous antibiotics | 816
responded to antibiotic treatment | 816
MOF improved | 816
CT-guided drainage performed | 1272
culture of drainage specimen no bacteria | 1272
drainage tube removed | 1968
follow-up abdominal CT confirmed shrinkage of IPA | 1968
began rehabilitation | 1968
discharged | 1968
ongoing follow-up | 1968
excellent results in activities of daily living | 1968
