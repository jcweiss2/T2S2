85 years old | 0
    female | 0
    visited emergency room | 0
    painful swelling on bilateral submandibular | 0
    painful swelling on submental | 0
    painful swelling on upper neck areas | 0
    overlying skin was edematous | 0
    overlying skin was reddish | 0
    ill-defined reddish border | 0
    extreme pain in upper neck area | 0
    underwent endodontic treatment on lower central incisor | -168
    symptoms persisted | -168
    swelling developed suddenly | -168
    febrile | 0
    body temperature 39℃ | 0
    medical history of steroid due to arthralgia | 0
    WBC 10.26×103/µL | 0
    ESR 3 mm/hr | 0
    neutrophil 93.1% | 0
    aPTT 45.9 seconds | 0
    CRP 202.96 mg/L | 0
    CT showed disseminated deep neck abscess | 0
    abscess extended into upper mediastinum | 0
    abscess extended to supraclavicular area | 0
    abscess extended to axillary areas | 0
    initial diagnosis odontogenic abscess | 0
    drained abscess | 0
    incised submental area | 0
    incised submandibular areas | 0
    dissected with fingers | 0
    dissected with mesenbaum scissors | 0
    underlying fascia opened | 0
    small amount of pus discharged | 0
    fascia discolored grayish | 0
    suggested fasciitis | 0
    incised skin along anterior border of sternocleidomastoid muscle | 0
    fascia along anterior neck discolored grayish | 0
    fascia along carotid sheath discolored grayish | 0
    detached diseased fascia from submental area to upper mediastinum | 0
    incised supraclavicular area | 0
    incised anterior border of trapezius muscle | 0
    explored infected areas | 0
    inserted silicon drains | 0
    administered triple antibiotic regimen | 0
    penicillin | 0
    aminoglycoside | 0
    metronidazole | 0
    microscopic examination acute infection | 0
    microscopic examination chronic infection | 0
    lymphocyte infiltration in necrotic fascia | 0
    diagnosed necrotizing fasciitis | 0
    pus culture betahemolytic streptococcal infection | 0
    sensitive to most antibiotics | 0
    condition not improved | 96
    CT showed infection spread under trapezius muscle | 96
    skin over shoulder area intense hot | 96
    skin over shoulder area reddish | 96
    airway obstruction expected | 96
    WBC 13.18×103/µL | 96
    ESR 15 mm/hr | 96
    neutrophil 87.7% | 96
    aPTT 46.3 seconds | 96
    CRP 151.46 mg/L | 96
    drained area under trapezius muscle | 96
    obtained artificial airway | 96
    tracheostomy | 96
    incised anterior border of trapezius muscle to greater extent | 96
    incised suprascapular area | 96
    inserted drain through and through | 96
    changed old drain | 96
    sent to intensive care unit | 96
    administered ventilator therapy | 96
    skin infection extended to upper chest | 240
    skin infection extended to shoulder area | 240
    CT showed multifocal abscess around left chest wall | 240
    CT showed multifocal abscess around shoulder area | 240
    CT showed multifocal abscess around carotid area | 240
    CT showed further deterioration | 240
    WBC 12.21×103/µL | 240
    ESR 11 mm/hr | 240
    neutrophil 75.7% | 240
    aPTT 38.6 seconds | 240
    CRP 14.2 mg/L | 240
    suspected uncontrolled necrotizing fasciitis | 240
    performed third operation | 240
    incised skin on chest over healthy area | 240
    dissected infected skin | 240
    elevated skin | 240
    subcutaneous fat necrotized | 240
    superficial fascia necrotized | 240
    dissected carotid space with finger | 240
    dissected necrotic tissue around upper chest | 240
    dissected necrotic tissue around trapezius area | 240
    pus culture Actinibacter baumanni | 240
    resistant to cabepenem | 240
    resistant to most antibiotics | 240
    changed antibiotic regimen to vancomycin | 240
    fasciotomy | 240
    skin loosely sutured | 240
    inserted drains | 240
    infection decreased gradually | 240
    skin over distal clavicular area not salvaged | 888
    closed skin with bilobed rotational flap | 888
    removed tracheostomy tube | 960
    discharged | 1344
    WBC 10.08×103/µL | 1344
    ESR 5 mm/hr | 1344
    neutrophil 71.3% | 1344
    aPTT 25.7 seconds | 1344
    CRP 20.4 mg/L | 1344