25 years old | 0
female | 0
nausea | -2
vomiting | -2
dizziness | -2
abdominal pain | -2
altered sensorium | -2
ingestion of mosquito repellent | -2
conscious | 0
pupils bilaterally semi constricted | 0
pupils sluggishly reactive to light | 0
crepitations present bilaterally | 0
respiratory rate 28/min | 0
blood pressure 110/70 mmHg | 0
gastric lavage | 0
gastric aspiration | 0
oral syrup charcoal | 0
atropine | 0
pantoprazole | 0
ondansetron | 0
tonic-clonic convulsions | 1
injection phenytoin | 1
injection diazepam | 1
injection hydrocortisone | 1
injection frusemide | 1
oxygen enrichment | 1
uncontrolled convulsions | 1
shifted to intensive care unit | 1
midazolam | 1
propofol | 1
endotracheal intubation | 1
oxygen enrichment | 1
midazolam infusion | 1
propofol infusion | 1
SpO2 maintained at 100% | 1
blood pressure 94/62 mmHg | 1
pulse rate 74/min | 1
arterial blood gas reports normal | 1
IV mannitol | 1
IV phenobarbitone | 1
seizure free for few hours | 2
seizures started again | 2
blood pressure 80/40 mmHg | 2
respiratory rate 35/min | 2
pulse rate 190/min | 2
SpO2 95% | 2
serum potassium 2.98 mmol/L | 2
serum calcium 2.5 mmol/L | 2
serum sodium 129 mmol/L | 2
injection dopamine | 2
potassium chloride | 2
hypertonic saline | 2
elective ventilation | 2
muscle paralysis | 2
controlled mechanical ventilation | 2
vecuronium | 2
dopamine dose increased | 2
propofol infusion stopped | 2
ABG reports no changes | 2
computed tomography scan of brain normal | 2
chest X-ray normal | 2
input/output charting for fluids | 2
central venous pressure 5-8 cm H2O | 2
ventilator for 48 h | 48
weaning started | 48
vecuronium and midazolam infusion stopped | 48
mode of ventilation changed to SIMV | 48
airway pressure support set | 48
positive end expiratory pressure set | 48
pulse rate 102 beats/min | 48
blood pressure 132/82 mmHg | 48
SpO2 above 96% | 48
total leucocyte count 7200/mm3 | 24
total leucocyte count 22,000/mm3 | 48
total leucocyte count 32,000/mm3 | 72
total leucocyte count 13,000/mm3 | 96
total leucocyte count 4000/mm3 | 144
dopamine infusion tapered down | 54
dopamine infusion stopped | 60
spontaneous respiration noticed | 60
muscle relaxation reversed | 60
neostigmine | 60
glycopyrrolate | 60
patient extubated | 60
oxygen through mask | 60
respiratory rate 25 breaths/min | 60
blood pressure 108/72 mmHg | 60
pulse rate 119/min | 60
pupils normally reacting to light | 60
nebulised with mistabron | 60
referred to psychiatrist | 96
shifted to ward | 96
discharged from hospital | 168