65 years old | 0
male | 0
admitted to the hospital | 0
chest pain | 0
radiated to left and right arms | 0
electrocardiogram showed anterolateral ischemia | 0
acute myocardial injury | -336
coronary angiography showed 90% stenosis of the circumflex artery | -336
percutaneous transluminal coronary angioplasty | -336
stent placement on left main, left anterior descending, and left circumflex | -336
dual antiplatelet therapy | -252
discharged from the hospital | -252
positive for Coronavirus-19 | -252
new ischemic episode | -144
uncompliant with DAPT therapy | -144
cardiac arrest | 0
ventricular fibrillation | 0
femoro-femoral VA-ECMO support | 0
second coronary angiography | 0
stent placement | 0
intra-aortic balloon pump placement | 0
trans-esophageal echocardiography | 0
severe LV dysfunction | 0
interventricular septum hypokinesia | 0
left atrial smoke | 0
minimal aortic valve opening | 0
mild aortic insufficiency | 0
severe reduction of right ventricle longitudinal and concentric function | 0
transeptal left atrial cannulation | 480
VA-ECMO converted to LAVA-ECMO | 480
TEE demonstrated improvement in right ventricle movement | 504
Levosimendan infusion | 504
transferred to cardiothoracic ICU | 528
progressive weaning from VA-ECMO | 528
oxygenator removed from the circuit | 528
LVAD | 528
vasopressor and inotropic support decreased | 528
platelet count reduced | 528
bleeding | 528
sepsis | 528
anticoagulation monitored | 528
activated coagulation time monitored | 528
activated partial thromboplastin time monitored | 528
pneumonia diagnosed | 528
antibiotics started | 528
fibro-bronchoscopies done | 528
renal failure | 528
continuous renal replacement therapy | 528
uncontrolled airway bleed | 936
death | 936