obesity | -20 years
psoriatic arthritis | -20 years
surgical hypoparathyroidism | -20 years
hypothyroidism | -20 years
total thyroidectomy | -20 years
multinodular goitre | -20 years
elective sleeve gastrectomy | 0
gastric perforations | 0
abdominal sepsis | 4
transfer to intensive care | 4
critically low calcium level | 4
continuous intravenous calcium gluconate infusion | 4
maintenance intermittent IV calcium boluses | 4
prolonged ICU admission | 4
weight loss 14 kg | 6 months
endocrinology advice | 14
TSH 5.83 mU/L | 14
intravenous triiodothyronine 10 µg BD | 14
euthyroidism | 14
high dose intravenous calcium | 14
ionised calcium measured daily | 14
serum phosphate level 1.07 | 14
intravenous calcitriol 1 µg alternate daily | 20
intravenous calcitriol ceased | 25
intramuscular cholecalciferol 150 000 units | 42
low 1,25(OH)vitamin D3 level | 42
normal renal function | 42
intravenous calcitriol recommenced | 84
intravenous thyroxine 200 µg alternate daily | 88
maintenance schedule established | 120
discharge from hospital | 240
normocalcaemia on review | 240
weight 71.8 kg | 240
BMI 29 kg/m2 | 240
follow-up 6 weeks | 276
follow-up 12 weeks | 300
follow-up 4 months | 336