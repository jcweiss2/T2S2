32 weeks pregnant | -672
decreased fetal movement | -672
fetal ultrasound | -672
fetal ascites | -672
edematous bowel loops | -672
antenatal scan | -672
TORCH | -672
emergency cesarean section | 0
abdominal distention | 0
mass felt on the right umbilicus | 0
shifted to the neonatal intensive care unit | 0
upper gastrointestinal contrast study | 0
normal C-loop | 0
ruled out malrotation | 0
altered nasogastric aspirates | 0
serial X-ray | 0
absence of flow of dye | 0
obstruction | 0
hemoglobin of 6 gm% | 0
clinical suspicion of bowel gangrene | 0
clinical suspicion of volvulus | 0
emergency laparotomy | 6
volvulus | 6
gangrene of 45 cm of the distal ileum | 6
herniating through mesenteric defect | 6
resection of gangrenous segment | 6
ileostomy | 6
ileocecal junction preserved | 6
elective stoma closure | 1800
uneventful hospital course | 1800
child is 5-year-old | 43800
growing well | 43800
no sequel of her disease | 43800