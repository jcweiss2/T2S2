49 years old | 0
female | 0
fell whilst bathing | -2
struck her face on the bath tap faucet | -2
5 cm partial thickness laceration below her left eye | -2
attended A&E department | -2
laceration was debrided, irrigated and sutured | -2
Elhers–Danlos syndrome | 0
ischaemic heart disease | 0
previous anaphylaxis to penicillin | 0
returned to A&E | -24
complaining of pain and swelling below the left eye | -24
eye was partially closed secondary to lower lid swelling | -24
eye examination was normal | -24
no deficit in visual acuity recorded | -24
discharged with oral clarithromycin | -24
re-attended A&E | -48
pyrexial | -48
tachycardic | -48
evidence of rigors | -48
confusion | -48
extensive left-sided facial swelling | -48
complete closure of the left eye | -48
involvement of the soft tissues of the left neck | -48
reduction in left visual acuity | -48
marked neutrophilia | -48
raised C-reactive protein | -48
laceration was opened | -48
necrotic skin edges | -48
absence of bleeding | -48
severe facial necrotizing fasciitis | -48
admitted | -48
underwent immediate widespread local excision of necrotic tissue | 0
peri-operative and post-operative IV clindamycin and gentamicin | 0
transferred to ICU | 0
reviewed the following morning | 24
clinically septic | 24
clear extension of necrotic tissue | 24
left eye involvement suspected | 24
urgent CT scan | 24
tissue features in keeping with a left retro-orbital necrosis | 24
further surgical excision of necrotic tissue | 48
exenteration of left orbital contents | 48
blood and tissue samples sent to microbiology laboratory | 48
cultured a florid growth of a Group A beta-haemolytic Streptococci | 48
confirmed the clinical suspicion of facial necrotizing fasciitis | 48
2-week period in ICU | 168
transferred for 3 weeks of ward-based care | 336
continued on oral clindamycin | 336
initial reconstruction with a split thickness skin graft | 504
second graft required | 504
current appearance | 1296