52 years old | 0
female | 0
abdominal pain | -48
nausea | -48
vomiting | -48
diarrhea | -24
increased liver enzyme alanine aminotransferase | -840
positive autoimmune antibody | -840
elevated immunoglobulin G | -840
coarse liver surface | -840
liver biopsy | -840
overlap syndrome | -840
autoimmune hepatitis | -840
ursodeoxycholic acid | -840
prednisolone | -840
mild heartburn | -48
abdominal tenderness | 0
mild fever | 0
tachycardia | 0
tachypnea | 0
abdominal hardness | 0
reduced white blood cells | 0
reduced platelets | 0
decreased neutrophil level | 0
elevated C-reactive protein level | 0
elevated aspartate aminotransferase | 0
elevated ALT | 0
elevated gamma glutamyl transferase | 0
prothrombin time international normalized ratio | 0
necrotizing gastritis | 0
septic shock | 0
intravenous hydration | 0.5
antibiotic treatment | 0.5
inotropics | 2
fluid treatment | 2
increased blood pressure | 2
severe stress-induced cardiomyopathy | 3
extracorporeal membrane oxygenation | 3
cardiac arrest | 3
death | 3
azathioprine | -336
reduced prednisolone | -144
discharge | -144 
admitted to the emergency room | 0 
admitted to the intensive care unit | 0.5 
discharged | -840