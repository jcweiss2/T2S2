10 weeks old|0
male|0
admitted to the hospital|0
abdominal distension|-24
lethargy|-24
fever|-72
poor feeding|-72
vomiting|-72
cessation of bowel movements|-24
progressive abdominal distension|-24
irritability|-24
small for gestational age|0
delayed in passing meconium at birth|0
constipation|0
up to date vaccination schedule|0
no family history of Hirschsprung's disease|0
no congenital disorders|0
height <3 percentile|0
weight <3 percentile|0
afebrile|0
tachycardia|0
tachypnea|0
hypotension|0
oxygen saturation 97%|0
unwell appearance|0
lethargy|0
marked dehydration|0
pale mottled skin|0
distended abdomen|0
tense abdomen|0
tender abdomen|0
reduced bowel sounds|0
agitation|0
crying|0
high leukocyte count|0
neutrophilia|0
thrombocytosis|0
elevated C-reactive protein|0
hyponatremia|0
hyperglycemia|0
elevated SGOT|0
elevated SGPT|0
compensated metabolic acidosis|0
multiple air fluid levels|0
distended loops of small intestine|0
no pneumoperitoneum|0
clinical sepsis|0
fluid resuscitation|0
broad-spectrum antibiotics|0
complicated intestinal obstruction|0
urgent laparotomy|0
ileal dilatation|0
ileal perforation|0
primary repair of ileal perforation|0
totally collapsed microcolon|0
Hirschsprung's disease diagnosis|0
transition zone at ileocecal valve|0
full thickness biopsies|0
appendectomy|0
protective ileostomy|0
absence of ganglion cells|0
enterocolitis|0
progressive deterioration post-surgery|0
intubation|0
monitoring in neonatal ICU|0
cardiopulmonary arrest|0
unsuccessful resuscitation|0
final diagnosis of ileal perforation|0
sepsis|0
septic shock|0
total colonic aganglionosis|0
death|24
