72-year-old-man | 0
hemodialysis | -149448
diabetic nephropathy | -149448
admitted to the emergency room | 0
fever | 0
penile pain | 0
vomiting | 0
diarrhea | 0
percutaneous transluminal angioplasty of the lower extremities | -149448
lanthanum carbonate hydrate | -149448
calcium carbonate | -149448
cilostazol | -149448
lansoprazole | -149448
cinacalcet | -149448
amlodipine | -149448
enalapril maleate | -149448
carvedilol | -149448
non-smoker | -149448
no alcohol consumption | -149448
good general condition | 0
physical examination | 0
penile pain worsened | -9
revisited the emergency room | -9
lost consciousness | -9
Glasgow Coma Scale score of 3 | 0
blood pressure 84/58 mmHg | 0
respiratory rate 28 breaths per minute | 0
heart rate 102 beats per minute | 0
temperature 37.6°C | 0
oxygen saturation 100% | 0
cold sweat | 0
swelling at the glans | 0
dark brownish changes at the glans | 0
white blood cell count 5,600 /μL | 0
hemoglobin 10.2 g/dL | 0
platelets 81,000 /μL | 0
sodium 141 mmol/L | 0
potassium 5.3 mmol/L | 0
chloride 103 mmol/L | 0
creatinine 9.71 mg/dL | 0
blood urea nitrogen 47.7 mg/dL | 0
albumin 3.3 g/dL | 0
calcium 9.4 mg/dL | 0
phosphorus 5.8 mg/dL | 0
parathyroid hormone 280 pg/mL | 0
C-reactive protein 129.8 mg/L | 0
total bilirubin 1.5 mg/dL | 0
aspartate aminotransferase 34 IU/L | 0
alanine aminotransferase 10 IU/L | 0
pH 7.031 | 0
PaCO2 62.4 Torr | 0
PaO2 80.6 Torr | 0
HCO3 15.7 mEq/L | 0
anion gap 25.0 mmol/L | 0
respiratory condition deteriorated | 0
worsening metabolic acidosis | 0
worsening respiratory acidosis | 0
hyperkalemia | 0
intubated | 0
admitted to the intensive care unit | 0
blackish changes on the entire penis | 3
blackish changes on the scrotum | 3
test incision in the perineum | 3
test incision in the penis | 3
test incision in the scrotum | 3
no effusion detected | 3
contrast-enhanced computed tomography | 3
no intestinal necrosis | 3
poor contrast enhancement of the penis | 3
no abscess | 3
no gas in the penis | 3
antibiotics | 3
vancomycin | 3
meropenem | 3
vasoactive agents | 3
noradrenaline | 3
vasopressin | 3
hydrocortisone | 3
continuous hemodiafiltration dialysis | 3
metabolic acidosis progressed | 3
hyperkalemia progressed | 3
died | 12
postmortem blood culture showed Streptococcus dysgalactiae subsp. equisimilis | 12
diagnosis of STSS | 12
antimicrobial susceptibility sensitive to β-lactam antibiotics | 12
calcification of the aorta | 12
ischemic necrosis of the stomach | 12
ischemic necrosis of the lower gastrointestinal tract | 12
calcified lesions | 12
infected thrombi in the subcutaneous tissue of the penis | 12
infected thrombi in the scrotum | 12
infected thrombi in the arterioles of the bladder wall | 12
