70 years old | 0
male | 0
emergency esophageal diversion | -720
injury to the cervical esophagus | -720
spinal surgery | -720
gastric pull-up procedure | -168
postoperative anastomotic leakage | -168
endoscopy | -168
esophageal stent | -168
discharged | -126
local cervical infection | -126
sepsis | -126
admitted to hospital | 0
malnutrition | 0
systemic inflammation | 0
jugular and cervical phlegmon | 0
hemoglobin level of 6.7 g/dL | 0
white blood cell count of 6400 cells/μL | 0
platelet count of 210 × 10^3/μL | 0
creatinine level of 0.76 mg/dL | 0
albumin level of 2.8 g/dL | 0
chest computed tomography scan | 0
endoscopy | 0
dislodged esophageal stent | 0
esophageal perforation | 0
infected cavity | 0
stenosis of the remaining esophagus | 0
stent removal | 0
endoscopic vacuum therapy | 24
EsoSponge system | 24
jugular and cervical phlegmon resolved | 168
repeated endoscopic balloon dilatation | 168
subtotal esophageal resection | 336
reconstruction using a free-jejunal graft interposition | 336
CT angiography | 336
partial sternotomy | 336
laparotomy | 336
jejunal segment harvested | 336
left carotid artery and left jugular vein used as recipient vessels | 336
graft implanted in an isoperistaltic position | 336
cervical anastomosis performed in an end-to-end fashion | 336
upper mediastinal gastro-jejunostomy performed in a side-to-side fashion | 336
upper sternum resected | 336
soft tissue defect covered with a sternocleidomastoid muscle flap | 336
abdominal reconstruction achieved by an end-to-end jejunojejunostomy | 336
postoperative course uneventful | 408
oral alimentation reestablished | 408
daily speech therapy | 408
anastomotic healing confirmed radiologically and endoscopically | 408
transferred to a rehabilitation clinic | 408
arterial hypertonus | -10080
non-active smoking status | -10080
ischemic stroke with incomplete senso-motoric hemiparesis | -10080
thyroidectomy | -10080
open prostatectomy due to prostate cancer | -10080
family history not related to present illness | 0
percutaneous jejunal feeding catheter inserted | 24
stent slippage | 48
stent position corrected | 48
stent dislocated again | 72
endoscopic management switched to EVT | 72
EVT performed | 96
fistula cavity cleaned | 120
cervical phlegmon resolved | 168
esophageal stenosis resolved | 168
salvage surgery planned | 168
esophageal reconstruction | 336
free jejunal graft interposition | 336
esophago-jejunostomy performed | 336
jejuno-gastrostomy performed | 336