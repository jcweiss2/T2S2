33 years old | 0
female | 0
abnormal uterine bleeding | -120
endometrial ablation | -720
dysuria | -72
grayish, malodorous vaginal discharge | -72
prescribed levofloxacin | -72
syncopal events | -72
admitted to the hospital | 0
blood pressure 74/24 mmHg | 0
afebrile | 0
no rash | 0
extremities were cool | 0
obesity | 0
abdominal exam benign | 0
pelvic examination normal | 0
urine β-human chorionic gonadotropin negative | 0
white blood cell count 60 × 10^3 cells/mm^3 | 0
hematocrit 42% | 0
platelets 38 × 10^3 cells/mm^3 | 0
lactate 6.5 mmol/L | 0
ascites | 0
pelvic ultrasound unremarkable | 0
empiric antibiotic therapy with vancomycin, cefepime, and metronidazole | 0
transferred to the intensive care unit | 0
white blood cell count 113 × 10^3 cells/mm^3 | 12
hematocrit 58% | 12
lactate 13.5 mmol/L | 12
tobramycin, clindamycin, and doxycycline added | 12
vasopressor support | 12
massive IV fluid resuscitation | 12
signs of disseminated intravascular coagulation | 12
received 46 units of blood product | 72
transthoracic echocardiogram showed large pericardial effusion | 24
cardiac tamponade | 24
pericardial drain placement | 24
bilateral pleural effusions | 24
bilateral chest tube placement | 24
exploratory laparotomy | 48
massive ascites | 48
uterus hyperemic | 48
vaginal swabs negative | 48
cervical swabs negative | 48
blood smear showed marked neutrophilia | 48
bone marrow biopsy negative | 48
human immunodeficiency virus-1 antibody negative | 48
blood, urine, pleural fluid, pericardial fluid, peritoneal fluid, and sputum cultures negative | 48
profound anasarca | 72
empiric plasmapheresis | 72
improvement in hemodynamics | 72
fluid removed with continuous venovenous hemofiltration | 72
edema improved | 96
pupils fixed and dilated | 96
CT head scan showed diffuse cerebral edema | 96
tonsillar herniation | 96
life support withdrawn | 96
died | 96
autopsy demonstrated diffuse edema | 120
evidence of DIC in all organs | 120
diffuse endometrial necrosis | 120
Clostridium bifermentans in endometrial tissue | 120