60 years old | 0
male | 0
admitted to the hospital | 0
biopsy proven PAN | -8760
on prednisone | -8760
on cyclophosphamide | -8760
prior failure on cyclophosphamide alone | -8760
paroxysmal atrial fibrillation | 0
hypertension | 0
not on calcium channels blocker | 0
dyslipidemia | 0
non-insulin dependent diabetes mellitus | 0
multiple prior admissions for PAN flares | -8760
history of an admission for septic shock | -17520
scrotal pain | 0
fever of 103°F | 0
fatigue | 0
tachycardic to 130 beats per minute | 0
hypotensive to 103/40 mm Hg | 0
broad-spectrum antibiotics | 0
vancomycin | 0
Zosyn (piperacillin/tazobactam) | 0
kidney function worsened | 24
switch in antibiotics to meropenem | 24
creatinine level continued to rise | 48
suspicion of acute interstitial nephritis less likely | 48
continued to spike fevers | 48
no specific source of an infection found | 48
no focus found on the CT chest, abdomen, and pelvis | 48
stopping all antibiotics | 48
macular rash | 168
rash progressed slowly | 168
involved axillary area | 168
involved chest, head, neck, and abdomen | 168
decline of mental status | 168
worsening of skin lesions | 168
element of bullae and vesicles | 168
dermatology team involved | 216
biopsy obtained | 216
initiating local steroid cream | 216
diagnosis of AGEP | 216
kidney injury | 216
neutrophilia | 216
cyclic fevers | 216
rash became pustular | 264
high grade fever of 109°F | 264
transfer to the intensive care unit | 264
protocol of cooling | 264
pulse steroids | 264
fever subsided | 312
improvement of the initial rash | 312
decreased progression of sloughing | 312
complete resolution of acute kidney injury | 312
taper in steroids | 312
skin biopsy | 0
urine analysis | 0
CT chest/abdomen/pelvis | 0
CBC/BMP/coagulation | 0
differential diagnosis | 0
Generalized acute pustular psoriasis (von Zumbusch type) | 0
Acute generalized exanthematous pustulosis (AGEP) | 0
Drug reaction with eosinophilia and systemic manifestation (DRESS) | 0
Steven Johnson syndrome | 0
Leukocytoclastic vasculitis | 0
Subcorneal pustular dermatosis (Sneddon–Wilkinson disease) | 0
Cutaneous candidiasis | 0
intra- and subcorneal spongiform | 216
superficial, interstitial, mid-dermal infiltrate rich in neutrophils | 216
dermal edema | 216
discharged | 720