55 years old | 0
male | 0
admitted to the hospital | 0
dyspnea | -720
dry cough | -720
joint pain | -720
bilateral distribution in the fingers | -720
hands | -720
wrists | -720
elbows | -720
shoulders | -720
hips | -720
knees | -720
ankles | -720
ibuprofen | -384
oxycodone-acetaminophen | -384
methylprednisolone | -384
joint pain worsened | -720
developed dyspnea | -720
negative SARS-CoV-2 tests | -24
presented to emergency department | -24
shortness of breath with exertion | -24
joint pain | -24
dry cough | -24
unintentional weight loss | -24
denied fever | -24
denied headache | -24
denied sore throat | -24
denied chest pain | -24
denied hemoptysis | -24
denied gastrointestinal symptoms | -24
denied calf swelling | -24
denied calf pain | -24
former smoker | -24000
no recent travel | 0
no sick contacts | 0
no exposure to toxic fume | 0
received Moderna SARS-CoV-2 vaccine | -720
blood pressure 98/63 mm Hg | 0
heart rate 93 beats/min | 0
respirations 18/min | 0
temperature 36.8 °C | 0
oxygen saturation 93% | 0
placed on 2 L oxygen | 0
oxygen saturation 98% | 0
bibasilar rales | 0
tenderness | 0
swelling of the fingers | 0
hands | 0
wrists | 0
elbows | 0
shoulders | 0
hips | 0
knees | 0
ankles | 0
erythematous papules on dorsum of left hand | 0
erythematous macules on fingers of left hand | 0
left elbow | 0
left knee | 0
no muscle tenderness | 0
D-dimer 1,702 ng/mL | 0
aspartate aminotransferase 86 U/L | 0
alanine aminotransferase 65 U/L | 0
CRP 3.70 mg/dL | 0
ESR 52 mm/h |7 0
normal complete blood count | 0
normal electrolytes | 0
normal total creatinine kinase | 0
normal procalcitonin | 0
negative blood cultures | 0
negative sputum cultures | 0
negative respiratory pathogen panel | 0
chest X-ray patchy atelectatic changes | 0
CTPA negative for pulmonary embolism | 0
nonspecific patchy atelectasis | 0
increased interstitial markings | 0
admitted to hospital | 0
rheumatology consult | 0
pulmonology consult | 0
infectious workup | 0
rheumatologic workup | 0
treated for community acquired pneumonia | 72
treated for autoimmune inflammatory arthropathy | 72
ILD | 72
azithromycin | 72
ceftriaxone | 72
fluticasone-vilanterol inhaler | 72
tiotropium bromide | 72
prednisone | 72
transitioned to cefuroxime | 144
prednisone 40 mg | 144
discharged | 144
followed up with rheumatology | 168
diagnosed CADM | 168
ILD | 168
anti-MDA5 antibody titers 72 | 168
started mycophenolate mofetil | 168
prednisone 60 mg | 168
follow-up pulmonology | 168
normal 6-min walk test | 168
PFT consistent with mild asthma | 168
diagnosed asthma | 168
mild ILD | 168
started fluticasone-salmeterol | 168
tiotropium bromide | 168
prescription for repeat chest X-ray | 168
new cough | 840
foamy sputum production | 840
bronchoscopy | 840
BAL | 840
transbronchial biopsy | 840
fever 40.3 °C | 840
readmitted | 840
concern for infection | 840
blood cultures | 840
sputum cultures | 840
(1,3)-beta-D-glucan | 840
BAL studies | 840
started vancomycin | 840
piperacillin-tazobactam | 840
sulfamethoxazole/trimethoprim | 840
methylprednisone | 840
high resolution CT scan | 840
traction bronchiectasis | 840
worsening bilateral infiltrates | 840
ground glass opacities | 840
septal thickening | 840
clinical status deteriorated | 840
increasing oxygen requirements | 840
hypoxia | 840
oxygen saturation 82-95% | 840
transbronchial biopsy normal | 840
BAL positive for Pneumocystis jirovecii | 840
diagnosed PCP | 840
transferred to ICU | 840
trimethoprim-sulfamethoxazole IV | 840
plasma exchange therapy | 840
hypoxia worsened | 840
bilevel positive airway pressure | 840
intubation | 840
pneumothorax | 840
pneumomediastinum | 840
cardiothoracic surgery consult | 840
no chest tube placement | 840
ventilator support | 840
norepinephrine | 840
PEA arrest | 840
death | 840
