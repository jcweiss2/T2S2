59 years old | 0
male | 0
presented with gross hematuria | 0
gross hematuria | 0
heavy smoker | 0
lower urinary tract symptoms | -26280
α1 blocker medication | -26280
mild pale | 0
blood pressure 120/60 mm/Hg | 0
pulse 70 | 0
mild tenderness in lower abdominal region | 0
hemoglobin 9 g/dl |8
white blood cell count 13 × 10^9/l | 0
platelet count 390 × 10^9/l | 0
normal creatinine | 0
normal urea | 0
normal electrolytes | 0
excess RBC/HPF | 0
30_50 WBC/HPF | 0
4–5 epithelial cells/HPF | 0
ultrasound showing grade 3 right renal hydronephrosis | 0
simple cyst (right renal) | 0
simple cyst (left renal) | 0
bladder diverticulum (right bladder wall) | 0
mass in bladder diverticulum | 0
CT confirmation of bladder diverticulum with mass | 0
cystoscopy | 24
enlarged prostate | 24
severe bladder trabeculation | 24
TUR-BT not feasible | 24
TUR-P performed | 24
partial cystectomy | 168
free visible margins | 168
para-aortic lymph node dissection | 168
foley catheter insertion | 168
transitional cell carcinoma (high grade) PT3 | 168
lymph nodes involvement | 168
cardiac arrhythmia | 168
right pleural effusion | 168
sepsis | 240
passed away | 240
