56 years old| 0
    man| 0
    diagnosed with nodular sclerosing CD30+ HL| -8640
    CD15+ HL| -8640
    stage IV disease| -8640
    diffuse involvement of lymph nodes| -8640
    bone marrow involvement| -8640
    liver involvement| -8640
    power-injectable port inserted| -8640
    six cycles of ABVD chemotherapy initiated| -8640
    adriamycin| -8640
    bleomycin| -8640
    vinblastine| -8640
    dacarbazine| -8640
    partial response achieved| -8640
    two other lines of chemotherapy| -8640
    poor clinical response| -8640
    evaluated for autologous HSCT| -8640
    pretransplant TTE revealed RA mass| -24
    2.2 × 1.8 cm RA mass| -24
    normal cardiac function| -24
    sent to emergency room| 0
    hemodynamically stable| 0
    asymptomatic| 0
    unremarkable physical examination| 0
    leukocytosis of 15,000 cells/mm3| 0
    hemoglobin of 7.5 mg/dL| 0
    normal platelet count| 0
    CT imaging showed RA mass| 0
    unclear etiology| 0
    extra-cardiac findings consistent with diffuse HL| 0
    TEE showed RA mass attached to posterior atrial wall| 0
    RA mass attached to CVC at SVC/RA junction| 0
    question of differentiating metastatic lesion vs thrombus| 0
    CMR obtained| 0
    no enhancement of RA mass with gadolinium| 0
    diagnosis of CRAT confirmed| 0
    started on heparin| 0
    anticoagulation initiated| 0
    cardiac thoracic surgery consulted| 0
    possible thrombectomy| 0
    developed fever| 0
    hypotension| 0
    pancytopenia| 0
    managed in ICU| 0
    broad spectrum antibiotics| 0
    vasopressors| 0
    rapid deterioration| 0
    succumbed to disease| 0
    <|eot_id|>