59 years old | 0
female | 0
laparoscopic adjustable band insertion | -7920
central abdominal pain | -336
abdominal distention | -336
nausea | -336
vomiting | -336
denied dysphagia | -336
denied odynophagia | -336
denied change in bowel habit | -336
afebrile | -336
tachycardic | -336
diffuse abdominal tenderness | -336
guarding | -336
inflammatory markers mildly elevated | -336
white cell count 13.7 × 10^9/L | -336
C-reactive protein 105 mg/L | -336
moderate hyperlactatemia | -336
lactate 2.4 mmol/L | -336
distended, air-filled stomach | -336
intragastric band erosion | -336
internalization of the entire gastric band and distal connector tubing within the gastric lumen | -336
moderate free fluid | -336
ascites | -336
mesenteric inflammatory fat stranding | -336
portal vein non-opacified | -336
possible portal vein thrombosis | -336
exploratory laparotomy | 0
ischemic small bowel segment resected | 0
engorged mesentery | 0
blood clots extruding out of the mesenteric vascular arcade | 0
on-table OGD | 0
deformed shaped stomach | 0
gastric band completely eroded through the wall of the stomach | 0
biofilm formed around the band device | 0
biofilm tracked to the stomach externally | 0
stomach opened | 0
device retrieved | 0
stomach closed in two layers | 0
abdominal drains inserted | 0
monitored in the intensive care unit | 0
focused hepatic ultrasound | 24
portal vein almost completely thrombosed | 24
commenced on therapeutic dose of tinzaparin sodium | 24
intensive gastroenterology input | 24
dietician input | 24
physiotherapy input | 24
hematology input | 24
barium meal | 504
normal gastric contours | 504
no filling defects | 504
no gastric outlet emptying | 504
discharged | 504