78 years old|0
woman|0
revised left total hip arthroplasty|0
presented to the emergency department|-504
abdominal pain|-504
hypotension|-504
placement of an antiprotrusio cage|-504
initial left total hip arthroplasty in 1998|-141120
osteoarthritis|-141120
progressive left hip pain|-141120
protrusio of the acetabular component|-141120
central bone weakening|-141120
revision of the left total hip arthroplasty|-141120
acetabuloplasty|-141120
medial acetabular bone grafting|-141120
placement of a unipolar hemiarthroplasty|-141120
left hip pain|-141120
radiographs showed progressive superomedial migration of the unipolar head|-141120
antiprotrusio cage placed|-141120
cervical squamous-cell carcinoma (stage IB; limited to the cervix)|0
treated with total hysterectomy in 1993|-217680
lymphoma treated with chemotherapy|0
splenectomy|0
not received pelvic irradiation|0
not on immunosuppressive medications (including steroids)|0
presented to the emergency department with abdominal pain|0
hypotensive|0
leukocytosis|0
pyuria|0
no symptoms of increased left hip pain|0
no edema|0
no erythema surrounding the left hip|0
CT scan of the abdomen and pelvis showed small bowel dilatation|0
severe left hip protrusio|0
medial migration of the acetabular hardware|0
hardware penetration of the sigmoid colon wall|0
large amount of fluid and gas surrounding the left hip and greater trochanter|0
sigmoid colon perforation|0
fistula to the left hip joint|0
fistula to periarticular soft tissues|0
CT-guided aspiration of the fluid collection lateral to the left greater trochanter|0
fecal material|0
culture grew Escherichia coli|0
culture grew Streptococcus viridans|0
culture grew Clostridium perfringens|0
surgery revealed 1-cm titanium flange of the acetabular cage perforating the sigmoid colon|0
proximal small bowel dilatation due to ileus|0
no findings of diverticulitis|0
bowel normally positioned|0
sigmoidectomy|0
Hartmann procedure|0
end-sigmoid colostomy|0
omental coverage of the hardware|0
lateral incision over the left hip|0
large pockets of brown fluid in the subcutaneous tissues|0
involved vastus lateralis muscle|0
involved left hip|0
debridement performed|0
cultures from the left hip grew Escherichia coli|0
cultures from the left hip grew Streptococcus viridans|0
cultures from the left hip grew Clostridium perfringens|0
removal of hardware initially not attempted due to risk of injury|0
seven left hip joint irrigations/debridements|336
hip disarticulation|336
femoral hardware removal|336
partial acetabular hardware removal|336
emergent femoral-femoral arterial bypass|336
left-lower-extremity ischemia|336
two-month hospitalization|1440
septicemia|0
two-week course in the intensive care unit|336
readmitted two weeks following initial discharge|720
gastrointestinal bleeding|720
infected left pelvic hematoma|720
osteomyelitis of the proximal left femur|720
decompression of the hematoma|720
serial irrigation and debridements of the left hip|720
removal of remaining acetabulum hardware (cemented cup, cage, four screws)|720
exacerbation of congestive heart failure|720
aspiration|720
became hypotensive|2160
died during her second hospitalization|2160
