69 years old | 0
male | 0
prostate cancer (cT4N0M1b) | -1008
chemotherapy | -1008
prednisolone 10 mg per day | -1008
proton pump inhibitor | -1008
Cabazitaxel Acetonate every two months | -1008
fever | -20
altered consciousness | 0
transferred to the hospital | 0
Glasgow Coma Scale E3V3M5 | 0
temperature 40.6 °C | 0
blood pressure 142/80 mmHg | 0
pulse rate 126/min | 0
respiratory rate 30/min | 0
SpO2 98 % | 0
pale conjunctive | 0
no icterus | 0
no abnormal chest findings | 0
median surgical scar | 0
no other remarkable abdominal findings | 0
mildly edematous lower extremities | 0
no palpable lymph nodes | 0
no rash | 0
no neck stiffness | 0
elevated white blood cell count | 0
anemia | 0
cytoplasmic vacuolation of white blood cells | 0
anisocytosis | 0
spherocytes | 0
high lactate dehydrogenase | 0
high creatine kinase | 0
severe hemolysis on first specimen | 0
severe hemolysis on re-drawn sample | 0
severe hemolysis six hours after arrival | 6
anemia progression | 6
hemolysis progression | 6
DIC progression | 6
plain chest X-ray no abnormalities | 0
chest CT no abscess | 0
abdominal CT no abscess | 0
sepsis treatment initiated | 0
blood cultures obtained | 0
sputum cultures obtained | 0
urinary cultures obtained | 0
piperacillin/tazobactam administered | 0
blood pressure drop two hours after arrival | 2
cardiopulmonary arrest | 2
cardiopulmonary resuscitation | 2
circulation recovered | 2
blood cell transfusion | 2
vasopressors initiated | 2
hypothermia treatment initiated | 2
worsening hemolysis | 2
difficulty maintaining blood pressure | 2
death | 30
Clostridium perfringens detected in blood cultures | 30
Gram-positive bacilli identified | 30
bacilli phagocytized by white blood cells | 30
serotype TW62 | 30
non-enterotoxin producing | 30
α toxin-producing type A | 30
susceptible to penicillins | 30
susceptible to β-lactams | 30
no postmortem examination | 30
