62 years old | 0
male | 0
prediabetes | 0
heavy smoker | 0
admitted with central chest pain | 0
ECG performed | 0
no ST elevation | 0
well perfused | 0
normotensive | 0
sinus rhythm | 0
chest auscultation | 0
normal heart sounds | 0
no added sounds | 0
no murmurs | 0
clear chest | 0
no arm claudication | 0
good pulses in both upper limbs | 0
normal full blood count | 0
raised fibrinogen | 0
raised troponin T | 0
raised brain natriuretic peptide | 0
coronary angiogram performed | 0
significant left main coronary artery disease | 0
three-vessel disease | 0
patent right brachiocephalic artery | 0
echocardiogram | 0
left ventricular ejection fraction 30% | 0
hypokinesia in inferior segments | 0
hypokinesia in anterior segments | 0
carotid arteries not imaged | 0
became unstable during anaesthetic induction | 0
ST-elevation | 0
urgent initiation of surgery | 0
surgical revascularization | 0
LIMA to LAD | 0
SVG to intermediate | 0
SVG to posterior descending artery | 0
off cardiopulmonary bypass easily | 0
minimal inotropic support | 0
stable echocardiographic appearances | 0
graft assessment | 0
patent grafts | 0
satisfactory diastolic Doppler flows | 0
developed mixed cardiogenic shock | 48
developed distributive shock | 48
intra-aortic balloon pump | 48
high doses of inotropes | 48
echocardiographic assessment | 48
no new regional wall motion abnormalities | 48
no dynamic ECG changes | 48
downward troponin trend | 48
inotropic support weaned | 168
IABP weaned | 168
deteriorated after becoming septic | 168
inotropic support restarted | 168
adrenaline | 168
noradrenaline | 168
milrinone | 168
empiric antibiotic coverage initiated | 168
meropenem | 168
repeat echocardiogram | 168
profound hypokinesia in mid-distal LAD territory | 168
no dynamic ECG changes | 168
down-trending troponin values | 168
deteriorating echocardiographic picture | 168
stunned anterior wall myocardium | 168
transferred to catheterization laboratory | 168
chronic total occlusion of left subclavian artery | 168
patent SVGs | 168
LIMA retrograde filling | 168
peak systolic gradient 60 mmHg | 168
PCI performed | 168
sirolimus-eluting stent implanted | 168
paclitaxel-eluting balloon inflation | 168
comprehensive invasive functional assessment | 168
FFR measured | 168
AF measured | 168
positive FFR | 168
AF increased by 14% | 168
LIMA occluded with coils | 168
Micro Vascular Plug implanted | 168
complete occlusion of LIMA | 168
improved significantly | 168
weaned from inotropic support | 168
weaned from ventilator | 168
discharged to ward | 168
minimal motor function impact | 168
discharged home | 720
good functional status | 720
EF 40% | 4320
hypokinesia of inferior wall | 4320
normalization of anterior wall contractility | 4320
