59 years old | 0
male | 0
acute disseminated encephalomyelitis (ADEM) | -1032
severe COVID-19 | -1032
encephalopathy | -1032
generalized motor weakness | -1032
multifocal magnetic resonance (MR) imaging findings | -1032
septic shock | -1032
inotropic support | -1032
acute kidney injury | -1032
haemodialysis | -1032
deranged liver function | -1032
provoked segmental pulmonary embolism | -1032
polyarticular gout flare | -1032
polyarticular gout | -1032
transferred out of intensive care | -1032
minimal neurological recovery | -1032
Glasgow Coma Scale (GCS) score of E4VTM1 | -1032
no consistent visual pursuit | -1032
no vocalizations | -1032
no functional communication | -1032
encephalopathy improved | -1032
Coma Recovery Scale-Revised (CRS-R) score 9/23 | -1032
followed instructions inconsistently | -1032
CRS-R score 10/23 | -1032
axonal sensorimotor polyneuropathy | -1032
critical illness polyneuropathy | -1032
transferred to inpatient rehabilitation facility | 0
GCS of E4V4M6 | 0
physiatrist-led transdisciplinary rehabilitation programme | 0
rehabilitation therapies | 0
physiotherapy | 0
occupational therapy | 0
speech therapy | 0
psychology reviews | 0
fortnightly dietician reviews | 0
weekly multidisciplinary conferences | 0
Functional Independence Measure (FIM) | 0
cognitive deficits | 0
sustained attention for 10–15 minutes | 0
disoriented | 0
slow information processing speed | 0
followed one-step commands | 0
impaired immediate information recall | 0
Abbreviated Mental Test (AMT) score 1/10 | 0
participation limited | 0
attentional deficits | 0
impaired short-term memory | 0
therapy in quiet environment | 0
coaxing required | 0
task simplification | 0
increased time for information processing | 0
irritability | 0
agitation | 0
time-out-on-the-spot techniques | 0
redirection | 0
unable to use cognitive remediation strategies | 0
daily reality orientation | 0
flexibility of therapy timings | 0
sleep wake regulation | 0
AMT improved to 3/10 | 0
quadriparesis | 0
spastic weakness in lower limbs | 0
Medical Research Council (MRC) grade 2/5 (left) | 0
MRC grade 1/5 (right) | 0
upper limbs MRC scale 3/5 | 0
periventricular lesions | 0
motor recovery complicated by CIP and steroid myopathy | 0
dependent in bed mobility | 0
poor sitting balance | 0
maximum assistance for ADLs | 0
sitting balance training | 0
sitting tolerance training | 0
verticalisation via tilt table | 0
task-specific training for ADLs | 0
mirror visual feedback | 0
orthostatic hypotension | 0
blood pressure drop from 135/92 mmHg to 112/87 mmHg | 0
scheduled fluid intake | 0
fluid boluses before therapy | 0
elastic compression stockings | 0
abdominal binders | 0
tolerated sitting at edge of bed | 0
mobilised in tilt-in-space wheelchair | 0
mild oropharyngeal dysphagia | 0
nasogastric tube feeding cessation | 0
blended diet | 0
video fluoroscopic swallowing study | 0
no aspiration | 0
normal diet | 0
functional communicative ability | 0
expressive speech | 0
receptive speech | 0
weight loss | 0
BMI 21.6 kg/m² | 0
nadir albumin level 24 g/L | 0
albumin improved to 30 g/L | 0
high caloric diet | 0
oral nutritional supplements | 0
nadir anaemia 6.3 mg/L | 0
anaemia improved to 10.2 mg/L | 0
immobilisation-related hypercalcemia | 0
hypercalcemia normalised | 0
decubitus ulcer | 0
Grade 3 sacral ulcer | 0
limited mobilisation efforts | 0
contraindicated Lokomat® | 0
bed-turning | 0
pressure relief mattresses | 0
pressure offloading | 0
sitting duration increased | 0
wound healing | 0
urinary incontinence | 0
indwelling urinary catheter | 0
spontaneous voiding | 0
dependent on diapers | 0
catheter-associated urinary tract infections | 0
Clostridium difficile diarrhoea | 0
recurrent polyarticular gout flares | 0
left hip aspiration | 0
right knee aspiration | 0
turbid straw-colored fluid | 0
negatively birefringent crystals | 0
no septic arthritis | 0
oral prednisolone | 0
febuxostat | 0
serum uric acid decreased from 903 µM/L to 483 µM/L | 0
gentle joint mobilisation | 0
acute lower body pain | 0
chronic lower body pain | 0
impaired sensory discrimination | 0
multifactorial pain | 0
acute pain flares | 0
chronic pain | 0
joint stiffness | 0
axonal sensorimotor polyneuropathy (CIP) | 0
central neuropathic pain | 0
spinal-thalamic-cortical pathway dysfunction | 0
adductor spasticity | 0
restricted hip abduction | 0
restricted hip flexion | 0
pain managed by acetaminophen | 0
pain managed by NSAIDs | 0
pain managed by gabapentin | 0
contraindicated physical modalities | 0
FIM scores improvement | 0
diagnostic delays | 0
normal computed tomography on Day 16 | 0
MR imaging on Day 34 | 0
early rehabilitation considerations | 0
decubitus ulcerations | 0
steroid-induced skin atrophy | 0
preventive nursing care | 0
nutrition | 0
neurocognitive sequelae | 0
persistent fatigue | 0
anxiety | 0
depression | 0
delayed neuroplastic mechanisms | 0
indeterminate prognosis | 0
chronic impairments | 0
hampered societal participation | 0
vocational cessation | 0
rehabilitation recommendations | 0
family engagement | 0
videoconferencing | 0
digital communication | 0
multiple organ dysfunction | 0
psychological interventions | 0
long-term morbidity | 0
physical disability | 0
cognitive disability | 0
long-term healthcare costs | 0
socioeconomic burden | 0
long COVID-19 | 0
intravenous immunoglobulin on Day 43 | -1032
intravenous immunoglobulin on Day 67 | -1032
intravenous immunoglobulin on Day 95 | -1032
intravenous immunoglobulin on Day 146 | -1032
nerve conduction study on Day 89 | -1032
transfer to ICU | -1032
intensive care unit (ICU) stay | -1032
FIM scores on Day 186 | 0
FIM scores on Day 223 | 0
FIM scores on Day 277 | 0
right knee and left hip aspiration | 0
Day 46 aspiration | -1032
Day 174 aspiration | -1032
Day 258 AMT improvement | 0
Day 258 wound healing | 0
Day 266 mobilisation | 0
Day 70 CRS-R score 9/23 | -1032
Day 72 follow instructions | -1032
Day 83 CRS-R score 10/23 | -1032
Day 108 nadir albumin | -1032
Day 53 hypercalcemia | -1032
Day 133 decubitus ulcer | -1032
Day 186 transfer to rehabilitation | 0
Day 189 swallowing study | 0
Day 258 events | 0
eight months into admission | 0
peak uric acid 903 µM/L | -1032
current uric acid 483 µM/L | 0
initial FIM score 26 | 0
FIM score 29 | 0
FIM score 34 | 0
motor sub-scores | 0
cognitive sub-scores | 0
self-care improvement | 0
sphincter control | 0
locomotion | 0
transfers | 0
communication improvement | 0
social cognition improvement | 0
no specific rehabilitation service | 0
detailed functional assessment | 0
family engagement challenges | 0
cross-border restrictions | 0
holistic rehabilitation approach | 0
long-term complications | 0
nil financial support | 0
no conflicts of interest | 0
