29 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
cardiogenic shock | -720 | -720 | Factual
biventricular failure | -720 | -720 | Factual
ejection fraction 5-10% | -720 | -720 | Factual
myopericarditis | -720 | -720 | Factual
constrictive physiology | -720 | -720 | Factual
PICC line placed | -720 | -720 | Factual
discharged on milrinone | -720 | -720 | Factual
fever | -24 | 0 | Factual
chills | -24 | 0 | Factual
septic shock | 0 | 0 | Factual
PICC line removed | 0 | 0 | Factual
IV vancomycin | 0 | 24 | Factual
piperacillin/tazobactam | 0 | 24 | Factual
vasopressor support | 0 | 24 | Factual
Chryseobacterium indologenes | 48 | 48 | Factual
ciprofloxacin | 48 | 336 | Factual
piperacillin/tazobactam | 48 | 336 | Factual
weaned off vasopressor support | 48 | 48 | Factual
pericardiectomy | 168 | 168 | Factual
discharged | 336 | 336 | Factual
inotrope independent | 336 | 336 | Factual
follow-up | 744 | 744 | Factual
no evidence of recurrent infection | 744 | 744 | Factual
NYHA Class I | 744 | 744 | Factual
improved functional status | 744 | 744 | Factual
furosemide | 0 | 744 | Factual
metoprolol succinate | 0 | 744 | Factual
sacubitril-valsartan | 336 | 744 | Factual
cardiomegaly | -720 | -720 | Factual
dilated right atrium | -720 | -720 | Factual
passive hepatic congestion | -720 | -720 | Factual
right ventricular failure | -720 | -720 | Factual
pericardial calcification | -720 | -720 | Factual
biventricular failure | -720 | -720 | Factual
constrictive pericarditis | -720 | -720 | Factual
left ventricular ejection fraction 23% | -720 | -720 | Factual
right ventricular ejection fraction 36% | -720 | -720 | Factual
delayed gadolinium enhancement | -720 | -720 | Factual
diastolic septal bounce | -720 | -720 | Factual
concentrically thickened pericardium | -720 | -720 | Factual
atrial flutter | -720 | -720 | Factual
rapid ventricular response | -720 | -720 | Factual
radiofrequency ablation | -720 | -720 | Factual
inotrope therapy | -720 | 0 | Factual
home milrinone infusion | -720 | 0 | Factual
elective pericardiectomy | -24 | -24 | Factual
fever 38.7°C | -24 | 0 | Factual
tachycardia | -24 | 0 | Factual
hypotension | 0 | 0 | Factual
elevated lactate level | 0 | 0 | Factual
severe rigours | 0 | 0 | Factual
blood cultures | 0 | 0 | Factual
Gram-negative rods | 48 | 48 | Factual
Chryseobacterium indologenes | 48 | 48 | Factual
ciprofloxacin | 48 | 336 | Factual
piperacillin/tazobactam | 48 | 336 | Factual
susceptibility testing | 48 | 48 | Factual
sensitive to ciprofloxacin | 48 | 48 | Factual
sensitive to piperacillin | 48 | 48 | Factual
sensitive to trimethoprim/sulfamethoxazole | 48 | 48 | Factual
resistant to meropenem | 48 | 48 | Factual
improved clinically | 48 | 336 | Factual
afebrile | 48 | 336 | Factual
weaned off vasopressor support | 48 | 48 | Factual
negative blood cultures | 48 | 336 | Factual
interval echocardiogram | 168 | 168 | Factual
left ventricular EF 50-55% | 168 | 168 | Factual
right ventricular systolic dysfunction | 168 | 168 | Factual
pericardiectomy | 168 | 168 | Factual
dense areas of adhesions | 168 | 168 | Factual
calcium | 168 | 168 | Factual
complete removal of pericardium | 168 | 168 | Factual
follow-up transthoracic echocardiogram | 336 | 336 | Factual
left ventricular EF 50-55% | 336 | 336 | Factual
right ventricular systolic dysfunction | 336 | 336 | Factual
discharged | 336 | 336 | Factual
inotrope independent | 336 | 336 | Factual
guideline-directed medical therapy | 336 | 744 | Factual
furosemide | 336 | 744 | Factual
metoprolol succinate | 336 | 744 | Factual
sacubitril-valsartan | 336 | 744 | Factual
follow-up | 744 | 744 | Factual
no evidence of recurrent infection | 744 | 744 | Factual
NYHA Class I | 744 | 744 | Factual
improved functional status | 744 | 744 | Factual