60 years old | 0
male | 0
admitted to the hospital | 0
fever | -24
working on farms | -672
close contact with swine | -672
stable vital signs | 0
no defining abnormal findings | 0
no specific findings in laboratory data | 0
no specific findings in urinalysis | 0
no active lung lesion | 0
mild gas accumulation | 0
discharged from the hospital | 24
revisited the emergency department | 24
persistent fever | 24
dizziness | 24
vomiting | 24
acutely ill | 24
drowsy | 24
low blood pressure | 24
low heart rate | 24
respiratory rate | 24
low body temperature | 24
clear lung sounds | 24
decreased bowel sounds | 24
leukopenia | 24
thrombocytopenia | 24
higher urea nitrogen | 24
higher creatinine | 24
hyperbilirubinemia | 24
metabolic acidosis | 24
meropenem administration | 24
vancomycin administration | 24
admitted to the intensive care unit | 24
vital signs at 6 hours of admission | 6
inotropics administration | 6
corticosteroid administration | 6
generalized tonic-clonic seizure | 14
low peripheral oxygen saturation | 14
endotracheal intubation | 14
mechanical ventilator application | 14
peripheral oxygen saturation at 16 hours of admission | 16
zero urine output | 16
continuous renal replacement therapy | 16
bacterial growth in blood cultures | 12
gram-positive cocci in blood cultures | 48
S. suis identification | 96
antibiotic susceptibility testing | 96
vancomycin and meropenem replacement with ampicillin/sulbactam | 96
vital signs stabilization | 96
dopamine and norepinephrine tapering | 96
hydrocortisone change to dexamethasone | 96
ventilator weaning and extubation | 168
continuous renal replacement therapy stop | 168
mental status improvement | 168
difficulty in hearing | 168
otoscopic examination | 168
tuning fork examination | 168
bilateral sensorineural hearing loss | 168
spinal tap | 168
cerebrospinal fluid analysis | 168
dexamethasone treatment continuation | 168
back pain | 240
magnetic resonance imaging of the lumbar spine | 240
infective spondylitis | 240
intramuscular abscess formation | 240
medical treatment continuation | 240
transfer to another hospital | 240
prolonged antibiotic treatment | 240
back pain improvement | 432
hearing difficulty persistence | 8760