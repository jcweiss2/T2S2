30 years old | 0
male | 0
Saethre-Chotzen syndrome | 0
admitted to the hospital | 0
shortness of breath | 0
abdominal pain | 0
nausea | 0
vomiting | 0
prior history of open surgical pulmonic valvotomy | -6720
prior history of pulmonary outflow homograft patch | -6720
gastric bypass for morbid obesity | -6720
recent treatment for bilateral lower extremity swelling | -168
antibiotics | -168
steroids | -168
admission BMI | 0
HR of 90 | 0
BP of 140/80 | 0
RR 27 breaths per minute | 0
Pulse Oximetry of 92% | 0
initiated on antibiotics | 0
nasal cannula oxygen | 0
intravenous fluids | 0
low lung volumes on chest x-ray | 0
acute left lower extremity superficial thrombophlebitis | 0
no evidence of acute pulmonary embolism | 0
cardiomegaly | 0
central pulmonary artery enlargement | 0
cholelithiasis | 0
nephrolithiasis | 0
left intrarenal calculus | 0
wedge-shaped infarct in the lower pole of the right kidney | 0
small cerebellar infarct | 0
transferred to the intensive care unit | 24
non-invasive ventilation with BiPAP | 24
intubated and placed on mechanical ventilation | 168
lung protective ventilation | 168
high PEEP strategy | 168
norepinephrine | 168
vasopressin | 168
failure of mechanical ventilation to improve hypoxemic respiratory failure | 168
initiation of veno-venous extracorporeal membrane oxygenation | 168
inhaled nitric oxide therapy | 192
transesophageal echocardiogram | 216
large intra-atrial bidirectional shunt | 216
right-to-left flow during systole | 216
left-to-right flow during diastole | 216
severe pulmonary regurgitation | 216
enlarged pulmonary artery | 216
absent left main and separate ostial connections of the left anterior descending and left circumflex coronary arteries | 216
bronchoscopy | 240
significant secretions in the right bronchial lower lobe | 240
influenza B | 240
pulmonary artery catheter | 240
hemodynamic and arterial blood gas profile changes | 240
pulmonary regurgitation and IAS required correction | 240
sepsis | 240
vasopressors | 240
judicious diuresis | 240
vasopressor wean | 240
drop in MAP | 240
increased hypoxemia | 240
CardioSeal patent foramen ovale closure device | 336
oxygen saturation improved | 336
balloon occlusion of the IAS | 336
oxygen saturation improved acutely | 336
30 mm cribriform ASD occluder device | 336
oxygen saturations and arterial oxygen pressure initially decreased | 336
improved modestly subsequent to the procedure | 336
weaned off inhaled nitric oxide | 480
interval echocardiography | 480
residual R-L shunt | 480
continued severe pulmonary regurgitation | 480
tracheostomy | 576
ventilator wean | 576
weaning of PEEP and FiO2 | 576
follow-up CT scans | 720
persistence of left cerebellar vermis infarct | 720
improved interstitial edema of the lung | 720
migration of the CardioSeal device | 720
angiographic removal | 720
mechanical ventilation discontinued | 912
supplemental oxygen delivery via a tracheostomy collar | 912
discharged to an acute rehabilitation unit | 912
primary closure of left atrial septal defect | 4320
pulmonic valve replacement | 4320
pulmonary outflow patch graft reconstruction | 4320
bovine pericardial patch | 4320
porcine heart valve Medtronic Hancock II | 4320
intraoperative pressure and oxygenation measurements | 4320
normal prosthetic pulmonary valve function | 4320
atrial septal defect closed | 4320
negative bubble study | 4320
outpatient cardiology clinic | 4752