8.75 years old | 0
male | 0
neutered | 0
Burmese | 0
5.6 kg | 0
admitted to the hospital | 0
lethargy | -72
anorexia | -72
tachypnoea | -72
restrictive breathing pattern | -72
pyrexia | -72
bright | 0
alert | 0
responsive | 0
respiratory rate 40 breaths/min | 0
mild increase in respiratory effort | 0
heart rate 170 bpm | 0
grade II/VI systolic murmur | 0
rectal temperature 38.1ºC | 0
midazolam administration | 0
butorphanol administration | 0
alfaxalone administration | 0
thoracocentesis | 0
pleural effusion | 0
bupivacaine administration | 0
thoracic drainage | 0
lavage | 0
amoxicillin-clavulanate administration | 0
buprenorphine administration | 0
IV fluid therapy | 0
oxygen therapy | 2
elevated respiratory effort | 12
mydriasis | 36
hypersalivation | 36
tonic–clonic seizure activity | 36
loss of consciousness | 36
stuporous | 36
sinus bradycardia | 36
hypotension | 36
intravenous lipid emulsion administration | 36.33
mentation improvement | 36.5
ambulatory | 36.5
mildly obtunded | 36.5
bradycardic | 36.5
hypersalivation | 36.5
thoracic lavage | 37
intrapleural bupivacaine discontinuation | 37
repeat venous blood gas analysis | 39
acidaemia | 39
hypokalaemia | 39
hyperglycaemia | 39
hyperlactataemia | 39
azotaemia | 39
decline in mental status | 46
relapse bradycardia | 46
repeat intravenous lipid emulsion administration | 46
improved mental status | 46.5
normotensive | 46.5
bradycardia | 46.5
general anaesthesia | 60
CT | 60
right middle lung lobe abscess | 60
median sternotomy | 60
hypotension | 60
noradrenaline CRI | 60
respiratory distress | 60
laryngeal oedema | 60
dexmedetomidine CRI | 60
re-intubation | 60
analgesia tapering | 72
discharged | 144