7 years old | 0
male | 0
admitted to the hospital | 0
high fever | -672
coughing | -672
pain in the legs | -672
dysesthesia | -672
waddling gait | -672
sister had flu-like syndrome | -168
symptomatic treatment | -672
deterioration of general state | -504
abdominal pain | -504
food intolerance | -504
acute respiratory failure | -504
tachycardia | 0
normal blood pressure | 0
respiratory retraction | 0
abdominal breathing | 0
diffuse rhonchi | 0
severe hypoxemia | 0
no hypercapnia | 0
chest X-ray showed bilateral interstitial pneumonia | 0
transferred to pediatric intensive care unit | 0
noninvasive ventilation | 0
chest X-ray control showed right basal consolidation | 24
dribble with probable aspiration | 24
agitation | 48
bilateral mydriasis | 48
intubation | 48
sedation | 48
mechanical ventilation | 48
neurological manifestations progressed to bulbar and peripheral motor deficit | 96
respiratory stabilization | 96
sedation released | 96
no seizures | 96
normal consciousness | 96
inability to speak | 96
communication via eye movements and blinking | 96
no spontaneous movements of arms and legs | 96
facial diplegia | 96
bilateral ptosis | 96
mydriasis without ophthalmoplegia | 96
severe swallowing disorders | 96
absence of cough | 96
tetraparesia predominant on upper limb | 96
brief hyperreflexia | 96
no Babinski reflex | 96
areflexia | 120
dysautonomia not diagnosed | 120
required vascular fillings | 120
hemodynamic stabilization | 120
no hypertension | 120
no heart rate lability | 120
Mycoplasma pneumonia identified | 0
Haemophilus influenza identified | 0
increased C-reactive protein | 0
increased procalcitonin | 0
toxicology studies negative | 0
other microbiological tests normal | 0
immune tests normal | 0
cerebrospinal fluid examinations normal | 0
no oligoclonal bands | 0
nonspecific anti-GM4 detected | 48
negative antiganglioside and antigalactocerebroside antibodies | 624
cerebral tomography scan normal | 48
cerebromedullar magnetic resonances normal | 120
no enhancements of nerve roots | 120
ultrasonography showed phrenic paresia | 504
electroencephalogram normal | 48
sensitive evoked potentials normal | 456
electromyogram decreased amplitude on upper limb | 192
axonal affection confirmed | 432
first course intravenous immunoglobulin | 120
no clinical improvement | 120
second course intravenous immunoglobulin | 504
recovery started | 504
treated with acyclovir | 0
treated with clarithromycin | 0
treated with ceftriaxone | 0
treated with cotrimoxazole | 0
treated with oseltamivir | 0
clarithromycin administered for 21 days | 0
amoxicillin–clavulanate associated for 8 days | 0
mechanical ventilation for 48 days | 0
oxygen requirement decreased | 0
muscle weakness | 0
swallowing troubles | 0
tracheostomy performed | 696
enteral feeding for 18 weeks | 0
gastrostomy | 1320
speech and oral intake improved | 0
intensive rehabilitation started | 0
left the hospital | 1848
proximal weakness | 1848
decreased upper limb deep tendon reflexes | 1848
fluid walking | 1848
no breathing troubles | 1848
no swallowing troubles | 1848
electromyogram control showed improvements | 4368
tracheostomy removed | 3024
gastrostomy removed | 3024
discrete hypotonia | 8760
fine motor skill difficulties | 8760
fatigability | 8760
intermittent hand tremors | 8760
normal deep tendon reflexes | 8760
electromyogram improving | 8760
discrete neurogenic involvement | 8760
