35 years old | 0 | 0 
female | 0 | 0 
pregnant | 0 | 0 
admitted to the hospital | 0 | 0 
fever | -240 | 0 
cough | -240 | 0 
dyspnoea | -120 | 0 
aggravated dyspnoea | -120 | 0 
yellow viscous sputum | -240 | 0 
chest distress | -240 | 0 
shortness of breath | -240 | 0 
cyanosis of the lip | 0 | 0 
thick breathing sounds in both lungs | 0 | 0 
dry and wet rales in the right lower lung | 0 | 0 
tachycardia | 0 | 0 
gestational age 34 + 4 weeks | 0 | 0 
G2P1 | 0 | 0 
pre-pregnancy weight 46.5 kg | 0 | 0 
body mass index 16.87 | 0 | 0 
weight gain 8.8 kg during pregnancy | 0 | 0 
uterine height 34 cm | 0 | 0 
abdominal circumference 89 cm | 0 | 0 
contractions sporadic and weak | 0 | 0 
head presentation | 0 | 0 
foetal heart sounds 142 beats/min | 0 | 0 
intrapelvic and extrapelvic measurements normal | 0 | 0 
increased CRP | 0 | 0 
increased erythrocyte sedimentation rate | 0 | 0 
increased procalcitonin | 0 | 0 
leukocytosis | 0 | 0 
neutrophilia | 0 | 0 
lymphopenia | 0 | 0 
abnormal liver enzymes | 0 | 0 
chest CT showed multiple plaques, miliary foci, nodular foci with partial consolidation and cavities | 0 | 0 
obstetric ultrasound showed a single viable foetus, head presentation, and oligohydramnios | 0 | 0 
cardiac ultrasound and lower extremity vascular ultrasound showed no significant abnormalities | 0 | 0 
S. aureus infection | 0 | 0 
COVID-19 infection | 0 | 0 
respiratory failure | 0 | 0 
caesarean section | 24 | 24 
oxyhemoglobin saturation decreased | 0 | 24 
oxyhemoglobin saturation increased | 24 | 48 
foetal distress | 0 | 24 
discharged | 264 | 264 
antibiotic therapy | 0 | 264 
antiviral therapy | 0 | 264 
glucocorticoids | 0 | 264 
acetaminophen | 0 | 264 
anticoagulant therapy | 0 | 264 
mNGS testing | 24 | 24 
S. aureus identified | 24 | 24 
COVID-19 identified | 24 | 24 
vancomycin | 24 | 264 
meropenem | 24 | 264 
sitafloxacin | 216 | 264 
chest CT showed improvement | 216 | 264 
pleural effusion absorbed | 216 | 264 
inflammatory lesions improved | 216 | 264 
electrolyte disturbance | 0 | 0 
hypoproteinaemia | 0 | 0 
oligohydramnion | 0 | 0 
premature live baby | 24 | 24 
maternal lower weight | 0 | 0 
elderly second parturient women | 0 | 0 
late pregnancy | 0 | 0 
G2P1 left occiput anterior | 0 | 0 
pregnancy combined with severe pneumonia | 0 | 0 
novel coronavirus infection | 0 | 0 
S. aureus infection | 0 | 0 
respiratory failure | 0 | 0 
treated with cefoperazone sodium and sulbactam sodium | 0 | 24 
treated with dexamethasone | 0 | 24 
high-flow nasal cannula oxygen therapy | 24 | 48 
assisted ventilation by endotracheal intubation | 24 | 48 
symptomatic treatment | 24 | 264 
fluid and ALB infusion | 24 | 264 
irrigation solution collected and tested for mNGS | 24 | 24 
bedside tracheoscopy | 24 | 24 
acid-fast bacilli in the sputum tuberculosis smear negative | 24 | 24 
tubercle bacillus-polymerase chain reaction negative | 24 | 24 
nontuberculosis mycobacterium-PCR negative | 24 | 24 
galactomannan experiments normal | 24 | 24 
bacterial resistance gene test | 24 | 24 
S. aureus resistant to macrolide and lincosamide antibiotics | 24 | 24 
chest CT showed multiple areas of inflammation in both lungs | 96 | 96 
mildly enlarged mediastinal lymph nodes | 96 | 96 
small amount of bilateral pleural effusion | 96 | 96 
CRP decreased | 96 | 96 
WBC count decreased | 96 | 96 
PCT decreased | 96 | 96 
potassium normal | 96 | 96 
D-dimer decreased | 96 | 96 
TB-PCR negative | 96 | 96 
chest CT showed inflammatory lesions improved | 216 | 216 
pleural effusion absorbed | 216 | 216 
antibiotics adjusted to sitafloxacin | 216 | 264 
patient condition stable | 264 | 264 
discharged from hospital | 264 | 264 
follow-up chest CT showed multiple lung inflammation absorbed | 336 | 336 
follow-up chest CT showed multiple lung inflammation apparently absorbed | 432 | 432 
mNGS results showed S. aureus and COVID-19 | 24 | 24 
S. aureus coverage 93.1785% | 24 | 24 
COVID-19 coverage 5.8690% | 24 | 24 
bacterial resistance gene test results showed S. aureus resistant to macrolide and lincosamide antibiotics | 24 | 24 
S. aureus sequence number 43700 | 24 | 24 
COVID-19 sequence number 10 | 24 | 24 
caesarean section performed | 24 | 24 
foetus transferred to neonatal ICU | 24 | 24 
patient transferred to respiratory ICU | 24 | 24 
patient received assisted ventilation by endotracheal intubation | 24 | 48 
patient received empirical antibiotic therapy | 24 | 264 
patient received symptomatic treatment | 24 | 264 
patient received fluid and ALB infusion | 24 | 264 
patient received high-flow nasal cannula oxygen therapy | 24 | 48 
patient received anticoagulant therapy | 24 | 264 
patient received treatments to relieve cough and reduce sputum | 24 | 264 
patient received other symptomatic treatment | 24 | 264 
patient condition improved | 96 | 264 
patient discharged from hospital | 264 | 264 
follow-up patient condition stable | 336 | 432 
follow-up patient discharged from hospital | 432 | 432