16 years old | 0
female | 0
admitted to the hospital | 0
syncope | -144
malaise | -144
fever | -144
fatigue | -144
chest pain | -144
shortness of breath | -144
presyncopal episode | -144
dizziness | -144
vision changes | -144
sweating | -144
true syncopal episode | -144
afebrile | 0
blood pressure 93/72 mmHg | 0
pulse rate 90s–100 beats per minute | 0
respiratory rate 16 | 0
oxygen saturation 100% | 0
mild pain from fall | 0
no head/facial bruising | 0
tachycardic | 0
normal heart sounds | 0
no murmurs | 0
lungs clear to auscultation | 0
no hepatosplenomegaly | 0
normal sinus rhythm | 0
low-voltage QRS complexes | 0
T-wave inversions | 0
normal electrolytes | 0
normal complete blood counts | 0
normal inflammatory markers | 0
mildly depressed left ventricular function | 0
ejection fraction 50% | 0
small pericardial effusion | 0
moderate-to-severe concentric LV hypertrophy | 0
LV diastolic septal and posterior wall thickness 1.4 cm | 0
hypertrophic cardiomyopathy suspected | 0
myocarditis suspected | 0
admitted for close monitoring | 0
initial troponin I 0.977 ng/mL | 0
fluid refractory hypotension | 24
sinus tachycardia | 24
tachypnea | 24
transferred to cardiac intensive care unit | 24
vasopressor support started | 24
dopamine started | 24
milrinone started | 24
viral polymerase chain reactions obtained | 24
influenza A positive | 24
peramivir started | 24
repeat echocardiogram | 48
increased pericardial effusion | 48
pericardiocentesis performed | 48
pericardial drain placement | 48
biphasic positive airway pressure started | 48
intravenous immunoglobulin given | 48
gradually improved | 120
weaned from intravenous infusions | 120
weaned from supplemental oxygen | 120
repeat TTE | 120
ejection fraction >70% | 120
persistent concentric LVH | 120
all symptoms resolved | 168
TTE revealed resolving LVH | 168
discharged | 168
cMRI showed normal biventricular chamber sizes | 3360
cMRI showed normal biventricular systolic function | 3360
cMRI showed normal LV mass | 3360
cMRI showed no LVH | 3360
cMRI showed no late gadolinium enhancement | 3360
echocardiogram showed resolution of LVH | 3360