49 years old | 0
female | 0
generalized weakness | -720
abdominal pain | -720
back pain | -720
abdominal fullness | -8760
marked splenomegaly | 0
hemoglobin 9 | 0
platelet count 40 | 0
white blood cell count 45 | 0
17% blasts | 0
bone marrow core biopsy 100% cellular | 0
myeloid predominance | 0
30% to 40% blasts | 0
complex 4-way rearrangement | 0
BCR-ABL rearrangement | 0
deletion in the long arm of chromosome 14 | 0
translocation between the short arm of chromosomes 7 and 12 | 0
BCR-ABL1 gene rearrangement | 0
next-generation sequencing negative for ASXL1, DNMT3A, FLT3, IDH1, IDH2, NPM1, RUNX1, TET2, TP53, and Wt1 | 0
CML-BC | 0
induction chemotherapy with cytarabine plus daunorubicin | 0
dasatinib 140 mg twice daily | 0
follow-up bone marrow biopsy | 168
complete morphologic remission | 168
normal female karyotype | 168
FISH negative for BCR-ABL translocation | 168
complete cytogenetic remission | 168
allogeneic hematopoietic stem cell transplant | 168
myeloablative conditioning with fludarabine and busulfan | 168
stable course | 1944
new leukocytosis | 1944
increased blast count | 1944
hemoglobin 11.7 | 1944
platelet count 20 | 1944
WBC 39 | 1944
10% peripheral blasts | 1944
prothrombin time 18 | 1944
internationalized normal ratio 1.6 | 1944
activated partial thromboplastin time 26 | 1944
fibrinogen 456 | 1944
negative soluble fibrin monomers | 1944
fever 38.4 | 1946
hypotension | 1946
sepsis | 1946
blood cultures showed no growth | 1946
CT scan of the abdomen and pelvis showed evidence of colitis | 1946
stool testing positive for Clostridioides difficile | 1946
peripheral blast count increased to 41% | 1948
bone marrow aspirate and core biopsy | 1947
nearly 100% cellular marrow | 1947
absent erythroids and megakaryocytes | 1947
85% to 90% blasts | 1947
relapse of CML-BC | 1947
fluorescence in situ hybridization analysis of peripheral blood confirmed BCR-ABL1 fusion | 1947
worsening coagulopathy | 1947
anemia | 1947
thrombocytopenia | 1947
hemoglobin 6.4 | 1947
hematocrit 19.2 | 1947
platelet count 9 | 1947
internationalized normal ratio increased to 4.1 | 1948
prothrombin time 52.7 | 1948
factor VII activity 3% | 1948
factor II activity 55% | 1948
factor X activity 57% | 1948
factor V activity 77% | 1948
oral vitamin K 5 mg | 1948
decreased level of responsiveness | 1948
transfer to intensive care unit | 1948
CT scan of the head ruled out intracranial hemorrhage | 1948
no evidence of bleeding | 1948
chemotherapy regimen for relapsed disease | 1950
cladribine 5 mg/m2 IV | 1950
cytarabine 20 mg subcutaneous twice daily | 1950
venetoclax for 21 days | 1950
clinical improvement | 1952
transferred back to the hematology ward | 1952
concerns for vision loss | 1952
dilated fundus exam showed severe bilateral retinal hemorrhages | 1952
coagulopathy improved | 1952
peripheral blast count decreased | 1952
FVII activity improved to 63% | 1980
hospital discharge | 1980
improvement of blurry vision | 1980
bone marrow aspirate and biopsy showed persistent disease | 4032
70% blasts | 4032
FVII activity decreased to 14% | 4032
INR 2.2 | 4032
decitabine and venetoclax for refractory disease | 4032
FVII level activity remained low at 15% | 4042
no bleeding | 4042
remission after 1 cycle of therapy | 4042
poor functional status | 4042
not a candidate for a second allogeneic hematopoietic stem cell transplantation | 4042