62 years old | 0
female | 0
alcohol abuse | -672
hypertension | -672
family history of seizure disorder | -672
daily alcohol intake | -672
admitted to the hospital | 0
dental pain | -72
facial swelling | -72
altered mental status | -72
Glasgow Coma Scale 13 | 0
not oriented to time or place | 0
febrile | 0
temperature 40° Celsius | 0
heart rate 160 beats per minute | 0
pupils 1 mm in diameter | 0
minimally reactive to light | 0
no afferent pupillary defect | 0
visual acuity at least hand motion | 0
orthotropic in primary gaze | 0
full ocular motility | 0
intraocular pressures 19 and 14 mm Hg | 0
right periorbital and temporal edema | 0
right periorbital and temporal erythema | 0
inferior chemosis of the right conjunctiva | 0
no conjunctival erythema | 0
septic shock | 0
serum anion gap 23 mEq/L | 0
lactic acid 4.8 mmol/L | 0
white blood cell count 15,000/mm3 | 0
started on intravenous vancomycin | 0
started on piperacillin/tazobactam | 0
started on metronidazole | 0
urinalysis unremarkable | 0
chest radiograph showed 2.7 cm right upper lung opacity | 0
chest radiograph showed heterogeneous basilar opacities | 0
CT of the chest without contrast showed bilateral lung masses and nodules | 0
CT of the chest without contrast showed septic emboli | 0
CT of the face with contrast showed multi-fascial space abscesses | 0
CT of the face with contrast showed phlegmon | 0
CT of the face with contrast showed gas extending to the right lateral supraorbital soft tissues | 0
CT of the face with contrast showed thrombophlebitic right retromandibular vein | 0
CT of the face with contrast showed thrombophlebitic superior temporal vein | 0
CT of the face with contrast showed periorbital cellulitis | 0
CT of the face with contrast showed thrombophlebitis of the right infraorbital facial vein | 0
CT of the face with contrast showed thrombophlebitis of the right internal jugular vein | 0
incision and drainage of facial abscesses | 24
extraction of five carious teeth | 24
blood cultures grew viridans group streptococci | 72
abscess cultures grew viridans group streptococci | 72
tracheal aspirate cultures negative | 72
urine cultures negative | 72
blood culture susceptibilities showed minimal inhibitory concentration of <0.1 μg/mL to penicillin | 72
discontinued vancomycin | 72
discontinued clindamycin | 72
discontinued piperacillin/tazobactam | 72
started on ampicillin/sulbactam | 72
considered anticoagulation for thrombophlebitis | 72
anticoagulation held due to eradication of bacteremia | 72
transferred out of the intensive care unit | 120
complained of binocular diplopia | 168
noted to have large right incomitant esotropia | 168
noted to have −4 abduction | 168
consistent with lateral rectus paralysis | 168
consistent with right sixth nerve palsy | 168
cranial nerve function intact | 168
extraocular movements intact | 168
no signs of nystagmus | 168
intraocular pressures 16 mm Hg | 168
visual acuities 20/30 bilaterally | 168
mild chemosis | 168
no conjunctival erythema | 168
CT angiogram of the head showed hypoenhancement of the right greater than left cavernous sinuses | 168
CT angiogram of the head showed concern for CST | 168
CT of the face with contrast showed persistence of multifascial abscesses | 168
repeat incision and drainage | 192
considered anticoagulation | 192
anticoagulation avoided due to upper gastrointestinal bleed | 192
discharged | 240
switched to ertapenem | 240
completed six weeks of treatment | 480
follow-up showed no improvement of sixth nerve palsy | 480