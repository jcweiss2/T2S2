53 years old | 0
male | 0
diagnosed with grade II follicular lymphoma | 0
autologous bone marrow transplant | 0
recurrence to initial chemotherapy | -672
treated with eight cycles of R-CVP | -2016
Rituximab | -2016
Cyclophosphamide | -2016
Vincristine | -2016
prednisone | -2016
treated with three cycles of R-ICE | -1344
Iphosphamide | -1344
Carboplatin | -1344
Etoposide | -1344
treated with two cycles of R-DA=EPOCH | -1008
dose-adjusted etoposide | -1008
prednisone | -1008
vincristine | -1008
cyclophosphamide | -1008
doxorubicin | -1008
rituximab | -1008
conditioning regimen prescribed with BEAM | 0
carmustine | 0
etoposide | 0
cytosine arabinoside | 0
melphalan | 0
prophylactic antimicrobial treatment prescribed with fluconazole | 0
neutropenia | 24
fever | 72
intense myalgia | 72
papular skin lesion | 72
papular skin lesion with rapid dissemination | 72
papular lesions progressed with central ischemia | 72
papular lesions progressed with necrosis | 72
empiric antimicrobial treatment with meropenen | 72
vancomycin | 72
liposomal amphotericin | 72
baseline total leukocyte count | 72
skin biopsy revealed abundant hyphae structures | 72
blood cultures identified Fusarium solani | 72
transferred to intensive care unit | 72
voriconazole added to antifungal therapy | 72
ophthalmologic evaluation revealed no signs of endophthalmitis | 72
radiographic images were unremarkable | 72
heavy myoglobinuria | 72
normal creatine phosphokinase | 72
worsened renal function | 72
increased blood lactate | 72
elevation of C-reactive protein | 72
elevation of pro-calcitonin | 72
serum (1-3)-β-d-glucan not assessed | 72
granulocyte transfused | 72
no significant improvement of clinical condition | 72
refractory septic shock | 72
intensive care support | 72
renal replacement therapy | 72
mechanical ventilation | 72
unresponsive cardiac arrest | 96
no previous history of fungal diseases | 0
no skin lesion observed prior to terminal event | 0
no nail lesion observed prior to terminal event | 0
fungal susceptibility testing revealed resistance to fluconazole | 72
fungal susceptibility testing revealed susceptibility to voriconazole | 72
fungal susceptibility testing revealed susceptibility to amphotericin | 72
investigation regarding potential source of infection conducted | 72
cultures of tap water negative for fungal growth | 72
cultures of shower bath water negative for fungal growth | 72
no skin lesion at hospital admission | -96
no nail lesion at hospital admission | -96
no skin lesion at post-transplant period | 0
no nail lesion at post-transplant period | 0
autologous BMT recipient | 0
neutropenia duration | 24
disseminated fusariosis | 72
fatal outcome | 96
negative hospital environmental cultures | 72
negative shower bath water cultures | 72
negative tap water cultures | 72
no prophylactic voriconazole | 0
increasing incidence of invasive mold infections | 0
hematological malignancies | 0
hematopoietic cell transplant recipients | 0
widespread use of rituximab | 0
treatment with amphotericin B | 72
treatment with voriconazole | 72
granulocyte transfusion | 72
lethal disseminated Fusarium infection | 96
pre-engraftment phase | 0
careful clinical evaluation of BMT candidates | 0
exhaustive vigilance of environmental cleansing procedures | 0
antifungal prophylaxis selection | 0
need for antifungal prophylaxis studies | 0
treated with three cycles of R&ndash;ICE | -1344
treated with two cycles of R-DA-EPOCH | -1008
