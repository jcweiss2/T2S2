63 years old | 0
    male | 0
    history of smoking (20 packs/year) | 0
    DVT in the left leg | -432
    rivaroxaban anticoagulant therapy | -432
    hospitalized due to abrupt onset of dyspnea | -168
    thoracic CT scan confirmed pulmonary thromboembolism | -168
    mass in the lower lobe of the right lung | -168
    ipsilateral ilo(mediastinal pathological lymph nodes | -168
    infra-clavear pathological lymph nodes | -168
    abdominal CT scan demonstrated splenic infarction | -168
    abdominal CT scan demonstrated renal infarction | -168
    developed right cerebellar signs | -144
    confusion | -144
    nystagmus | -144
    ataxia | -144
    dysmetria | -144
    adiadochokinesia | -144
    MRI of the brain revealed multiple cerebral and cerebellar areas | -144
    hyperintense in fluid-attenuated inversion recovery/fast spin echo sequences | -144
    diffusion restriction | -144
    moderate patchy and gyriform enhancement | -144
    ischemic lesions on an embolic basis | -144
    miliary brain metastases | -144
    transthoracic echocardiogram (TTE) | -144
    transesophageal echocardiogram (TEE) not performed | -144
    spontaneous rapid improvement of neurological state | -144
    complete resolution of confusion | -144
    complete resolution of cerebellar symptoms | -144
    cardio embolic origin of brain lesions suspected | -144
    TEE carried out | -144
    revealed PFO | -144
    paradoxical arterial embolisms | -144
    no surgical correction of PFO | -144
    discharged | -144
    prescribed subcutaneous LMWH | -144
    lung cancer diagnosis | 0
    locally advanced non-small cell lung cancer (NSCLC) | 0
    PET scan confirmed locally advanced extension | 0
    EBUS-guided transbronchial needle aspiration performed | 0
    diagnosis of large-cell carcinoma of the lung | 0
    immunohistochemistry (IHC) | 0
    positive for cytokeratin pool | 0
    lacked expression of TTF-1 | 0
    lacked expression of p40 | 0
    lacked expression of chromogranin A | 0
    lacked expression of synaptophysin | 0
    positivity for cytokeratin CAM5.2 | 0
    excluded lymphoma | 0
    no EGFR mutations | 0
    no ALK gene rearrangements | 0
    PD-L1 tumor proportion score 55% | 0
    candidate for immunotherapy with pembrolizumab | 0
    onset of diplopia | 0
    gait impairment | 0
    hospitalization (University Hospital of Parma, Italy) | 0
    CT scan documented evolution of the lesion | 0
    developed substernal chest pain | 24
    dyspnea | 24
    body temperature regular | 24
    blood pressure regular | 24
    heart rate regular | 24
    diastolic murmur consistent with aortic regurgitation | 24
    sinus tachycardia (90 beats/min) | 24
    ST segment elevation in DII-DIII-aVF derivations | 24
    elevated serum troponin I | 24
    peak value 22.91 ng/ml | 24
    TTE showed reduced LVEF 45% | 24
    mobile mass on anterior leaflet of mitral valve | 24
    moderate aortic insufficiency | 24
    acute pulmonary edema | 24
    respiratory failure | 24
    noninvasive ventilation | 24
    coronary angiography showed reduced flow (TIMI score=2) | 24
    embolus appearance | 24
    no atherosclerotic lesions | 24
    admitted to intensive care unit | 24
    therapy with aspirin | 24
    therapy with β-blockers | 24
    maintained LMWH treatment | 24
    suspicion of infective endocarditis | 24
    blood culture tests | 24
    empiric intravenous antibiotic therapy | 24
    linezolid 600 mg twice daily | 24
    daptomycin 6 mg/kg once daily | 24
    piperacillin/tazobactam 4.5 g three times daily | 24
    petechiae on the skin of lower limbs | 24
    abdominal CT scan performed | 24
    abdominal pain | 24
    loss of blood in the stool | 24
    occlusion of distal branch of superior mesenteric artery | 24
    thinning of corresponding ileal loop | 24
    emergency segmental ileo-cecal resection | 24
    histological diagnosis of bowel infarction | 24
    remained intubated | 24
    TEE performed | 24
    mobile echogenic mass 0.8×0.6 cm on mitral valve | 24
    moderate aortic insufficiency | 24
    reduced LVEF 40% | 24
    no signs of PFO | 24
    negativity of blood cultures | 24
    normal procalcitonin | 24
    diffuse embolic manifestations | 24
    diagnosis of NBTE | 24
    coma | 24
    brain CT scan documented increased infarct lesions | 24
    progression of cerebral ischemic events | 24
    onset of novel interested foci | 24
    multi-organ failure | 24
    passed away | 24
    ~70 days after lung cancer diagnosis | 1680

    
