Here is the table of events and timestamps:

pregnancy diagnosis | 0
37.6 weeks of gestation | 0
viable intrauterine pregnancy | 0
fetal heart rate 143 beats per minute | 0
fetus situated longitudinally with cephalic presentation, back to the left | 0
cervix 6 cm dilated | 0
70% effaced | 0
station +1 | 0
intact membranes | 0
mild edema of the extremities | 0
normal osteotendinous reflexes | 0
obstetrical ultrasound | -5
pregnancy of 37+0 weeks of gestation | -5
posterior body placenta maturation grade III | -5
amniotic fluid index of 8.7 cm | -5
5th percentile of 50 for gestational age | -5
biophysical profile of 8/8 | -5
Hadlock of 34.2% | -5
weight of 3033 grams | -5
spontaneous rupture of the membranes | -4
7 cm dilation | -4
effective labor | -4
4 contractions every 10 minutes that lasted 40 to 45 seconds | -4
no uterotonic agents | -4
fully dilated | -4
100% clearance | -4
station of +3 | -4
fetus in left occiput anterior position | -4
live newborn | -4
Apgar scores of 7 and 9 | -4
gestational age of 40 weeks | -4
height 48 cm | -4
weight of 2650 grams | -4
Schultze mechanism | -4
placenta came out with normal characteristics | -4
grade III uterine inversion | -4
manual reinversion | -4
no success | -4
total blood loss of 1200 mL | -4
UA | -4
oxytocin | -4
carbetocin | -4
misoprostol | -4
exploratory laparotomy | -4
uterine inversion evaluated | -4
reinversion was successful | -4
UA persisted | -4
PPH | -4
Hayman hemostatic suture | -4
no response | -4
bilateral ligation of the anterior trunk of the hypogastric artery | -4
immediate recovery of uterine tone | -4
cessation of PPH | -4
uterus regained tone in approximately 5 minutes | -4
postligation bleeding was only 50 mL | -4
2 bags of packed red blood cells transfused | -4
hemoglobin level of 7 g | -4
transferred to the recovery room | -4
transferred to the medical intensive care unit | -4
transferred to a hospital room | -4
normal diet | -4
ambulation | -4
spontaneous uresis | -4
normal peristalsis | -4
breastfeeding | -4
discharged on the second day | -4
description of the technique of bilateral ligation of the hypogastric artery in its anterior trunk | -4
initial anatomic reference from where the retroperitoneum is incised | -4
bifurcation of the common iliac artery identified | -4
correct identification of the decussation of the ureter above the artery | -4
retroperitoneum dissected parallel to the entire course of the hypogastric artery | -4
anterior trunk is carefully dissected until it is completely freed and ligated with absorbable catgut suture 1-0 | -4
hemostasis is checked | -4
same procedure is performed contralaterally | -4
ligation of the anterior trunk of the hypogastric artery bilaterally | -4
no complications | -4
effective, safe, and fertility-preserving surgical procedure | -4