56 years old | 0
male | 0
admitted to the hospital | 0
severe anal pain | 0
bleeding | 0
history of external hemorrhoids | -7200
denied any systemic diseases | 0
thrombosed external protruding hemorrhoid | 0
surgery suggested | 0
preoperative blood pressure 108/96 mmHg | 0
pulse 59 beats per minute | 0
oxygen saturation 100% | 0
other examination results were normal | 0
routine laboratory examinations were within normal limits | 0
routine chest X-ray examination was normal | 0
hemorrhoidectomy | 0
vital signs were similar to those from preoperative examination | 24
temperature 36.4 oC | 24
blood pressure 85/50 mmHg | 24
pulse 83 beats per minute | 24
good spirits | 24
fair activity | 24
moderate wound pain | 24
mild swelling | 24
no pus or bloody discharge | 24
Mefenamic acid 250mg QID PO | 24
Pethidine 50mg PRN | 24
increased pulse rates to 108 beats per minute | 48
persistent hypotension | 48
denied having dizziness | 48
denied chills | 48
denied weakness | 48
denied poor appetite | 48
denied low urine output | 48
sepsis considered | 48
stress ulcer induced gastrointestinal bleeding considered | 48
dehydration considered | 48
denied tarry stool | 48
denied epigastric discomfort | 48
planned to give intravenous fluid | 48
refused to establish an intravenous line | 48
water intake encouraged | 48
vital signs closely monitored | 48
fever to 38.6 oC | 72
chills | 72
blood pressure 70/42 mmHg | 72
pulse 124 beats per minute | 72
oxygen saturation 97% | 72
two sets of blood cultures | 72
laboratory tests | 72
leukocytosis | 72
elevated C-reactive protein | 72
blood urea nitrogen 40.6 mg/dL | 72
creatinine 2.6 mg/dL | 72
decreased platelets | 72
intravenous fluid | 72
antibiotics | 72
Cefmetazole 1g Q8H | 72
rechecked vital signs | 74
blood pressure 155/110 mmHg | 74
pulse 88 beats per minute | 74
oxygen saturation 95% | 74
general soreness | 74
discomfort | 74
consciousness change | 80
body temperature 36.1 oC | 80
blood pressure 68/51 mmHg | 80
pulse 144 beats per minute | 80
respiratory rate 27 per minute | 80
oxygen saturation 95% | 80
immediate intravenous fluid resuscitation | 80
artery blood gas analysis | 80
pH 7.32 | 80
pCO2 16.9 mmHg | 80
pO2 118.9 mmHg | 80
HCO3 8.5 mmol/L | 80
sent to the intensive care unit | 80
endotracheal tube put in place | 80
Sodium bicarbonate given | 80
persistent metabolic acidosis | 80
continuous venous-venous hemofiltration | 80
sudden cardiac arrest | 80
cardiopulmonary resuscitation | 80
emergent extracorporeal membrane oxygenation | 80
ECMO applied | 80
cardiac arrest again | 82
expired | 82
blood culture yielded Streptococcus pyogenes | 82
wound culture yielded Streptococcus pyogenes | 82