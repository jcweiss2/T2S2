23 years old | 0
male | 0
admitted to the hospital | 0
abdominal pain | 0
jaundice | 0
biliary cirrhosis | -3456
abnormal liver function tests | -3456
alcohol consumption | -3456
visited the emergency room | -168
abdominal pain | -168
discharged | -168
visited the emergency room | -24
abdominal pain | -24
discharged | -24
hepatosplenomegaly | 0
collateral vessels | 0
esophageal varices | 0
total bilirubin | 0
direct bilirubin | 0
aspartate aminotransferase | 0
alanine aminotransferase | 0
proximal limb pain | 0
skin sensitivity | 0
family history of multiple skin blisters | 0
porphyria | 0
increased coproporphyrin | 0
uroporphyrin | 0
acute liver failure | 0
hypovolemic shock | 0
intra-abdominal bleeding | 0
renal function deteriorated | 0
continuous renal replacement therapy | 0
listed for liver transplantation | 696
sinus tachycardia | 696
echocardiogram | 696
pulmonary edema | 696
pulmonary effusion | 696
model for end-stage liver disease score | 696
intubated | 696
norepinephrine | 696
Bispectral Index monitor | 696
ventilator care | 696
arterial cannulation | 696
central venous cannulation | 696
multifunction Swan-Ganz catheter | 696
endotracheal tube | 696
general anesthesia | 696
propofol | 696
remifentanil | 696
atracuronium | 696
hypovolemic acute renal failure | 696
dopamine | 696
liver transplantation operation | 771
crystalloid | 771
colloid | 771
albumin | 771
packed red blood cells | 771
fresh frozen plasma | 771
platelet concentrate | 771
cryoprecipitate | 771
calcium gluconate | 771
anuric | 771
acute renal failure | 771
transferred to ICU | 1071
alert | 72
renal function improved | 72
continuous renal replacement therapy discontinued | 72
motor function weak | 72
extubation delayed | 72
motor power grade 2 | 216
severe sensory and motor polyneuropathy | 216
tracheostomy | 312
liver function tests improved | 216
liver function worsened | 744
fever | 744
antibiotics | 744
multi-organ failure | 2496
expired | 2496