68 years old | 0
male | 0
admitted to the hospital | 0
chief complaint of subjective fever | 0
bilateral leg pain | 0
worsening blistering | 0
bleeding from BP lesions | 0
history of chronic lymphocytic leukemia | -8760
history of bullous pemphigoid | -1460
hospital admission 2 weeks prior | -336
treated with prednisone | -336
treated with doxycycline | -336
shave biopsy of the bullous skin lesions | -336
diagnosed with refractory CLL | -8760
treated with rituximab | -8760
treated with cyclophosphamide | -8760
treated with vincristine | -8760
treated with prednisone | -8760
treated with fludarabine | -8760
started on ibrutinib | -2628
treated with apixaban | -2628
diagnosed with deep vein thrombosis | -2628
diagnosed with chronic obstructive pulmonary disease | -2628
diagnosed with diastolic heart failure | -2628
diagnosed with non-insulin dependent diabetes mellitus | -2628
treated with intravenous immunoglobulin | -2628
developed sepsis | 24
developed atrial fibrillation | 24
developed hypotension | 24
transferred to the intensive care unit | 24
started on broad spectrum antibiotics | 24
started on vancomycin | 24
started on meropenem | 24
held ibrutinib | 24
continued prophylactic acyclovir | 24
tapered prednisone | 24
shave biopsy results showed trophozoites | 48
started on intravenous fluconazole | 48
stabilized in the intensive care unit | 72
discontinued vancomycin | 72
discontinued meropenem | 72
consulted with dermatology | 72
repeat punch biopsies performed | 72
switched to intravenous liposomal amphotericin B | 72
negative blood cultures | 72
negative cryptococcal antigen | 72
negative urine histoplasma antigen | 72
negative urine blastomycosis antigen | 72
negative serum coccidioides antibody | 72
computed tomography of the chest, abdomen and pelvis | 72
hiatal hernia | 72
splenomegaly | 72
transferred out of the intensive care unit | 120
continued on intravenous liposomal amphotericin B | 120
punch biopsies showed clusters of septate hyphae | 120
X-rays of the bilateral tibia and fibula | 120
subcutaneous skin thickening | 120
fungal cultures from punch biopsies returned positive for mucormycosis | 336
developed foul smelling drainage | 480
white blood cell count increased | 480
started on daptomycin | 480
started on meropenem | 480
wound cultures grew Pseudomonas | 480
wound cultures grew E. coli | 480
completed 7-day course of antibiotics | 544
transitioned to posaconazole | 672
discharged to a skilled nursing facility | 1440