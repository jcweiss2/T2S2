15 years old | 0
    male | 0
    mild infrequent asthma | 0
    road traffic accident | -120
    suspected intracranial involvement | -120
    not wearing a helmet | -120
    collision with a car | -120
    incident on bright daylight | -120
    hill side location | -120
    possible inhalation of water or soil | -120
    Glasgow Coma Scale 6 | -120
    oxygen saturation 75% | -120
    intubated | -120
    respiratory failure | -120
    chest xray reveals massive right haemothorax | -120
    segmented fracture of 6th posterior rib | -120
    ipsilateral chest tube inserted | -120
    300 ml blood drained | -120
    transferred to tertiary hospital | -120
    CT brain reveals subarachnoid haemorrhage | -120
    punctate intracerebral haemorrhage | -120
    burr hole done | -120
    intracranial pressure monitoring attached | -120
    transferred to ICU | -120
    ventilator support | 0
    minimal inotropic support (0.1-0.2 mcg/kg/min Noradrenaline) | 0
    extubation attempted after 72 hours | 72
    improvement in neurological status | 72
    minimal inotropic support | 72
    low ventilator settings | 72
    reintubation after 8 hours | 80
    moderate ventilator settings | 80
    significant secretions | 80
    fever (38-40°C) | 80
    bronchoscopy performed | 80
    purulent secretions | 80
    blood cultures positive for Burkholderia pseudomallei | 80
    tracheal secretions cultures positive | 80
    bronchoalveolar lavage cultures positive | 80
    gram negative bacilli with safety-pin appearance | 80
    sensitivity to amoxicillin-clavulanate | 80
    sensitivity to ceftazidime | 80
    sensitivity to doxycycline | 80
    sensitivity to imipenem | 80
    sensitivity to trimethoprim-sulfamethoxazole | 80
    Hepatitis B negative | 80
    Hepatitis C negative | 80
    HIV negative | 80
    syphilis negative | 80
    CXR shows right hemithorax consolidation | 80
    low to moderate ventilator support | 80
    minimal inotropic support | 80
    extubated after 168 hours | 168
    discharged to general ward after 504 hours | 504
    IV Meropenem started after 168 hours | 168
    IV Ceftazidime deescalated after 168 hours | 168
    oral trimethoprim-sulfamethoxazole planned | 504
    no commercial conflicts | 0
    