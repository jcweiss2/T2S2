22 years old | 0
female | 0
admitted to the hospital | 0
swallowing difficulties | 0
throat pain | 0
local inflammation of the tonsils | 0
tonsillitis | 0
symptomatic therapy with ibubrufen | 0
discharged | 0
paresis of the abducens nerve | 144
paresis of the oculomotor nerve | 144
mydriasis of the right eye | 144
impairment in function of the musculus levator | 144
impairment in motion of the right eye | 144
prism cover test | 144
exophthalmos on the right side | 216
paralysis of the abducens nerve on the left eye | 216
photophobia | 216
incomplete trismus | 216
signs of meningism | 216
fever | 216
leucocytosis | 216
thrombocytopenia | 216
activated coagulation | 216
international normalized ratio | 216
magnetic resonance imaging | 216
thromboses in the cavernous sinus | 216
thrombosis of the superior ophthalmic vein | 216
abscess in the right temporal lobe | 216
computed tomography of the neck | 216
abscess in the left tonsil | 216
thrombus in the right internal jugular vein | 216
computed tomography of the lung | 216
septic emboli | 216
starting abscesses | 216
diagnosis of Lemierre's syndrome | 216
high-dose intravenous antibiotic therapy | 216
anticoagulation therapy | 216
blood cultures | 216
anaerobic cultures | 216
Fusobacterium necrophorum | 240
operative drainage of the left tonsillary abscess | 288
progressive brain abscess | 288
switched to ceftriaxon and metronidazole | 288
mycotic aneurysm in the right internal carotid artery | 288
transferred to a neurosurgical intensive care unit | 288
discharged from the hospital | 2160
residual sign of an abducens nerve paralysis | 2160
oculomotor nerve paralysis | 2160