42 years old | 0
female | 0
admitted to the hospital | 0
altered mental status | 0
low grade fevers | -120
sudden deterioration in mental status | 0
history of intravenous drug use | -8760
extraction of all maxillary teeth | -2160
mandibular dental infection | -720
treated with oral amoxicillin | -720
temperature was 36.7 °C | 0
heart rate was 98 beats/min | 0
respiratory rate was 17 breaths/min | 0
blood pressure was 131/66 mm Hg | 0
oxygen saturation of 99% on room air | 0
denies fevers | 0
denies chills | 0
denies chest pain | 0
denies dyspnea | 0
denies nausea | 0
denies vomiting | 0
denies diarrhea | 0
denies skin lesions | 0
denies numbness | 0
denies tingling | 0
denies weakness of the lower extremities | 0
prominent holosystolic murmur at the apex | 0
petechial rash scattered on the abdomen | 0
petechial rash scattered on the palms | 0
petechial rash scattered on the soles of the feet | 0
encephalopathy | 0
facial droop | 0
slurred speech | 0
admitted to the intensive care unit | 0
started on empiric antibiotic treatment with vancomycin | 0
started on empiric antibiotic treatment with meropenem | 0
became unresponsive to voice | 24
minimally responsive to pain | 24
left hemi-neglect | 24
right gaze deviation | 24
Glasgow Coma Scale (GCS) was 6 | 24
intubated for airway protection | 24
leukocytosis of 24.7 × 10^9/L | 24
87.6% neutrophils | 24
platelet count of 17 × 10^9/L | 24
liver and kidney functions were within normal | 24
declined a HIV test | 24
innumerable acute to subacute embolic infarcts in both cerebral and cerebellar hemispheres | 24
proximal right internal carotid artery T-shaped acute thrombus | 24
occlusion of the right middle cerebral artery | 24
subarachnoid hemorrhage in the right parietal region | 24
subarachnoid hemorrhage around the posterior aspect of the midbrain | 24
echo densities on the tricuspid valve | 24
echo densities on the aortic valve | 24
echo densities on the mitral valve | 24
blood culture grew S. marcescens | 48
antibiotic changed to cefepime | 72
cardiothoracic surgery consulted | 72
patient was a poor candidate for surgery | 72
neurological status continued to deteriorate | 120
no cough or gag reflex | 144
pupils were fixed and mid-dilated | 144
family decided to withdraw care | 144
discharged to hospice care | 144