39 years old | 0
male | 0
admitted to the hospital | 0
ulcerative colitis | -8760
sclerosing cholangitis | -8760
azathioprine | 0
ursacol | 0
prednisone | 0
simvastatin | 0
spironolactone | 0
folic acid | 0
calcium carbonate | 0
good general condition | 0
healthy skin tone | 0
well hydrated | 0
feverless | 0
jaundiced | 0
stable vital signs | 0
target painless hepatomegaly | 0
spider veins | 0
lower limb edema | 0
high fever | 12
tachycardia | 12
myalgia | 12
anuria | 12
ceftriaxone | 12
lesions resembling purplish erythematous plaques | 12
recent trip to the coastal area | -24
samples for leptospirosis | 0
samples for dengue | 0
samples for yellow fever | 0
samples for spotted fever | 0
samples for meningococcemia | 0
negative results for leptospirosis | 0
negative results for dengue | 0
negative results for yellow fever | 0
negative results for spotted fever | 0
negative results for meningococcemia | 0
unresponsive to volume | 24
dyspnea | 24
respiratory distress | 24
transferred to the ICU | 24
vasoactive drugs | 24
mechanical ventilation | 24
skin lesions became confluent | 24
blisters | 24
discharge of sero-sanguineous fluids | 24
therapy with ceftriaxone changed to meropenem | 24
therapy with ceftriaxone changed to oxacillin | 24
blood cultures revealed growth of gram-negative bacillus | 24
Vibriovulnificus identified | 48
death | 32
sepsis | 12
septic shock | 24
disseminated intravascular coagulation | 24
necrotizing fasciitis | 24
leukocytosis | 24
alteration in renal function | 24
edema | 24
accumulation of fluid in the affected tissues | 24
elevated levels of ferritin | 0
elevated transferrin saturation | 0
immunodeficiencies | -8760
liver disease | -8760
diseases of iron accumulation | -8760
diabetes mellitus | 0
use of steroids | 0
chronic renal failure | 0
raw seafood ingestion | -24
doxycycline | 0
prophylactic measures | 0
microbial surveillance | 0
warning to consumers | 0 
culture result available | 72 
post-mortem | 72 
septicemia | 24 
refractory septic shock | 24 
intensive care unit support | 24 
antibiotic therapy | 24 
death | 32 
V. vulnificus-induced illness in Southern Brazil | 0 
water temperature | 0 
global climate change | 0 
microbial surveillance | 0 
warning to consumers | 0 
education about the risk associated with the consumption of raw seafood | 0