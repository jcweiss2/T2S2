28 years old | 0
nonpregnant | 0
female | 0
no known comorbidities | 0
fever | -120
epistaxis | -120
high grade fever | 0
tachycardia | 0
blood pressure of 80/50 mmHg | 0
mild icterus | 0
no organomegaly | 0
chest was clear | 0
hemoglobin of 13.3 g/dL | 0
total leukocyte count of 15,200/cu.mm | 0
platelets 30,000/cumm | 0
prerenal acute kidney injury | 0
total bilirubin of 3.2 mg/dL | 0
mild serum transaminitis | 0
peripheral smear showed trophozoites of Plasmodium vivax malaria | 0
peripheral smear showed schizonts of Plasmodium vivax malaria | 0
complicated vivax malaria | 0
sepsis | 0
multi-organ dysfunction | 0
treated with fluids | 0
inotropic support | 0
parenteral anti-malarials | 0
platelet transfusion | 0
hemoptysis | 48
tachypnea | 48
bilateral diffuse coarse crepitations | 48
chest-X-ray showed bilateral diffuse opacities | 48
arterial blood gas pH of 7.44 | 48
HCO3 of 15 mEq/l | 48
PaO2 of 44.5 mmHg | 48
PaCO2 of 16 mmHg | 48
hemoglobin decreased to 10.5 mg/dL | 48
shifted to intensive care unit | 48
provisional diagnosis of diffuse alveolar hemorrhage | 48
oxygen inhalation | 48
illness worsened | 72
mechanical ventilation | 72
intravenous steroids | 72
blood culture negative | 72
urine culture negative | 72
ultrasonography of abdomen suggestive of polyserositis | 72
moderate ascites | 72
minimal bilateral pleural effusion | 72
Dengue NS1ag positive | 72
Chikungunya IgM positive | 72
confirmed by reverse transcription polymerase chain reaction for Dengue | 72
confirmed by reverse transcription polymerase chain reaction for Chikungunya | 72
succumbed to co-infection with malaria | 96
succumbed to co-infection with dengue | 96
succumbed to co-infection with chikungunya | 96
