49 years old | 0
    woman | 0
    hepatocellular carcinoma | 0
    end-stage hepatitis B liver cirrhosis | 0
    MELD score 14 | 0
    Child-Pugh class B | 0
    hypertension | 0
    well controlled with medications | 0
    blood type A, Rh+ | 0
    ABO compatible donor | 0
    anesthesia induced with fentanyl | 0
    anesthesia induced with thiopental sodium | 0
    anesthesia induced with vecuronium | 0
    anesthesia maintained with oxygen, air, desflurane | 0
    neuromuscular block maintained with atracurium | 0
    hemodynamic monitoring | 0
    piggyback technique | 0
    preservation of caval flow | 0
    reperfusion of graft liver | 0
    right posterior sectionectomy | 0
    decreased right hepatic venous flow | 0
    relatively large size of graft liver | 0
    morbid obesity | 0
    graft blood flow did not improve | 0
    intractable bleeding occurred | 0
    rapid volume resuscitation | 0
    hypovolemia aggravated | 0
    cardiac arrest occurred | 0
    chest compression started | 0
    epinephrine 1 mg injected 4 times | 0
    aggressive volume resuscitation continued | 0
    spontaneous circulation recovered | 8
    normal sinus rhythm | 8
    serum potassium level elevated | 8
    serum calcium level decreased | 8
    hematocrit level decreased | 8
    significant oozing continued | 8
    surgical hemostasis | 8
    operator decided to stop surgery | 8
    intensive medical treatment | 8
    planned second operation | 8
    gauze packing | 8
    transferred to surgical ICU | 8
    crystalloid infused | 0
    5% albumin infused | 0
    colloid infused | 0
    leukocyte depleted red blood cell infused | 0
    leukocyte depleted platelet concentrate infused | 0
    cell saver blood infused | 0
    fresh frozen plasma infused | 0
    cryoprecipitate infused | 0
    urine output | 0
    estimated blood loss | 0
    metabolic acidosis | 24
    pH < 7.2 | 24
    azotemia | 24
    creatinine level over 2.0 mg/dl | 24
    ongoing graft failure | 24
    intractable bleeding | 24
    severe hypoxemia | 24
    mechanical ventilation | 24
    tidal volume 6 ml/kg | 24
    respiratory rate 30 breaths/minute | 24
    PEEP up to 10 cmH2O | 24
    chest radiography revealed pulmonary congestion | 24
    echocardiography | 24
    anuria developed | 7
    continuous renal replacement therapy started | 7
    brain tomography | 7
    no definite abnormal finding | 7
    failure of conventional ventilatory support | 24
    decision to initiate VV ECMO | 24
    normal heart function | 24
    no need of cardiac support with ECMO | 24
    existing central cannula removed | 24
    Swan-Ganz catheter removed | 24
    drainage cannula placed in right femoral vein | 24
    return cannula placed in right internal jugular vein | 24
    CAPIOX emergent bypass system primed | 24
    CRRT continued through ECMO circuit | 24
    VV ECMO circulation maintained | 24
    heparin not used | 24
    antithrombin injected | 24
    ACT measured | 24
    ACT maintained between 120-180 s | 24
    SpO2 95% | 24
    FiO2 0.3-0.4 at ventilator | 24
    FiO2 1.0 at ECMO | 24
    transferred to operating room for deceased donor LT | 24
    warm ischemic time 41 minutes | 24
    cold ischemic time 446 minutes | 24
    preoperative chest radiograph showed pulmonary congestion | 24
    bilateral pleural effusions | 24
    MELD score 30 | 24
    high risk of massive bleeding | 24
    decided to discontinue CRRT during operation | 24
    planned ECMO application | 24
    intubated | 24
    body temperature monitored | 24
    administered fluid heated | 24
    warm blanket | 24
    humidifier applied | 24
    limbs covered | 24
    room temperature maintained | 24
    SpO2 stable 97-100% | 24
    FiO2 0.5 at ventilator | 24
    ECMO flow 4-5 L/min | 24
    gas sweep 57-6 L/min | 24
    body temperature maintained | 24
    compartment syndrome concern | 24
    surgery finished without suturing abdominal wall | 24
    crystalloid administered | 24
    colloid administered | 24
    dextrose water administered | 24
    cell saver autotransfusion | 24
    leukocyte-depleted red blood cell infused | 24
    fresh frozen plasma infused | 24
    plateletpheresis infused | 24
    cryoprecipitate infused | 24
    no severe oozing | 24
    no acute massive bleeding | 24
    hematocrit level maintained over 24% | 24
    no rapid volume resuscitation | 24
    no hypotensive episode | 24
    no urine excreted | 24
    sedation maintained | 24
    CRRT restarted | 24
    ECMO continued | 24
    body temperature maintained | 24
    Glasgow coma scale tested | 24
    pupil size checked | 24
    light reflex checked | 24
    limb movement checked | 24
    orientation checked | 24
    pupil dilatation did not occur | 24
    light reflex normal | 24
    continuous sedation | 24
    muscular relaxation therapy with cisatracurium | 24
    arterial oxygen saturation improved | 64
    chest roentgenogram improved | 64
    sonography | 64
    improved coagulopathy | 64
    graft functional | 64
    hemodynamic stability achieved | 64
    norepinephrine tapered | 64
    recovery from hepatic failure | 64
    ECMO flow reduced to 3.0 L/min | 64
    oxygen flow reduced to zero | 64
    FiO2 increased to 0.6 | 64
    ABGAs showed appropriate oxygenation | 64
    ECMO removed | 64
    PaO2/FiO2 ratio improved | 64
    PaCO2 level similar | 64
    ventilatory demand decreased | 64
    PaO2/FiO2 stabilized | 64
    laparotomy wound closure | 120
    liver congestion noted | 120
    hepatic drainage failed | 120
    surgical decompression performed | 120
    stenosis at intrahepatic IVC developed | 120
    stenting performed | 168
    graft failure not improved | 168
    leg necrosis | 168
    sepsis | 168
    fentanyl stopped | 168
    cisatracurium stopped | 168
    continuous eye opening | 168
    low grade motor responses | 168
    no improvement of consciousness | 168
    expired | 576
    multi-organ failure | 576
    uncontrolled sepsis | 576
    