69 years old | 0
female | 0
breast cancer | -2520
radical surgery | -2520
high fever | -96
pain in right upper limb | -96
swelling in right upper limb | -96
admitted to hospital | 0
septic shock | 0
confused | 0
blood pressure 80/40 mmHg | 0
heart rate 105 beats/min | 0
breathing frequency 25 breaths/min | 0
armpit temperature 39°C | 0
peripheral oxygen saturation 94% | 0
WBC count 1.17×10^9/L | 0
platelet count 70×10^9/L | 0
hemoglobin 94 g/L | 0
neutrophils 85.5% | 0
IL-6 > 5000 pg/mL | 0
CRP 164.0 mg/L | 0
serum creatinine 158 µmol/L | 0
mild edema of upper arm and forearm | 0
vascular color ultrasound of extremities normal | 0
empirical meropenem | 0
vancomycin | 0
norepinephrine | 0
rehydration | 0
low-molecular-weight heparin | 0
drugs for raising platelets | 0
topical magnesium sulfate | 0
procalcitonin decreased to 9.47 pg/mL | 24
mNGS results indicated SDSE | 24
cyanosis of fingers and toes | 48
large purpura on skin | 48
large blisters | 48
liver function tests showed steep rise in transaminases | 72
progression of limb end ischemia | 72
blood cultures showed SDSE | 72
Streptococcus isolated from blood | 72
hypotension | 72
multiple organ dysfunction | 72
coagulation dysfunction | 72
liver function dysfunction | 72
renal function dysfunction | 72
blister formation | 72
limb gangrene | 72
STSS diagnosed | 72
drug sensitivity results | 72
ceftriaxone | 72
anisodamine | 72
transferred from ICU to general ward | 240
ischemia at extremities worsened | 240
amputation performed | 240
SPG developed | 240