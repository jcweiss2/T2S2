79 years old| 0
    male | 0
    acute abdominal pain | -72
    HPVG detected by abdominal CT | -24
    transferred to our hospital | -24
    no remarkable past medical history | 0
    body temperature: 37.2°C | 0
    blood pressure: 112/74 mmHg | 0
    pulse rate: 68 beats/min | 0
    abdominal distention | 0
    rebound tenderness | 0
    abdominal guarding | 0
    peritoneal irritation | 0
    white blood cell count of 18,400/μL | 0
    C-reactive protein concentration of 17.7 mg/dL | 0
    dehydration | 0
    metabolic acidosis | 0
    base excess of −7.0 mmol/L | 0
    creatine kinase elevated (28,327 IU/L) | 0
    distention of the small intestine | 0
    subileus | 0
    contrast defect in a region of the small intestine | 0
    small amount of ascites around the intestine | 0
    no thrombus in any artery | 0
    wall of the appendix moderately thickened | 0
    urgent laparotomy | 0
    generalized peritonitis caused by intestinal necrosis | 0
    small amount of turbid ascites | 0
    dilated small intestine | 0
    no intestinal ischemia detected | 0
    discoloration of the appendix with wall thickening | 0
    gangrenous appendicitis | 0
    no macroscopic perforation observed | 0
    appendectomy | 0
    abdominal drainage | 0
    pathological diagnosis of gangrenous appendicitis | 0
    no evidence of malignancy | 0
    Escherichia coli in ascitic culture | 0
    intravenous antibiotic treatment (meropenem) | 0
    septic shock | 24
    DIC | 24
    admitted to ICU | 24
    blood purification therapy | 24
    HPVG disappeared | 168
    left ICU | 168
    discharged from hospital | 312
    
    