63 years old | 0
male | 0
170cm tall | 0
69kg | 0
admitted to the hospital | 0
epigastric bloating | 0
discomfort | 0
history of extensive smoking | -672
hypertension | -672
chronic kidney disease | -672
Child C liver disease | -672
portal hypertension | -672
ascites | -672
oesophageal varices | -672
gastropathy | -672
treated with antibiotics | 0
ascitic drainage | 0
culture-negative neutrocystic ascites | 0
developed acute severe abdominal pain | 624
computed-tomography abdominal and pelvis investigation | 624
perforated duodenal ulcer | 624
exploratory laparotomy | 624
roux loop mucosal patch | 624
transferred to the surgical intensive care unit (ICU) | 624
ventilatory and haemodynamic support | 624
high intra-abdominal pressure | 672
oliguric acute kidney impairment | 672
abdominal compartment syndrome | 672
managed medically with paralysis | 672
renal replacement therapy | 672
duodeno-jejunal anastomotic leak | 840
second exploratory laparotomy | 840
tube diversion | 840
primary repair of the wound dehiscence pedicled omentoplasty | 840
definitive surgery | 960
primary exclusion | 960
roux loop gastrojejunostomy | 960
significant blood loss | 960
received packed red cells | 960
received pooled platelets | 960
received fresh frozen plasma | 960
noradrenaline infusion | 960
ventilatory support | 960
difficult ventilation | 962
peak pressure rose | 962
end-tidal carbon dioxide rose | 962
paralysed with atracurium | 962
sedated with propofol | 962
ventilator pressure-time curve demonstrated increased peak and plateau pressures | 962
chest was clear bilaterally | 962
generalised poor air entry throughout | 962
multiple endotracheal tube suctioning | 962
arterial blood gas | 962
pH 6.99 | 962
pCO2 106mmHg | 962
pO2 125mmHg | 962
base excess -6 | 962
chest X-ray | 962
intra-abdominal pressure 31mmHg | 962
noradrenaline increased | 962
vasopressin started | 962
haemoglobin dropping | 962
intra-abdominal haemorrhage suspected | 962
abdominal compartment syndrome suspected | 962
fourth exploratory laparotomy | 984
small amount of intra-abdominal bleeding | 984
blood clots | 984
moderate generalised bowel oedema | 984
opening of the peritoneum | 984
improvement in ventilation | 984
improvement in haemodynamics | 984
Ppeak improved | 984
tidal volume improved | 984
vasopressin stopped | 984
noradrenaline weaned | 984
post-operatively improved | 984
Ppeak remained high | 984
respiratory acidosis persisted | 984
intra-abdominal pressure improved | 984
arterial blood gas | 984
pH 7.164 | 984
pCO2 72.8mmHg | 984
pO2 152mmHg | 984
BE -4 | 984
bedside bronchoscopy | 984
large mucus plug found | 984
endotracheal tube exchanged | 984
immediate improvement in Ppeak | 984
noradrenaline stopped | 984
arterial blood gases | 985
pH 7.42 | 985
pCO2 39.1mmHg | 985
pO2 76.1mmHg | 985
BE 0.5 | 985
gastrointestinal bleeding | 1200
breakdown of the surgical anastomosis | 1200
overwhelming sepsis | 1200
multiorgan failure | 1200
died | 1200