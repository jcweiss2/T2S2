53 years old | 0
male | 0
admitted to the hospital | 0
altered mental status | 0
hypotension | 0
fever | 0
respiratory distress | 0
diabetic nephropathy | -672
renal replacement therapy | -672
diabetic retinopathy | -672
bilateral amaurosis | -672
cardiac arrest | 0
acute respiratory failure | 0
cardiopulmonary resuscitation | 0
return to spontaneous blood circulation | 0
orotracheal intubation | 0
normocytic normochromic anemia | 0
mixed hyperbilirubinemia | 0
conserved renal function | 0
no electrolyte disorders | 0
CT angiography negative for pulmonary embolism | 0
positive polymerase chain reaction for SARS-CoV-2 | 0
respiratory distress | 0
fever | 0
no vaccination | 0
unknown COVID-19 variant | 0
somnolent but alertable | 1
obeying simple orders | 1
intact brainstem reflexes | 1
normal motor function | 1
normal sensitive function | 1
brain CT | 1
supratentorial bilateral frontal leukoencephalopathy | 1
small vessel disease | 1
calcified atheromatous plaques | 1
no other abnormalities | 1
deterioration of mental status | 24
stupor | 24
severe hypoglycemia | 24
glucose levels of 18 mg/dl | 24
MRI | 24
symmetric focal high intensity signals in T2-weighted images | 24
symmetric focal high intensity signals in FLAIR | 24
symmetric focal high intensity signals in DWI | 24
bilateral middle cerebellar peduncles | 24
hypoglycemic encephalopathy | 24
glucose level normalization | 48
improvement of mental status | 48
multiple comorbidities | 72
worsen respiratory status | 72
stop all invasive interventions | 72
end-of-life symptom management order protocol | 72
death | 96