73 years old | 0
woman | 0
vaginal vault cancer stage 4 | 0
received 10 fractions of palliative RT to the vagina | 0
received 1 cycle of chemotherapy | 0
doing well at home until one week before her admission | -168
presented to the emergency room | 0
complaints of shortness of breath | 0
fever | 0
constipation | 0
generalized weakness | 0
unresponsiveness | 0
oxygen saturation was 89% on room air | 0
temperature 101.9F | 0
respiratory rate of 24 | 0
heart rate of 140 | 0
blood pressure measuring 110/65 | 0
purple urinary bag in one of the PCN stents | 0
PCN stents placed 4 months ago | -2928
history of bilateral hydroureteronephrosis | -2928
chronic kidney disease | -2928
impingement of vaginal vault mass on both the ureters | -2928
history of acute renal failure | -2928
underlying tumour (post-renal acute kidney failure) | -2928
catheter bag with <50 mL of urine output | 0
Karnofsky performance status 40 | 0
family noticed a colour change 3 days ago | -72
provisional diagnosis of PUBS | 0
purple colour throughout the bag on visual examination | 0
high white blood cell count of 16,760/mm3 | 0
urinary pH 7.5 | 0
moderate leukocytes in the urine | 0
tested positive for nitrates | 0
tested positive for leucocyte esterase |B0
no trace of ingestion of medications/food items | 0
no trace of poisonous materials | 0
no haematuria | 0
no porphyria | 0
started on empirical IV cefoperazone and sulbactam combination | 0
started on levofloxacin 500 mg | 0
other supportive medications | 0
urine culture grew Escherichia coli >105 CFU/mL | 0
urine culture grew Klebsiella spp. | 0
gram-negative bacteremia | 0
urine discolouration subsided | 120
no clinical improvement | 120
disease burden | 120
ongoing sepsis | 120
multi-organ failure | 120
advanced nature of the disease | 120
poor prognosis | 120
decision for no aggressive treatment | 120
preferred palliative intent | 120
delirious | 120
increased breathlessness | 120
fever spikes | 120
condition gradually deteriorated | 120
expired | 144
discharged | 144
