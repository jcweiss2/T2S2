65 years old | 0
    male | 0
    presented to the emergency | 0
    multiple blisters | 0
    erosions all over body | 0
    oral mucosa involvement | 0
    scalp involvement | 0
    superadded maggot infection | -4320
    previous episodes of lesions | -8640
    lesions subsided | -8640
    treatment with steroids | -8640
    unknown generic medications | -8640
    lesions developed over 6 months | -4320
    lesions worsened | -4320
    brought to tertiary hospital | 0
    febrile | 0
    numerous flaccid blisters | 0
    erosions covering >85% body surface area | 0
    slough present | 0
    maggots present | 0
    Nikolsky sign positive | 0
    PV diagnosis confirmed by skin biopsy | 0
    PV diagnosis confirmed by Tzanck smear | 0
    intravenous dexamethasone pulse (120 mg) | 0
    supportive care (fluids) | 0
    supportive care (FFP) | 0
    supportive care (dressings) | 0
    routine blood investigation normal | 0
    blood culture sterile | 0
    urine culture sterile | 0
    intravenous antibiotics (Piperacillin/Tazobactam) | 0
    intravenous antibiotics (Teicoplanin) | 0
    pus culture sensitivity | 0
    adjuvant immunosuppressors held back due to infection | 0
    extensive lesions | 0
    high susceptibility to infections | 0
    shifted to isolation ICU | 0
    oozing from skin ulcerations | 0
    hemorrhagic excoriation | 0
    peeling of skin | 0
    oral methyl prednisolone (1 mg/kg) | 0
    no improvement in skin lesions | 0
    general condition worsened | 168
    hypoproteinemia | 168
    pleural effusion | 168
    blood culture showed enterobacter | 168
    pus culture showed Staphylococcus aureus | 168
    pus culture showed Proteus mirabilis | 168
    intravenous Tigecycline | 168
    intravenous Vancomycin | 168
    erosions persisted | 168
    no re-epithelialization | 168
    perilesional Nikolsky sign positive | 168
    new blisters developed | 168
    sepsis | 168
    persistent high grade fever | 168
    albumin levels fell to 2.1 mg | 168
    hold IV methyl prednisolone pulse therapy | 168
    hold cyclophosphamide | 168
    TPE cycle planned | 168
    TPE performed | 168
    plasma exchange with cell separator | 168
    femoral access with dialysis catheter | 168
    TPE scheduled alternate-day intervals | 168
    five sessions over 10 days | 168
    anticoagulation with citrate (ACD) | 168
    replacement with isotonic saline | 168
    replacement with 4% human albumin | 168
    replacement with FFP | 168
    monitoring hemodynamic parameters | 168
    complications monitored and reverted | 168
    calcium gluconate administered | 168
    hemogram monitored | 168
    serum electrolytes monitored | 168
    total protein monitored | 168
    albumin monitored | 168
    Nikolsky sign negative after third TPE | 264
    no new lesions after third TPE | 264
    exudation reduced | 264
    dressings remained dry | 264
    60-70% re-epithelialization | 264
    90% healing after last TPE | 408
    oral lesions healed completely | 408
    erosions on back persisted | 408
    erosions on anterior thigh persisted | 408
    erosions on buttocks persisted | 408
    IV methyl prednisolone (1 g/day) | 408
    cyclophosphamide (500 mg/day) | 408
    Pulse therapy for three days | 408
    further improvement in lesions | 408
    clinically stable | 408
    plan for more TPE cycles | 408
    cost restraint prevented TPE | 408
    discharged | 408
    monthly IV dexamethasone pulse | 408
    oral prednisolone (60 mg/day) | 408

    