55 years old|0
    male|0
    experienced a trivial fall|0
    severe back pain|0
    analgesics|-48
    bed rest|-48
    pain relieved|-48
    back pain gradually increased|0
    incapacitated from routine activities|0
    persistent back pain|0
    restriction of movements|0
    gibbus at thoracolumbar junction|0
    spasm of para-spinal muscles|0
    restricted spine movements|0
    painful spine movements|0
    normal motor power|0
    normal sensation distally|0
    intact reflexes|0
    normal bladder function|0
    normal bowel function|0
    anorexia|0
    loss of weight|0
    well-controlled type-2 diabetes|0
    surgical fixation of humerus fracture|0
    no smoking|0
    no alcohol use|0
    no childhood illnesses|0
    raised CRP|0
    raised ESR|0
    high normal white cell count|0
    normal bone profile|0
    normal renal function|0
    normal liver function|0
    T12 compression fracture|0
    marrow edema|0
    fluid in fracture site|0
    prevertebral soft-tissue swelling|0
    epidural soft-tissue component|0
    differential diagnosis of tumor|0
    pseudoarthrosis|0
    infection|0
    osteopenic|0
    T-score -2|0
    intact posterior cortex|0
    severe unremitting pain|0
    osteoporotic fracture|0
    metastasis|0
    transpedicular biopsy|0
    kyphoplasty|0
    general anesthesia|0
    prone position|0
    transpedicular biopsy needles inserted|0
    minimal resistance|0
    no initial aspiration material|0
    saline injected|0
    sero-sanguineous material|0
    pus|0
    microbiology sent|0
    cytology sent|0
    fluid analysis sent|0
    infection suspected|0
    kyphoplasty deferred|0
    extubation|0
    severe bronchospasm|0
    decreased saturation|0
    inability to maintain tidal volume|0
    intubation|0
    respiratory acidosis|0
    pH 7.16|0
    PaCO2 72 mm Hg|0
    PaO2 82 mm Hg|0
    bilateral lung infiltrates|0
    mechanical ventilation|0
    PaO2/FiO2 205|0
    progression of pulmonary edema|0
    multifocal infiltrates|0
    pleural fluid|0
    intravenous vancomycin|0
    improved after 24 hours|24
    ventilator weaning|24
    endo-tracheal tube detached|48
    high dependency unit|48
    chest clear|72
    infiltrates resolved|72
    Staphylococcus aureus culture|72
    imipenum sensitive|72
    linezolid sensitive|72
    bronchial lavage culture|72
    pleural fluid culture|72
    endotracheal tube culture|72
    negative blood culture|72
    septic pulmonary emboli|72
    intravenous linezolid|72
    oral linezolid|72
    thoracolumbar orthosis|72
    CRP normalization|72
    ESR normalization|72
    symptom free|432
    uneventful recovery|432
    