57 years old | 0
Hispanic | 0
male | 0
admitted to the hospital | 0
history of coronary artery disease | -3024
history of myocardial infarction | -3024
history of ischemic dilated cardiomyopathy | -3024
pocket infection of cardiac resynchronization therapy defibrillator | 0
initial device and leads implanted | -7776
generator change | -432
2-month history of erythema | -1440
discomfort around left upper chest implant site | -1440
edema | -1440
serosanguinous drainage | -1440
oral amoxicillin treatment | -1440
nonbacteremic | 0
afebrile | 0
laboratory investigations within normal limits | 0
echocardiography revealed severely reduced left ventricular systolic function | 0
ejection fraction of 20%–25% | 0
global hypokinesis of the left ventricle | 0
no evidence of vegetations | 0
preoperative computed tomography revealed leads scarred to lateral wall of superior vena cava | 0
transvenous lead extraction | 0
cardiac resynchronization therapy defibrillator pocket capsule dissected out | 0
device removed | 0
coronary sinus and right atrial leads extracted | 0
right ventricular lead extracted with laser assistance | 0
patient became hypotensive | 0
transesophageal echocardiography revealed large pericardial effusion | 0
emergency midsternotomy performed | 0
pericardium opened | 0
significant amount of blood seen | 0
bleeding manually controlled with pressure | 0
cardiopulmonary bypass instituted | 0
5-mm tear in superior cavoatrial junction located | 0
perforation in right atrium located | 0
oozing hematoma at level of innominate vein located | 0
lesions repaired with multiple 4-0 polypropylene sutures | 0
right ventricular lead capped and abandoned | 0
intra-aortic balloon pump placed | 0
multiple blood transfusions | 0
coagulopathy developed | 0
transfusions of cryoprecipitate, platelets, fresh frozen plasma, and factor VII | 0
chest closed | 0
transferred to intensive care unit | 0
severe cardiogenic shock | 0
multiorgan failure | 0
hypotensive | 0
required large doses of vasopressin, epinephrine, and norepinephrine | 0
hypoxic respiratory failure | 0
mechanical ventilation | 0
liver failure | 0
albumin and multiple blood products given | 0
broad-spectrum antibiotics adjusted | 0
oliguric | 0
continuous venovenous hemodialysis for acute renal failure | 24
bilateral, symmetrical cyanotic changes to all 5 digits of upper and lower extremities | 48
vasopressor administration stopped | 48
upper- and lower-digit ischemia progressed to dry gangrene | 216
dull pain | 216
no ability to move fingers and toes | 216
bilateral stiffness | 216
2+ pitting edema | 216
nonexistent capillary refill time | 216
palpable 2+ peripheral pulses | 216
Doppler study showed flat waveforms on all digits and toes bilaterally | 216
intra-aortic balloon pump removed | 168
endotracheal tube removed | 168
albumin discontinued | 264
liver enzymes returned to normal limits | 264
kidney function gradually improved | 984
hemodialysis stopped | 984
mental status improved | 984
necrotic lesions treated conservatively with povidone-iodine dressings | 648
debridement | 648
negative-pressure wound therapy | 648
purulent, foul-smelling material drained from left infraclavicular operative site | 1296
transferred to facility for further management of pocket infection | 1296
preoperative transesophageal echocardiography revealed diminished ejection fraction | 1296
laser extraction of retained lead | 1308
pus drained from subfascial area | 1308
antibiotic regimen started | 1308
microbial cultures grew Enterobacter cloacae and Staphylococcus epidermidis | 1308
transvenous implantable cardioverter-defibrillator system implanted | 1312
evaluation of hands and feet revealed no signs of local infection or wet gangrene | 1312
black skin changes and demarcation lines clearly defined | 1312
frank mummification of digits and toes | 1312
discharged to home health services | 1848
amputation and debridement of necrotic feet | 2544
amputation of fingers scheduled | 2544