61 years old | 0
male | 0
admitted to the hospital | -120
acute abdominal pain | -120
fever | -120
perforated duodenal ulcer | -120
sepsis | -120
primary surgical closure | -120
right internal jugular vein catheterization | -120
intensive care unit treatment | -120
transferred to general ward | -96
CVC removal | 0
shortness of breath | 0
chest discomfort | 0
unconscious | 0
cardiopulmonary resuscitation | 0
return of spontaneous circulation | 5
transthoracic echocardiogram | 5
multiple air bubbles in right and left ventricles | 5
ostium secundum atrial septal defect | 5
right-to-left shunt | 5
brain computed tomography | 5
gas within centrum semiovale | 5
gas within cerebral sulci | 5
gas within cavernous sinuses | 5
free air in neck | 5
free air in jugular vein | 5
free air in left ventricle | 5
transferred to our hospital | 6
blood pressure 107/75 mmHg | 6
heart rate 134 beats/min | 6
respiratory rate 30 breaths/min | 6
temperature 35.8°C | 6
Glasgow coma scale 3/15 | 6
no brain stem reflex | 6
chest X-ray | 6
extensive bilateral infiltrates | 6
pulmonary edema | 6
arterial blood gas analysis | 6
pH 7.141 | 6
PaCO2 52.3 mmHg | 6
PaO2 53.6 mmHg | 6
HCO3 14.8 mEq/L | 6
SaO2 74% | 6
venovenous ECMO support | 6
mechanical ventilation | 6
FiO2 1.0 | 6
pulmonary edema ameliorated | 120
lung injury ameliorated | 120
weaned off ECMO support | 168
ejection fraction of left ventricle preserved | 72
no regional wall motion abnormalities | 72
apical left ventricle thrombus | 72
anticoagulation therapy | 72
acute renal failure | 6
improved without hemodialysis | 168
diffuse cerebral ischemia | 168
brain magnetic resonance imaging | 168
tracheostomy | 168
transferred to general ward | 168