89 years old|0
female|0
referred to medical center with loss of consciousness|0
sudden LOC|0
admitted to emergency department via ambulance|0
loss of consciousness|-0.5
dry cough|-48
body aches|-48
no comorbidity|0
no drug history|0
no alcohol history|0
no smoking history|0
no allergy|0
vaccinated twice with Sinopharm vaccine|0
GCS score three|0
oral temperature 36.5°C|0
normal vital signs|0
oxygen saturation 98%|0
elevated lactate dehydrogenase|0
elevated C-reactive protein|0
elevated ESR|0
elevated CPK|0
elevated urea|
