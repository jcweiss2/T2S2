52 years old | 0
male | 0
admitted to the hospital | 0
general weakness | -240
right upper quadrant pain | -96
diagnosed with PC-type MCD | -4380
computed tomography (CT) scans | -4380
right axillary lymph node biopsy | -4380
chemotherapy | -4380
loss to follow-up | -4380
smoking history | -4380
contrast-enhanced CT scan | 0
acute calculous cholecystitis | 0
lymphadenopathy | 0
splenomegaly | 0
bilateral pleural effusion | 0
ascites | 0
anemia | 0
thrombocytopenia | 0
lymphopenia | 0
azotemia | 0
stress-induced cardiomyopathy | 0
percutaneous transhepatic gallbladder drainage | 0
serum immunofixation electrophoresis | 0
polyclonal hypergammaglobulinemia | 0
bone marrow study | 0
plasmacytosis | 0
reductions in platelet count | 0
reductions in hemoglobin (Hgb) | 0
reductions in lymphocyte | 0
reductions in total cholesterol | 0
reductions in albumin | 0
increases in international normalized ratio (INR) | 0
increases in blood urea nitrogen | 0
increases in creatinine | 0
increases in C-reactive protein (CRP) | 0
increases in erythrocyte sedimentation rate (ESR) | 0
increases in vascular endothelial growth factor (VEGF) | 0
chemotherapy | 0
pulmonary edema | 168
dyspnea | 168
oliguria | 168
aggressive treatment | 168
intensive care unit (ICU) | 168
echocardiography | 552
normalization of left ventricular systolic function | 552
improvements in pulmonary edema | 552
improvements in azotemia | 552
transfusions of leukocyte-poor and irradiated packed red blood cells (RBC) | 552
transfusions of platelets | 552
transfusions of fresh frozen plasma (FFP) | 552
elective laparoscopic cholecystectomy | 720
preanesthetic evaluation | 720
blood transfusion | 720
physical examination | 720
abdominal distension | 720
chest X-ray | 720
pulmonary function test | 720
electrocardiogram (ECG) | 720
thoracic CT scan | 720
modified Allen's test | 720
arterial pressure monitoring | 720
arterial blood gas sampling | 720
FloTrac/Vigileo monitor | 720
preoxygenation | 720
general anesthesia | 720
tracheal tube insertion | 720
sevoflurane | 720
remifentanil | 720
central venous oximetry catheter | 720
surgery | 720
Calot's triangle | 720
inflammation | 720
adhesion | 720
open cholecystectomy | 720
perioperative drainage of ascites | 720
cisatracurium | 720
ephedrine | 720
vital signs monitoring | 720
Vigileo monitor | 720
bispectral index | 720
arterial blood gas analysis (ABGA) | 720
surgery completion | 750
anesthesia termination | 750
tracheal tube removal | 750
ICU | 750
postoperative vital signs | 750
postoperative laboratory findings | 750
general ward | 750
chemotherapy | 750
cough | 4320
sputum | 4320
fungal pneumonia | 4320
treatment | 4320
deterioration | 4320
ventilator care | 4320
ICU | 4320
expiration | 4320