88 years old | 0
male | 0
admitted to the hospital | 0
skin color change in the right scrotal area | 0
right scrotal pain | -168
right scrotal swelling | -168
red skin color change in the right scrotal area | -24
skin color changed from red to black with foul-smelling | -24
voiding dysfunction | -6048
benign prostatic hyperplasia | -6048
a-blocker | -6048
5 alpha reductase inhibitor | -6048
Memokath 028 implantation | -6048
refractory to medical therapy for LUTS with BOO | -6048
TURP | -6048
high ASA score | -6048
NSTEMI | -6048
cerebrovascular accident | -6048
poor-controlled COPD | -6048
spinal stenosis | -6048
MIS under local anesthesia | -6048
intraurethral lidocaine injection | -6048
analgesic injection intravenously | -6048
Qmax improved | -1304
residual urine volume decreased | -1304
suprapubic cystostomy | -2880
acute urinary retention | -2880
Memokath 028 not working | -2880
broad-spectrum antibiotics | 0
meropenem | 0
vancomycin | 0
clindamycin | 0
necrotic tissues excised | 24
right orchiectomy | 24
necrotic change of right spermatic cord and epididymis | 24
Memokath 028 stent removed | 24
culture swab in open wound | 24
erythematous change of prostatic urethra | 24
mechanical ventilation | 24
total parenteral nutrition | 24
hemodialysis | 48
incomplete surgical debridement | 48
necrotic tissues debrided | 72
elevated liver enzyme and bilirubin level | 288
total platelet count decreased | 312
prothrombin time and international normalized ratio prolonged | 312
died | 336
Fournier’s gangrene | 0
acute prostatitis | 0
sepsis | 0
multiorgan failure | 0
Enterobacter cloacae isolated | 0
urine analysis | 0
pyuria | 0
procalcitonin level elevated | 0
serum lactate level elevated | 0
serum creatinine level elevated | 0
serum glucose level elevated | 0
abdominal-pelvic enhanced computed tomography | 0
emphysematous changes | 0
inflammatory infiltration | 0
prostatic urethral stent observed | 0
necrotic skin lesion | 0
tenderness and heat of entire prostate | 0
white blood cell count elevated | 0
C-reactive protein level elevated | 0
digital rectal examination | 0
Fournier’s gangrene severity index | 0
broad-spectrum antibiotics administration | 0
surgical debridement | 24
necrotic tissues with foul-smelling fluid excised | 24
right orchiectomy performed | 24
Memokath 028 stent removed | 24
culture swab in prostatic stent | 24
antibiotics susceptibility | 24
incomplete surgical debridement | 48
necrotic tissues debrided | 72
elevated liver enzyme and bilirubin level | 288
total platelet count decreased | 312
prothrombin time and international normalized ratio prolonged | 312
died | 336