60 years old | 0
woman | 0
admitted to the hospital | 0
epilepsy | -120
unwitnessed fall | -120
3-cm laceration on the medial aspect of her forehead | -120
CT of the head without contrast | -120
nausea | -96
vomiting | -96
diarrhea | -96
generalized weakness | -96
severe fatigue | -96
seizure-like activities | -96
altered mental status | -96
diffuse shaking movements | -96
non-specific headaches | -168
low back pain | -168
neck pain | -168
hearing loss | -168
hallucinations | -96
chronic obstructive pulmonary disease | 0
hypertension | 0
hyperlipidemia | 0
depression | 0
anxiety | 0
migraines | 0
multiple sclerosis | 0
immunosuppressive therapy with fingolimod | 0
temperature of 37.6 °C | 0
heart rate of 110 bpm | 0
blood pressure of 191/84 mm Hg | 0
respiratory rate of 16 breaths per minute | 0
oxygen saturation of 97% | 0
bilateral periorbital ecchymosis | 0
small forehead laceration with sutures | 0
surrounding ecchymosis and bruising | 0
tachycardia | 0
regular rhythm | 0
no murmurs | 0
no rubs | 0
no gallops | 0
lungs clear | 0
no wheezing | 0
no rales | 0
no rhonchi | 0
fluent speech | 0
no aphasia | 0
cranial nerves II-XII intact | 0
5/5 muscle strength | 0
intact sensation | 0
normal reflexes | 0
negative Babinski sign | 0
no dysmetria | 0
no nuchal rigidity | 0
negative Kernig maneuver | 0
negative Brudzinski maneuver | 0
hemoglobin 11.4 g/dL | 0
hematocrit 32.7% | 0
white blood cell 20.8 × 103/µL | 0
platelets 141 × 103/µL | 0
sodium 128 mEq/L | 0
potassium 2.5 mEq/L | 0
chloride 88 mEq/L | 0
creatinine 0.64 mg/dL | 0
blood urea nitrogen 12 mg/dL | 0
calcium 8.9 mg/dL | 0
glucose 200 mg/dL | 0
lactic acid 2.2 mmol/L | 0
cardiac high-sensitivity troponin T 0.03 ng/mL | 0
ECG sinus tachycardia | 0
diffuse non-specific ST-segment depression | 0
CT scan of the head without contrast | 0
small frontal scalp hematoma | 0
MRI of brain and brainstem | 0
progressive periventricular white matter lesions | 0
blood cultures obtained | 0
back pain | 24
nausea | 24
vomiting | 24
photosensitivity | 24
EEG diffuse slowing | 24
encephalopathy | 24
obtunded | 48
unable to follow commands | 48
repeat head and neck images unremarkable | 48
blood cultures heavy growth of yeast | 48
concern for cryptococcal meningitis | 48
lumbar puncture performed | 48
started on amphotericin | 48
CSF WBC count 0 | 48
CSF RBC count 2434 cells | 48
CSF total protein 58 mg/dL | 48
CSF glucose 3 mg/dL | 48
CSF Cryptococcus antigen positive | 48
blood cultures confirmed Cryptococcus neoformans | 48
flucytosine added | 48
unresponsive | 96
hypoxic | 96
endotracheal intubation | 96
bradycardic | 96
cardiac arrest | 96
advance cardiac life support initiated | 96
ROS achieved | 96
troponin 1.43 ng/mL | 96
ECG Q waves anteriorly | 96
poor R wave progression | 96
ST-segment elevations in leads V1 to V4 | 96
echocardiogram ejection fraction 20-25% | 96
hypokinesis of anterior, anteroseptal, and apical segments | 96
basal hyperkinesis | 96
Takotsubo cardiomyopathy | 96
CT angiogram of the chest | 96
no significant coronary calcifications | 96
hemodynamic instability | 96
dual vasopressor support | 96
norepinephrine | 96
epinephrine | 96
continued clinical decline | 96
increasing vasopressors | 96
significant ventilator support | 96
no cough reflexes | 96
no corneal reflexes | 96
no pharyngeal reflexes | 96
decision for comfort care | 96
patient passed away | 96
