33 years old | 0
female | 0
admitted to the hospital | 0
history of headache | -1200
history of myalgia | -1200
history of nausea | -1200
history of vomiting | -1200
evaluated elsewhere | -1200
treated for migraine | -1200
intermittent episodes of hypotension | -720
persistent leucocytosis | -720
treated with multiple courses of empirical broad-spectrum antibiotics | -720
developed anasarca | -720
no history of hematuria | 0
no reduction in urine output | 0
afebrile | 0
blood pressure 110/70 mmHg | 0
no postural hypotension | 0
systemic examination unremarkable | 0
nephrotic range proteinuria | 0
microscopic hematuria | 0
hypoalbuminemia | 0
hypercholesterolemia | 0
hypertriglyceridemia | 0
serum creatinine 1.08 mg/dl | 0
leucocytosis | 0
neutrophil 71% | 0
lymphocyte 19% | 0
eosinophil 3% | 0
monocyte 6% | 0
basophil 1% | 0
anti-nuclear antibody negative | 0
anti-double stranded deoxyribonucleic acid antibody negative | 0
Complement C3c and C4 levels normal | 0
started on diuretics | 0
started on intravenous albumin | 0
blood culture did not grow any pathogen | 0
renal biopsy | 0
mild increase in mesangial matrix | 0
mesangial hypercellularity | 0
immunofluorescence study negative | 0
diagnosis of idiopathic unsampled focal and segmental glomerulosclerosis | 0
started on prednisolone | 0
electron microscopy | 0
mesangial proliferative glomerulonephritis | 0
mesangial electron dense deposits | 0
discharged | 0
myalgia | 120
giddiness | 120
weakness | 120
tachycardia | 120
tachypnea | 120
hypotension | 120
worsening leucocytosis | 120
neutrophilic predominance | 120
elevated serum procalcitonin levels | 120
broad-spectrum antibiotic coverage | 120
intravenous meropenem | 120
total leucocyte count increased | 144
imaging of chest and abdomen | 144
no focus of sepsis | 144
managed in the intensive care unit | 144
meropenem | 144
inotropic support | 144
clinical improvement | 216
reduction of inotropic requirement | 216
normalization of the total leucocyte count | 216
blood culture grew non-O1, non-O139 V. cholerae | 216
sensitive to ampicillin | 216
sensitive to tetracycline | 216
sensitive to cotrimoxazole | 216
sensitive to cefotaxime | 216
sensitive to ofloxacin | 216
sensitive to meropenem | 216
stool culture did not grow any pathogen | 216
visited a beach for swimming and bathing | -1344
exposure to sea-water | -1344
consumed no sea-food | -1344
completed 2 weeks of meropenem | 336
repeat blood culture documented to be sterile | 336
discharged in stable condition | 336
advice to continue prednisolone | 336