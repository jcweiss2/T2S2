101 years old | 0
male | 0
admitted to the hospital | 0
cough | -24
productive sputum | -24
wheezing | -24
hypertension | 0
coronary artery disease | 0
old cerebral infarction |>0
diabetes mellitus | 0
WBC 9.28×109/L | 0
neutrophils 80.4% | 0
lymphocytes 11.3% | 0
CRP 2.67 mg/dl | 0
Procalcitonin <0.05 ng/mL | 0
CT scan showed new patchy ground glass opacities in the right upper lung and right middle lobe | 0
community acquired pneumonia | 0
flomoxef | 0
levofloxacin | 0
fever 38.3°C | 48
adenovirus IgM positive | 48
adenovirus | 48
meropenem | 48
tigecycline | 48
persistent fever | 0
lethargy | 0
thrombocytopenia | 0
elevated creatinine | 0
elevated transaminase levels | 0
PCT peak at 1.78 ng/mL | 0
vancomycin | 0
piperacillin/tazobactam | 0
respiratory failure | 864
CT scan showed new bilateral patchy infiltrates | 864
CT scan showed lung cavity (7 mm × 8 mm) in the anterior segment of the left upper lobe | 864
bronchoscopy | 864
yellowish-white secretion in left main bronchus | 864
edematous and congested mucosa | 864
bronchoalveolar lavage | 864
mNGS revealed E. faecium | 864
BALF culture confirmed E. faecium | 864
vancomycin-resistant | 864
linezolid-sensitive | 864
linezolid 600 mg IV q12d | 864
clinical improvement | 864
thrombocytopenia (platelets 44 ×109/L) | 864
linezolid discontinued | 864
contezolid 400 mg PO q12d | 864
thrombopoietin | 864
platelet counts returning to normal | 864
cavitary lesion resolved | 864
decreased patchy infiltrations in the left upper lobe | 864
nearly 4-month course of contezolid therapy | 864
follow-up CT scan showed disappearance of lung cavity lesion and patchy infiltrations | 864
discharged | 0
