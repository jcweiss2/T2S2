68 years old | 0
male | 0
diabetes mellitus type II | -672
hypertension | -672
chronic kidney disease stage 5 | -672
heart failure with preserved ejection fraction | -672
admitted to the hospital | 0
shortness of breath | 0
generalized body aches | 0
worsening of kidney function | 0
diuretic therapy | 0
hemodialysis | 264
hypotensive | 528
lethargic | 528
decrease in urine output | 528
shifted to the MICU | 528
bolus of crystalloids | 528
norepinephrine infusion | 528
echo | 528
moderate pericardial effusion | 528
subcostal approach | 528
coagulopathy | 528
hepatomegaly | 528
apical approach | 528
INR 1.7 | 528
Fresh Frozen Plasma (FFP) | 528
increased vasopressors requirements | 552
lactate 8 mmol/L | 552
anuric | 552
continuous renal replacement therapy | 552
liver enzymes increased | 552
alanine aminotransferase 1729 U/L | 552
aspartate aminotransferase 1772 U/L | 552
INR 2 | 552
diagnosed with acute ischemic hepatitis | 552
coagulopathy | 552
emergency pericardiocentesis | 552
FFP | 552
vitamin K | 552
advanced cardiac monitoring device | 552
cardiac index 0.9 L/min/m2 | 552
systemic vascular resistance > 4000 dynes/sec/cm5 | 552
cardiogenic shock | 552
cardiac tamponade | 552
repeated coagulation profile | 552
INR 2.3 | 552
activated prothrombin complex concentrate (FEIBA) | 552
coagulation profile repeated | 556
INR 1.9 | 556
pre-pericardiocentesis echo | 556
pericardiocentesis | 556
60 mL of fluid drained | 556
asystole cardiac arrest | 580
cardiopulmonary resuscitation | 580
death | 596