56 years old | 0
    African American female | 0
    presented to the Emergency Department | -144
    swelling over left labia | -144
    swelling opened and began to drain | -48
    temperature 36.8°C | 0
    blood pressure 100/60 mmHg | 0
    pulse 96-100 beats per minute | 0
    respiratory rate 20 breaths per minute | 0
    arterial oxygen saturation 98% | 0
    white blood cell count 17.4×10^9 per liter | 0
    started on vancomycin | 0
    started on piperacillin/tazobactam | 0
    surgery consult requested | 0
    pelvic CT scan obtained | 0
    CT showed cutaneous ulceration over left labia | 0
    CT showed air in subcutaneous fat of left groin | 0
    CT showed air in subcutaneous fat of left lower abdominal wall | 0
    inflammatory fat stranding along left lateral abdominal wall | 0
    LRINEC score 3 | 0
    LRINEC score potential 7 | 0
    decision for immediate explorative surgery | 0
    gynecology team involved | 0
    explorative surgery of pelvic and abdominal regions | 0
    diagnosis of necrotizing soft tissue infection confirmed | 0
    infection originating at left vulva | 0
    infection spreading to abdominal wall | 0
    first aggressive debridement performed | 0
    second look exploration surgery | 24
    further debridement of vulvar area | 24
    additional pockets of necrosis in abdominal wall discovered | 24
    additional debridement of necrosis | 24
    three surgeries for debridement and closure | 24
    stay in surgical intensive care unit | 120
    microbiology samples determined Clostridium clostridiforme | 120
    microbiology samples determined Bacteroides | 120
    Jackson-Pratt drain placed | 0
    drain removed during follow-up | 720
    healed well with no complications | 720
    proper bowel function | 720
    favorable cosmetic outcome | 720
    hemodynamic instability | 0
    tachycardia | 0
    hypotension | 0
    initial misdiagnosis with cellulitis | -24
    delay in surgical consultation | -24
    sepsis upon presentation | 0
    suspicion of NF raised | 0
    surgical intervention performed | 0
    <|eot_id|>
    56 years old | 0
African American female | 0
presented to the Emergency Department | -144
swelling over left labia | -144
swelling opened and began to drain | -48
temperature 36.8°C | 0
blood pressure 100/60 mmHg | 0
pulse 96-100 beats per minute | 0
respiratory rate 20 breaths per minute | 0
arterial oxygen saturation 98% | 0
white blood cell count 17.4×10^9 per liter | 0
started on vancomycin | 0
started on piperacillin/tazobactam | 0
surgery consult requested |A 0
pelvic CT scan obtained | 0
CT showed cutaneous ulceration over left labia | 0
CT showed air in subcutaneous fat of left groin | 0
CT showed air in subcutaneous fat of left lower abdominal wall | 0
inflammatory fat stranding along left lateral abdominal wall | 0
LRINEC score 3 | 0
LRINEC score potential 7 | 0
decision for immediate explorative surgery | 0
gynecology team involved | 0
explorative surgery of pelvic and abdominal regions | 0
diagnosis of necrotizing soft tissue infection confirmed | 0
infection originating at left vulva | 0
infection spreading to abdominal wall | 0
first aggressive debridement performed | 0
second look exploration surgery | 24
further debridement of vulvar area | 24
additional pockets of necrosis in abdominal wall discovered | 24
additional debridement of necrosis | 24
three surgeries for debridement and closure | 24
stay in surgical intensive care unit | 120
microbiology samples determined Clostridium clostridiforme | 120
microbiology samples determined Bacteroides | 120
Jackson-Pratt drain placed | 0
drain removed during follow-up | 720
healed well with no complications | 720
proper bowel function | 720
favorable cosmetic outcome | 720
hemodynamic instability | 0
tachycardia | 0
hypotension | 0
initial misdiagnosis with cellulitis | -24
delay in surgical consultation | -24
sepsis upon presentation | 0
suspicion of NF raised | 0
surgical intervention performed | 0