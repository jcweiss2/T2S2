52 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
right upper quadrant pain | -168 | 0 | Factual
abdominal fullness and distention | -168 | 0 | Factual
paroxysmal pain | -168 | 0 | Factual
worsened after meals | -168 | 0 | Factual
no nausea | 0 | 0 | Negated
no vomiting | 0 | 0 | Negated
no stiffness | 0 | 0 | Negated
no fever | -168 | 0 | Negated
hepatic abscess | -24 | 0 | Factual
treated with hepatic puncture and drainage | -24 | 0 | Factual
afebrile | 0 | 0 | Factual
pulse rate of 80 beats/minute | 0 | 0 | Factual
blood pressure of 118/73 mmHg | 0 | 0 | Factual
respiratory rate of 26 breaths/minute | 0 | 0 | Factual
leukocyte count of 16.4×10^9/L | 0 | 0 | Factual
neutrophil 94.5% | 0 | 0 | Factual
haemoglobin level of 85 g/L | 0 | 0 | Factual
platelet count of 240×10^9/L | 0 | 0 | Factual
procalcitonin level of 2.3 ng/mL | 0 | 0 | Factual
plasma fibrinogen level of 7.48 g/L | 0 | 0 | Factual
liver and renal function tests slightly abnormal | 0 | 0 | Factual
serum glutamic oxalacetic transaminase level of 67 U/L | 0 | 0 | Factual
glutamic-pyruvic transaminase level of 83 U/L | 0 | 0 | Factual
cholinesterase level of 1360 U/L | 0 | 0 | Factual
total protein and albumin levels of 50.8 and 21.5 g/L | 0 | 0 | Factual
blood urea nitrogen level of 10.8 mmol/L | 0 | 0 | Factual
creatinine level of 51.3 umol/L | 0 | 0 | Factual
negative for HIV | 0 | 0 | Negated
negative for syphilis | 0 | 0 | Negated
abdominal distension | 48 | 48 | Factual
mild bellyache | 48 | 48 | Factual
extreme thirst | 48 | 48 | Factual
right abdominal tenderness | 48 | 48 | Factual
no rebound or guarding | 48 | 48 | Negated
temperature of 36.8 °C | 48 | 48 | Factual
drainage catheter yield of 150 mL of fulvous fluid | 48 | 48 | Factual
abdominal and pelvic computed tomography (CT) scan | 48 | 48 | Factual
irregular, slightly low-density lesion in the right posterior hepatic lobe | 48 | 48 | Factual
gas density shadow inside | 48 | 48 | Factual
liquid density shadow and high-density drainage tube shadow | 48 | 48 | Factual
round-like low-density lesion of about 0.8 cm in diameter | 48 | 48 | Factual
appendix thickened to about 20 mm in diameter | 48 | 48 | Factual
structure of the ascending colon near the ileocecal region became disorganised | 48 | 48 | Factual
multiple gas accumulation and dilation in the bowel | 48 | 48 | Factual
air-fluid levels inside the abdomen | 48 | 48 | Factual
hepatic abscesses | 48 | 48 | Factual
ileus | 48 | 48 | Factual
mild ascites | 48 | 48 | Factual
abdominal infection | 48 | 48 | Factual
peritonitis | 48 | 48 | Factual
pre-shock | 72 | 72 | Factual
insufficient blood pressure of 93/59 mmHg | 72 | 72 | Factual
exploratory laparotomy | 72 | 72 | Factual
fulvous purulent exudate and necrotic tissue | 72 | 72 | Factual
partial postnecrotic defect in the peritoneum | 72 | 72 | Factual
massive epiploon adhesion in the right upper abdomen | 72 | 72 | Factual
two perforations | 72 | 72 | Factual
ileocecal resection | 72 | 72 | Factual
partial resection of the ascending colon | 72 | 72 | Factual
ileostomy | 72 | 72 | Factual
drainage of hepatic, abdominal and extraperitoneal abscesses | 72 | 72 | Factual
orotracheal intubation | 96 | 96 | Factual
hypotension | 96 | 96 | Factual
anemia | 96 | 96 | Factual
fever | 96 | 96 | Factual
transferred to the intensive care unit (ICU) | 96 | 96 | Factual
noradrenaline | 96 | 168 | Factual
ventilator | 96 | 168 | Factual
intravenous hydration | 96 | 168 | Factual
nutritional support therapy | 96 | 168 | Factual
blood transfusion | 96 | 168 | Factual
intravenous tigecycline | 96 | 120 | Factual
piperacillin/tazobactam | 96 | 120 | Factual
body temperature monitoring | 96 | 168 | Factual
routine blood count monitoring | 96 | 168 | Factual
procalcitonin level monitoring | 96 | 168 | Factual
C-reactive protein (CRP) level monitoring | 96 | 168 | Factual
temperature of 39.3°C | 120 | 120 | Factual
pulse rate of 130 beats/minute | 120 | 120 | Factual
leukocyte count of 35.9×10^9/L | 120 | 120 | Factual
neutrophils 92.4% | 120 | 120 | Factual
procalcitonin level of 8.15 ng/mL | 120 | 120 | Factual
CRP level of 174 mg/L | 120 | 120 | Factual
anaerobic blood culture positive | 120 | 120 | Factual
Gram stain revealed short Gram-positive bacillus | 120 | 120 | Factual
matrix-assisted laser desorption/ionization time-of-flight mass spectrometry (MALDI-TOF MS) | 120 | 120 | Factual
identified as E. lenta | 120 | 120 | Factual
plasma fibrinogen fell to 1.0 g/L | 144 | 144 | Factual
tigecycline replaced by teicoplanin | 144 | 144 | Factual
piperacillin/tazobactam discontinued | 144 | 144 | Factual
ertapenem added | 144 | 144 | Factual
cultures of the drainage fluid | 144 | 144 | Factual
Escherichia coli isolated | 144 | 144 | Factual
ertapenem and teicoplanin | 144 | 168 | Factual
fever improved | 168 | 168 | Factual
leukocytosis improved | 168 | 168 | Factual
procalcitonin level improved | 168 | 168 | Factual
CRP level improved | 168 | 168 | Factual
transferred to the general ward | 168 | 168 | Factual
ertapenem and teicoplanin for another 14 days | 168 | 336 | Factual
debridement | 168 | 336 | Factual
dressing change | 168 | 336 | Factual
symptomatic supportive treatment | 168 | 336 | Factual
repeated blood cultures negative | 336 | 336 | Factual
CT scan showed improvement | 336 | 336 | Factual
discharged | 504 | 504 | Factual
oral antibiotics (clindamycin) | 504 | 504 | Factual
follow-up | 672 | 672 | Factual
complete resolution of the abscess | 672 | 672 | Factual