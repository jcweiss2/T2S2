12-month-old|0
female|0
premature birth|0
vaginal delivery|0
low birth weight|0
neonatal sepsis|-672
parenteral antibiotics|-672
no surgical drainage|-672
no ultrasound-guided repeated aspiration|-672
referred to department|0
painless limping|0
right hip pain|0
walking on tiptoe|0
pelvic obliquity|0
Trendelenburg-Duchenne gait|0
limited right hip abduction|0
limited internal rotation|0
lower-extremity length discrepancy|0
shortening of right femur|0
plain anteroposterior radiographs|0
viable femoral head|0
decreased neck-shaft angle|0
relative overgrowth of greater trochanter|0
proximally migration|0
shortening of femoral neck|0
severe coxa vara|0
femoral neck pseudoarthrosis|0
vertical orientation of the capital physis|0
preoperative Hilgenreiner-epiphyseal angle|0
Choi Type IIIB|0
Johari Group V|0
proximal femoral valgus osteotomy|0
adductor tenotomy|0
adductor soft tissue release|0
correction of neck shaft angle|0
lateral approach|0
subperiosteal detachment of vastus lateralis|0
closing wedge valgus osteotomy|0
130° angled blade plate|0
internal fixation|0
postoperative partial weight bearing|0
postoperative Trendelenburg gait correction|0
restored right lower extremity alignment|0
corrected lower-extremity length discrepancy|0
intertrochanteric osteotomy|0
valgisation|0
transfer of greater trochanter|0
postoperative Hilgenreiner-epiphyseal angle|0
acetabular depth improvement|0
consolidation of osteotomy|0
hardware removal|0
no hip pain|0
better hip range of motion|0
hip flexion|0
hip extension|0
hip abduction|0
hip adduction|0
internal rotation|0
external rotation|0
no difficulties with recreational activities|0
osteotomy healed|0
able to squat|0
able to run|0
able to climb stairs|0
able to walk without limp|0
shortening reduced|0
x-ray showed neck shaft angle|0
union of pseudoarthrosis|0
