28 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
farmer | 0 | 0 | Factual
ingestion of two fresh tablets of Celphos | -4 | -4 | Factual
vomiting | -4 | 0 | Factual
abdominal pain | -4 | 0 | Factual
agitated | 0 | 0 | Factual
anxious | 0 | 0 | Factual
irritable | 0 | 0 | Factual
pulse rate not palpable | 0 | 0 | Factual
blood pressure not recordable | 0 | 0 | Factual
heart rate 110/min | 0 | 0 | Factual
respiratory rate 28/min | 0 | 0 | Factual
oxygen saturation 95% | 0 | 0 | Factual
sinus tachycardia | 0 | 0 | Factual
T wave inversion in lead 3 | 0 | 0 | Factual
intravenous crystalloids | 0 | 24 | Factual
intravenous magnesium sulphate | 0 | 24 | Factual
intravenous calcium gluconate | 0 | 24 | Factual
intravenous hydrocortisone | 0 | 24 | Factual
intravenous dopamine | 0 | 24 | Factual
intravenous noradrenaline | 0 | 24 | Factual
gastric lavage with potassium permanganate | 0 | 0 | Factual
activated charcoal | 0 | 24 | Factual
arterial blood gas analysis | 0 | 0 | Factual
metabolic acidosis | 0 | 24 | Factual
intubation | 0 | 0 | Factual
shifted to intensive care unit | 0 | 0 | Factual
blood pressure 60-80 mmHg | 6 | 6 | Factual
pulse rate 120/min | 6 | 6 | Factual
respiratory rate 20/min | 6 | 6 | Factual
input/output 3L/300 ml | 6 | 24 | Factual
monomorphic ventricular tachycardia | 48 | 48 | Factual
DC cardio-version | 48 | 48 | Factual
intravenous amiodarone | 48 | 96 | Factual
cardiac bio-markers raised | 48 | 48 | Factual
cardiac bio-markers normalised | 336 | 336 | Factual
arterial blood gas analysis | 96 | 96 | Factual
blood urea 100 mg/dl | 96 | 96 | Factual
serum creatinine 4.5 mg/dl | 96 | 96 | Factual
urine output 400 ml/24 hours | 96 | 96 | Factual
aspartate amino-transferase/alanine amino-transferase 80/90 IU/L | 96 | 96 | Factual
alkaline phosphatase 200 U/L | 96 | 96 | Factual
S bilirubin 2.5 mg/dl | 96 | 96 | Factual
liver and kidney involvement | 96 | 96 | Factual
blood pressure 100/70 mmHg | 120 | 120 | Factual
pulse rate 110/min | 120 | 120 | Factual
respiratory rate 22/min | 120 | 120 | Factual
total leucocyte count 14000/mm3 | 120 | 120 | Factual
polymorphonuclear leucocytosis | 120 | 120 | Factual
urea 200 mg/dl | 120 | 120 | Factual
S. creatinine 7.5 mg/dl | 120 | 120 | Factual
urine output 400 ml/24 hours | 120 | 120 | Factual
arterial blood gas analysis | 120 | 120 | Factual
re-appearance of acidosis | 120 | 120 | Factual
haemodialysis | 120 | 120 | Factual
haemodialysis | 168 | 168 | Factual
blood urea 70 mg/dl | 168 | 168 | Factual
creatinine 4.0 mg/dl | 168 | 168 | Factual
urine output 1200 ml/24 hours | 168 | 168 | Factual
extubation | 144 | 144 | Factual
shifted to step down unit | 192 | 192 | Factual
vitals normal | 192 | 192 | Factual
liver and kidney functions improving | 192 | 336 | Factual
discharge | 336 | 336 | Factual