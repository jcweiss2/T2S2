45 years old | 0
    male | 0
    received yellow fever vaccine | 0
    fever | 168
    myalgia | 168
    headache | 168
    vomiting | 168
    jaundice | 216
    abdominal pain | 216
    conjunctival suffusion | 216
    altered mental status | 216
    respiratory failure | 216
    hemodynamic instability | 216
    admitted to Intensive Care Unit | 216
    leukocytosis | 216
    thrombocytopenia | 216
    elevated alanine aminotransferase | 216
    elevated aspartate aminotransferase | 216
    elevated total bilirubin | 216
    elevated creatinine | 216
    elevated creatine phosphokinase | 216
    elevated prothrombin-time international normalized ratio | 216
    started ceftriaxone | 216
    switched to piperacillin-tazobactam | 216
    started methylprednisolone | 216
    received hemoderivatives transfusion | 216
    hemodialysis | 216
    negative blood cultures | 216
    negative dengue fever serology | 216
    negative leptospirosis serology | 216
    abdominal CT without significant findings | 216
    moderate free fluid in abdominal cavity | 216
    persistent altered mental status | 336
    frontal lobe bleeding | 336
    severe diffuse brain dysfunction | 336
    death | 480
    confirmed yellow fever infection | 480
    liver steatosis | 480
    hepatocytic necrosis | 480
    perivascular lymphocyte encephalitis | 480
    angioinvasive hyalohyphomycosis | 480
    fungal embolism | 480
    thrombosis of vessels | 480
    endomyocarditis | 480
    cardiomyocyte necrosis | 480
    fungal brain abscesses | 480
    necrotizing encephalitis | 480
    rough kidney surface | 480
    hyalinized glomeruli | 480
    tubular atrophy | 480
    benign nephrosclerosis | 480
    hematogenic acute pyelonephritis | 480
    renal papillary neoplasm | 480
    clear cell renal adenocarcinoma | 480
    pancreatic fat necrosis | 480
    fungal thrombosis | 480
    Aspergillus spp. infection | 480
    yellow fever vaccine virus confirmed | 480
    