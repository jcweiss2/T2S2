44 years old | 0
female | 0
Caucasian | 0
facial paralysis | -672
acoustic neuroma removal | -672
lagophthalmos | -672
keratopathy | -672
gold weight implantation | 0
right upper eyelid swelling | 264
erythema | 264
limitation of abduction | 264
orbital cellulitis | 264
intravenous cefuroxime | 264
complete limitation of gaze | 268
afferent pupillary defect | 268
necrosis of lower eyelid | 268
necrosis of upper eyelid margins | 268
necrosis of anterior ocular segment | 268
computed tomography scan | 268
gold weight removal | 272
necrosis of upper eyelid tarsus | 272
necrosis of lower eyelid | 272
necrosis of limbus | 272
necrosis of conjunctiva | 272
corneal opacity | 272
dense cataract | 272
full thickness biopsy | 272
necrotic conjunctiva | 272
necrotic skin | 272
diffuse acute inflammatory reaction | 272
gram-positive cocci | 272
Staphylococcus capitis | 272
intravenous vancomycin | 272
piperacillin/tazobactam | 272
visual acuity light perception | 272
transcranial Doppler | 276
normal flow in ophthalmic arteries | 276
fever | 296
chills | 296
tachycardia | 296
restlessness | 296
systemic involvement | 296
scleral necrosis | 296
worsening eyelid swelling | 296
worsening necrosis | 296
axial computed tomography scan | 296
air bubbles under eyelid | 296
intraconal fat haziness | 296
evisceration | 300
debridement of necrotic tissue | 300
acute nonspecific necrotizing panophthalmitis | 300
gram-positive cocci | 300
Staphylococcus epidermidis | 300
Candida albicans | 300
Candida glabrata | 300
Clindamycin | 300
voriconazole | 300
systemic condition deterioration | 304
fever | 304
urinary retention | 304
desaturation | 304
acidosis | 304
intensive care unit admission | 304
vancomycin | 304
meropenem | 304
fluconazole | 304
condition improvement | 312
ocular condition stabilization | 312
severe contracted socket | 8760
nonhealing third-degree chemical burn | 8760
right anterior thigh | 8760
wound debridement | 8760
local anesthesia | 8760
lack of patient cooperation | 8760
second operation | 8760
complete debridement | 8760
general anesthesia | 8760
split thickness skin graft | 8760
negative pressure dressing | 8760
dressing tear | 8784
partial skin graft take | 8784
Sulfamylon wet-to-dry dressing | 8784
tenderness | 8784
itching | 8784
unrest | 8784
full thickness third degree burn | 8808
no signs of infection | 8808
further operation | 8816
debridement | 8816
partial thickness skin graft | 8816
dressing and skin graft removal | 8816
full length cast | 8816
self-induced damage suspicion | 8816
factitious disorder suspicion | 8816
psychiatric consult | 8816
no factitious disorder diagnosis | 8816