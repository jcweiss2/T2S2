41 years old | 0
female | 0
smoker | 0
15 pack-year history | 0
admitted to the hospital | 0
endoscopic resection of a submucous uterine myoma | 0
general anesthesia | 0
fentanyl | 0
propofol | 0
I-gel laryngeal mask No. 4 | 0
desflurane | 0
lithotomy position | 0
hysteroscopy | 0
bipolar 9-mm resectoscope | 0
0.9% saline | 0
end-tidal CO2 dropped | -50
pulse oximetry dropped | -50
crackling sounds from the base of the lungs | -50
pulmonary oedema suspected | -50
irrigated saline checked | -50
9000 mL of saline used | -50
4000 mL of saline collected | -50
surgery stopped | -50
generalized oedema noticed | -50
distended abdomen | -50
cervical oedema | -50
inspired fraction of oxygen increased | -50
arterial blood analysis | -50
pH 7.09 | -50
PaCO2 41 mmHg | -50
PO2 70 mmHg | -50
HCO3+ 12.4 mEq/L | -50
Na+ 145 mEq/L | -50
K+ 2.3 mEq/L | -50
Ca2+ 0.76 mEq/L | -50
hemoglobin 5.9 g/dL | -50
O2 sat 89% | -50
blood glucose level 50 mg/dL | -50
sodium bicarbonate administered | -40
furosemide administered | -40
laryngeal mask replaced by tracheal tube | -40
airway oedema observed | -40
arytenoid region oedema | -40
intubation of 6.5-mm tracheal tube | -40
arterial and central lines put | -40
potassium chloride administered | -40
calcium chloride administered | -40
magnesium sulfate administered | -40
dextrose administered | -40
laparoscopy performed | -30
no uterine rupture | -30
intestinal loops oedema | -30
peritoneal free fluid observed | -30
bladder catheter inserted | -30
auricular temperature 33°C | -30
admitted to ICU | 0
postoperative chest X-ray | 2
bilateral pulmonary oedema | 2
electrolyte disturbances corrected | 2
acidosis corrected | 2
hemoglobin increased | 6
temperature returned to normal | 6
generalized oedema resolved | 6
urine output 3000 mL | 6
extubation | 6
oxygen supplementation | 12
transferred to general ward | 24
discharged | 48