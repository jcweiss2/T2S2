57 years old | 0
male | 0
admitted to the hospital | 0
acute abdomen | 0
nausea | 0
vomiting | 0
supra=umbilical incarcerated incisional hernia | 0
body mass index 38.3 kg/m2 | 0
elevated white cell count | 0
elevated CRP | 0
elevated interleukins | 0
elevated creatinine | 0
elevated urea | 0
amiodarone | 0
pantoprazole | 0
bisoprolol | 0
eplerenone | 0
sacubitril/valsartan | 0
eliquis | 0
l-thyroxin | 0
dilated cardiomyopathy | 0
ejection fraction 15-20% | 0
atrial fibrillation | 0
left atrial thrombus | 0
implantable cardioverter defibrillator | 0
radioiodine therapy | 0
laparoscopic appendectomy | 0
perforated appendicitis | 0
peritonitis | 0
emergency laparotomy | 0
incarcerated ischaemic ileum | 0
tinny pale intramural lesions | 0
resected ileum | 0
end-to-end ileo-ileostomy | 0
sepsis | 0
cardiopulmonary instability | 0
intensive care for 4 days | 0
discharged home on postoperative day 11 | 264
resected ileum histology: hemorrhagic mucosa | 0
resected ileum histology: mural necrosis | 0
three foci of well-differentiated NET | 0
immunohistochemistry positivity: CK AE 1/3 | 0
immunohistochemistry positivity: synaptophysin | 0
immunohistochemistry positivity: chromogranin | 0
immunohistochemistry positivity: CD56 | 0
NET grade 1 (Ki67 < 1%) | 0
NET mitotic activity 1 mitosis/10 HPF | 0
staging pT2m | 0
staging pN0 | 0
staging pL0 | 0
staging pV0 | 0
resection margins R0 | 0
six-week post-surgery NET workup | 432
CT thorax, abdomen, pelvis: no neuroendocrine disease | 432
no increased DOTATATE avidity on 68Ga PET/CT | 432
plasma chromogranin A elevated | 432
5-HIAA normal | 432
denied carcinoid syndrome symptoms | 432
suspected residual neuroendocrine disease | 432
repeat laparotomy | 432
palpation of entire small bowel | 432
ileum resection with multiple intramural deposits | 432
end-to-end ileo-ileostomy | 432
remaining 280 cm small intestine | 432
postoperative course uneventful | 432
histology: 25 well-differentiated NET | 432
immunohistochemistry positivity: chromogranin | 432
immunohistochemistry positivity: synaptophysin | 432
immunohistochemistry positivity: SSTR 2A | 432
Ki67 <2% (G1) | 432
staging pT1m | 432
staging pN1 | 432
staging pL0 | 432
staging pV0 | 432
resection margins R0 | 432
last follow-up 9 months post-surgery | 6480
no evidence of disease | 6480
alive | 6480
