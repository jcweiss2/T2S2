61 years old | 0
male | 0
admitted to the intensive care unit | 0
acute respiratory distress | 0
shock | 0
unconscious | 0
Glasgow Coma Scale score of 10/15 | 0
tachycardic at 145 bpm | 0
hypotensive at 86/51 mm Hg | 0
polypneic at 32 cpm | 0
desaturated at 40% at room air | 0
desaturated at 78% under high mask concentration 15 L/mn | 0
body temperature 38.5°C | 0
diffuse subcrackling rales | 0
ulcerative lesions of the nasal cavity | 0
ulcerative lesions of the oral cavity | 0
blood gas lactate level 3.24 | 0
blood gas PaO2/FiO2 ratio of 105 | 0
elevated white blood cells to 14,600/µL | 0
elevated C-reactive protein level to 230 mg/L | 0
procalcitonin positive at 2.32 g/L | 0
lymphopenia at 180/µL | 0
anemia at 8.4 g/dL | 0
prothombin time at 51% | 0
high level of D-dimers 2.76 mg/L | 0
normal renal function | 0
normal hepatic function | 0
sinus tachycardia | 0
CT scan bilateral infectious bronchopneumonia | 0
CT scan moderate bilateral pleurisy | 0
CT scan no signs of pulmonary embolism | 0
transthoracic echocardiogram normal | 0
pneumonia caused by Klebsiella rhinoscleromatis | 0
ARDS | 0
septic shock | 0
intubated | 0
vasoactive drugs noradrenaline at rate 0.25 mcg/kg/min | 0
intravenous Triaxon 2 g/d | 0
intravenous ciprofloxacin 200 mg twice a day | 0
bacterium detected in distal pulmonary swab | 0
bacterium detected in blood culture | 0
organ dysfunction failure | 240
passed away | 240
nasal cavity rhinoscleroma | -672 (assuming nasal cavity rhinoscleroma was diagnosed prior to admission, approximated to 4 weeks earlier)
