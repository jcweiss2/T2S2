69 years old | 0
female | 0
paraplegic | -18000
public road accident | -18000
implanted for intrathecal therapy | -4320
Ascenda catheter | -4320
Synchromed II pump | -4320
baclofen | -4320
morphine | -4320
doses unchanged | -4320
daily administration of 300 μg of baclofen | -4320
daily administration of 400 μg of morphine | -4320
fillings scheduled every 10 weeks | -4320
pump replacement | -2160
lymphatic collection | -2160
regular aspirations | -2160
diffusion dried up | -840
fever | -24
chills | -24
fatigue | -24
presented to the Emergency Department | 0
Glasgow Coma Scale score of 15/15 | 0
nausea | 0
cloudy liquid issuing from a small hole | 0
indurated zone surrounding the pump | 0
elevated C-reactive protein | 0
antibiotherapy begun | 0
vancomycin | 0
cefotaxime | 0
local surgical cleaning of the site of the pump | 24
cerebrospinal fluid sample collected | 24
elevated white blood cell count | 24
elevated protein concentration | 24
low glycorrhachia | 24
Gram-positive cocci | 24
Streptococcus dysgalactiae | 24
antibiotics switched to amoxicillin | 48
rifampicin | 48
hospitalized in the intensive care unit | 0
transferred to the infectious diseases department | 72
ablation of the pump and intrathecal catheter | 216
new intrathecal catheter placed | 216
tunnelled to the right hypochondrium | 216
linked to an implanted port | 216
external pump connected to the port | 216
continuous administration of the intrathecal therapy | 216
replacement of the implanted port by a new Synchromed II pump | 408
discharged for outpatient follow up | 432
antibiotic therapy prolonged at home | 432
cured of this acute episode | 2592