12 years old | 0
    female | 0
    steroid-resistant nephrotic syndrome | 0
    presented to the emergency department | 0
    fever | 0
    shortness of breath | 0
    cough | 0
    tachycardic | 0
    tachypneic | 0
    supplemental oxygen | 0
    normal saline bolus | 0
    chest X-ray bilateral pulmonary edema | 0
    sepsis | 0
    vancomycin | 0
    cefotaxime | 0
    admitted to pediatric intensive care unit | 0
    nephrotic syndrome | -6264
    steroid-responsive | -6264
    relapses when steroid dose tapered | -6264
    renal biopsy minimal change disease | -6312
    genetic testing heterozygous non-coding mutation in TRPC6 | -6312
    cyclophosphamide | -6312
    1.5-year remission | -6312
    tacrolimus | -8760
    partial clinical response | -8760
    improved edema | -8760
    persistent proteinuria | -8760
    concern for FSGS | -8760
    repeat biopsy interstitial nephritis | -8760
    Acthar Gel | -1440
    tacrolimus continued | -1440
    S. pneumoniae blood culture | 8
    nasopharyngeal swab PCR positive for parainfluenza type 2 | 8
    oliguria | 8
    creatinine increased from 1.4 to 2.4 mg/dL | 8
    hemoglobin decreased from 11.4 to 7.4 g/dL | 8
    Acthar discontinued | 8
    tacrolimus discontinued | 8
    unwashed packed red blood cells transfusion | 8
    continuous veno-venous hemodiafiltration | 8
    respiratory failure | 96
    intubation | 96
    chest CT bilateral patchy consolidation | 96
    bilateral pleural effusions | 96
    high-dose hydrocortisone | 96
    platelet count decreased | 96
    clinical condition worsened | 96
    intravenous vasoactive support | 96
    plasma exchange started | 120
    FFP replacement | 120
    pHUS considered | 120
    direct Coombs test negative | 120
    plasma exchange completed | 168
    direct Coombs test positive | 168
    platelet count nadir 36 | 312
    platelet count improved | 312
    supportive care | 0
    antibiotics | 0
    temporary KRT | 0
    creatinine returned to baseline 0.6 mg/dL | 936
    discharged home | 936
    angiotensin-converting enzyme inhibitor therapy | 936
    persistent nephrotic syndrome | 936
    