42 years old | 0
man | 0
renal failure secondary to adult polycystic kidney disease | 0
recurrent urinary tract infections following renal transplantation 7 months earlier | -5040
admitted with dysuria | 0
right-sided loin pain | 0
blood pressure 140/80 mmHg | 0
pulse 80 beats/minute | 0
temperature 38.5°C | 0
white cell count 12.5 × 103/mm3 | 0
haemoglobin 9.5 g/L | 0
platelet count 568 × 103/mm3 | 0
