28 years old | 0
male | 0
thermal burn | -1
improper handling of a gasoline can | -1
superficial, deep partial-thickness burns | -1
full-thickness burns | -1
total body surface area lesions | -1
chest and abdominal debridement | 0
decompression incisions | 0
protective tracheal intubation | 0
increased C-reactive protein | 0
moderately elevated procalcitonin | 0
severe hypoproteinemia | 0
ABSI | 0
Baux | 0
R-Baux | 0
local conservative nonsurgical treatment | 48
lavage | 48
dressing with silver-containing products | 48
admission to the Intensive Care Unit | 48
respiratory support using mechanical ventilation | 48
signs of an extremely aggressive burn-induced inflammatory reaction | 48
increased CRP | 48
decreased albumin | 48
increased presepsin | 48
decreased serum iron | 48
extubation | 72
conservative local treatment methods | 72
removing devitalized tissue | 72
application of special topical antimicrobial agents | 72
excision and grafting with expanded meshed autografts | 72
proton-pump inhibitor | 72
thromboprophylaxis with enoxaparin | 72
analgesics | 72
antioxidants | 72
oligoelements | 72
enteral and parenteral nutrition | 72
normal feeding | 72
adequate tissue perfusion | 72
mean arterial pressure | 72
diuresis | 72
lactate | 72
central venous oxygen saturation | 72
colonization of the wound with Pseudomonas aeruginosa | 192
increased presepsin value | 192
antibiotic therapy with colistin | 192
antibiotic therapy with cefoperazone/sulbactam | 192
swab cultures | 192
decrease in presepsin | 336
excision and grafting with expanded meshed autograft | 840
discharge | 1056