41 years old | 0
premenopausal woman | 0
re-presented to the metropolitan hospital emergency department | 0
worsening abdominal pain | 0
vomiting | 0
non-bloody diarrhoea | 0
fever | 0
inpatient treatment for bilateral Escherichia coli pyelonephritis | -240
reported 3 weeks of intermittent abdominal pain | -504
returning from overseas travel to Indonesia | -504
Stage 4 endometriosis | -34560
bilateral endometriomas | -34560
rectal nodule | -34560
obliterated pouch of Douglas | -34560
fixed anterior uterus | -34560
diagnosed on ultrasound | -34560
no previous laparoscopies | -34560
one previous caesarean section | -34560
well controlled asthma | -34560
denied any recent sexual intercourse | 0
no uterine instrumentation | 0
no history of PID | 0
no history of sexually transmitted infections | 0
not taking any regular medication | 0
not on any contraceptives | 0
had regular menstrual cycles | 0
tachycardic | 0
hypotensive | 0
febrile | 0
right renal angle tenderness | 0
generalised lower abdominal tenderness | 0
rebound | 0
guarding | 0
right adnexal tenderness on bimanual exam | 0
no palpable masses | 0
no cervical motion tenderness | 0
speculum examination unremarkable | 0
normal cervix visualised macroscopically | 0
no abnormal vaginal discharge | 0
elevated lactate (3.1 mmol/L) | 0
in shock | 0
elevated inflammatory parameters | 0
leucocytosis of 16.9 × 109/L | 0
93% neutrophilia | 0
rise in C-reactive protein (CRP) 315 mg/L | 0
acute kidney injury | 0
elevated creatinine 100 μmol/L | 0
reduced estimated glomerular filtration rate (eGFR) 60 mL/min/1.73m2 | 0
quantitative beta hCG negative | 0
urinalysis negative | 0
microscopy negative | 0
urine culture negative | 0
endocervical swabs negative for Chlamydia trachomatis | 0
endocervical swabs negative for Neisseria gonorrhoea | 0
blood cultures negative | 0
stool culture positive for Campylobacter jejuni | 0
CT abdomen showed bilateral enlarged ovaries | 0
septated cysts | 0
low-density mass in the presacral space | 0
fat stranding | 0
transvaginal deep infiltrating endometriosis ultrasound demonstrated multiple endometriomas | 0
right ovarian cyst 54 mm × 31 mm × 32 mm | 0
three left ovarian cysts | 0
largest left ovarian cyst 39 mm × 33 mm × 38 mm | 0
ovaries fixed in the pelvis | 0
kissing ovaries sign | 0
sliding sign negative | 0
bowel adherent to the posterior wall of the uterus | 0
two bowel nodules | 0
differential diagnoses included colitis | 0
differential diagnoses included urosepsis | 0
differential diagnoses included appendicitis | 0
differential diagnoses included tuboBovarian abscesses | 0
tuboBovarian abscess less likely given stable appearance compared with previous imaging | 0
managed empirically for sepsis | 0
adult sepsis pathway | 0
fluid resuscitation | 0
broadBspectrum intravenous antibiotics (ceftriaxone and metronidazole) | 0
condition deteriorated over the next 24B36 h | 24
ongoing fever | 24
tachycardia | 24
hypotension | 24
required transfer to the intensive care unit | 24
inotropic support | 24
changed to intravenous amoxicillin with clavulanic acid | 24
commenced on azithromycin for Campylobacteriosis | 24
day 5 of hospital admission | 120
ongoing pain | 120
infective signs | 120
repeat CT abdomen pelvis | 120
interval increase in left multiloculated adnexal mass | 120
increased surrounding fat stranding | 120
free fluid in the pelvis | 120
bowel wall thickening of the sigmoid | 120
bowel wall thickening of the descending colon | 120
bowel wall thickening of the transverse colon | 120
possible inflammatory or infective nature | 120
decision made for exploratory laparoscopy | 120
underwent urgent laparoscopic washout | 120
drainage of tuboBovarian abscesses | 120
source control of infection | 120
sterile abscess culture fluid positive for Escherichia coli | 120
right adnexal tissue histopathology showed abscess formation | 120
no evidence of endometriosis | 120
managed with intravenous antibiotics | 120
intravenous fluids | 120
condition greatly improved | 120
discharged from hospital | 168
plan for outpatient followBup | 168
repeat pelvic scan | 168
