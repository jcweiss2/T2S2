26 years old | 0
    woman | 0
    rural area of Peru | 0
    two vaginal deliveries without complications | 0
    complete prenatal care during current pregnancy | 0
    three doses of tetanus, diphtheria, and pertussis (DTaP) during childhood | 0
    one dose of tetanus and diphtheria (Tdap) vaccine during each pregnancy | 0
    last dose of Tdap on June 14, 2020 at 27 weeks of gestation | -1104
    presented to hospital in active phase of labor at 38 weeks of gestation | 0
    vaginal delivery | 0
    child weighing 3.7 kg | 0
    postpartum hemorrhage two days after delivery | 48
    hypotension | 48
    tachycardia | 48
    altered sensorium | 48
    flaccid uterus | 48
    pelvic ultrasound demonstrated retention of placental tissue | 48
    uterine curettage performed | 48
    discharged four days later | 96
    headache 14 days after discharge | 336
    nausea | 336
    general malaise | 336
    fever | 336
    vital signs within normal ranges | 336
    scant lochia without bad odor | 336
    absence of vaginal bleeding | 336
    hematocrit 24% | 336
    hemoglobin 7.3 g/dL | 336
    white blood cells 14,000 m/mm3 | 336
    creatinine 104 μmol/L | 336
    urinalysis: 12 white blood cells per high power field | 336
    urinalysis: eight epithelial cells per high power field | 336
    positive urine culture for E. coli sensitive to ceftriaxone | 336
    hospitalized with presumptive diagnosis of urinary tract infection | 336
    severe anemia | 336
    treatment with ceftriaxone 2 g IV daily | 336
    iron saccharate | 336
    hydration | 336
    altered mental status on day two of hospitalization | 384
    no response to external stimuli | 384
    Glasgow Coma Scale score of seven | 384
    nuchal stiffness | 384
    limb stiffness | 384
    intubation performed for airway protection | 384
    transferred to more equipped hospital | 384
    laboratory exam unremarkable | 384
    non-contrast cerebral computed tomography unremarkable | 384
    lumbar puncture performed | 384
    white cell count: 30/mm3 | 384
    glucose: 42 mg/dl | 384
    proteins: 70 g/L | 384
    CSF culture showed no growth | 384
    blood cultures showed no growth | 384
    admitted to intensive care unit (ICU) | 384
    empiric treatment for meningitis with ceftriaxone | 384
    vancomycin | 384
    acyclovir | 384
    severe trismus on second day of hospitalization in ICU | 432
    increased respiratory rate | 432
    spasms of upper and lower extremities | 432
    trunk spasms | 432
    passive motion of limbs caused diffuse spasms | 432
    clinical diagnosis of severe tetanus | 432
    vaginal cultures obtained | 432
    vaginal cultures showed no growth | 432
    treatment with penicillin G four million units IV every four hours for seven days | 432
    two doses of 500 units of IM anti-tetanus immunoglobulin | 432
    extubated on sixth day of hospitalization | 528
    clinical improvement observed | 528
    discharged on 27th day of hospitalization | 648
    gait disorder | 648
    mild long-term memory impairment | 648
    