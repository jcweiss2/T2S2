75 years old | 0 | 0 
male | 0 | 0 
admitted to the hospital | 0 | 0 
fever | -168 | 0 
chills | -168 | 0 
dizziness | -168 | 0 
remission after fever | -168 | 0 
no headache | -168 | 0 
no abdominal pain | -168 | 0 
no diarrhea | -168 | 0 
no sputum | -168 | 0 
no nasal congestion | -168 | 0 
no runny nose | -168 | 0 
hypertension | -6720 | 0 
body temperature 39.0 °C | -168 | 0 
levofloxacin 0.5 g qd | 0 | 72 
body temperature above 39.0 °C | 0 | 72 
blood culture indicated penicillin-resistant Staphylococcus | 72 | 72 
Vancomycin injection 500000 U q6h | 72 | 168 
body temperature returned to normal | 168 | 168 
discharged from the hospital | 168 | 168 
high fever again | 192 | 192 
maximum body temperature 39.7 °C | 192 | 192 
chills | 192 | 192 
cough | 192 | 192 
sputum | 192 | 192 
no chest pain | 192 | 192 
no limb twitching | 192 | 192 
pupils sluggish in light reflection | 192 | 192 
confused | 192 | 192 
mentally soft | 192 | 192 
could only communicate briefly | 192 | 192 
muscle strength test could not cooperate | 192 | 192 
voluntary activities were seen | 192 | 192 
diarrhea | 192 | 192 
high-frequency oxygen inhalation | 192 | 192 
piperacillin and tazobactam 4.5 g q8h | 192 | 240 
methylprednisolone injection 40 mg | 192 | 192 
body temperature above 38.3 °C | 192 | 240 
levofloxacin 0.5 g qd | 240 | 288 
body temperature returned to normal | 288 | 288 
consciousness became clear | 288 | 288 
CRP dropped to 76.4 mmol/L | 288 | 288 
transferred to the general ward of the Department of Respiratory Medicine | 288 | 288 
atrial fibrillation | 288 | 288 
unresponsiveness | 288 | 288 
slurred speech | 288 | 288 
shortness of breath | 288 | 288 
slow light reflexes | 288 | 288 
stiff neck | 288 | 288 
increased muscle tone | 288 | 288 
wet rales in both lungs | 288 | 288 
repeated fever | 288 | 336 
body temperature fluctuating around 38.7 °C | 288 | 336 
sudden blood pressure drops | 288 | 336 
septic shock | 288 | 336 
active rehydration | 288 | 336 
norepinephrine micropump | 288 | 336 
vancomycin injection 1 million units q12h | 288 | 336 
meropenem injection 1.0 g q8h | 288 | 336 
methylprednisolone reduced to 20 mg | 288 | 336 
methylprednisolone stopped | 336 | 336 
unconscious | 336 | 336 
base of the tongue fell back | 336 | 336 
shortness of breath | 336 | 336 
stiff neck | 336 | 336 
tremor of the limbs | 336 | 336 
heart rate dropped to 40 beats per minute | 336 | 336 
trachea intubated | 336 | 336 
breathing assisted by a ventilator | 336 | 336 
condition continued to deteriorate rapidly | 336 | 336 
multiple organ failure | 336 | 336 
family decided to discontinue further treatment | 336 | 336 
died | 336 | 336