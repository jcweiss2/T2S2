85 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
farmer | 0 | 0 | Factual
active lifestyle | 0 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
atrial fibrillation | -6720 | 0 | Factual
benign prostatic hypertrophy | -6720 | 0 | Factual
trismus | -144 | 0 | Factual
hypertonia | -144 | 0 | Factual
injured his leg | -144 | -144 | Factual
C. tetani infection | -144 | 0 | Factual
immunoglobulins | -144 | -120 | Factual
tetanus vaccination | -144 | -120 | Factual
metronidazole | -144 | -134 | Factual
transferred to ICU | -120 | -120 | Factual
tracheostomy | -120 | -120 | Factual
mechanical ventilation | -120 | 0 | Factual
vasoactive support | -120 | 0 | Factual
seizures | -120 | 0 | Factual
baclofen | -120 | 0 | Factual
midazolam | -120 | 0 | Factual
diazepam | -120 | 0 | Factual
electroencephalography | -120 | -120 | Factual
slow cerebral activity | -120 | 0 | Factual
respiratory failure | -120 | 0 | Factual
opacity on chest radiography | -120 | 0 | Factual
peripheral leukocytosis | -120 | 0 | Factual
ventilator-associated pneumonia | -120 | 0 | Factual
blood cultures | -120 | -120 | Factual
tracheal secretion samples | -120 | -120 | Factual
Klebsiella pneumoniae | -120 | 0 | Factual
methicillin-sensitive Staphylococcus aureus | -120 | 0 | Factual
piperacillin-tazobactam | -120 | -100 | Factual
transferred to geriatric unit | -100 | -100 | Factual
coma | -100 | 0 | Factual
spontaneous breathing | -100 | 0 | Factual
supplemental oxygen | -100 | 0 | Factual
tracheal cannula | -100 | 0 | Factual
antibiotic therapy switched to linezolid | -96 | -82 | Factual
septic shock | -96 | 0 | Factual
meropenem | -96 | -79 | Factual
awoke | -79 | -79 | Factual
feeding tube removed | -79 | -79 | Factual
cholestasis | -79 | 0 | Factual
acute edematous pancreatitis | -79 | 0 | Factual
endoscopic treatment postponed | -79 | -79 | Factual
urinary tract infection | -72 | -65 | Factual
multidrug-resistant organisms | -72 | 0 | Factual
K. pneumoniae | -72 | 0 | Factual
Acinetobacter baumannii | -72 | 0 | Factual
Enterococcus faecalis | -72 | 0 | Factual
colistin | -72 | -65 | Factual
amoxicillin-clavulanate | -72 | -65 | Factual
clinical condition improved | -65 | -65 | Factual
transferred to rehabilitation unit | -65 | -65 | Factual
MDRO isolation | -65 | 0 | Factual
tracheal supplemental oxygen | -65 | 0 | Factual
bladder catheter | -65 | 0 | Factual
pressure ulcers | -65 | 0 | Factual
sarcopenic | -65 | 0 | Factual
low handgrip strength | -65 | 0 | Factual
low appendicular skeletal mass | -65 | 0 | Factual
rehabilitation | -65 | 0 | Factual
Clostridioides difficile infection | -60 | -50 | Factual
oral vancomycin | -60 | -50 | Factual
atrial fibrillation with third-degree atrioventricular block | -57 | -57 | Factual
single-chamber pacemaker implantation | -57 | -57 | Factual
hyperkinetic delirium | -55 | -55 | Factual
Pseudomonas aeruginosa bloodstream infection | -55 | -48 | Factual
ceftazidime-avibactam | -55 | -48 | Factual
amikacin | -55 | -48 | Factual
SARS-CoV-2 | -53 | -53 | Factual
remdesivir | -53 | -50 | Factual
droplet isolation | -53 | 0 | Factual
recurrence of C. difficile | -50 | -40 | Factual
fidaxomicin | -50 | -40 | Factual
transferred to geriatric medicine unit | -40 | -40 | Factual
bloodstream infection due to Candida parapsilosis | -38 | -21 | Factual
caspofungin | -38 | -21 | Factual
cefazolin | -38 | -21 | Factual
bloodstream infection due to P. aeruginosa | -28 | -18 | Factual
piperacillin-tazobactam | -28 | -21 | Factual
aztreonam | -21 | -14 | Factual
ceftazidime-avibactam | -21 | -14 | Factual
cefepime | -14 | 0 | Factual
tracheostomy closure | -7 | -7 | Factual
nutritional supplementation | -7 | 0 | Factual
discharge | 0 | 0 | Factual
postural transition with assistance | 0 | 0 | Factual
motor and respiratory reconditioning | 0 | 0 | Factual
rehabilitation follow-up | 0 | 0 | Factual
ENT follow-up | 0 | 0 | Factual
geriatric follow-up | 0 | 0 | Factual