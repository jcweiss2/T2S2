18 years old | 0
female | 0
history of untreated hypertension | 0
history of morbid obesity | 0
history of chronic back pain | 0
history of IVDU | 0
presented with worsening low back pain | -144
presented with diffuse abdominal pain | -144
presented with lower extremity weakness | -144
presented with anorexia | -144
presented with fever | -144
presented with chills | -144
presented with shortness of breath | -144
presented with dizziness | -144
presented with constipation | -144
reported recent use of acetaminophen | -144
reported recent use of gabapentin | -144
reported recent use of hydrocodone | -144
reported recent use of methamphetamines | -144
reported recent use of marijuana | -144
admitted to the hospital | 0
blood pressure of 79/53 mmHg | 0
heart rate of 149 bpm | 0
lactic acid of 4.2 mg dl−1 | 0
WBC 37 500 u l−1 | 0
erythrocyte sedimentation rate 75 mm h−1 | 0
urine toxicology positive for cannabis and amphetamines | 0
midline tenderness of the lumbar spine | 0
3/5 strength in bilateral lower extremities | 0
bilateral shoulder warmth, erythema and tenderness | 0
limited range of motion | 0
multiple needle puncture sites on the antecubital fossas bilaterally | 0
smaller puncture wounds between the toes of the right foot | 0
blood cultures collected | 0
empirically started on vancomycin, metronidazole, aztreonam and IV fluids | 0
MRSA with sensitivities to vancomycin, rifampin, levofloxacin, clindamycin, daptomycin, and linezolid | 0
bilateral shoulder plain radiographs showed no abnormalities | 0
arthrocentesis of the acromioclavicular (AC) joints | 0
WBC of 93 137 u l–1 in one shoulder and 32 043 u l–1 in the other | 0
aspirates were cultured and grew MRSA | 0
taken for emergent surgical debridement of the shoulders | 0
intubated | 0
MRI of the lumbar spine showed L3–L5 osteomyelitis with facet septic arthritis, dorsal paraspinous myositis, L2–L5 epidural abscess, and bilateral psoas myositis and abscesses | 0
MRI of the bilateral shoulders after debridement showed septic arthritis of the AC joints, right distal trapezius abscess, and left supraclavicular abscess | 0
MRI of the brain showed no acute intracranial processes | 0
transthoracic echocardiogram (TTE) was negative for any valvular vegetations | 0
repeat surgical debridement of the shoulders was performed | 0
neurosurgery evaluated the patient for possible debridement of the epidural abscess | 0
leukocytosis continued to rise and peaked at 52 100 u l–1 | 0
trough levels of vancomycin were being monitored | 0
repeat blood cultures continued to be positive for MRSA | 0
antibiotics were escalated to daptomycin and ceftaroline | 0
blood cultures became negative on day 14 | 14
rifampin was added to the current antibiotic regimen | 14
repeat MRI of the lumbar spine showed worsening epidural abscess | 14
neurosurgery took the patient for surgical drainage with drain placement | 18
intraoperative wound cultures were positive for MRSA and Proteus mirabilis | 18
improved clinically, all drains were removed | 24
discharged on day 28 | 28
prescribed oral levofloxacin and rifampin for an additional 52 days | 28