8 years old | 0
female | 0
born in Guyana | -4 years * 8760 = -35040
living in France | -4 years * 8760 = -35040
unremarkable familial history | 0
unremarkable medical history | 0
admitted to the hospital | 0
severe bilateral optic neuritis | 0
longitudinally extensive transverse myelitis (LETM) | 0
methylprednisolone | 0
oral tapering steroids | 0
fully recovered | 24 * 3 = 72
another LETM occurred | 5 * 30 * 24 = 3600
AQP4-Ab in the serum | 3600
diagnosis of NMOSD | 3600
immunoadsorptions/plasma exchanges | 3600
mycophenolate mofetil | 3600
RTX | 3600
9 severe relapses | 3600
permanent visual disability | 3600
right amblyopia | 3600
visual acuity | 3600
Expanded Disability Status Scale = 3 | 3600
RTX infusion-related reaction | 6 * 30 * 24 = 4320
anaphylactic-like reaction | 7 * 30 * 24 = 5040
hospitalization in an intensive care unit | 5040
B-cells detected | 5040
severe sepsis | 5040
infection of a central catheter | 5040
subcutaneous OFA | 9 * 12 * 30 * 24 = 77760
one injection of 20 mg every week | 77760
one injection of 20 mg every 4 weeks | 77760 + 4 * 7 * 24 = 78144
detection of antibodies against RTX | 9 * 12 * 30 * 24 + 1 * 12 * 30 * 24 = 90720
no further relapse | 2 * 12 * 30 * 24 = 90720
clinical examination was normal | 11 * 12 * 30 * 24 = 95040
visual disability | 95040
Expanded Disability Status Scale = 3 | 95040
MRI revealed no radiologic activity | 12 * 30 * 24 = 95040
atrophy of optic nerves | 95040
persistent spinal cord lesion | 95040
tolerance was perfect | 95040
no anaphylactic-like nor infectious event | 95040
complete B-cell depletion | 95040
no lymphopenia | 95040
no hypogammaglobulinemia | 95040