16 years old | 0
    primigravida | 0
    admitted to the emergency room | 0
    pregnancy diagnosis of 37.6 weeks | 0
    viable intrauterine pregnancy | 0
    fetal heart rate of 143 beats per minute | 0
    fetus situated longitudinally | 0
    cephalic presentation | 0
    back to the left | 0
    cervix 6 cm dilated | 0
    70% effaced | 0
    station +1 | 0
    intact membranes | 0
    mild edema of the extremities | 0
    normal osteotendinous reflexes | 0
    obstetrical ultrasound performed | 0
    pregnancy of 37+0 weeks | 0
    posterior body placenta | 0
    maturation grade III | 0
    amniotic fluid index of 8.7 cm | 0
    biophysical profile of 8/8 | 0
    Hadlock of 34.2% | 0
    weight of 3033 grams | 0
    decided to continue labor monitoring | 0
    spontaneous rupture of the membranes | -5
    labor progressed over 5 hours | -5
    effective labor | -5
    4 contractions every 10 minutes | -5
    contractions lasted 40 to 45 seconds | -5
    no need for uterotonic agents | -5
    moved to the labor room | -5
    fully dilated | -5
    100% clearance | -5
    station of +3 | -5
    fetus in left occiput anterior position | -5
    live newborn delivered | 0
    Apgar scores of 7 and 9 | 0
    gestational age of 40 weeks | 0
    height 48 cm | 0
    weight of 2650 grams | 0
    placenta came out with Schultze mechanism | 0
    placenta with normal characteristics | 0
    grade III uterine inversion | 0
    maneuvers for manual reinversion performed | 0
    manual reinversion unsuccessful | 0
    total blood loss of 1200 mL | 0
    uterine atony | 0
    use of oxytocin | 0
    use of carbetocin | 0
    use of misoprostol | 0
    persistent uterine inversion | 0
    decided to perform exploratory laparotomy | 0
    under general anesthesia | 0
    evaluated uterine inversion | 0
    reinversion successful | 0
    uterine atony persisted | 0
    postpartum hemorrhage persisted | 0
    decided to place Hayman hemostatic suture | 0
    no response to Hayman suture | 0
    bilateral ligation of anterior trunk of hypogastric artery | 0
    immediate recovery of uterine tone | 0
    cessation of postpartum hemorrhage | 0
    uterus regained tone in 5 minutes | 0
    postligation bleeding of 50 mL | 0
    transfused 2 bags of packed red blood cells | 24
    hemoglobin level of 7 g | 24
    transferred to recovery room | 24
    transferred to medical intensive care unit | 24
    transferred to hospital room | 48
    normal diet | 48
    ambulation | 48
    spontaneous uresis | 48
    normal peristalsis | 48
    breastfeeding | 48
    discharged on the second day | 48
    no postoperative complications | 48
    <|eot_id|>
    
    16 years old | 0
primigravida | 0
admitted to the emergency room | 0
pregnancy diagnosis of 37.6 weeks | 0
viable intrauterine pregnancy |"0
fetal heart rate of 143 beats per minute | 0
fetus situated longitudinally | 0
cephalic presentation | 0
back to the left | 0
cervix 6 cm dilated | 0
70% effaced | 0
station +1 | 0
intact membranes | 0
mild edema of the extremities | 0
normal osteotendinous reflexes | 0
obstetrical ultrasound performed | 0
pregnancy of 37+0 weeks | 0
posterior body placenta | 0
maturation grade III | 0
amniotic fluid index of 8.7 cm | 0
biophysical profile of 8/8 | 0
Hadlock of 34.2% | 0
weight of 3033 grams | 0
decided to continue labor monitoring | 0
spontaneous rupture of the membranes | -5
labor progressed over 5 hours | -5
effective labor | -5
4 contractions every 10 minutes | -5
contractions lasted 40 to 45 seconds | -5
no need for uterotonic agents | -5
moved to the labor room | -5
fully dilated | -5
100% clearance | -5
station of +3 | -5
fetus in left occiput anterior position | -5
live newborn delivered | 0
Apgar scores of 7 and 9 | 0
gestational age of 40 weeks | 0
height 48 cm | 0
weight of 2650 grams | 0
placenta came out with Schultze mechanism | 0
placenta with normal characteristics | 0
grade III uterine inversion | 0
maneuvers for manual reinversion performed | 0
manual reinversion unsuccessful | 0
total blood loss of 1200 mL | 0
uterine atony | 0
use of oxytocin | 0
use of carbetocin | 0
use of misoprostol | 0
persistent uterine inversion | 0
decided to perform exploratory laparotomy | 0
under general anesthesia | 0
evaluated uterine inversion | 0
reinversion successful | 0
uterine atony persisted | 0
postpartum hemorrhage persisted | 0
decided to place Hayman hemostatic suture | 0
no response to Hayman suture | 0
bilateral ligation of anterior trunk of hypogastric artery | 0
immediate recovery of uterine tone | 0
cessation of postpartum hemorrhage | 0
uterus regained tone in 5 minutes | 0
postligation bleeding of 50 mL | 0
transfused 2 bags of packed red blood cells | 24
hemoglobin level of 7 g | 24
transferred to recovery room | 24
transferred to medical intensive care unit | 24
transferred to hospital room | 48
normal diet | 48
ambulation | 48
spontaneous uresis | 48
normal peristalsis | 48
breastfeeding | 48
discharged on the second day | 48
no postoperative complications | 48