55 years old | 0
female | 0
admitted to the hospital | 0
fever | -168
malaise | -168
fatigue | -168
decreased appetite | -168
productive cough | -144
abdominal pain | -144
watery diarrhea | -144
mental status changes | -168
nonresponsive to her name | -168
visual hallucinations | -168
denies headache | 0
denies loss of consciousness | 0
denies neck rigidity | 0
denies seizure | 0
denies focal neurological symptoms | 0
denies chest pain | 0
denies hemoptysis | 0
denies difficulty breathing | 0
allergy to penicillin | 0
returned from Ghana | -432
traveled to California | -168
denies receiving malaria prophylaxis | 0
denies vaccination against yellow fever | 0
denies vaccination against hepatitis A virus | 0
developed symptoms in California | -168
visited a hospital in California | -168
discharged from hospital in California | -168
lethargic | 2
respiratory distress | 2
oral temperature 38.6°C | 2
heart rate 121 beats/min | 2
blood pressure 100/51 mmHg | 2
respiratory rate 45 breaths/min | 2
SpO2 93% | 2
dry mucous membranes | 2
decreased bilateral breath sounds | 2
tenderness to palpation of the left lower quadrant abdomen | 2
no obvious jaundice | 2
no enlarged lymph nodes | 2
no splenomegaly | 2
lethargic and confused | 2
Glasgow coma scale score 14 | 2
pupils equal, round, and reactive to light | 2
no cranial nerve or sensory deficit | 2
neck supple | 2
Brudzinski’s sign negative | 2
Kernig’s sign negative | 2
leukocytosis | 2
white cell count 19 800/µL | 2
neutrophils 44% | 2
lymphocytes 22% | 2
eosinophil 1% | 2
platelets 51 000/µL | 2
hemoglobin 11.8 g/dL | 2
hematocrit 35.3% | 2
red blood cell distribution width 16.9% | 2
lactate dehydrogenase 2714 U/L | 2
haptoglobin <8 mg/dL | 2
prothrombin time/international normalized ratio 14.9/1.4 | 2
troponin 0.161 ng/mL | 2
blood glucose 26 mg/dL | 2
blood urea nitrogen 157 mg/dL | 2
creatinine 7.52 mg/dL | 2
estimated glomerular filtration rate 6 mL/min | 2
bicarbonate 5 mmol/L | 2
anion gap 36 | 2
lactic acid 16.2 mmol/L | 2
sodium 131 mmol/L | 2
potassium 5.5 mmol/L | 2
chloride 91 mmol/L | 2
alanine transaminase 542 U/L | 2
aspartate transaminase 1328 U/L | 2
total bilirubin 14.5 mg/dL | 2
albumin 2.2 mg/dL | 2
malaria smear positive | 2
parasitemia 25% | 2
ring forms/trophozoites | 2
developing gametocytes | 2
arterial blood gas pH 7.03 | 2
pCO2 20 | 2
HCO3 0 | 2
intubated and mechanically ventilated | 5
transferred to ICU | 5
severe malaria diagnosed | 5
Plasmodium falciparum malaria | 5
multi-organ failure | 5
respiratory failure | 5
renal failure | 5
hepatic failure | 5
septic shock | 5
disseminated intravascular coagulation | 5
cerebral malaria | 5
acute toxic-metabolic encephalopathy | 5
acute hypoxemic respiratory failure | 5
acute respiratory distress syndrome | 5
vasopressors started | 5
steroids started | 5
infectious disease consultation | 5
IV quinidine started | 5
IV doxycycline started | 5
CDC contacted | 5
empiric broad-spectrum antibiotic coverage started | 5
IV meropenem started | 5
IV vancomycin started | 5
QTc prolongation | 24
quinidine switched to IV artesunate | 24
parasitemia improved | 24
acidosis improved | 24
positive end-expiratory pressure decreased | 24
FiO2 requirements decreased | 24
computed tomography of the brain unremarkable | 48
lumbar puncture | 48
white blood cells 3 per high-power field | 48
neutrophils 12% | 48
lymphocytes 48% | 48
monocytes 38% | 48
no organisms on gram stain | 48
vancomycin discontinued | 48
meropenem discontinued | 48
parasitemia 0.3% | 120
parasitemia negative | 144
multi-organ failure treated | 144
septic shock treated | 144
disseminated intravascular coagulation treated | 144
renal replacement therapy | 144
platelet transfusions | 144
patient clinically improving | 144
IV artesunate completed | 120
oral doxycycline started | 120
discharged to rehabilitation facility | 168