30 years old | 0
male | 0
Saethre-Chotzen syndrome | 0
open surgical pulmonic valvotomy | -672
pulmonary outflow homograft patch | -672
presented to a community hospital | 0
shortness of breath | 0
abdominal pain | 0
nausea | 0
vomiting | 0
gastric bypass | -672
morbid obesity | -672
BMI 42 | -672
bilateral lower extremity swelling | -672
antibiotics | -672
steroids | -672
admission HR 90 | 0
BP 140/80 mmHg | 0
RR 27 breaths per minute | 0
pulse oximetry 92% | 0
antibiotics initiated | 0
nasal cannula oxygen | 0
intravenous fluids | 0
chest x-ray low lung volumes | 0
acute left lower extremity superficial thrombophlebitis | 0
CT angiography no acute pulmonary embolism | 0
significant cardiomegaly | 0
central pulmonary artery enlargement | 0
cholelithiasis | 0
nephrolithiasis | 0
left intrarenal calculus | 0
right kidney wedge-shaped infarct | 0
small cerebellar infarct | 0
transferred to intensive care unit | 24
BiPAP initiated | 24
intubated | 168
mechanical ventilation initiated | 168
lung protective ventilation | 168
ARDS diagnosis | 168
high PEEP strategy | 168
MAP <60 mmHg | 168
norepinephrine initiated | 168
vasopressin initiated | 168
FiO2 1.0 | 168
PEEP 16 | 168
ABG pH 7.4 | 168
ABG pCO2 41 | 168
ABG paO2 42 | 168
ECMO activation | 168
CT scan no bilateral opacities | 168
no echocardiography | 168
inhaled nitric oxide initiated | 168
iNO 40 ppm | 168
oxygen saturation improved to 94% | 168
paO2 65.9 | 168
transferred to our institution | 168
transesophageal echocardiogram performed | 168
large intra-atrial bidirectional shunt | 168
severe pulmonary regurgitation | 168
enlarged pulmonary artery 4.9 cm | 168
absent left main coronary artery | 168
separate ostial connections | 168
bronchoscopy performed | 168
significant secretions right bronchial lower lobe | 168
influenza B positive | 168
pulmonary artery catheter placed | 168
pulmonary regurgitation | 168
IAS correction deferred | 168
concern for sepsis | 168
continued iNO | 168
diuresis | 168
vasopressor wean | 168
hypoxemia | 168
day four after admission | 96
cardiac catheterization laboratory | 96
PFO closure device placed | 96
oxygen saturation improved acutely | 96
residual R-L shunt | 96
severe pulmonary regurgitation | 96
weaned off iNO | 240
day twelve | 288
tracheostomy performed | 288
ventilator weaning | 288
ICU day fifteen | 360
CT scans | 360
left cerebellar vermis infarct | 360
improved interstitial edema | 360
device migration | 360
angiographic removal | 360
hospital day nineteen | 456
mechanical ventilation discontinued | 456
supplemental oxygen via tracheostomy collar | 456
discharged to acute rehabilitation unit | 456
home oxygen 2-4L | 456
six months post-discharge | 4320
atrial septal defect closure | 4320
pulmonic valve replacement | 4320
pulmonary artery patch graft | 4320
normal prosthetic pulmonary valve function | 4320
ASD closed | 4320
negative bubble study | 4320
