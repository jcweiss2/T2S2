74 years old | 0
male | 0
admitted to the hospital | 0
lower abdominal pain | -96
signs of infection | -96
deterioration in overall well-being | -96
uncontrolled diabetes mellitus | -6720
metformin | -6720
right femur fracture | -17280
sequela of stroke | -17280
motor aphasia | -17280
facial paralysis | -17280
urethral stenosis | -6720
recurrent urinary tract infections | -6720
intravenous antibiotics | -144
dysuria | -96
fever | -96
pneumaturia | -96
lower abdominal tenderness | 0
hyperglycemia | 0
elevated inflammatory markers | 0
C-reactive protein | 0
lactate levels | 0
leukocytes in urine | 0
nitrites in urine | 0
diffuse thickening of the bladder wall | 0
air bubbles in the bladder wall | 0
intraparenchymal air bubbles | 0
intrluminal gas in the bladder | 0
white blood cells in urine | 0
red blood cells in urine | 0
emphysematous cystitis | 0
broad-spectrum antimicrobial therapy | 0
ceftriaxone | 0
metronidazole | 0
gentamicin | 0
urinary catheter insertion | 0
cloudy urine | 0
gas in urine | 0
polymorphic flora | 0
intensive care unit | 0
close clinical and biochemical monitoring | 0
vigilant surveillance strategy | 0
bladder necrosis | 0
abscess formation | 0
bladder perforation | 0
intravenous antibiotics | 0
insulin therapy | 0
improvement in overall condition | 336
discharged from the hospital | 480