64 years old | 0
female | 0
admitted to the hospital | 0
severe headache | 0
right periorbital and mid-facial swelling | 0
fever | -336
headache | -336
light pain in the right ear | -336
purulent secretion from the ear | -336
swelling and redness of the skin behind the right ear | -336
tinnitus | -336
hearing disorder | -336
right acute mastoiditis | -336
Amoxicillin | -336
painkillers | -336
anti-inflammatory drugs | -336
improved slightly | -192
severe headache | -192
anorexia | -192
high fever | -192
confusion | -192
arterial hypertension | 0
angiotensin-converting enzyme inhibitors | 0
right facial and periorbital swelling | 0
right blepharoptosis | 0
chemosis | 0
proptosis | 0
visual acuity of 7/12 on her right eye | 0
no visual fields abnormalities | 0
intraocular pressures in both eyes were normal | 0
no relative afferent pupillary defect | 0
color vision was normal | 0
no signs of optic disc swelling | 0
febrile | 0
conscious, but somnolent | 0
no other neurological deficits | 0
inflammatory parameters were significantly elevated | 0
renal and liver functions within normal limits | 0
prothrombin G20210A mutation | 0
coagulation profile and urinalysis were both normal | 0
non-opacification of the right cavernous sinus | 0
Ceftriaxone | 0
Enoxaparin | 0
shortness of breath | 96
reduced oxygen saturation | 96
unilateral homogeneous opacification on right lobar lung | 96
air bronchograms | 96
right lobar pneumonia | 96
non-invasive mechanical ventilation | 96
Amikacin | 96
Piperacillin–Tazobactam | 96
improved | 168
symptoms resolved | 168
control contrast-enhanced magnetic resonance angiography | 168
persistence of the lacunar image in the right cavernous sinus | 168
ophthalmological symptoms improved | 168
periorbital swelling has diminished | 168
discharged | 336
oral anticoagulant – Acenocoumarol | 336
follow-up CT venogram | 504
full recovery | 504