74 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
hypertension | 0 | 0 | Factual
insulin-dependent diabetes mellitus type 2 | 0 | 0 | Factual
diabetic retinopathy | 0 | 0 | Factual
weight loss | -168 | 0 | Factual
iron deficiency anemia | -168 | 0 | Factual
tumor in the colon ascendens | -168 | 0 | Factual
liver metastases | -168 | 0 | Factual
right hemicolectomy | 0 | 0 | Factual
low-grade pT3cN0 adenocarcinoma | 0 | 0 | Factual
absence of metastases in 24 excised lymph nodes | 0 | 0 | Factual
lymphovascular growth | 0 | 0 | Factual
no vascular or perineural growth | 0 | 0 | Factual
activated BRAF mutation | 0 | 0 | Factual
loss of expression of MLH1 and PMS2 | 0 | 0 | Factual
mismatch repair-deficient (MMR-D)/microsatellite-instable (MSI) tumor | 0 | 0 | Factual
pembrolizumab therapy | 0 | 336 | Factual
symptoms of a cold | 168 | 168 | Factual
leukocytosis | 168 | 168 | Factual
slight increase in C-reactive protein | 168 | 168 | Factual
dry coughing | 528 | 528 | Factual
no fever | 528 | 528 | Factual
increase in AST and ALT | 528 | 528 | Factual
ICI-induced hepatitis grade 2 | 528 | 528 | Factual
prednisolone therapy | 528 | 1008 | Factual
decrease in C-reactive protein and AST | 528 | 1008 | Factual
increase in white blood cells and neutrophils | 528 | 1008 | Factual
dyspnea | 696 | 696 | Factual
myocardial infarction suspected | 696 | 696 | Factual
elevation of troponin T | 696 | 696 | Factual
septal hypokinesia | 696 | 696 | Factual
no dynamic change in troponin T | 696 | 696 | Factual
somnolence | 720 | 720 | Factual
difficulty walking | 720 | 720 | Factual
dysarthria | 720 | 720 | Factual
hoarseness | 720 | 720 | Factual
pain in neck and right leg | 720 | 720 | Factual
difficulty raising right leg | 720 | 720 | Factual
increase in prednisolone dose | 720 | 720 | Factual
no signs of stroke | 720 | 720 | Factual
increase in creatine kinase and myoglobin levels | 720 | 720 | Factual
ICI-induced myositis suspected | 720 | 720 | Factual
gradual decrease in creatinine levels | 720 | 1008 | Factual
antibodies against acetylcholine receptor and titin | 720 | 720 | Factual
myasthenia gravis (MG) | 720 | 720 | Factual
albumin in cerebrospinal fluid | 720 | 720 | Factual
inability to sit up | 1008 | 1008 | Factual
severe dysarthria and dysphagia | 1008 | 1008 | Factual
need for oxygen | 1008 | 1008 | Factual
absent reflexes | 1008 | 1008 | Factual
transfer to intensive care unit | 1008 | 1008 | Factual
intubation | 1032 | 1032 | Factual
methylprednisolone therapy | 1032 | 1064 | Factual
intravenous immunoglobulins | 1032 | 1032 | Factual
infliximab therapy | 1104 | 1104 | Factual
improvement in muscle strength | 1128 | 1128 | Factual
carbon dioxide retention | 1164 | 1164 | Factual
noninvasive ventilation | 1164 | 1164 | Factual
sinus bradycardia | 1164 | 1164 | Factual
death | 1164 | 1164 | Factual
respiratory insufficiency | 1164 | 1164 | Factual
polymyositis | 1164 | 1164 | Factual
autopsy | 1164 | 1164 | Factual
significant stenosis of right coronary artery | 1164 | 1164 | Factual
no fibrosis or signs of recent myocardial infarction | 1164 | 1164 | Factual
softened tongue | 1164 | 1164 | Factual
no surgical complication after hemicolectomy | 1164 | 1164 | Factual
liver metastasis | 1164 | 1164 | Factual
hepatocellular cancer (HCC) | 1164 | 1164 | Factual
response to pembrolizumab therapy | 1164 | 1164 | Factual
inflammatory infiltration of lymphocytes | 1164 | 1164 | Factual
fibrosis | 1164 | 1164 | Factual
myocardial infarction | 1164 | 1164 | Factual
inflammatory infiltrate | 1164 | 1164 | Factual