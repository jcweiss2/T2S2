admitted to the emergency room | 0
pregnancy diagnosis of 37.6 weeks of gestation | 0
viable intrauterine pregnancy | 0
fetal heart rate of 143 beats per minute | 0
fetus situated longitudinally with cephalic presentation | 0
cervix 6 cm dilated | 0
70% effaced | 0
station +1 | 0
intact membranes | 0
mild edema of the extremities | 0
normal osteotendinous reflexes | 0
obstetrical ultrasound | 0
pregnancy of 37+0 weeks of gestation | 0
posterior body placenta maturation grade III | 0
amniotic fluid index of 8.7 cm | 0
biophysical profile of 8/8 | 0
Hadlock of 34.2% | 0
weight of 3033 grams | 0
continue labor monitoring | 0
spontaneous rupture of the membranes | -5
7 cm dilation | -5
labor progressed over 5 hours | -5
effective labor | -5
4 contractions every 10 minutes | -5
contractions lasted 40 to 45 seconds | -5
no need for uterotonic agents | -5
moved to the labor room | -5
fully dilated | -5
100% clearance | -5
station of +3 | -5
fetus in left occiput anterior position | -5
live newborn delivered | 0
Apgar scores of 7 and 9 | 0
gestational age of 40 weeks | 0
height 48 cm | 0
weight of 2650 grams | 0
placenta came out with normal characteristics | 0
grade III uterine inversion | 0
manual reinversion maneuvers performed | 0
total blood loss of 1200 mL | 0
UA | 0
oxytocin used | 0
carbetocin used | 0
misoprostol used | 0
persistent uterine inversion | 0
exploratory laparotomy | 1
utrine inversion evaluated | 1
reinversion successful | 1
UA persisted | 1
PPH | 1
Hayman hemostatic suture placed | 1
no response to Hayman suture | 1
bilateral ligation of the anterior trunk of the hypogastric artery | 2
immediate recovery of uterine tone | 2
cessation of PPH | 2
uterus regained tone in approximately 5 minutes | 2
postligation bleeding of 50 mL | 2
2 bags of packed red blood cells transfused | 2
gasometry showed a hemoglobin level of 7 g | 2
transferred to the recovery room | 3
transferred to the medical intensive care unit | 3
transferred to a hospital room | 24
normal diet | 24
ambulation | 24
spontaneous uresis | 24
normal peristalsis | 24
breastfeeding | 24
discharged on the second day | 48
no postoperative complications | 48