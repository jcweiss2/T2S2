71 years old | 0
female | 0
arthritis | -8760
central serous retinopathy | -8760
deep vein thrombosis | -8760
hyperlipidemia | -8760
osteoporosis | -8760
fatigue | -216
abdominal pain | -216
loss of appetite | -216
anemia | 0
mild thrombocytopenia | 0
abnormal liver function tests | 0
hemoglobin 10.7 g/dL | 0
Na+ 128 mmol/L | 0
AST 110 U/L | 0
ALT 73 U/L | 0
GGTP 94 U/L | 0
albumin 2.6 gm/dL | 0
hepatic and portal vein thrombosis | 0
hepatitis | 0
pancreatitis | 0
colitis | 0
right hepatic vein thrombosis | 0
pancreatic tail mass | 0
pancreatic carcinoma | 0
pancreatic neuro-endocrine tumor | 0
CT-guided needle core biopsy | 0
diffuse large B-cell lymphoma | 0
cell block | 0
CD20 positive | 0
CD79a positive | 0
CD45 positive | 0
PAX-5 positive | 0
MUM-1 non-contributory | 0
Ki-67 high | 0
bone marrow aspirate | 0
bone marrow biopsy | 0
no bone marrow involvement | 0
Weisella confusa bacteremia | 24
Enterococcus faecalis bacteremia | 24
piperacillin-tazobactam | 24
up-trending creatinine | 48
elevated lactate dehydrogenase | 48
diastolic blood pressure fluctuating | 48
up-trending liver function tests | 48
vancomycin | 72
meropenem | 72
metronidazole | 96
septic shock | 96
intubated | 120
norepinephrine drip | 120
stress dose steroids | 120
disseminated intravascular coagulopathy | 144
pulmonary emboli | 144
multi-organ failure | 168
death | 312
autopsy | 312
pancreatic mass | 312
lymphoma cells | 312
intravascular lymphomatous proliferation | 312
CD20 positive | 312
MUM1 weak | 312
Pax-5 weak | 312
CD5 positive | 312
CD3 negative | 312
CD10 negative | 312
Ki-67 high | 312
Epstein-Barr encoding region negative | 312