45 years old | 0
female | 0
admitted to the hospital | 0
severe lower abdominal | -12
bright red per rectal bleeding | -12
diagnosed with right-sided colon cancer | - months 
pelvic side wall lymph node metastases | - months 
surgery | - months 
R0 resection | - months 
radiotherapy | - weeks 
adjuvant FOLFOX chemotherapy | -168
nausea | -168
abdominal discomfort | -168
constipation | -168
schizophrenia | 0
Clozapine | 0
tachycardia | 0
high-grade fevers | 0
worsening pain | 0
pneumoperitoneum | 0
sigmoid faecaloma | 0
stercoral perforation | 0
ischaemic changes | 0
emergency laparotomy | 0
grossly dilated sigmoid colon | 0
redundant sigmoid colon | 0
inspissated faecaloma | 0
necrosis of the wall | 0
Hartmann’s procedure | 0
extensive washout | 0
vasopressor support | 0
septic shock | 0
granulocyte colony stimulating factor (G-CSF) | 0
febrile neutropaenia | 0
suspended Clozapine | 0
recovered well post-operatively | 240
discharged to rehabilitation | 240
full thickness perforation | 0
ischaemic necrosis | 0
massive faecaloma | 0
stercoral perforation | 0