29 years old | 0
female | 0
native mitral and aortic valve endocarditis | 0
active IVDU | 0
mother of two young children | 0
poor social support network | 0
admitted to Emergency Department | 0
underplayed severity of cardiac condition | 0
unwilling to quit IVDU | 0
initial decision to treat conservatively | 0
antibiotic therapy | 0
developed severe cardiogenic shock | 24
severe aortic and mitral valve regurgitation | 24
referred for emergency inpatient cardiac surgery | 24
obtained mother's consent | 24
aortic valve replacement | 24
complex mitral valve repair | 24
could not be weaned off cardiopulmonary bypass machine | 24
severe biventricular dysfunction | 24
postcardiotomy venoarterial ECMO | 24
five days of clinical progress | 120
one failed attempt to wean off ECMO | 120
successfully discontinued ECMO | 168
remained in ICU | 168
total of 75 days in hospital | 1800
discharged to local convalescence center | 1800
continuation of rehabilitation | 1800
COVID-19 pandemic | -1000
peak of COVID-19 pandemic | 0
limited resources | 0
shortage of ICU beds | 0
shortage of nurses | 0
shortage of cardiac surgical operating rooms | 0
shortage of ECMO machines | 0
shortage of perfusionists | 0
high-risk cardiac surgical procedure | 24
high possibility of developing prosthetic valve endocarditis | 24
postoperative complications | 24
high mortality rates | 24
prolonged postoperative hospital stays | 168
massive consumption of resources | 168
ethical principle of stewardship | 0
decision to perform surgery | 24
contingency plan of rehabilitation | 24
close community follow-up | 24
organization support from Street Health | 24
protect patient's children | 24
use of ECMO for patients with active endocarditis and IVDU | 24
limited experience with percutaneous ECMO | 0
longer hospital stays | 168
higher rates of complications | 168
moral distress | 24
allocation of scarce resources | 0
rationing of ECMO | 0
stringent eligibility criteria | 0
patient's ability to appreciate harm of IVDU | 0
choice to pursue ECMO | 24
patient's survival | 24
future rehabilitation | 1800
long-term mechanical circulatory support | 168
limited evidence to guide patient selection | 0
expert opinion against long-term support | 0
social support and ventricular device care programs | 1800
heart transplantation | 1800
high-risk procedure | 1800
intense immunosuppression | 1800
satisfactory social support network | 1800
no reports of heart transplants in patients with infective endocarditis due to active IVDU | 0
patient's options slim | 168
ability to refrain from IVDU | 1800
potential LVAD or cardiac transplantation | 1800
healthcare team's wish to avoid | 168
allocation of scarce resources amidst COVID-19 pandemic | 0
main ethical dilemma | 0
rapid rise in cases | 0
elevated needs for life support systems | 0
stringent eligibility criteria | 0
patient eligible for ECMO | 24
no other co-morbidities | 0
vast limitation in resources | 0
decision difficult to pursue ECMO | 24
patient tolerated ECMO | 168
slowly weaned off | 168
long recovery | 1800
multidisciplinary team approach | 168
postoperative abstinence from IVDU | 1800
education on dangers of IVDU | 168
intensive counseling | 168
critical need for patient to abstain from IVDU | 168
patient's mind changed | 1800
promised to never use intravenous drugs again | 1800
one-month follow-up appointment | 720
close follow-up throughout care | 1800