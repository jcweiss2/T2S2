60 years old | 0
male | 0
admitted to the hospital | 0
fever | -2
hypotension | -2
altered mental status | -2
low back pain | -2
epigastric pain | -2
chills | -2
vomiting | -2
disoriented | -2
dusky discoloration of face and extremities | -2
splenectomy | -44160
cholecystectomy | -7300
multiple laparotomies | -7300
dog bites | -168
scratches from dog | -168
intravenous fluids | 0
packed red blood cells | 0
levofloxacin | 0
CT scan of chest, abdomen, and pelvis | 0
acute respiratory distress syndrome | 0
intubated | 2
worsening confusion | 2
hypoxemia | 2
transferred to hospital | 2
heavily sedated | 2
mechanically ventilated | 2
blood pressure 80/58 mmHg | 2
heart rate 111 beats per minute | 2
temperature 38.5°C | 2
coarse breath sounds | 2
absent peripheral pulses | 2
cold, dusky extremities | 2
mottling of skin | 2
violaceous purpura on thighs | 2
superficial linear scratches | 2
erythema | 2
intravenous fluids | 2
vasopressors | 2
blood cultures collected | 2
white blood cell count 18.0 × 10^9/L | 2
platelet count 14 × 10^9/L | 2
international normalized ratio 1.7 | 2
fibrinogen 178 mg/dL | 2
creatinine 3.8 mg/dL | 2
lactate 5.6 mmol/L | 2
PaO2 60 mmHg | 2
urinalysis | 2
erythrocytes and leukocytes in urine | 2
protein in urine | 2
bilirubin in urine | 2
bacteria in urine | 2
empiric broad-spectrum antibiotics | 2
vancomycin | 2
cefepime | 2
ampicillin | 2
doxycycline | 2
acyclovir | 2
CT scan of head | 4
lumbar puncture | 4
cerebrospinal fluid analysis | 4
Gram stain | 4
herpes simplex virus PCR | 4
ampicillin discontinued | 4
acyclovir discontinued | 4
continuous renal replacement therapy | 4
peripheral blood Wright's stain | 6
neutrophils with blue inclusions | 6
buffy coat Gram stain | 6
Gram-negative rods | 6
cefepime changed to piperacillin-tazobactam | 6
ciprofloxacin | 6
NGS assay | 96
plasma sample sent for analysis | 96
microbial DNA detected | 120
Capnocytophaga canimorsus identified | 120
antibiotic regimen narrowed | 120
piperacillin-tazobactam monotherapy | 120
blood culture grew Gram-negative rods | 120
Gram stain morphology | 120
MALDI-TOF attempted | 120
16S ribosomal ribonucleic acid PCR sequencing attempted | 120
Clostridium difficile colitis | 600
Candida tropicalis fungemia | 600
recurrent sepsis | 624
gangrene of upper and lower extremities | 624
comfort care only | 624
patient died | 960
postmortem analysis | 960
16S sequencing confirmed Capnocytophaga canimorsus | 960