74 years old | 0
male | 0
admitted to the hospital | 0
altered mental status | 0
fever | -48
cough with mucopurulent sputum | -48
abdominal pain | -48
hypertension | -6720
gastroesophageal reflux | -6720
moderate alcohol consumption | -6720
lansoprazole | -6720
perindopril | -6720
amlodipine | -6720
disoriented | 0
uncooperative | 0
blood pressure 135/85 mmHg | 0
heart rate 103 beats/min | 0
respiratory frequency 18 breaths/min | 0
peripheral oxygen saturation 85% | 0
tympanic temperature 39.6 °C | 0
livedo reticularis | 0
increased capillary refill time | 0
bilateral rhonchi | 0
intense epigastric and right hypochondrium pain | 0
muscle guarding | 0
hypoxic respiratory failure | 0
leukocytosis with neutrophilia | 0
altered liver profile | 0
aspartate aminotransferase 1896 U/L | 0
alanine aminotransferase 640 U/L | 0
lactate dehydrogenase 2499 U/L | 0
alkaline phosphatase 230 U/L | 0
total bilirubin 4.78 mg/dL | 0
increased blood lactate level | 12
C-reactive protein increased | 12
procalcitonin 83.86 ng/mL | 12
blood cultures sent | 12
piperacillin/tazobactam started | 12
abdominal CT scan | 12
diffuse heterogeneous structure with hypodensity within the right lobe of the liver | 12
areas with gas within the right lobe of the liver | 12
emphysematous hepatitis diagnosed | 12
acute liver failure diagnosed | 12
severe metabolic acidosis | 24
distributive shock | 24
vasopressor support started | 24
vancomycin started | 48
metronidazole started | 48
fluconazole started | 48
multiorgan failure | 72
died | 72
blood cultures grew Escherichia coli | 72
autopsy decision deterred | 72