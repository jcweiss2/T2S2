58 years old | 0
female | 0
hypertension | -8760
generalized anxiety disorder | -8760
depression | -8760
hepatitis C | -8760
diagnosed with retroperitoneal leiomyosarcoma | -720
radical resection of the tumor | -720
segmental duodenectomy | -720
inferior vena cava closure | -720
nausea | -48
vomiting | -48
right upper quadrant abdominal pain | -48
biopsy confirmed recurrent disease | -48
started on chemotherapy | -48
AIM75/10 | -48
doxorubicin | -48
ifosfamide | -48
mesna | -48
neutropenic fever | -24
thiamine | -24
bisacodyl | -24
docusate-senna | -24
clonidine | -24
losartan | -24
nifedipine | -24
ondansetron | -24
dexamethasone | -24
metoclopramide | -24
oxycodone | -24
fluconazole | -24
paroxetine | -24
altered mental status | 0
confusion | 0
memory impairment | 0
inability to follow commands | 0
inability to form coherent speech | 0
total delirium observation score 10 | 0
increased thiamine dose | 0
methylene blue | 0
discontinued paroxetine | 0
worsening confusion | 6
total delirium observation score 13 | 6
severe sinus tachycardia | 6
hypertension | 6
diaphoresis | 6
fever | 6
combativeness | 6
hyperreflexia | 6
ocular clonus | 6
spontaneous muscular clonus | 6
facial tremors | 6
discontinued methylene blue | 6
discontinued ondansetron | 6
IV lorazepam | 6
metoprolol | 6
acetaminophen | 6
hydromorphone | 6
transferred to critical care unit | 6
intubation | 6
elevated measures of care | 6
normal laboratory tests | 6
workup for sepsis | 6
computed tomography | 6
magnetic resonance imaging | 6
continued thiamine | 6
supportive care | 6
mentation improved | 144
extubated | 144
discharged from hospital | 360
follow-up appointment | 720
surgical resection | 2160
no evidence of disease | 2880