10 years old| 0
    male | 0
    papulovesicular skin lesions | -240
    fever | -96
    lesions over hands | -240
    lesions over lower abdomen | -240
    lesions over perineal areas | -240
    lesions over buttocks | -240
    altered sensorium | -24
    malena | -24
    respiratory rate 32/min | 0
    heart rate 173/min | 0
    capillary refill time 4 seconds | 0
    blood pressure 90/50 mm Hg | 0
    SpO2 93% in room air | 0
    poor peripheral pulses | 0
    severe pallor | 0
    crusted pus discharging lesions over hands | 0
    crusted pus discharging lesions over lower abdomen | 0
    crusted pus discharging lesions over perineal area | 0
    crusted pus discharging lesions over buttocks | 0
    Glasgow Coma Scale score E4M4V4 | 0
    generalized hypotonia | 0
    elicitable deep tendon reflexes | 0
    flexor plantar reflex | 0
    no cranial nerve palsies | 0
    absent meningeal signs | 0
    normal systemic examinations | 0
    infected scabies considered | 0
    septic shock considered | 0
    disseminated intravascular coagulation considered | 0
    upper gastrointestinal bleeding considered | 0
    normal saline boluses resuscitation | 0
    intravenous adrenaline infusion | 0
    intravenous noradrenaline infusion | 0
    intravenous vasopressin infusion | 0
    intravenous dobutamine infusion | 0
    packed red blood cells transfusion | 0
    intravenous antibiotics administration | 0
    mechanical ventilation | 0
    shifted to pediatric intensive care unit | 6
    acute kidney injury | 48
    peritoneal dialysis | 48
    deranged liver function tests | 0
    inotropes tapered | 96
    inotropes stopped | 96
    extubated | 144
    severe anemia | 168
    hypotensive shock | 168
    multiple episodes of massive malena | 168
    fluid boluses resuscitation | 168
    PRBCs transfusions | 168
    vasoactive drugs administration | 168
    upper gastrointestinal endoscopy | 168
    bleeding lesion in first part of duodenum | 168
    computed tomography angiography | 168
    gastroduodenal artery pseudoaneurysm | 168
    digital subtraction angiography guided coil embolization | 168
    transiently controlled bleeding | 168
    massive episodes of malena | 180
    PRBC transfusion | 180
    second endovascular cyanoacrylate glue embolization | 192
    life-threatening upper gastrointestinal bleeding | 192
    massive PRBC transfusion | 192
    fresh frozen plasma transfusion | 192
    platelet concentrates transfusion | 192
    normal amylase levels | 192
    normal ANA | 192
    normal ANCA | 192
    normal HBsAg | 192
    normal HCV | 192
    normal HIV reports | 192
    laparotomy | 216
    duodenostomy | 216
    ligation of gastroduodenal artery aneurysm | 216
    upper gastrointestinal bleeding stopped | 216
    inotropes tapered | 264
    respiratory support tapered | 264
    extubated | 264
    critical illness neuromyopathy | 264
    discharged | 600
    ambulatory at 6 months follow-up | 0
    no recurrence of symptoms | 0
    