42 years old|0
female|0
admitted to the hospital|0
JIA|-108000
anakinra|-108000
hydroxychloroquine|-108000
chronic adrenal insufficiency|-108000
hydrocortisone|-108000
seizure disorder|-108000
culture negative infective endocarditis|-108000
cardioembolic stroke|-108000
mechanical fall|-168
C7 vertebral fracture|-168
cervical collar|0
pain control|0
acute on chronic hypoxic respiratory failure|0
hypercapnic respiratory failure|0
rescue BiPAP|0
encephalopathic|0
respiratory acidosis|0
carbon dioxide retention (>105 mm Hg)|0
intubated|0
computed tomography thorax|0
left-sided opacification|0
left-sided pneumonia|0
adequate antibiotic therapy|0
failed spontaneous breathing trials|0
neuromuscular weakness|0
left-sided diaphragmatic weakness|0
tracheotomy|312
percutaneous endoscopic gastrostomy|312
subarachnoid hemorrhage|0
comminuted fracture of the distal left tibia|0
progressive weakness|-8760
progressive muscular weakness (worsening over past year)|-8760
mechanical ventilation|0
nonverbal status|0
serum aldolase elevated (11.8 U/L)|0
serum aldolase normalized (4.6 U/L)|96
creatine kinase normal (70 U/L)|0
thyroid-stimulating hormone elevated (8.15 IU/mL)|0
free thyroxine normal (0.98 ng/dL)|0
alanine aminotransferase elevated (36 U/L)|0
aspartate aminotransferase elevated (62 U/L)|0
bilirubin normal|0
creatinine low (0.2-0.4 mg/dL)|0
wheelchair use|0
hematuria (past)|-108000
secondary systemic lupus erythematosus|-108000
synovitis (both hands)|0
Enterococcus faecalis urinary tract infection|0
septic shock|0
muscle weakness (all extremities)|0
proximal muscles affected (⅗ strength)|0
distal muscles affected (⅘ strength)|0
hyporeflexic|0
clonus (both ankles)|0
brain MRI consistent with prior stroke|0
bilateral encephalomalacia|0
spinal MRI unremarkable|0
EMG suggested myopathy|0
decreased motor unit recruitment (proximal extremities)|0
myopathic changes (proximal muscles)|0
irritability (proximal and distal arm muscles)|0
myositis panel negative|0
muscle biopsy|0
granular myopathy|0
rimmed vacuoles|0
type II fiber atrophy|0
scattered inflammation|0
electron microscopy (autophagosomes)|0
curvilinear bodies|0
CD3 positive (T-lymphocytes)|0
CD68 positive (histiocytes)|0
hydroxychloroquine-induced myopathy|0
continued hydroxychloroquine|0
inpatient physical therapy|0
hydroxychloroquine level (763 ng/mL)|0
hydrocortisone continued|0
discontinuation of hydroxychloroquine|0
respiratory failure reversed|0
