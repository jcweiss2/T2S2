40 years old|0
female|0
obesity|0
confusion|0
dysuria|0
CT scan showing left EPN|0
transferred to tertiary care center|0
admitted to Medical ICU|0
awake|0
oriented|0
denied hematuria|0
denied flank pain|0
denied chest pain|0
denied shortness of breath|0
denied history of nephrolithiasis|0
afebrile|0
tachycardic|0
normotensive|0
tachypneic|0
saturating well on room air|0
WBC of 34|0
platelet count 66|0
lactate 5.8|0
BUN 56|0
creatinine 3.22|0
glucose 485|0
alkaline phosphatase 498|0
AST 39|0
ALT 43|0
Hemoglobin A1C 7.6|0
urine cultures grew E. coli|0
blood cultures grew E. coli|0
suprapubic tenderness|0
CT imaging revealed gas within left kidney parenchyma|0
4 mm stone within proximal left ureter|0
no hydronephrosis|0
air in collecting systems of both kidneys|0
no definite parenchymal gas on right|0
CT revealed heterogenous liver with cirrhotic nodules|0
moderate abdominal ascites|0
no drainable collection|0
diagnosed with Child Class C cirrhosis|0
started on rifaximin|0
started on lactulose|0
workup not completed|0
nonalcoholic fatty liver disease considered|0
MELD-Na score 31|0
guarded prognosis|0
initial management included intravenous fluids|0
insulin drip|0
Zosyn|0
insertion of bilateral double J stents|0
retrograde pyelogram showed no hydroureteronephrosis|0
foley left in place|0
worsening acidosis|0
required continued intubation|0
returned to ICU in stable condition|0
required dialysis|72
required bicarbonate drip|72
required pressors|72
tachypnea|72
low volumes prevented extubation|72
family updated|72
wish to proceed with surgery only if percutaneous drainage not possible|72
repeat CT scan obtained|72
CT showed worsening left EPN|72
near complete necrosis of left renal upper pole|72
new right EPN|72
new right colon pneumatosis|72
new portal venous gas|72
planning for definitive surgical intervention|72
emergent left nephrectomy|72
general surgery consulted|72
bowel resection considered|72
concern surgery would be fatal|72
decision for comfort measures|72
terminally extubated|96
died|96
