39 years old | 0
male | 0
untreated arterial hypertension | 0
admitted to the Institute of Cardiology | 0
suspected acute coronary syndrome | 0
atypical chest pain | 0
blood pressure 180/110 mm Hg | 0
heart rate of 74 beats per minute | 0
loud systolic murmur | 0
no symptoms of heart failure | 0
ECG sinus rhythm 73 beats per minute | 0
left ventricle hypertrophy | 0
negative T waves in II, III, aVF | 0
coronary angiography | 0
atherosclerotic lesions | 0
maximum luminal diameter stenosis 30–40% in the right coronary artery | 0
troponin I level 0.03 ng/ml | 0
troponin I level 0.07 ng/ml | 0
D-dimer level elevated 1.0 µg/ml | 0
ACS excluded | 0
echocardiography | 0
bicuspid aortic valve | 0
degenerative changes | 0
calcifications | 0
aortic stenosis | 0
mean pressure gradient 45 mm Hg | 0
mild aortic regurgitation | 0
disproportionate concentric left ventricle hypertrophy | 0
maximum wall thickness 1.7 cm | 0
normal left ventricle systolic function | 0
LVEF 65% | 0
ascending aorta diameter 5.6 cm | 0
indexed for body surface area 2.6 cm/m² | 0
Z-score 9.23 | 0
thoracic aortic aneurysm | 0
computed tomography confirmed BAV | 0
dilatation of the ascending aorta 5.5 cm | 0
aortic dissection not discovered | 0
chronic pancreatitis | 0
recurrent exacerbations | 0
alcohol overuse | 0
type C chronic viral hepatitis | 0
hyperlipidemia | 0
offered cardiothoracic surgery | 0
refused surgery | 0
pharmacological treatment | 0
β-blocker | 0
angiotensin-converting enzyme inhibitor | 0
diuretic | 0
atorvastatin | 0
acetylsalicylic acid | 0
blood pressure control unknown | 0
cerebrovascular event | -8760
aphasia | -8760
hospitalization in Department of Neurology | -8760
echocardiography repeated | -8760
ultrasonography of cervical arteries | -8760
calcified cervical arteries | -8760
admitted to emergency room | -2160
abrupt onset of chest pain | -2160
chest pain persisted for 3 hours | -2160
severe retrosternal pain | -2160
pain radiated to left upper limb | -2160
loud systolic murmur | -2160
blood pressure 163/98 mm Hg right arm | -2160
blood pressure 135/93 mm Hg left arm | -2160
heart rate 65 beats per minute | -2160
ECG sinus rhythm 72/min | -2160
LVH features | -2160
negative T waves in II, III, aVF | -2160
negative T waves in V3–V6 | -2160
new findings in ECG | -2160
troponin I level 0.34 ng/ml | -2160
medical history BAV | -2160
medical history TAA | -2160
medical history arterial hypertension | -2160
coronary angiography 3 years prior | -2160
acute aortic dissection suspected | -2160
bedside transthoracic echocardiography | -2160
dissection flap in ascending aorta | -2160
computed tomography confirmed | -2160
ascending aorta dilatation 6.3 cm | -2160
aortic dissection | -2160
intimal tear 2.5 cm above aortic valve | -2160
dissection flap extended from right coronary artery ostium to aortic arch | -2160
right subclavian artery aberrant | -2160
right common carotid artery involved | -2160
left subclavian artery proximal segment involved | -2160
pharmacological treatment administered | -2160
referred for surgery | -2160
Bentall procedure performed | 0
total aortic root replacement | 0
St Jude Medical 29 mm conduit | 0
re-implantation of coronary arteries | 0
distal ascending aorta replaced with Datascope 22 mm prosthesis | 0
postoperative course typical | 24
conscious | 24
respiratory sufficient | 24
circulation supported with dobutamine | 24
LVEF 50% | 24
extubated on 1st postoperative day | 24
stable condition for 2 days | 24
postoperative day 4 | 96
excited and restless | 96
fever 39°C | 96
postoperative day 6 | 144
symptoms of septic shock | 144
multiorgan failure | 144
mediastinum drained | 144
empiric antibiotic therapy | 144
intensive care treatment | 144
died on 8th postoperative day | 192
cardiopulmonary insufficiency | 192
