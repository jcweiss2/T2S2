45 years old | 0
female | 0
admitted to the hospital | 0
shortness of breath | -48
malaise | -1344
lethargy | -1344
slow speech | -1344
edema of the face and extremities | -1344
progressive weight gain | -1344
no history of medical illness | 0
no drug history | 0
temperature 36°C | 0
blood pressure 90/52 mmHg | 0
heart rate 74 beats/min | 0
obese | 0
hypothermic | 0
pulsus paradoxus | 0
facial edema | 0
coarse hair | 0
dry skin | 0
engorged jugular vein | 0
mild pallor | 0
non-pitting edema of the extremities | 0
oxygen saturation 84% | 0
cardiac apical impulse not visible | 0
apex beat not felt | 0
heart sounds soft and distant | 0
bilateral basal rales | 0
mild hepatomegaly | 0
delayed relaxation of deep reflexes | 0
cardiomegaly | 0
globular enlargement of the cardiac silhouette | 0
pericardial effusion | 0
electrical alternans | 0
low voltage pattern | 0
right ventricular diastolic collapse | 0
pericardiocentesis | 1
pericardial fluid tapping | 1
450 ml pericardial fluid tapped | 1
improvement in cardiopulmonary status | 2
reduction of tachycardia and tachypnea | 2
oxygen saturation increased to 94% | 2
reduction of cardiomegaly | 2
minimal pericardial effusion | 2
no evidence of tamponade | 2
primary hypothyroidism | 0
high TSH | 0
low T3 and T4 levels | 0
thyroxine 100 μg daily | 2
thyroxine increased to 200 μg daily | 4
discharged | 336
follow-up echocardiogram | 2160
near total resolution of pericardial effusion | 2160
resolution of symptoms and signs | 2160
Hemoglobin 11.5 g% | 0
erythrocyte sedimentation rate 24 | 0
total leukocyte count 9850 mm3 | 0
platelet count 2.1 lac | 0
blood urea level 24 mg% | 0
serum creatinine level 1.1 mg% | 0
liver function test within normal limits | 0
serum TSH 84 mU/ml | 0
T3 26.2 ng/dl | 0
T4 0.56 μg/dl | 0
lipid profile | 0
total cholesterol 317 mg/dl | 0
high-density lipoprotein cholesterol 52 mg/dl | 0
triglyceride 214 mg/dl | 0
serum sodium 136 mEq/l | 0
serum potassium 4.2 mEq/l | 0
HIV negative | 0
HbSAg negative | 0
pericardial fluid analysis | 1
golden yellow pericardial fluid | 1
lymphocytes 8-10/mm3 | 1
proteins 4.7 g% | 1
sugar 80 mg% | 1
cholesterol 192 mg% | 1
no organisms grown on culture | 1