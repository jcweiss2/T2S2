45 years old | 0
female | 0
admitted to the hospital | 0
intermittent pain abdomen | -72
loss of appetite | -168
mild breathlessness | -72
no history of jaundice | 0
no history of hematemesis | 0
no history of malena | 0
no history of nausea and vomiting | 0
no history of chest pain | 0
no history of systemic medical disease | 0
history of previous exposure to general anesthesia | -10080
delayed emergence from anesthesia | -10080
heart rate 86/min | 0
occasional missed beats | 0
blood pressure 118/72 mmHg | 0
decreased air entry over left lower zones | 0
abnormal ventricular complexes on ECG | 0
tenderness over left hypochondrium and epigastric region | 0
no associated organomegalies | 0
Mallampatti Score grade II | 0
cystic lesion with air and fluid level at left lower zones on chest X-ray | 0
hydatid cyst of liver and lower lobe of left lung | 0
cyst in close proximity to the heart | 0
tab albendazole 400 mg twice daily started | -336
incentive spirometry taught | -336
premedication with tab ranitidine 150 mg | -12
premedication with tab metoclopramide | -12
premedication with tab alprazolam 0.25 mg | -12
general anesthesia and double lumen tube intubation planned | 0
thoracic epidural analgesia planned | 0
monitors attached for ECG, NIBP, ETCO2, and SpO2 | 0
IV access secured | 0
inj hydrocortisone 100 mg IV injected | 0
inj chlorpheniramine 25 mg IV injected | 0
inj adrenaline and inj theophylline kept ready | 0
epidural catheter inserted | 0
test dose of 3 mL of 2% lignocaine with 15 μg adrenaline injected | 0
8 mL of 0.75% ropivacaine injected into epidural space | 0
inj midazolam 1 mg IV administered | 0
inj glycopyrollate 0.2 mg IV administered | 0
inj fentanyl 50 μg IV administered | 0
induction of anesthesia with inj thiopentone sodium 250 mg | 0
complete muscle relaxation with inj suxamethonium 100 mg | 0
trachea intubated with 35 Fr left-sided double lumen tube | 0
bilateral equal air entry checked | 0
ventilation for each lung checked individually | 0
position of double lumen tube checked and confirmed by fiberoptic bronchoscopy | 0
anesthesia maintained with O2, N2O, and isoflurane | 0
muscle relaxation maintained with inj vecuronium bromide | 0
thoracoscopy done in right lateral decubitus position | 0
clamping bronchial lumen and ventilating only the right lung | 0
surgical procedure stopped and both lungs ventilated for 5 min every 30 min | 0
bradyarrhythmias observed on ECG monitor | 40
surgery stopped | 40
bradyarrhythmias subsided spontaneously | 40
inj lignocaine 60 mg given stat IV | 80
inj amiodarone 150 mg administered as bolus | 85
inj amiodarone infusion started | 85
surgical procedure accomplished uneventfully | 120
drainage and excision of lung cyst | 120
patient made supine | 120
laparoscopic drainage and excision of liver cyst | 120
ventilation of both lungs carried out simultaneously | 120
continuous monitoring of HR, ECG, NIBP, SpO2, and ETCO2 | 0
intermittent ABG done | 0
fluid intake and urine output remained within normal limits | 0
residual neuromuscular blockade reversed with inj neostigmine 2.5 mg and inj glycopyrrolate 0.05 mg | 240
trachea extubated | 240
patient shifted to ICU | 240
pain relief managed by epidural top-up of 8 mL of 0.25% ropivacaine | 240
postoperative ECG and echocardiography carried out | 288
patient shifted to surgical ICU | 288
recovery uneventful | 288