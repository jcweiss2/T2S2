46 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
arterial hypertension | -10080 | 0 | Factual
obesity | -10080 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
fever | -336 | 0 | Factual
hypotension | -336 | 0 | Factual
asthenia | -336 | 0 | Factual
cardiological examination | -672 | -672 | Factual
electrocardiogram (ECG) | -672 | -672 | Factual
transthoracic echocardiography (TTE) | -672 | -672 | Factual
COVID-19 infection | -336 | -336 | Factual
rhinitis | -336 | -336 | Factual
mild cough | -336 | -336 | Factual
alert | 0 | 0 | Factual
oriented | 0 | 0 | Factual
cooperative | 0 | 0 | Factual
asthenic | 0 | 0 | Factual
blood pressure (BP) 85/55 mmHg | 0 | 0 | Factual
heart rate (HR) 120 bpm | 0 | 0 | Factual
arterial oxygen saturation 85% | 0 | 0 | Factual
fever 38.3 C° | 0 | 0 | Factual
femoral central venous catheter (CVC) | 0 | 0 | Factual
sinus tachycardia | 0 | 0 | Factual
diffuse low voltages | 0 | 0 | Factual
absence of significant repolarization abnormalities | 0 | 0 | Factual
neutrophilic leukocytosis | 0 | 0 | Factual
C-reactive protein (CRP) elevation | 0 | 0 | Factual
Procalcitonin elevation | 0 | 0 | Factual
high sensitivity Troponin (hs-Tn) elevation | 0 | 0 | Factual
brain natriuretic peptide (BNP) elevation | 0 | 0 | Factual
creatinine elevation | 0 | 0 | Factual
transaminases elevation | 0 | 0 | Factual
total bilirubin elevation | 0 | 0 | Factual
reverse transcription-polymerase chain reaction (RT-PCR) nasopharyngeal swab negative | 0 | 0 | Factual
COVID-19 IgM antibody test positive | 0 | 0 | Factual
normal left ventricular (LV) cavitary dimensions | 0 | 0 | Factual
diffuse LV parietal thickening | 0 | 0 | Factual
increased myocardial echogenicity | 0 | 0 | Factual
severely reduced LV global systolic function | 0 | 0 | Factual
ejection fraction (EF) 26% | 0 | 0 | Factual
dP/dT ratio 672 mmHg/sec | 0 | 0 | Factual
indexed stroke volume (SVi) 11 ml/m2 | 0 | 0 | Factual
cardiac index (CI) 1.3 l/min/m2 | 0 | 0 | Factual
grade II LV diastolic dysfunction | 0 | 0 | Factual
normal cavitary dimensions | 0 | 0 | Factual
reduced global right ventricular (RV) systolic function | 0 | 0 | Factual
basal end-diastolic diameter (EDD) 37 mm | 0 | 0 | Factual
mean diameter 28 mm | 0 | 0 | Factual
TAPSE 14 mm | 0 | 0 | Factual
tricuspid S-wave velocity at tissue doppler imaging (TDI) 7.3 cm/sec | 0 | 0 | Factual
inferior vena cava (IVC) dilated | 0 | 0 | Factual
right ventricular systolic pressure (RVSP) 41 mmHg | 0 | 0 | Factual
absence of hemodynamically significant valvulopathy | 0 | 0 | Factual
pericardial effusion | 0 | 0 | Factual
blood cultures | 0 | 0 | Factual
broad-spectrum antibiotic therapy | 0 | 24 | Factual
INN-daptomycin | 0 | 24 | Factual
piperacillin/tazobactam | 0 | 24 | Factual
crystalloid hydration | 0 | 24 | Factual
nasal cannula ventilatory therapy | 0 | 24 | Factual
norepinephrine | 0 | 12 | Factual
poor hemodynamic response | 12 | 12 | Factual
levosimendan | 12 | 36 | Factual
bolus administration avoided | 12 | 12 | Factual
continuous maintenance intravenous infusion | 12 | 36 | Factual
BP increased to 100/60 mmHg | 12 | 12 | Factual
HR decreased to 110 bpm | 12 | 12 | Factual
further hemodynamic improvement | 24 | 24 | Factual
BP 125/70 mmHg | 24 | 24 | Factual
HR 95 bpm | 24 | 24 | Factual
diuresis 1800 ml | 12 | 24 | Factual
control TTE | 12 | 24 | Factual
improvement of systolic performance indices | 12 | 24 | Factual
LV EF 66% | 24 | 24 | Factual
dP/dT ratio 1275 mmHg/sec | 24 | 24 | Factual
TAPSE 23 mm | 24 | 24 | Factual
tricuspid S-wave velocity at TDI 11.2 cm/sec | 24 | 24 | Factual
SVi 27 ml/m2 | 24 | 24 | Factual
CI 2.5 l/min/m2 | 24 | 24 | Factual
LV diastolic function improvement | 24 | 24 | Factual
IVC diameter 18 mm | 24 | 24 | Factual
IVC collapse 100% | 24 | 24 | Factual
RVSP 28 mmHg | 24 | 24 | Factual
cardiac magnetic resonance imaging (CMR) | 24 | 24 | Factual
endomyocardial biopsy | 48 | 48 | Factual
lymphocytic myocarditis | 48 | 48 | Factual
coronary arteriography | 48 | 48 | Factual
normal coronary circulation | 48 | 48 | Factual
discharged | 504 | 504 | Factual
excellent hemodynamic compensation | 504 | 504 | Factual
normal laboratory findings | 504 | 504 | Factual
normal electrocardiographic findings | 504 | 504 | Factual
normal echocardiographic findings | 504 | 504 | Factual
TTE at 1 month | 744 | 744 | Factual
TTE at 3 months | 2232 | 2232 | Factual
normal LV and RV systolic and diastolic function | 744 | 2232 | Factual