43 years old | 0
    woman | 0
    Chron’s disease | 0
    infliximab | 0
    azathioprine | 0
    fever | 0
    thoracic pain | 0
    elevated inflammatory parameters | 0
    nasopharyngeal swab for SARS-CoV-2 negative | 0
    bilateral community-acquired pneumonia | 0
    chest radiograph | 0
    discharged | 0
    cefuroxime | 0
    same symptoms | -72
    organ dysfunction negative | -72
    Streptococcus pneumoniae urinary antigen test negative | -72
    Legionella pneumophila urinary antigen test negative | -72
    nasopharyngeal swab for SARS-CoV-2 negative | -72
    blood samples collected | -72
    sputum samples collected | -72
    admitted to the hospital | -72
    piperacillin-tazobactam | -72
    acute rapidly progressive respiratory failure | -48
    admitted to the intensive care unit | -48
    invasive mechanical ventilation | -48
    normal cardiac function | -48
    no signs of pulmonary embolism | -48
    significant consolidation of both lungs | -48
    suspicion of organizing pneumonia | -48
    vancomycin | -48
    methylprednisolone | -48
    mixed acidaemia | -24
    refractory hypoxemia | -24
    extracorporeal membrane oxygenation | -24
    transferred to Infectious Diseases ICU | -24
    blood samples negative | -24
    sputum samples negative | -24
    blood collected | 0
    bronchial lavage collected | 0
    bronchoalveolar lavage collected | 0
    urine collected | 0
    etiological investigation | 0
    meropenem | 0
    vancomycin | 0
    liposomal amphotericin | 0
    cardiovascular failure | 24
    hypoperfusion | 24
    hypotension | 24
    anasarca | 24
    hyperlacticaemia | 24
    anuric acute kidney injury | 24
    liver failure | 24
    worsening pancytopenia | 24
    blood transfusions | 24
    vasopressor therapy | 24
    continuous renal replacement therapy | 24
    sodium bicarbonate | 24
    albumin supplementation | 24
    plasmapheresis | 24
    yeast growing in blood bottle | 72
    Saprochaete clavata identified | 96
    Saprochaete clavata isolated again | 96
    died | 120
    Legionella pneumophila PCR positive | 120
    <|eot_id|>