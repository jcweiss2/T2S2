18 years old | 0
male | 0
history of methicillin-resistant Staphylococcus aureus (MRSA) impetigo | -8760
right tibia fracture | -8760
intramedullary fixation (IMN) | -8760
interlocking screws removed | -8760
skin irritation | -8760
pain | -8760
redness and swelling at the surgical site | -730
stitch abscess | -730
MRSA | -730
oral antibiotic treatment | -730
fever | -672
right groin pain | -672
viral infection | -672
systemic fever | -644
myalgia | -644
difficult and painful ambulation | -644
right forearm cellulitis | -644
right sudden onset uveitis | -644
systemic rash | -644
right hip lymphadenopathy | -644
increased CRP | -644
increased WBC count | -644
elevated hepatic enzymes | -644
elevated lactic dehydrogenase (LDH) | -644
elevated creatine phosphokinase (CPK) levels | -644
intravenous (IV) antibiotics | -644
hemodynamic deterioration | -576
fulminant MRSA sepsis | -576
ultrasound-guided drainage | -576
further enlargement of the abscesses diameter | -552
persistent fever | -552
CRP level of 36 mg/dL | -552
WBC count of 20,000 | -552
surgical intervention | -528
combined approach of Smith-Peterson and modified Stoppa | -528
general anaesthesia with muscle relaxant | -528
supine position with a bump and the knee to flex the thigh | -528
contralateral pelvic elevation to 20 degrees | -528
Stoppa approach | -528
medial side of the abscess | -528
lateral sides of the abscess | -528
anterior approach of the hip (Smith-Peterson) | -528
rectus abdominis muscles split vertically | -528
rectus and the femoral neurovascular structures retracted | -528
iliopectineal fascia released | -528
iliopsoas visualized and elevated | -528
obturator neurovascular bundle exposed and protected | -528
quadrilateral surface and posterior column dissected | -528
obturator internus muscle and adductor brevis muscle debridement and lavage | -528
Smith-Peterson approach | -528
rectus femoris detached from its both origins | -528
rectus femoris and iliopsoas retracted medially | -528
gluteus medius retracted laterally | -528
hip capsule exposed | -528
abscess drainage and debridement | -528
almost complete recovery | -504
normal ambulation without any pain or functional limitations | -504
return to daily activities | -504