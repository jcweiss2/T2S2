74 years old | 0
female | 0
admitted to the hospital | 0
low-grade fever | -48
cough | -48
shortness of breath | -48
elective right total knee replacement | -168
pain in the right knee | -168
redness in the right knee | -168
swelling in the right knee | -168
essential hypertension | -168
obesity | -168
myasthenia gravis | -168
osteoarthritis | -168
body temperature of 37.3°C | 0
blood pressure of 121/82 | 0
pulse of 87 beats per minute | 0
respiratory rate of 16 breaths per minute | 0
oxygen saturation of 87% | 0
bilateral rhonchi with rales | 0
patchy air space opacity in the right upper lobe suspicious for pneumonia | 0
negative for influenza A and B | 0
nasopharyngeal swab specimen | 0
sent to the state laboratory for detection of SARS-CoV-2 | 0
admitted to the airborne-isolation unit | 0
broad-spectrum antibiotics with cefepime and levofloxacin | 0
2 L of supplemental oxygen | 0
mild diarrhea | 72
generalized weakness | 72
fatigue | 72
1 g/kg intravenous immunoglobulin | 72
mild MG exacerbation | 72
pending MG crises | 72
arterial blood gases | 72
complete blood count | 72
basic metabolic profile studies | 72
mild absolute lymphopenia | 72
anemia | 72
pH of 7.46 | 72
pCO2 of 44.6 mmHg | 72
pO2 of 94.7 mmHg | 72
bicarbonate of 31.4 mmol/L | 72
positive for SARS-CoV-2 | 96
oral hydroxychloroquine 400 mg once | 96
azithromycin 500 mg once a day intravenously | 96
zinc sulfate 220 mg 3 times a day | 96
oral vitamin C 1 g twice a day | 96
broad-spectrum antibiotics discontinued | 96
SOB worsened rapidly | 120
oxygen requirements went up to 15 L | 120
drowsy | 120
in moderate distress | 120
unable to protect the airways | 120
blood pressure of 78/56 mmHg | 120
heart rate of 112 beats per minute | 120
temperature 38°C | 120
respiratory rate of 28 breaths per minute | 120
bilateral alveolar infiltrates due to pneumonia and interstitial edema | 120
ARDS | 120
intubated on an emergent basis | 120
pressure-regulated volume-controlled mechanical ventilation | 120
norepinephrine 0.02 mcg/kg/min | 120
septic shock | 120
colchicine 0.6 mg twice a day | 120
elevated interleukin-6 levels | 120
high-dose vitamin C 11 g per 24 h | 168
clinical condition started to improve slowly | 168
norepinephrine support was stopped | 168
CXR showed significant improvement of the pneumonia and interstitial edema | 168
spontaneous breathing trial with CPAP/PS | 168
positive end-expiratory pressure (PEEP) of 7 mmHg | 168
PS above PEEP of 10 mmHg | 168
fraction of inspired oxygen of 40% | 168
ABGs revealed a pH of 7.49 mmHg | 168
pCO2 of 40.2 mmHg | 168
pO2 of 77.1 mmHg | 168
bicarbonate of 30.2 mmol/L | 168
extubated to 4 L of oxygen with a nasal cannula | 168
oxygen saturation of 92% | 168
CXR revealed almost complete resolution of the infiltrates | 168
discharged from the hospital | 168
still positive by RT-PCR for SARS-CoV-2 | 168
14 days of quarantine | 168