43 years old | 0
    Hispanic | 0
    female | 0
    no significant medical history | 0
    right upper quadrant abdominal pain | -168
    fever | -168
    nausea | -168
    vomiting | -168
    diarrhea | -168
    hypotensive | 0
    tachycardic | 0
    temperature of 38.0 °C | 0
    pulse of 138 beats per minute | 0
    respiratory rate of 18 per minute |5
    blood pressure of 90/54 mm Hg | 0
    pulse oximetry of 99% on room air | 0
    dry mucosal membranes | 0
    diffuse abdominal tenderness | 0
    transferred to intensive care unit | 0
    septic shock | 0
    white blood cell count of 5,620/µL | 0
    hemoglobin of 11.7 g/dL | 0
    sodium level of 130 mmol/L | 0
    potassium of 3.3 mmol/L | 0
    creatinine of 3.3 mg/dL | 0
    glomerular filtration rate of 15.26 mL/min | 0
    total bilirubin of 1.5 mg/dL | 0
    aspartate aminotransferase of 246 U/L | 0
    alanine aminotransferase of 185 U/L | 0
    alkaline phosphatase of 131 U/L | 0
    lipase of 35 U/L | 0
    lactic acid of 7.2 mmol/L | 0
    COVID-19 positive | 0
    no supplemental oxygen required | 0
    no specific treatment for COVID-19 | 0
    CT scan of abdomen | 0
    hypodense cystic structure in right liver lobe | 0
    follow-up ultrasound | 24
    9.9-cm mass in right lobe of liver | 24
    follow-up MRI scan of abdomen | 24
    heavily septated 13-cm hepatic abscess in posterior right hepatic lobe | 24
    fluid boluses | 0
    intravenous vancomycin | 0
    intravenous piperacillin/tazobactam | 0
    percutaneous drainage | 24
    1,110 mL of purulent fluid | 24
    CT scan for needle placement | 24
    small pneumoperitoneum | 24
    Streptococcus viridans culture | 24
    antibiotics switched to ampicillin/sulbactam | 24
    RUQ pain improved | 24
    discharge | 192
    antibiotic regimen changed to amoxicillin | 192
    left lower quadrant abdominal pain | 192
    repeat CT of abdomen | 192
    decreased size of liver lesion | 192
    pelvic abscess measuring 13.6 × 5 cm | 192
    unchanged pneumoperitoneum | 192
    perforated sigmoid diverticulum | 192
    CT-guided percutaneous drainage | 192
    mixed gram-positive and gram-negative flora culture | 192
    Candida albicans culture | 192
    discharged with drains | 192
    20-day course of amoxicillin | 192
    fluconazole | 192
    returned to hospital for drain removal | 240
    improvement of LLQ pain | 240
    no jaundice | 0
    no bacteremia | 0
    no venous thromboembolism | 0
    no history of diverticulitis | 0
    single hepatic abscess | 24
    no multiple hepatic abscesses | 24
    no portal vein thrombosis | 24
    no acute diverticulitis initially | 0
    no personal history of diverticulitis | 0
    no bacteremia | 0
    no Candida albicans in hepatic abscess | 24
    mixed flora in pelvic abscess | 192
    received antibiotics prior to pelvic aspiration | 192
    no colonoscopy reported | 0
    no weight loss | 0
    no jaundice | 0
    no acute cholangitis | 0
    no Streptococcus anginosus | 0
    no portal vein thrombosis | 0
    no venous thromboembolism | 0
    no surgical drainage required | 24
    no multiple abscesses | 24
    no loculated abscess | 24
    no complications from drainage | 24
    no recurrence of hepatic abscess | 240
    no mortality | 240
    no diabetes mellitus | 0
    no hypertension | 0
    no atrial fibrillation | 0
    no preexisting conditions | 0
    Hispanic female | 0
    younger than average patient | 0
    no initial LLQ pain | 0
    no initial pelvic abscess | 0
    no initial perforated diverticulitis | 0
    no bacteremia | 0
    no jaundice | 0
    no weight loss | 0
    no Streptococcus intermedius in pelvic abscess | 192
    no Candida albicans in hepatic abscess | 24
    no acute diverticulitis at presentation | 0
    no initial findings of diverticulitis | 0
    no colonoscopy reported | 0
    no specific treatment for COVID-19 | 0
    no oxygen required | 0
    no jaundice | 0
    no venous thromboembolism | 0
    no portal vein thrombosis | 0
    no bacteremia | 0
    no complications from antibiotics | 192
    no recurrence after discharge | 240
    no mortality | 240
    no diabetes mellitus | 0
    no hypertension | 0
    no atrial fibrillation | 0
    no preexisting comorbidities | 0
    no history of diverticulitis | 0
    no initial pelvic abscess | 0
    no initial perforated diverticulum | 0
    no bacteremia | 0
    no jaundice | 0
    no weight loss | 0
    no venous thromboembolism | 0
    no portal vein thrombosis | 0
    no surgical drainage required | 24
    no complications from drainage | 24
    no recurrence of abscess | 240
    no mortality | 240
    no diabetes | 0
    no hypertension | 0
    no atrial fibrillation | 0
    no comorbidities | 0
    no history of diverticulitis | 0
    no bacteremia | 0
    no jaundice | 0
    no weight loss | 0
    no venous thromboembolism | 0
    no portal vein thrombosis | 0
    no surgical intervention | 24
    no complications post-discharge | 240
    no mortality | 240