34 years old | 0
female | 0
admitted to the hospital | 0
epigastric pain | -48
dyspnea | -48
diaphoresis | -48
nausea | -48
vomiting | -48
weight loss | -4320
left flank pain | 0
mild abdominal tenderness | 0
ascites | 0
palpable painful mass in left upper abdomen | 0
hypotension | 0
blood pressure 90/50 mmHg | 0
heart rate 75 bpm | 0
moist rales | 0
ST-segment elevation in inferior limb leads | 0
dopamine infusion | 0
bolus saline replacement | 0
emergency coronary angiogram | 0
high thrombus burden in distal right coronary artery | 0
cardiac arrest during angiography | 0
ventricular fibrillation | 0
defibrillation with 360 J | 0
cardiopulmonary resuscitation | 0
asystole | 0
adrenaline administration | 0
sinus rhythm achieved | 0
predilatation with balloon | 0
tirofiban infusion | 0
no reflow after stent deployment | 0
drug-eluting stent implanted | 0
TIMI Grade 3 flow achieved | 48
regional wall motion abnormalities | 24
hypokinesia of inferior, posterior, and septal segments | 24
ejection fraction 40% | 24
right atrial mass adhering to inferior vena cava | 24
no paradoxical embolism | 24
intracardiac mass thought to be thrombus | 72
anticoagulation with rivaroxaban | 72
dual antiplatelet therapy | 72
normal haematological parameters | 72
normal biochemical parameters | 72
normal lipid profile | 72
normal tumour markers | 72
normal connective tissue markers | 72
normal thrombophilia panel | 72
cancer antigen 125 elevated | 72
possible cancer-induced thrombosis | 168
CT scan of abdomen and pelvis | 168
11.3 cm enhanced necrotic mass in left adrenal gland | 168
tumour thrombus in inferior vena cava | 168
normal twenty-four-hour urine analyses | 312
image-guided tissue sampling | 408
histopathological confirmation of PHEOs | 408
metastatic foci on PET and CT | 408
persistence of thrombus despite anticoagulation | 408
diagnosis of malignant PHEOs | 480
treatment with 177Lu-DOTATATE PRRT initiated | 480
discharged | 720
readmitted with ascites and dyspnea | 2160
septic shock | 2160
death due to nosocomial infections | 2160
