40 years old | 0 | 0 
African-American | 0 | 0 
female | 0 | 0 
admitted to the emergency department | 0 | 0 
history of chronic eczema | -720 | 0 
previous alcohol abuse | -720 | 0 
gout | -720 | 0 
hypothyroidism | -720 | 0 
cutaneous eruption | -336 | 0 
desquamation of the hands | -336 | 0 
desquamation of the feet | -336 | 0 
desquamation of the perioral skin | -336 | 0 
desquamation of the perineal skin | -336 | 0 
pain | -336 | 0 
swelling | -336 | 0 
hair loss | -336 | 0 
increasing weakness | -576 | 0 
fatigue | -576 | 0 
intermittent diarrhea | -576 | 0 
unintentional weight loss | -576 | 0 
70 pounds weight loss | -576 | 0 
psychosocial habits | -720 | 0 
1 to 2 glasses of wine a day | -720 | 0 
smoking | -720 | 0 
no significant family history | 0 | 0 
not on any medications | 0 | 0 
dermatologic examination | 0 | 0 
erythematous desquamative patches | 0 | 0 
erosions | 0 | 0 
crusted lesions | 0 | 0 
diffuse nonscarring alopecia | 0 | 0 
scaling patches on the vermillion lips | 0 | 0 
punch biopsy of the left medial thigh | 0 | 0 
psoriasiform epidermal spongiosis | 0 | 0 
superficial perivascular lymphohistiocytic infiltrate | 0 | 0 
diffuse hypogranulosis | 0 | 0 
broad overlying parakeratosis | 0 | 0 
ballooning degeneration of the spinous layer | 0 | 0 
methicillin-resistant Staphylococcus aureus sepsis | 0 | 48 
Escherichia coli sepsis | 0 | 48 
pneumonia | 0 | 48 
admitted to the intensive care unit | 0 | 48 
ventilator respiratory support | 0 | 48 
systemic antibiotics | 0 | 48 
laboratory and imaging studies | 0 | 48 
necrolytic acral erythema ruled out | 0 | 48 
pellagra ruled out | 0 | 48 
biotin deficiency ruled out | 0 | 48 
low zinc levels | 0 | 0 
antitransglutaminase antibodies positive | 0 | 0 
antiendomysium antibodies positive | 0 | 0 
diagnosis of celiac disease | 0 | 0 
zinc deficiency | 0 | 0 
history of excessive alcohol intake | -720 | 0 
chronic low zinc levels | -720 | 0 
deficiency dermatitis | -336 | 0 
distal duodenal biopsy | 0 | 48 
focal villi blunting | 0 | 48 
Brunner's gland hyperplasia | 0 | 48 
treated with a gluten-free diet | 48 | 336 
treated with zinc sulfate | 48 | 336 
resolution of gastrointestinal symptoms | 336 | 336 
resolution of cutaneous symptoms | 336 | 336