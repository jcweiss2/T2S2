10 years old | 0
male | 0
unrelated healthy parents | 0
first and only son | 0
refractory epilepsy | -120 months
insomnia | -120 months
born by cesarean section | -120 months
38 weeks gestation | -120 months
no intrauterine growth restriction | -120 months
weight 3200g | -120 months
length 52 cm | -120 months
APGAR score 9-9 | -120 months
perioral cyanosis | -120 months
transferred to intensive care unit | -120 months
probable diagnosis of neonatal sepsis | -120 months
echocardiogram reported patent ductus arteriosus | -120 months
patent ductus arteriosus closed spontaneously | -120 months
newborn screening normal | -120 months
discharged after 11 days | -119 months
recurrent pulmonary infections | -120 months
multiple hospital admissions | -120 months
severe gastroesophageal reflux | -120 months
breast milk intolerance | -120 months
Nissen fundoplication | -114 months
gastrostomy | -114 months
atonic seizures | -113 months
childhood spasms | -113 months
valproic acid | -113 months
Fanconi syndrome | -112 months
oxcarbazepine | -112 months
severe hyponatremia | -112 months
phenobarbital | -112 months
phenytoin | -112 months
atomoxetine | -112 months
aripiprazole | -112 months
quetiapine fumarate | -112 months
haloperidol | -112 months
sertraline | -112 months
pregabalin | -112 months
olanzapine | -112 months
topiramate | -112 months
levetiracetam | -112 months
mirtazapine | -112 months
ethyl loflazepate | -112 months
lacosamide | 0
clobazam | 0
brivaracetam | 0
acetazolamide | 0
hypokalemia | 0
potassium supplementation | 0
weight below third percentile | -120 months
height below third percentile | -120 months
head circumference below third percentile | -120 months
subclinical hypothyroidism | -108 months
selective immunodeficiency | -108 months
nephrocalcinosis | -108 months
microcephaly | -120 months
elongated eyelid fissures | -120 months
eversion of outer third of lower eyelid | -120 months
arched and broad eyebrows | -120 months
depressed nasal tip | -120 months
short columella | -120 months
small and spaced teeth | -120 months
micrognathia | -120 months
large cup-shaped ears | -120 months
low implantation | -120 months
bilateral retroauricular pits | -120 months
polydactyly of right hand | -120 months
polydactyly of left foot | -120 months
surgically treated | -114 months
bilateral palmar aberrant folds | -120 months
sacral dimple | -120 months
Kabuki syndrome suspected | -12 months
KMT2D gene sequencing | -12 months
exome sequencing | 0
homozygous variant in OTUD6B gene | 0
c.433C>T variant | 0
pathogenic variant | 0
weight 24 kg | 0
height 1.24 m | 0
delayed overall development | 0
head support delayed | 0
sitting with support delayed | 0
no gait development | 0
only emits sounds | 0
obeys simple commands | 0
solid foods orally | 0
liquids by gastrostomy | 0
levothyroxine | 0
gamma globulin | 0
insulin resistance | 0
allergic colitis | 0