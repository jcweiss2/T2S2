32 years old | 0
    female | 0
    dental abscess on left inferior 3rd molar | -672
    treated with oral amoxicillin/clavulanate | -672
    odynophagia | -144
    painful left submandibular edema | -144
    severe upper airway respiratory distress | 0
    trismus | 0
    extension of inflammatory signs to anterior cervical region | 0
    leukocytosis | 0
    elevated C-reactive protein | 0
    diffuse thickening of soft tissues with phlegmon and emphysema | 0
    abscess extension to submandibular, parapharyngeal, and retrosternal spaces | 0
    bulging of the walls of the airway at the base of the tongue | 0
    left internal jugular vein thrombosis | 0
    transferred to tertiary referral centre | 0
    fibreoptic nasotracheal intubation | 0
    surgical drainage of abscesses | 0
    admitted to Intensive Care Unit | 0
    daily bedside drainage of submandibular region | 0
    intravenous corticosteroids | 0
    empiric antibiotic therapy with ceftriaxone and metronidazole | 0
    extension of vein thrombosis to brachiocephalic vein | 48
    intravenous non-fractioned heparin initiated | 48
    Gram staining showed polymicrobial flora | 0
    abscess cultures grew Streptococcus anginosus | 0
    blood cultures sterile | 0
    HIV negative | 0
    normal serum immunoglobulins | 0
    clinical and imaging improvement | 192
    successful extubation | 192
    transferred to infirmary | 192
    persistence of left internal jugular vein thrombosis | 192
    defervescence | 192
    neck tenderness resolution | 192
    completed 24 days of ceftriaxone and metronidazole | 576
    discharged | 600
    anticoagulation with enoxaparin | 600
    
    