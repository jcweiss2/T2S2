26 years old | 0
male | 0
admitted to the hospital | 0
weakness of all four limbs | -24
addicted to multiple medicines | -6720
tramadol | -6720
diclofenac | -6720
pheniramine | -6720
dexamethasone | -6720
heparin | -6720
bronchial asthma | -8760
on and off steroids | -8760
conscious | 0
oriented | 0
hemodynamically stable | 0
heart rate of 112 beats/min | 0
non-invasive blood pressure of 130/80 mmHg | 0
respiratory rate of 24/min | 0
temperature of 99°F | 0
no pallor | 0
no signs of clubbing | 0
no lymphadenopathy | 0
oral thrush | 0
chest examination was grossly normal | 0
cardiovascular system examination was grossly normal | 0
per abdomen examination was grossly normal | 0
power was grade 3/5 in upper limbs | 0
power was grade 1/5 in lower limbs | 0
generalized areflexia | 0
planters were bilateral flexors | 0
sensory examination was normal | 0
arterial blood gas (ABG) at admission showed a normal pH | 0
hyperkalemia (K+ = 6.01) | 0
tachypnoeic | 1
respiratory rate of 36-40/min | 1
non-invasive ventilation | 1
heart rate went up to 130 beats/min | 1
pulses got feeble | 1
blood pressure dropped down to 100/56 mmHg | 1
invasive lines were put in | 1
central venous cannulation | 1
arterial line | 1
central venous pressure was 6 cm H2O | 1
mean arterial pressure (MAP) was 55 mmHg | 1
resuscitated with a fluid bolus of 1 litre normal saline | 1
blood pressure improved with MAP going up to 64 mmHg | 2
given 500 mL of normal saline | 2
started on normal saline 100 mL/h infusion | 2
urine output was >0.5 mL/kg | 2
chest X-ray showed a patch of consolidation | 2
echocardiography showed global hypokinesia | 2
severe left ventricular dysfunction | 2
ejection fraction of 30% | 2
repeat ABG after 6 h showed metabolic acidosis | 6
lactic acidosis | 6
hyperkalemia (pH = 7.257, pCO2 = 27.2, pO2 = 98.6, HCO3− = 13.8, Lactate = 7.1, K+ = 7.0) | 6
anti-hyperkalemia treatment was started | 6
calcium gluconate | 6
dextrose-insulin | 6
salbutamol nebulization | 6
slow low-efficiency dialysis (SLED) of 8 h | 6
episode of pulseless ventricular tachycardia | 6.33
defibrillated | 6.33
cardiopulmonary resuscitation (CPR) | 6.33
anti-hyperkalemia regimen was repeated | 6.33
urgent serum K+ levels done at the time of event were 9.1 mEq/L | 6.33
revived with normal sinus rhythm | 6.73
intubated | 6.73
put on invasive ventilatory support | 6.73
started on inotropes | 6.73
started on vasopressors | 6.73
subsequent ABG done before the end of planned duration of SLED still showed persistent hyperkalemia | 14
planned to extend the ongoing SLED | 14
after another 4 h of extended SLED | 18
blood gas still showed raised potassium values | 18
SLED was further extended | 18
total duration of 20 h | 20
post dialysis | 20
lab serum K+ level of 7.6 mEq/L | 20
developed blisters all over the body | 24
coagulopathy | 24
thrombocytopenia | 24
started empirically on ceftriaxone | 0
shifted to meropenem | 24
teicoplanin | 24
ampicillin | 24
deteriorating clinical condition | 24
taken up for SLED again | 24
dialyzed for more than 32 h | 32
refractory hyperkalemia remained | 40
fludrocortisone in the dose of 100 μg/day was also added | 48
correlating thrombocytopenia and coagulopathy with heparin | 48
activated clotting time was monitored | 48
protamine sulphate was also given | 48
episode of upper gastrointestinal bleed | 72
went into asystole | 72
CPR was done | 72
could not be revived | 72
declared dead | 72
blood cultures obtained after 72 h showed methicilin-resistant staphylococci | 72