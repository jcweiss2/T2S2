24 years old | 0
female | 0
pregnant | 0
admitted to the hospital | 0
abdominal pain | -120
abdominal distension | -120
constipation | -120
increasing severity of pain | -120
no significant past medical history | 0
no significant past surgical history | 0
uneventful menstrual history | 0
uneventful antenatal history | 0
dehydrated | 0
hypotension | 0
tachycardia | 0
tachypnea | 0
asymmetrically distended abdomen | 0
tenderness all over abdomen | 0
empty rectum on digital examination | 0
foetal viability assessed | 0
no threatened preterm labour | 0
elevated white cell count | 0
normal urine analysis | 0
distended bowel loop on ultrasound | 0
moderate amount of free fluid in peritoneal cavity | 0
single viable foetus on ultrasound | 0
clinical diagnosis of intestinal obstruction | 0
abdominal X-ray performed | 0
dilated large bowel on X-ray | 0
abnormal gas pattern on X-ray | 0
coffee bean appearance on X-ray | 0
sigmoidoscopy performed | 0
twisted sigmoid colon on sigmoidoscopy | 0
failure to negotiate obstruction | 0
foetal distress | 0
deceleration in heart rate | 0
decision to perform caesarean section | 0
concomitant caesarean section | 0
exploration of abdomen for intestinal obstruction | 0
initial resuscitation | 0
taken to emergency theatre | 0
midline laparotomy | 0
enormously distended sigmoid loop | 0
ischemic and gangrenous changes | 0
no signs of perforation | 0
necrotic colon | 0
posterior displacement by pregnant uterus | 0
lower segment caesarean section | 0
preterm infant delivered | 0
male infant | 0
infant weighed 750g | 0
infant admitted to neonatal ICU | 0
infant on mechanical ventilation | 0
gangrenous sigmoid colon resected | 0
Hartmann’s procedure | 0
end colostomy fashioned | 0
closure of rectal stump | 0
post-operative course uneventful | 0
discharged home on 9th post-operative day | 216
infant discharged home after 10 weeks in neonatal ICU | 720
reversal of Hartmann’s | 4320
bowel continuity restored | 4320
colo-rectal anastomosis | 4320