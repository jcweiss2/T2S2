term appropriate for gestational age male baby | 0
born to a 29-year-old mother | 0
elective lower segment cesarean section | 0
mother had high-grade fever | -48
mother had severe multiple joint pains | -48
mother developed diffuse hyperpigmentation of body | -44
baby developed high-grade fever | 72
baby admitted in neonatal intensive care unit | 72
baby started on antibiotics | 72
fever decreased in intensity | 120
baby developed generalized edema | 144
baby developed tenderness | 144
baby developed paradoxical cry | 144
baby developed decreased urine output | 168
features of acute renal failure | 168
dialysis started | 168
platelet transfusions given | 168
dialysis continued for 2 days | 192
platelet transfusions given for 3 days | 216
baby was relatively better | 288
urine output improved | 288
baby was relatively active | 360
feed was reintroduced | 360
baby tolerated feeds well | 360
platelet count remained low | 360
baby referred to our center | 432
persistent symptoms | 432
paradoxical cry | 432
significant thrombocytopenia | 432
mild bleeding manifestations | 432
baby was lethargic and inactive | 432
oral mucosal bleeds | 432
evidence of mucositis | 432
no hepatosplenomegaly | 432
C-reactive protein elevated | 432
hemoglobin 11 g/dL | 432
total leukocyte count 28,000/mm3 | 432
lymphocytosis | 432
platelet count 18,000/mm3 | 432
normal prothrombin and activated partial thromboplastin time | 432
serum sodium 129 mmol/L | 432
serum potassium 4.9 mmol/L | 432
plasma urea 112 mg/dL | 432
serum creatinine 1.8 mg/dL | 432
serum glutamic pyruvic transaminase elevated | 432
serum glutamic oxaloacetic transaminase elevated | 432
blood culture reported sterile | 432
TORCH screen normal | 432
cerebrospinal fluid study normal | 432
platelet transfusion given | 432
plasma urea and serum creatinine normalized | 480
other laboratory parameters normalized | 504
magnetic resonance imaging done | 504
focal areas of bleeds in the basal ganglia and subcortical areas | 504
mother tested for chikungunya IgM and IgG | 504
mother's chikungunya IgM and IgG reported positive | 504
baby's serology reported negative | 504
diagnosis of congenital chikungunya made | 504
baby improved with supportive management | 504
irritability and paradoxical cry persisted | 504
baby discharged | 756
baby kept under follow-up | 756
fixed flexion deformity of the right thumb | 1296