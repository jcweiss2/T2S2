75 years old | 0
female | 0
hypertension | 0
diabetes mellitus type II | 0
chronic kidney disease (CKD stage II) | 0
obesity (BMI 38.4 kg/m2) | 0
hyperlipidemia | 0
admitted to the hospital | 0
right upper quadrant abdominal pain | -336
nausea | -336
vomiting | -336
afebrile | 0
stable vital signs | 0
epigastric tenderness | 0
white blood cell count of 22,200/μL | 0
serum lipase of 804 U/L | 0
amylase level of 484 U/L | 0
gallstone in gallbladder | 0
pancreatic necrosis | 0
non-occlusive splenic vein thrombosis | 0
intravenous fluid | 0
IV antibacterials | 0
analgesics | 0
bowel rest | 0
persistent leukocytosis | 24
inability to tolerate oral intake | 24
hypoxemic respiratory failure | 24
intubation | 24
mechanical ventilation | 24
repeat CT scan abdomen/pelvis | 48
large collection | 48
pancreatic necrosectomy | 72
abdominal washout | 72
wide drainage | 72
vasopressor requirements | 72
ventilator support | 72
post-operative day (POD) 10 | 240
repeat CT scan of abdomen/pelvis | 240
posterior wall gastric perforation | 240
gastric perforation repair | 240
primary repair of gastric perforation | 240
one week after gastric perforation repair | 336
febrile episode | 336
elevated WBC count | 336
second posterior wall gastric perforation | 336
primary repair of second gastric perforation | 336
abdominal washout | 336
pancreatic necrosectomy | 336
twenty-eight days later from index operation | 672
third posterior wall gastric perforation | 672
CMV inclusion bodies | 672
HIV status negative | 672
intravenous ganciclovir | 672
CMV IgM titer negative | 672
CMV IgG titer positive | 672
CMV PCR 3,860,104 IU/mL | 672
ganciclovir treatment | 672
leukocytosis trending down | 696
weaned off vasopressors | 696
CMV PCR titer decreased | 696
total parenteral nutrition (TPN) | 696
tracheostomy | 696
jejunostomy feeding tube placement | 696
ganciclovir discontinued | 688
abdominal wound dehiscence | 720
debridement | 720
negative pressure wound therapy | 720
skin grafting | 720
urine and bronchoalveolar lavage cultures positive for Candida albicans and Pseudomonas aeruginosa | 720
treated with antifungals and antibiotics | 720
discharged to a rehabilitation center | 840
discharged home | 1008
tracheostomy decannulated | 1008
started on regular diet | 1008
follow up CT scans | 1008
no evidence of leak | 1008
outpatient esophagogastroduodenoscopy (EGD) | 2160
no malignancy | 2160
no Helicobacter pylori | 2160
no CMV infection | 2160