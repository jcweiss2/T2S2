65 years old | 0
male | 0
chest pain | -24
chest pain radiating to left arm | -24
chest pain radiating to right arm | -24
anterolateral ischemia on ECG | -24
emergency department admission | 0
acute myocardial injury | -336
cardiac arrest | 0
ventricular fibrillation on ECG | 0
coronary angiography (90% stenosis of circumflex artery) | -336
percutaneous transluminal coronary angioplasty | -336
stent placement on left main coronary artery | -336
stent placement on left anterior descending coronary artery | -336
stent placement on left circumflex coronary artery | -336
dual antiplatelet therapy (DAPT) initiation | -312
discharge from hospital | -312
Coronavirus-19 positive (asymptomatic) | -312
non-compliance with DAPT therapy | -288
new ischemic episode | -288
anterolateral ischemia on ECG | -288
femoro-femoral VA$ECMO support | 0
second coronary angiography | 0
stent placement on same vessels | 0
intra-aortic balloon pump (IABP) placement | 0
intensive care unit (ICU) admission | 0
trans-esophageal echocardiography (TEE) | 0
severe left ventricular dysfunction | 0
interventricular septum hypokinesia | 0
left atrial smoke | 0
minimal aortic valve opening | 0
mild aortic insufficiency | 0
severe reduction of right ventricle longitudinal function | 0
severe reduction of right ventricle concentric function | 0
transeptal left atrial cannulation | 480
VA$ECMO converted to LAVA$ECMO | 480
improvement in right ventricle movement | 480
improvement in anterior septum movement | 480
improvement in posterior wall movement | 480
persistent severe left ventricular dysfunction | 480
Levosimendan infusion | 504
progressive weaning from VA$ECMO | 528
conversion to LVAD | 528
vasopressor support decreased | 528
inotropic support decreased | 528
improved cardiac function | 528
reduced platelet count | 0
bleeding at cannula insertion sites | 0
airway bleeding | 0
packed red blood cell transfusions (4 units) | 0
strict coagulation monitoring | 0
pneumonia | 0
antibiotics initiation | 0
fibro-bronchoscopies | 0
renal failure (stage 3) | 0
continuous renal replacement therapy | 0
uncontrolled airway bleed | 936
death | 936
