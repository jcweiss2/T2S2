28 years old | 0
male | 0
near drowning | -120
ventilated | -120
acute respiratory distress syndrome | -120
ceftriaxone | -120
high-grade fever | 0
tachypnea | 0
oxygen saturation of 87% | 0
leukocytosis | 0
hemoglobin 11.1 g% | 0
normal electrolytes | 0
creatinine of 1.8 mg/dl | 0
endotracheal secretions sent for gram, fungal, acid-fast stain, and cultures | 0
blood samples sent for gram, fungal, acid-fast stain, and cultures | 0
urine samples sent for gram, fungal, acid-fast stain, and cultures | 0
antibiotic coverage changed to cefoperazone + sulbactam | 0
bilateral alveolar shadows on Chest X-ray | 0
cystic lesion in the lung parenchyma on Chest X-ray | 0
multiple ill-defined, round hypodense lesions in bilateral cerebral hemispheres with surrounding edema on CT brain | 0
multiple, well-defined, round, variable sized nodular lesions scattered in both lungs, with few of them showing central cavitation on CT chest | 0
patchy hypodensities in both kidneys on CT scan abdomen | 0
patchy hypodensities in the gluteal muscles bilaterally on CT scan abdomen | 0
normal echocardiography | 0
bronchoalveolar lavage (BAL) | 0
transbronchial biopsy | 0
antibiotic escalated to meropenem | 0
all microbiological laboratory reports negative on 2nd day of ICU admission | 48
serum galactomannan raised on 2nd day of ICU admission | 48
endotracheal aspirate for fungal stain showed Aspergillus species on 2nd day of ICU admission | 48
voriconazole and caspofungin combination started | 48
hemoptysis | 48
tachycardia | 48
desaturation | 48
fresh frozen plasma administered | 48
tranexamic acid administered | 48
septic shock | 72
vasopressors administered | 72
worsening respiratory acidosis | 72
leukopenia | 72
transbronchial biopsy report revealed neutrophilic exudates and foci of fungal broad hyphae, broad angle branching | 72
BAL specimen on culture revealed Aspergillus fumigatus growth | 96
patient expired | 120