36 years old | 0
female | 0
pregnant | 0
admitted to hospital | 0
recurrent vomiting | 0
epigastric pain | 0
diagnosed with uterine fibroid | -238
weight loss | -238
using iron tablets | -238
history of weight loss | -238
no change in bowel habits | -238
no hematemesis | -238
no rectal bleeding | -238
no hematuria | -238
no passing stones | -238
looked ill | 0
markedly dehydrated | 0
drowsy | 0
blood pressure 126/76 mmHg | 0
pulse rate 94 min–1 | 0
respiratory rate 30 min–1 | 0
temperature 36.6°C | 0
no lymphadenopathy | 0
no thyromegaly | 0
no edema | 0
uterus size of 40 weeks | 0
tender epigastric area | 0
drowsy and hypotonic | 0
brisk deep tendon reflexes | 0
no obvious focal neurological sign | 0
planter reflexes were down-going | 0
chest and cardiovascular systems were unremarkable | 0
hemoglobin 8.7 g/dl | 0
WBCs 7000 μl–1 | 0
platelets 445 000 μl–1 | 0
ESR 109 mm/h | 0
toxic granulation of WBCs | 0
BUN 4.4 mmol/l | 0
creatinine 59 μmol/l | 0
HCO3 22 mmol/l | 0
Na 138 mmol/l | 0
Ca 4.8 mmol/l | 0
uric acid 508 μmol/l | 0
lactic acid 1.2 mmol/l | 0
phosphorous 0.8 mmol/l | 0
HIV serology was negative | 0
calcium at 14 weeks’ gestation was 2.43 mmol/l | -238
ALT 4 u/l | 0
AST 11 u/l | 0
ALP 150 u/l | 0
total protein 72 g/l | 0
albumen 30 g/l | 0
cholesterol 4.05 mmol/l | 0
triglyceride 3.59 mmol/l | 0
PTH 3 pg/ml | 0
TSH 0.68 mIU/l | 0
free thyroxin 16.6 pmol/l | 0
cortisol 1849 nmol/l | 0
vitamin D 15 ng/ml | 0
given normal saline infusion | 0
given intramuscular calcitonin | 0
transferred to medical intensive care unit | 0
developed rupture membrane | 24
urgent cesarean section | 24
hypercalcemia | 0
hypotension | 24
blood transfusion | 24
delivered a baby girl | 24
removed uterine masses | 24
septicemia | 48
septic shock | 48
vasopressors | 48
broad-spectrum antibiotics | 48
postoperative laboratory test | 48
serum calcium 2.34 mmol/l | 48
phosphorus 1.1 mmol/l | 48
BUN 6.2 mmol/l | 48
Cr 75 mmol/l | 48
Na 143 mmol/l | 48
K 4.2 mmol/l | 48
HCO3 16 mEq/l | 48
chloride 113 mEq/l | 48
albumin 21 g/l | 48
serum lactate 5.19 | 48
serum PTH 155 pg/ml | 48
serum amylase 88 u/l | 48
serum lipase 73 u/l | 48
Hb 5.8 g/dl | 48
platelets 125 000 μl–1 | 48
CT scan of chest and pelvis | 72
MRI of brain | 72
MRA | 72
evidence of infarcts | 72
vasospasm of internal carotid | 72
middle and anterior carotid arteries | 72
diffuse ischemic changes | 72
condition began to improve | 96
discharged home | 168
final diagnosis of humoral hypercalcemia | 168
serum calcium remained within normal range | 432
diagnosed with hypercalcemic crisis | 0
hypercalcemia due to uterine fibroid | 0
humoral hypercalcemia of benignancy | 0
PTH-rP producing malignant tumors | -238
primary hyperparathyroidism | -238
hyperthyroidism | -238
immobilization | -238
vitamin D and vitamin A overdose | -238
familial hypocalciuric hypercalcemia | -238
diuretic phase of acute renal failure | -238
chronic renal failure | -238
thiazide diuretics | -238
sarcoidosis | -238
milk-alkali syndrome | -238
Addison's disease | -238
parathyroid hormone-related protein | -238
humoral hypercalcemia of malignancy | -238
breast cancer | -238
lung cancer | -238
ovarian cancer | -238
renal cell carcinoma | -238
lymphoma | -238
multiple myeloma | -238
calcitonin | 0
hemodialysis | 24
urgent hemodialysis | 24
physiotherapy | 168
generalized muscle weakness | 168
stiffness | 168