68 years old | 0
female | 0
residence in a long-term nursing facility | 0
dementia | 0
admitted to the hospital | 0
vomiting | -72
diarrhea | -72
bilateral leg swelling | -72
vague leg discomfort | -72
increased diuretic dose | -72
denied nausea | 0
denied abdominal pain | 0
denied bleeding | 0
denied fevers | 0
denied focal leg pain | 0
denied redness | 0
denied trauma | 0
denied rash | 0
denied shortness of breath | 0
denied chest pain | 0
nonalcoholic fatty liver disease | -672
cirrhosis | -672
chronic kidney disease stage III | -672
insulin-dependent type 2 diabetes | -672
never smoked cigarettes | 0
no history of alcohol | 0
no history of substance abuse | 0
afebrile | 0
heart rate of 55 | 0
BP of 96/43 mm Hg | 0
respiratory rate of 16 breaths/min | 0
oxygen saturation of 96 % | 0
BMI of 36 kg/m2 | 0
alert and conversant | 0
oriented to self and place only | 0
mucous membranes dry | 0
sclera anicteric | 0
regular heart rate | 0
no S3 | 0
normal JVP | 0
clear lungs | 0
abdomen benign | 0
stool hemoccult negative | 0
pitting lower extremity edema | 0
no focal tenderness | 0
no erythema | 0
hemoglobin level of 8.7 g/dL | 0
WBC count of 12,400/μL | 0
91 % segmental neutrophils | 0
no bands | 0
platelets of 77,000/μL | 0
sodium level of 138 mM | 0
potassium level of 4.4 mM | 0
bicarbonate level of 15 mM | 0
BUN level of 72 mg/dL | 0
creatinine level of 4.16 mg/dL | 0
total bilirubin of 1.9 mg/dL | 0
aspartate aminotransferase of 63 u/L | 0
alanine aminotransferase of 34 u/L | 0
INR of 2.1 | 0
ammonia of 94 umol/L | 0
venous lactate of 1.6 mmol/L | 0
sinus bradycardia | 0
multiple nodular densities | 0
ill-defined airspace opacities | 0
hypotensive | 2
BP of 78/34 mm Hg | 2
received fluid resuscitation | 2
received empiric broad spectrum antibacterials | 2
admitted to the hospital | 0
received additional IV fluids | 2
normal lactic acid level | 2
negative blood cultures | 2
negative urine cultures | 2
unable to produce sputum | 2
nasal swab for methicillin resistant Staphylococcus aureus negative | 2
vancomycin stopped | 50
liver enzymes elevated | 50
bedside portable ultrasound consistent with cirrhosis | 50
no evidence of biliary obstruction | 50
echocardiogram showed normal systolic and diastolic function | 50
progressive oliguric renal failure | 72
urinary sediment demonstrating acute tubular necrosis | 72
dialysis initiated | 72
hypoxic respiratory failure | 72
admitted to the Intensive Care Unit | 72
intubated | 72
follow up chest X-ray demonstrated worsening bilateral airspace disease | 96
supported with mechanical ventilation | 96
pressors | 96
dialysis | 96
intravenous piperacillin/tazobactam continued | 96
vancomycin resumed | 96
CVVHD initiated | 96
respiratory function stabilized | 240
unable to be weaned from the ventilator | 240
weakness | 240
waxing and waning encephalopathy | 240
hypervolemia | 240
pressor-dependent | 240
treated with stress-dose steroids | 240
hematologic abnormalities | 240
thrombocytopenia | 240
anemia | 240
coagulopathy | 240
transitioned to comfort care | 432
died | 432
autopsy demonstrated hepatic cirrhosis | 432
massive abdominal ascites | 432
esophageal varices | 432
intratubular oxylate crystals | 432
nodular glomerulosclerosis | 432
arterial and arteriolar nephrosclerosis | 432
mild to moderate aortocoronary atherosclerosis | 432
mild cardiomegaly | 432
myocyte hypertrophy | 432
acute and chronic pancreatitis | 432
heavy lungs | 432
ill-defined areas of consolidation | 432
septated hyphae with acute angle branching | 432
invasive pulmonary aspergillosis | 432
bilateral organizing pulmonary thromboemboli | 432