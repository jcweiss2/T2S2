48 years old| 0
    male| 0
    admitted to the hospital (outside hospital) | -1440
    diagnosed with multisystem sarcoidosis (bone marrow, liver, lymph nodes) | -1440
    progressive abdominal pain | -5760
    100-pound weight loss | -5760
    nausea | -5760
    vomiting | -5760
    paraplegia (due to motor vehicle accident) | -52560
    urinary retention | -52560
    asthma | 0
    type 2 diabetes mellitus | 0
    gastroesophageal reflux disease | 0
    hiatal hernia | 0
    hypertension | 0
    alcoholism | 0
    MRI thoracic spine (showing degenerative disc disease) | -26208
    MRI lumbar spine (showing disc bulging at L5–S1) | -26208
    albuterol | 0
    terazosin | 0
    oxybutynin | 0
    pantoprazole | 0
    leukopenia | -1440
    anemia | -1440
    CT abdomen and pelvis (revealing lymph node adenopathy, splenomegaly, liver parenchyma changes) | -1440
    liver biopsy | -1440
    bone marrow biopsy | -1440
    retroperitoneal lymph node biopsy | -1440
    diagnosed with sarcoidosis | -1440
    prednisone | -1440
    methotrexate | -1440
    admitted to the same hospital (3 days prior to transfer) | -72
    chest pain | -72
    anorexia | -72
    nausea | -72
    vomiting | -72
    continued abdominal pain | -72
    hypotension (blood pressure 85/63 mmHg) | 0
    temperature 98.6°F | 0
    pulse 117 bpm | 0
    respiratory rate 22 bpm | 0
    oxygen saturation 95% | 0
    CT thorax (negative for pulmonary embolism, moderate pleural effusions) | 0
    CT abdomen and pelvis (stable changes, new ascites) | 0
    negative urine and blood cultures | 0
    lactate 2.3 mmol/L | 0
    INR >12 | 0
    fibrinogen 50 mg/dL | 0
    ALT 86 IU/L | 0
    AST 204 IU/L | 0
    WBC 0.8 K/uL | 0
    hemoglobin 7.9 g/dL | 0
    platelets 92 K/uL | 0
    admitted to ICU | 0
    suspected sepsis | 0
    intravenous fluids | 0
    cefepime | 0
    vancomycin | 0
    vitamin K | 0
    hematology consultation | 0
    infectious disease consultation | 0
    rheumatology consultation | 0
    cefepime discontinued | 72
    vancomycin discontinued | 72
    methylprednisolone 1 gram for 3 days | 0
    transferred to our hospital | 0
    blood pressure 87/64 mmHg | 0
    pulse 104 bpm | 0
    respiratory rate 19 bpm | 0
    temperature 98.2°F | 0
    oxygen saturation 99% | 0
    soft, diffusely tender abdomen | 0
    rebound tenderness | 0
    bowel sounds | 0
    hepatosplenomegaly | 0
    pancytopenia (WBC 0.8 k/uL) | 0
    hemoglobin 9.3 g/dL | 0
    platelets 90 k/uL | 0
    ANC 0.76 K/uL | 0
    ALT 146 IU/L | 0
    AST 224 IU/L | 0
    INR 1.99 | 0
    PT 22 | 0
    PTT 43 | 0
    fibrinogen 106 mg/dL | 0
    D-Dimer 5.06 | 0
    lactic acid 5.0 mmol/L | 0
    ferritin 6,420 ng/mL | 0
    triglycerides 168 mg/dL |