61 years old | 0
    male | 0
    admitted to the emergency department | 0
    fever | -168
    dysphagia | -168
    cervical swelling | -168
    impacted fish bones in his throat | -168
    examined by the endoscopist | -168
    oral antibiotics | -168
    no improvement | -168
    dysphonia | 0
    cough | 0
    deterioration of general condition | 0
    body temperature 39 °C | 0
    white blood cell count 18,900/mm3 | 0
    hemoglobin level 11.3 g/dL | 0
    CRP 64 ng/ml | 0
    plasma glucose level 680 mg/dl | 0
    pH 7.4 | 0
    plasma osmolarity 320 mOsm/kg | 0
    nonketotic hyperosmolar coma | 0
    taken into the intensive care unit | 0
    intravenous insulin | 0
    0.9% NaCl administered | 0
    ceftriaxon 2 gr/day intravenously | 0
    fever remained high after three days | 72
    neck ultrasound examination | 72
    neck pain | 72
    abscess formation in the upper mediastinum | 72
    close relation to thyroid gland | 72
    cervicothoracic computed tomography (CT) | 72
    gas in upper mediastinum | 72
    pleural effusion in both hemithorax | 72
    gram stain of the needle aspiration | 72
    polymorphonuclear leukocytes existence | 72
    no bacteria | 72
    needle aspirat culture failed to show bacterial growth | 72
    ceftriaxon discontinued | 72
    meropenem 3 gr/day intravenously | 72
    symptoms resolved after five days of antibiotic treatment | 120
    control cervicothoracic CT on 10th day | 240
    abscess formation disappeared | 240
    pleural effusion disappeared | 240
    discharged after fifteen days | 360
    mediastinitis | 0
    diabetic patient | 0
    