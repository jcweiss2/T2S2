18 years old | 0
male | 0
hypertension | -672
diabetes | -672
fever | -144
rigors | -144
generalized headache | -144
altered mentation | -144
body malaise | -144
nausea | -144
vomiting | -144
history of malaria | -672
previous uncomplicated malarial infections | -672
febrile | 0
tachypneic | 0
disoriented | 0
splenomegaly | 0
normal vesicular breath sounds | 0
normal abdominal examination | 0
WBC count | 0
hemoglobin | 0
thrombocytopenia | 0
elevated creatinine | 0
elevated BUN | 0
low sodium | 0
normal serum electrolytes | 0
normal liver profile | 0
normal coagulation profile | 0
normal chest X-ray | 0
P. falciparum | 0
high parasitemia | 0
admitted to ICU | 0
intravenous artesunate-based regimen | 0
improved clinical status | 12
improved lab parameters | 12
shifted to general ward | 72
acute abdomen | 120
progressive abdominal pain | 120
nausea | 120
non-bilious vomiting | 120
low Hb | 120
urgent CBC | 120
grouping/crossmatch | 120
abdominal ultrasound | 120
contrast-enhanced CT scan | 120
hypoechoic nodular cystic area | 120
splenic laceration | 120
intraparenchymal hematoma | 120
intraparenchymal free fluid | 120
grade 3 splenic injury | 120
splenectomy | 120
evacuated 2.5 L of frank blood | 120
splenectomy done | 120
uneventful postoperative period | 168
discharged home | 168