32 years old | 0
male | 0
admitted to the hospital | 0
fracture of the right sacroiliac joint | 0
open wound of right tibial fracture | 0
elective surgery | 0
sacroiliac disruption | 0
pubic diastasis | 0
high-grade fever | 72
tachycardia | 72
hypotension | 72
increasing pain | 72
progressive swelling | 72
erythema | 72
crepitus | 72
severely swollen skin | 72
brownish skin | 72
necrotic wound | 72
foul smelling wound | 72
gas in the interfacial planes | 72
extensive gas formation | 72
increased total leukocyte counts | 72
erythrocyte sedimentation rate | 72
C-reactive-protein | 72
presumptive diagnosis of gas gangrene | 72
emergency surgical debridement | 72
wound debridement | 72
pus pockets removed | 72
necrosed medial gastrocnemius muscle debrided | 72
tissue and pus sample sent to microbiology laboratory | 72
gram-staining | 72
variable Gram-positive rods | 72
pus and tissue samples cultured | 72
anaerobic blood agar plate showed growth | 96
aerobic culture showed no growth | 96
colony identified as C. sordellii | 96
injection clindamycin started | 96
injection linezolid started | 96
antibiotics deescalated | 120
injection metronidazole started | 120
injection clindamycin continued | 120
patient clinical condition improved | 120
hyperbaric oxygen therapy | 144
wound healed | 240
repeated pus culture from the wound was sterile | 240
patient discharged | 480