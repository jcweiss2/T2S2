9 years old | 0
female | 0
Afghan | 0
admitted to the hospital | 0
car accident | -672
surgery at an Indian hospital | -672
external fixation | -672
femur nail | -672
dehydration | 0
undernourishment | 0
decreased serum concentration of total protein | 0
decreased creatinine | 0
anemia | 0
decubitus dorsal ulcers | 0
multiple wounds | 0
scab | 0
yellow pus | 0
fistula of her left hip joint | 0
methicillin resistant Staphylococcus aureus (MRSA) | 0
carbapenem resistant Pseudomonas aeruginosa | 0
Gram negative bacteria species with extended spectrum beta-lactamase activity (ESBL) | 0
Citrobacter sedlakii | 0
Escherichia coli | 0
Proteus mirabilis | 0
Klebsiella pneumoniae | 0
methicillin susceptible S. aureus | 0
P. mirabilis (non ESBL) | 0
Enterococcus faecalis | 0
Enterococcus hirae | 0
Bacteroides fragilis | 0
peptostreptococci | 0
initial treatment at the intensive care unit | 0
admitted to the pediatric surgery ward | 336
improved general condition | 336
16 surgeries | 336
60 dressing changes | 336
general anesthetics | 336
cefazoline | 0
imipenem | 0
meropenem | 0
ampicillin + clindamycin | 0
amoxicillin + clindamycin | 0
ceftazidime | 0
ceftaroline | 0
cefuroxime | 0
MRSA isolation | -168
decolonization cycle | -168
MRSA not found | -168
MRSA recolonization | 1344
biopsy sample | 1344
MRSA detection | 1344
amputation of her lower legs | 1440
knee disarticulation | 1440
systemic inflammatory response syndrome | 1440
increased heart rate | 1440
increased white blood cell count | 1440
decreased blood pressure | 1440
body temperature rose | 1440
C-reactive protein concentration increased | 1440
MRSA in blood culture | 1440
septic infection | 1440
antibiotic treatment with ceftaroline | 1440
improved general condition | 1464
final revision surgery | 1512
removal of the condylar cartilage | 1512
debridement of necrotic tissue | 1512
MRSA detection | 1512
inflammation parameters remained low | 1512
ceftaroline application stopped | 1512
discharged from the hospital | 2160
typing of MRSA isolates | 0
National Reference Centre for Staphylococci and Enterococci | 0
Robert Koch Institute | 0
informed consent | 0
ethics approval | 0
Institutional Review Board of Klinikum Ingolstadt | 0
standard treatment procedures | 0
no additional samples | 0
scientific purposes | 0
severe infection of both legs | 0
multiresistant bacteria | 0
bacteriologic analyses | 0
MRSA infection | 0
endogenous MRSA infection | 0
typing results | 0
screening results | 0
decolonization measures | 0
MRSA decolonization | 0
continuous MRSA monitoring | 0
infection treatment with ceftaroline | 1440
ceftaroline dosage | 1440
ceftaroline safety | 1440
ceftaroline efficacy | 1440
vancomycin | 0
linezolid | 0
daptomycin | 0
pediatric patients | 0
ceftaroline treatment | 1440
MRSA pneumonia | 0
body weight | 0
general condition | 0
initial therapy | 1440
low-dose treatment | 1440
postoperative course | 1440
satisfactory | 1440
circulation stabilized | 1440
body temperature decreased | 1440
C-reactive protein concentration | 1440
white blood cell count | 1440
extended wounds | 1440
inflammation parameters | 1512
ceftaroline MIC | 1440
reduced antibiotic susceptibility | 1440
clonal lineages | 0
ST228 | 0
ST239 | 0
CC8 | 0
ceftaroline resistance | 1440
MICs | 1440
treatment efficiency | 1440
susceptibility interpretive criteria | 0
pharmacokinetic | 0
pharmacodynamic | 0
in vitro analyses | 0
breakpoint | 0
treatment failure | 0
potent antibiotic | 0
broadly resistant MRSA | 0
speaker’s honorarium | 0
AstraZeneca | 0
conflicts of interest | 0
Figure 1 | 0
Microbiological results | 0
antibiotic treatment | 0
Figure 2 | 0
Vital signs | 1440
MRSA finding | 1440
MAP | 1440
mean arterial pressure | 1440
intensive care unit | 1440
Table 1 | 0
Characteristics of MRSA isolates | 0
spa type | 0
CC | 0
SCCmec | 0
PVL | 0
phenotypic resistance pattern | 0
MIC ceftaroline | 0
BMD | 0
Etest | 0
EUCAST guidelines | 0