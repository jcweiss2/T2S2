68 years old | 0
male | 0
Caucasian | 0
anterior mediastinal mass | -672
thymoma | -672
declined surgery | -672
gross hematuria | 0
oral mucosal bleeding | 0
generalized weakness | -720
fatigue | -720
subjective fever | -720
unintentional weight loss | -720
marked pancytopenia | 0
broad spectrum antibiotics | 0
transfused with red blood cells | 0
transfused with platelets | 0
severe thrombocytopenia | 0
neutropenia | 0
inappropriately low retic count | 0
admitted to the intensive care unit | 0
vancomycin | 0
piperacillin/tazobactam | 0
intravenous methylprednisolone | 0
bone marrow biopsy | 24
severe AA | 24
cyclosporine | 48
eltrombopag | 48
anti-thymocyte globulin | 48
thymoma resection | 48
platelets count improved | 72
absolute neutrophil count remained low | 72
posaconazole | 72
acyclovir | 72
transient sudden loss of consciousness | 120
hypotension | 120
oxygen desaturation | 120
stroke alert | 120
CT brain | 120
new maxillary swelling | 120
maxillary swelling increased | 144
intubated | 144
sedated | 144
self-tamponade | 144
blood cultures positive | 216
Gram-negative rods | 216
Fungemia | 216
cefepime | 216
micafungin | 216
multiorgan failure | 216
DNR | 216
cardiopulmonary arrest | 216
expired | 216
profound pancytopenia | 0
white blood cells low | 0
absolute neutrophil count low | 0
RBCs low | 0
platelets low | 0
hemoglobin low | 0
reticulate count low | 0
peripheral blood smear | 0
mild anisocytosis | 0
bone marrow biopsy | 24
profound hypocellularity | 24
decreased numbers in all hematopoietic lineages | 24
bone marrow aspirate | 24
no evidence of dysplasia | 24
residual cells | 24
HUS/TTP screening labs | 0
lactate dehydrogenase normal | 0
haptoglobin elevated | 0
fibrinogen elevated | 0
direct bilirubin elevated | 0
renal function test | 0
elevated creatinine | 0
elevated BUN | 0
electrolytes normal | 0
urine cultures negative | 0
blood cultures negative | 0
Lyme disease suspected | 0
Ehrlichia chaffeensis suspected | 0
antibodies screening negative | 0
complement C3 normal | 0
complement C4 elevated | 0
ANA negative | 0
ANCA negative | 0
myasthenia-related anti-Ach antibodies negative | 0
myeloperoxidase antibodies negative | 0
proteinase-3 antibodies negative | 0
Vitamin B12 normal | 0
chest X-ray | 0
CT chest | 0
interval enlargement of anterior mediastinal mass | 0
thymoma versus invasive thymoma | 0
differential diagnosis | 0
TR-AA | 0
HUS/TTP | 0
leukemia | 0
myelodysplasia | 0
multiple myeloma | 0
autoimmune conditions | 0
infective agents | 0
outcome | 216
fatal TR-AA | 216
optimal treatment | 0
high-dose systemic steroids | 0
cyclosporine | 48
eltrombopag | 48
anti-thymocyte globulin | 48
broad spectrum antibiotics | 0
RBCs transfusion | 0
platelets transfusion | 0
AA-related complications | 120
severe thrombocytopenia | 120
neutropenia | 120
rapidly expanding soft tissue neck swelling | 120
impeded respiration | 120
emergent endotracheal intubation | 144
mechanical ventilation | 144
bacteremia | 216
fungemia | 216
septic shock | 216
multiorgan failure | 216
cardiopulmonary arrest | 216
DNR | 216
expired | 216