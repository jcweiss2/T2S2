52 years old | 0
    female | 0
    admitted to the hospital | 0
    colicky | 0
    left flank pain | 0
    no chronic diseases | 0
    no immunodeficiency diseases | 0
    no urolithiasis | 0
    no urinary tract infections | 0
    vital signs stable | 0
    blood pressure 110/70 mmHg | 0
    respiratory rate 20/min | 0
    pulse rate 69/min | 0
    temperature 37.0℃ | 0
    left flank pain | 0
    left costovertebral angle tenderness | 0
    WBC 9,970/mm3 | 0
    neutrophils 84.4% | 0
    lymphocytes 6.4% | 0
    hemoglobin 10.6 g/dL | 0
    platelet count 142,000/mm3 | 0
    CRP 57.5 mg/dL | 0
    BUN 19 mg/dL | 0
    creatinine 0.8 mg/dL | 0
    total protein 6.5 g/dL | 0
    albumin 3.2 g/dL | 0
    total bilirubin 2.2 mg/dL | 0
    aspartate aminotransferase 34 IU/L | 0
    alanine aminotransferase 47 IU/L | 0
    no WBCs in urinalysis | 0
    RBCs over 100/HPF | 0
    urinary stone in left ureter | 0
    ESWL on 3rd day | 72
    ESWL on 4th day | 96
    received 8,000 shocks | 72
    flank pain aggravated | 72
    costovertebral angle tenderness aggravated | 72
    body temperature rose to 39.9℃ | 168
    blood pressure 70/50 mmHg | 168
    heart rate 125/min | 168
    respiratory rate 26/min | 168
    temperature 39.0℃ | 168
    oxygen saturation 80% | 168
    moved to ICU | 168
    mechanical ventilation | 168
    shock management | 168
    WBC 18,400/mm3 | 168
    neutrophils 90.4% | 168
    lymphocytes 5.5% | 168
    hemoglobin 11 g/dL | 168
    platelet count 92,000/mm3 | 168
    CRP 240 mg/dL | 168
    BUN 56 mg/dL | 168
    creatinine 2.4 mg/dL | 168
    cefepime administration | 168
    vancomycin administration | 168
    computed tomography showed ureter stone | 168
    hydroureteronephrosis | 168
    no WBCs in urine | 168
    no RBCs in urine | 168
    urine cultures negative | 168
    blood cultures positive for gram-negative bacilli | 168
    Achromobacter xylosoxidans identified | 168
    imipenem/cilastatin 4 µg/mL | 168
    meropenem 4 µg/mL | 168
    piperacillin-tazobactam 8 µg/mL | 168
    ampicillin 16 µg/mL | 168
    ciprofloxacin 2 µg/mL | 168
    amikacin 32 µg/mL | 168
    aztreonam 16 µg/mL | 168
    cefepime 16 µg/mL | 168
    cefepime resistant | 168
    antibiotics changed to imipenem | 168
    blood cultures negative for A. xylosoxidans on 14th day | 336
    renal function worsened | 336
    continuous renal replacement therapy | 336
    Burkholderia cepacia isolated on 16th day | 384
    B. cepacia susceptible to imipenem/cilastatin | 384
    central venous catheter removed | 384
    tip culture negative | 432
    repeated blood cultures negative after three days | 432
    respiratory failure | 504
    bilateral opacities on chest imaging | 504
    passed away | 696
    septic shock | 696
    multiple organ failure | 696
    16S rRNA sequencing identified isolate | 696
    primers 515FPL and 13B used | 696
    sequencing with Taq polymerase | 696
    GenBank comparison | 696
    100% sequence identity with A. xylosoxidans | 696