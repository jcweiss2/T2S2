69 years old | 0
male | 0
treated for high-grade B-cell non-Hodgkin lymphoma | 0
developed from advanced follicular lymphoma through Richter’s transformation | 0
comorbidities: severe chronic ischemic heart disease | 0
arterial hypertension | 0
chronic bronchitis | 0
type 2 diabetes mellitus | 0
intended for treatment with three cycles of salvage immunochemotherapy with rituximab, ifosfamide, carboplatin, and etoposide (RC-ICE) | 0
autologous haematopoietic stem cell transplantation | 0
second cycle complicated by oropharyngeal mucositis with candida superinfection | -672
treated by amikacin | -672
piperacillin/tazobactam | -672
fluconazole | -672
third cycle of R-ICE with pegfilgrastim support | -504
first episode of sepsis | -336
not participated in the telemonitoring project | -336
seventh day of the third cycle of R-ICE | -168
called emergency phone number | -168
not feeling well over the past 2 days | -168
weakness | -168
diarrhea | -168
fever | -168
dyspnea | -168
advised to go to the hospital immediately | -168
initial examination revealed signs of septic shock | -168
hypotensive with blood pressure 90/57 mm Hg | -168
tachycardic (120/min) | -168
dyspneic | -168
immediately admitted to the ICU | -168
laboratory findings: neutropenia – WBC count of 0.68 × 109/L | -168
absolute neutrophil count (ANC) of 0.6 × 109/L | -168
CRP concentration on admission was 120 mg/L | -168
kidney injury classified as 1st stage of acute kidney injury (KDIGO) | -168
lactate acidosis (4.32 mmol/L) | -168
base excess of −9.8 | -168
electrolyte imbalance: hyponatremia of 133 mmol/L | -168
hypokalemia of 3.2 mmol/L | -168
broad-spectrum antibiotics administered immediately (meropenem, linezolid) | -168
fluid resuscitation initiated | -168
hypotension progressed, necessitating continuous infusion of norepinephrine | -168
blood cultures revealed Escherichia coli sensitive to antibiotics | -168
stool samples: non-toxin-producing Clostridium difficile detected | -168
CRP peaked 2 days later at 286 mg/L | -144
kidney injury progressed into oligoanuric acute kidney insufficiency stage 3 (KDIGO) | -144
treated with continuous diuretic support | -144
chest X-ray showed bilateral opacities at the bases of the lungs | -144
differential diagnosis: co-infection combined with ischemic damage following septic shock | -144
treatment complicated by oral candidiasis | -144
herpes labialis | -144
necessitating additional antimicrobial treatment | -144
patient’s condition gradually improving until thirteenth day | -144
fever returned | -144
diarrhea returned | -144
E. coli cultivated from blood culture from peripherally inserted central catheter | -144
C. difficile detected in stool samples | -144
Clostridioides toxin detected | -144
peripherally inserted central catheter extracted | -144
catheter tip culture negative | -144
antibiotic treatment: piperacillin, tazobactam, amikacin, fidaxomicin | -144
patient finally recovered | -144
discharged after 27 days of ICU hospitalization | 0
therapy succeeded | 0
treatment strategy changed | 0
intended autologous stem cell transplantation replaced by chimeric antigen receptor-T cell therapy | 0
enrolled in telemedicine project | 0
lymphoma progressed before chimeric antigen receptor-T cell therapy initiated | 0
combination of rituximab, gemcitabine, oxaliplatin used as bridge therapy | 0
fifth day of the second cycle of regimen | 504
developed another infectious complication | 504
fever (38.4°C) detected during regular morning measurement | 504
contacted by phone | 504
advised to go to the hospital | 504
admitted within 3 hours from first occurrence of fever | 504
diarrhea | 504
vomiting | 504
blood pressure of 189/93 mm Hg | 504
irregular tachycardia with multiple ventricular extrasystoles | 504
immediately admitted to the ICU | 504
laboratory findings: WBC of 3.16 × 109/L | 504
neutrophils 2.95 × 109/L | 504
WBC decreased to 1.1 × 109/L the next day | 552
CRP level on admission was 32 mg/L | 504
peaking 2 days later at 271 mg/L | 552
serum electrolytes within normal range | 504
renal parameters within normal range | 504
intravenous hydration initiated | 504
antibiotic treatment: cefepime and amikacin | 504
granulocyte colony-stimulating factor administered | 504
blood culture revealed E. coli sensitive to antibiotics | 504
first-line therapy sufficient | 504
patient recovered after 10 days | 552
discharged from the hospital | 552
