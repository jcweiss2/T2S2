24 years old|0
male|0
weighing 80 kg|0
no co-morbidities|0
sore throat| -240
difficulty in swallowing| -240
pain on left side of the neck| -96
swelling on left side of the neck| -96
severe throbbing headache| -48
vomiting| -48
restlessness| -48
bulge in posterior pharyngeal wall|0
deviated uvula to the right|0
febrile|0
tachycardic|0
tender swelling on left side of the neck|0
Hb 13.3 gm%|0
total count 9800 cells/cumm|0
platelet count 282210 cells/cumm|0
ESR 37 mm/h|0
HIV negative|0
left parapharyngeal abscess|0
thrombosis of left IJV|0
reduced flow or stasis in left transverse and sigmoid sinuses|0
diagnosis of Lemierre's syndrome|0
parapharyngeal abscess drained|0
imepenem started|0
fondaparinux started|0
persistent hypotension|48
systolic pressures 70-90 mmHg|48
total count decreased to 3720 cells/cumm|48
platelet count dropped to 35000/cumm|48
activated partial thromboplastin time prolonged (84 s)|48
serum procalcitonin 1.4 ng/mL|48
diagnosis of septic shock|48
shifted to intensive care unit|48
imipenem stopped|48
vancomycin started|48
clindamycin started|48
metronidazole started|48
single donor platelet units transfused|48
central venous access via right femoral vein|48
fondaparinux stopped|48
noradrenaline infusion started|48
S. aureus sensitive to vancomycin and clindamycin|48
blood culture negative|48
no anaerobes isolated|48
progressively tachypneic|96
hypoxemic|96
bilateral lower zone opacities on chest X-ray|96
intubated|96
ventilated|96
gradual recovery|168
weaned off inotrope|168
weaned off ventilator support|168
platelet count improved to 379000/cumm|168
coagulation normalized|168
chest X-ray normalized|168
discharged to ward|240
Glasgow coma scale 15/15|0
no neurological deficits|0
discharged from hospital|504
oral linezolid continued for 3 weeks|504
