66 years old | 0
female | 0
admitted to the hospital | 0
fever | -72
systemic fatigue | -72
confusion | -72
restlessness | -72
depression | -100000
rectal cancer | -100000
osteoarthritis of the left knee | -100000
amitriptyline | -100000
trazodone | -100000
triazolam | -100000
flunitrazepam | -100000
duloxetine | -100000
aripiprazole | -100000
Glasgow Coma Scale, E3V4M5 | 0
blood pressure, 140/86 mmHg | 0
heart rate, 130 beats/min | 0
body temperature, 40.4 °C | 0
respiratory rate, 26/min | 0
SpO2, 94% | 0
costovertebral angle tenderness | 0
confusion | 0
C-reactive protein elevation | 0
creatine kinase elevation | 0
renal function tests elevation | 0
pyuria | 0
ureteral stone in the right urinary duct | 0
swelling of the right kidney | 0
septic shock | 0
obstructive pyelonephritis | 0
urolithiasis | 0
meropenem | 0
intraurethral catheter | 0
haloperidol | 0
improved hemodynamics | 48
noradrenaline administration ended | 48
lucid | 48
afebrile | 48
worsened consciousness | 48
Glasgow Coma Scale, E1VTM2 | 48
hyperthermia | 72
roving eye movement | 72
decreased tonus | 120
cogwheel rigidity | 120
clonic spasms | 120
elevated creatine kinase | 120
hepatitis virus antigens negative | 120
human immunodeficiency virus antigen negative | 120
autoantibodies negative | 120
vitamins normal | 120
trace elements normal | 120
improved pyelonephritis | 72
albuminocytologic dissociation | 96
bacterial culture negative | 96
herpes virus PCR negative | 96
cytomegalovirus antigen negative | 96
electroencephalography normal | 96
NMS diagnosis | 96
dantrolene | 96
bromocriptine | 96
renal replacement therapy | 96
tracheostomy | 120
MRI showed diffuse hyperintense signal in the cerebellar cortex | 240
MRI showed symmetrical hyperintense signals in the cerebellar dentate nucleus, superior cerebellar peduncle, and thalamus | 240
MRI showed hyperintense signals in the bilateral substantia nigra and bilateral globus pallidus | 648
improved brain MRI findings | 2160
transferred to another hospital for rehabilitation | 3564