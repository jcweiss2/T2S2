36 years old | 0
female | 0
admitted to the hospital | 0
abdominal pain | 0
constipation | 0
jaundice | 0
hypertension | -48
pre-eclamptic toxaemia | -48
emergency lower segment caesarean section (LSCS) | -48
delivered triplets | -48
elevated alanine amino transferase (ALT) | -24
elevated aspartate amino transferase (AST) | -24
hyperbilirubinaemia | -24
tachycardia | 0
heart rate of 140/minute | 0
blood pressure 176/100 mmHg | 0
peripheral oxygen saturation of 92% | 0
tachypnoea | 0
decreased air entry in bilateral lower lung fields | 0
abdomen was tender, distended and tense | 0
oliguria | 0
right-sided consolidation with pleural effusion | 0
massive intraperitoneal collection with thickened bowel loops | 0
severe thrombocytopenia | 0
haemoglobin of 10.2 g% | 0
white blood cells 11.2 × 10^9/L | 0
normal coagulation profile | 0
diagnostic ascites tapping | 0
bowel injury suspected | 0
exploratory laparotomy | 12
haemorrhagic liver parenchyma | 12
no bowel, uterus or abdominal organ injury | 12
received 12 units of platelets | 12
intubated | 12
shifted to the intensive care unit (ICU) | 12
metabolic acidosis | 12
cultures of urine, sputum and blood sent | 12
negative cultures | 24
hepatitis viral markers and HIV negative | 24
peripheral smear showed fragmented red cells | 24
anaemia with dimorphic cells | 24
polychromatic cells with burr cells | 24
thrombocytopenia | 24
leucocytosis with absolute neutrophilia | 24
microangiopathic haemolytic anaemia | 24
hyperbilirubinaemia | 24
elevated liver enzymes | 24
hypoalbuminaemia | 24
antineutrophilic cytoplasmic antibodies (ANCAs) negative | 24
antinuclear antibodies (ANAs) negative | 24
plasmapheresis initiated | 30
plasmapheresis done eight times | 30-216
haemodialysis done four times | 30-216
received five units of packed red cells | 48
thrombocytopenia improved | 240
liver function tests improved | 240
renal function improved | 240
lung condition improved | 240
extubated | 264
urine output increased | 312
shifted to the ward | 360
discharged home | 600