63 years old | 0
male | 0
admitted to the hospital | 0
productive cough | -72
dyspnea | -72
pulmonary tuberculosis | -8760
treated (pulmonary tuberculosis) | -8760
smoking 15 packs/year | -8760
sought medical care | -1344
treated with symptomatic medication | -1344
plain chest radiography | -1344
mild mediastinal enlargement | -1344
bulging on the right atrium contour | -1344
afebrile | 0
normal hemodynamic parameters | 0
no peripheral edema | 0
normal lung examination | 0
ejection murmur | 0
raised jugular venous pressure | 0
hepatomegaly | 0
normal remaining examination | 0
unremarkable laboratory workup | 0
pericardium thickening | 0
mild effusion | 0
left ventricular ejection fraction 60% | 0
mass infiltrating pericardium | 0
mass infiltrating anterior wall of the right atrium | 0
bilateral pulmonary nodules | 0
pulmonary nodules up to 2.6 cm | 0
mass diffusely involving pericardium | 0
compression of right ventricle’s outflow tract | 0
compression of pulmonary artery | 0
compression of superior vena cava | 0
pericardial biopsy | 0
no evidence of malignancy (pericardium) | 0
pulmonary nodule biopsy | 0
sinusoidal vascular channels | 0
atypical endothelial cells | 0
positivity for CD31 | 0
positivity for CD34 | 0
negativity for Desmin | 0
negativity for S100 Protein | 0
diagnosis of angiosarcoma | 0
metastatic angiosarcoma primary to the right atrium | 0
chemotherapy with doxorubicin | 0
chemotherapy with ifosfamide | 0
reduction in pulmonary nodules size | 504
pulmonary infection | 864
admitted to emergency department | 864
refractory septic shock | 864
death | 864
