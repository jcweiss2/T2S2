55 years old | 0
female | 0
Caucasian | 0
admitted to the hospital | 0
chest pain | 0
palpitations | 0
shortness of breath | 0
nausea | 0
blood pressure 182/87 mmHg | 0
heart rate 74 bpm | 0
temperature 98.3°F | 0
oxygen saturation 94% | 0
troponin 0.26 ng/mL | 0
creatinine 1.5 mg/dL | 0
white blood cell 21.6 K/uL | 0
blood glucose 497 mg/dL | 0
aspartate aminotransferase 110 U/L | 0
alanine aminotransferase 133 U/L | 0
lactic acid 6.9 mmol/L | 0
pro-BNP 926 pg/mL | 0
ST segment elevations in leads V1 and V2 | 0
CT pulmonary angiography with contrast | 0
incidental finding of 3.5 cm x 4.1 cm hypodense right adrenal mass | 0
admitted to the intensive care unit | 0
heparin drip at 12 Units/kg/hr | 0
metoprolol 12.5 mg two times daily | 0
cefepime 1 g | 0
lactated ringers bolus 30 ml/kg | 0
insulin drip at 0.1 Units/Kg/hr | 0
worsening chest pain | 12
worsening palpitations | 12
troponin rose to 1.00 ng/mL | 12
emergent echocardiogram | 12
ejection fraction 40-45% | 12
septal hypokinesis | 12
lateral hypokinesis | 12
anteroseptal hypokinesis | 12
posterolateral hypokinesis | 12
cardiac angiography | 24
normal coronary vessels | 24
myocarditis considered | 24
erythrocyte sedimentation rate 0 mm/hr | 24
improvement in chest pain | 48
oxygen requirement decreased | 48
lactic acid trended down to 2.0 mmol/L | 48
blood glucose decreased to 179 mg/dL | 48
AST improved to 39 U/L | 48
ALT improved to 41 U/L | 48
plasma metanephrine 2.13 nmol/L | 48
normetanephrine 4.15 nmol/L | 48
doxazosin 2 mg daily | 48
carvedilol 3.125 mg two times daily | 48
CT Adrenal with and without contrast | 72
complex right adrenal mass suspicious for pheochromocytoma | 72
robotic assisted laparoscopic right adrenalectomy | 168
histochemical features consistent with pheochromocytoma | 168
echocardiogram 2 months after adrenalectomy | 1440
resolution of cardiomyopathy | 1440