57 years old | 0 | 0 | Factual
Hispanic | 0 | 0 | Factual
male | 0 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
history of coronary artery disease | -0 | 0 | Factual
myocardial infarction | -0 | 0 | Factual
ischemic dilated cardiomyopathy | -0 | 0 | Factual
pocket infection of his cardiac resynchronization therapy defibrillator | -0 | 0 | Factual
initial device and leads implanted | -6480 | -6480 | Factual
generator change | -432 | -432 | Factual
2-month history of erythema | -720 | -0 | Factual
discomfort around his left upper chest implant site | -720 | -0 | Factual
edema | -0 | 0 | Factual
serosanguinous drainage | -0 | 0 | Factual
oral amoxicillin treatment | -720 | -0 | Factual
nonbacteremic | 0 | 0 | Factual
afebrile | 0 | 0 | Factual
laboratory investigations within normal limits | 0 | 0 | Factual
echocardiography revealed severely reduced left ventricular systolic function | 0 | 0 | Factual
ejection fraction of 20%–25% | 0 | 0 | Factual
global hypokinesis of the left ventricle | 0 | 0 | Factual
no evidence of vegetations | 0 | 0 | Factual
preoperative computed tomography revealed that his leads were scarred to the lateral wall of the superior vena cava | 0 | 0 | Factual
transvenous lead extraction | 0 | 0 | Factual
cardiac resynchronization therapy defibrillator pocket capsule was dissected out | 0 | 0 | Factual
device removed | 0 | 0 | Factual
coronary sinus and right atrial leads extracted | 0 | 0 | Factual
right ventricular lead extracted | 0 | 0 | Factual
patient suddenly became hypotensive | 0 | 0 | Factual
transesophageal echocardiography revealed a large pericardial effusion | 0 | 0 | Factual
emergency midsternotomy | 0 | 0 | Factual
pericardium opened | 0 | 0 | Factual
significant amount of blood seen | 0 | 0 | Factual
bleeding manually controlled with pressure | 0 | 0 | Factual
cardiopulmonary bypass instituted | 0 | 0 | Factual
5-mm tear in the superior cavoatrial junction | 0 | 0 | Factual
perforation in the right atrium | 0 | 0 | Factual
oozing hematoma at the level of the innominate vein | 0 | 0 | Factual
lesions repaired with multiple 4-0 polypropylene sutures | 0 | 0 | Factual
right ventricular lead capped and abandoned | 0 | 0 | Factual
intra-aortic balloon pump placed | 0 | 0 | Factual
coagulopathy developed | 0 | 0 | Factual
transfusions of cryoprecipitate, platelets, fresh frozen plasma, and factor VII | 0 | 0 | Factual
coagulopathy improved | 0 | 0 | Factual
chest closed | 0 | 0 | Factual
postoperatively transferred to the intensive care unit | 0 | 0 | Factual
severe cardiogenic shock | 0 | 24 | Factual
multiorgan failure | 0 | 24 | Factual
hypotensive | 0 | 24 | Factual
required large doses of vasopressin, epinephrine, and norepinephrine | 0 | 24 | Factual
hypoxic respiratory failure | 0 | 24 | Factual
mechanical ventilation | 0 | 168 | Factual
liver failure | 0 | 24 | Factual
albumin | 0 | 240 | Factual
blood products given | 0 | 240 | Factual
broad-spectrum antibiotics | 0 | 240 | Factual
oliguric | 0 | 24 | Factual
continuous venovenous hemodialysis | 24 | 984 | Factual
bilateral, symmetrical cyanotic changes | 48 | 216 | Factual
vasopressor administration stopped | 48 | 48 | Factual
upper- and lower-digit ischemia progressed to dry gangrene | 216 | 216 | Factual
dull pain | 216 | 216 | Factual
no ability to move his fingers and toes | 216 | 216 | Factual
bilateral stiffness | 216 | 216 | Factual
2+ pitting edema | 216 | 216 | Factual
nonexistent capillary refill time | 216 | 216 | Factual
palpable 2+ peripheral pulses | 216 | 216 | Factual
Doppler study showed flat waveforms | 216 | 216 | Factual
intra-aortic balloon pump removed | 168 | 168 | Factual
endotracheal tube removed | 168 | 168 | Factual
albumin discontinued | 240 | 240 | Factual
liver enzymes returned to normal limits | 240 | 240 | Factual
kidney function improved | 240 | 984 | Factual
hemodialysis stopped | 984 | 984 | Factual
mental status improved | 240 | 984 | Factual
sedation weaned off | 240 | 984 | Factual
necrotic lesions treated conservatively | 240 | 984 | Factual
povidone-iodine dressings | 240 | 984 | Factual
debridement | 648 | 648 | Factual
negative-pressure wound therapy | 648 | 984 | Factual
purulent, foul-smelling material drained | 648 | 984 | Factual
transferred to our facility | 1296 | 1296 | Factual
preoperative transesophageal echocardiography | 1296 | 1296 | Factual
ejection fraction of 10%–15% | 1296 | 1296 | Factual
laser extraction of his retained lead | 1392 | 1392 | Factual
pus drained from the subfascial area | 1392 | 1392 | Factual
antibiotic regimen started | 1392 | 1392 | Factual
microbial cultures grew Enterobacter cloacae and Staphylococcus epidermidis | 1392 | 1392 | Factual
transvenous implantable cardioverter-defibrillator system implanted | 1536 | 1536 | Factual
evaluation of his hands and feet | 1536 | 1536 | Factual
no signs of local infection or wet gangrene | 1536 | 1536 | Factual
black skin changes and demarcation lines | 1536 | 1536 | Factual
frank mummification of his digits and toes | 1536 | 1536 | Factual
discharged | 1848 | 1848 | Factual
amputation and debridement of his necrotic feet | 2544 | 2544 | Factual
amputation of his fingers scheduled | 2544 | 0 | Factual