51 years old | 0
male | 0
admitted to ICU | 0
acute circulatory failure | 0
diarrhea | -48
rigors | -48
chronic kidney disease | -10000
diabetes mellitus | -10000
sarcoidosis | -10000
hepatosplenic involvement | -10000
splenectomy | -5040
hydroxychloroquine treatment | -10000
no immunosuppressive drug | 0
vaccinated against Streptococcus pneumoniae | -10000
vaccinated against Neisseria meningitidis | -10000
no antibiotic prophylaxis | 0
one dog at home | -10000
central body temperature 34.4 °C | 0
heart rate 121/min | 0
arterial blood pressure 80/40 mmHg | 0
respiratory rate 20/min | 0
SpO2 99% | 0
Glasgow coma score 15 | 0
alert and oriented | 0
no neck stiffness | 0
lung auscultation irrelevant | 0
abdominal examination irrelevant | 0
no heart murmur | 0
extensive non-blanching rash | 0
lactic acidosis | 0
acute-on-chronic kidney failure | 0
disseminated intravascular coagulation | 0
biological inflammatory syndrome | 0
thoracic and abdominal CT-scan | 0
transthoracic echocardiography | 0
negative urinary sample examination | 0
negative pneumococcal urinary antigen test | 0
empirical antibiotic therapy with cefotaxime | 0
massive fluid loading | 0
renal replacement therapy | 0
invasive mechanical ventilation | 0
hydrocortisone | 0
vasopressor support with norepinephrine | 0
clinical condition deterioration | 5
death | 10
blood cultures drawn | 0
Enterococcus cecorum identification | 9
susceptible to ampicillin | 9
susceptible to vancomycin | 9
susceptible to linezolid | 9
susceptible to rifampicin | 9
susceptible to third-generation cephalosporin | 9
sterile blood cultures after cefotaxime | 6