71 years old | 0
    African American woman | 0
    type 2 diabetes mellitus | 0
    chronic kidney disease stage IV | 0
    hypertension | 0
    heart failure with preserved ejection fraction | 0
    chronic obstructive pulmonary disease | 0
    gout | 0
    admitted to the burn intensive care unit | 0
    worsening maculopapular rash | -168
    allopurinol | -168
    erosive rash | -168
    coverage of 25% total body surface area | -168
    ocular involvement | -168
    oropharyngeal involvement | -168
    skin biopsies consistent with SJS/TEN | 0
    SCORTEN score 4 | 0
    IV corticosteroids | 0
    IVIG therapy | 0
    respiratory failure | 0
    intubation | 0
    septic shock | 0
    ileus | 0
    oliguric renal failure | 0
    continuous renal replacement therapy | 0
    bloody diarrhea | 504
    drop in hemoglobin from 10.3 to 6.5 g/dL | 504
    Clostridium difficile assay negative | 504
    upper endoscopy showing antral gastritis | 504
    colonoscopy revealing perianal skin breakdown | 504
    cecum ulcers | 504
    ileocecal valve ulcers | 504
    ascending colon ulcerated, edematous mucosa | 504
    hematochezia | 504
    transfusion-dependent anemia | 504
    over 70 units of packed red blood cells | 504
    unsuccessful colonoscopy | 504
    unsuccessful radiologic guided embolization | 504
    ileocecectomy recommended | 504
    family declined surgical management | 504
    IV dexamethasone 100 mg daily | 504
    IV methylprednisolone 120 mg daily | 504
    prolonged prednisone taper | 504
    multidisciplinary conference discussed infliximab therapy | 504
    risks of further immunosuppression outweighed benefits | 504
    bleeding not slowed in response to corticosteroid therapy | 504
    death | 1728
    septic shock refractory to vasopressors | 1728
    