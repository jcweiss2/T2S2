51 years old | 0
male | 0
admitted to the hospital | 0
high-grade fever | -360
intermittent fever | -360
cough with expectoration | -360
breathlessness | -24
nebulized bronchodilators | -360
steroids | -360
quinolones | -360
hypertension | 0
childhood onset bronchial asthma | 0
chronic steroid therapy | 0
tachycardia | 0
tachypnea | 0
bilateral crepitations | 0
wheeze | 0
eschar on the left side of the chest | 0
azithromycin | 0
doxycycline | 0
oseltamivir | 0
throat swab for H1N1 | 0
sepsis workup | 0
intubated | 0
meropenem | 0
teicoplanin | 0
CT scan of the brain | 0
CT scan of the thorax | 0
CT scan of the abdomen | 0
bilateral multifocal patchy consolidation | 0
minimal right-sided pleural effusion | 0
collapse of left lung fields | 0
consolidation | 0
tracheal aspirate sent for Gram stain | 0
moderate polymorphonuclear neutrophils | 0
branching filamentous bacilli | 0
Nocardia species | 0
cotrimoxazole | 0
imipenem | 0
tracheal aspirates | 24
Gram stain findings | 24
dry chalky white colonies | 24
pitting on blood agar | 24
pitting on chocolate agar | 24
amikacin | 24
ciprofloxacin | 24
linezolid | 24
ceftriaxone | 24
resistant to cotrimoxazole | 24
resistant to amoxicillin-clavulanate | 24
Nocardia otitidiscaviarum | 24
MALDI-TOF MS | 24
acid-fast stain for Mycobacteria | 24
HIV 1 and 2 antibodies | 24
H1N1 RT-PCR | 24
white blood cell counts | 24
neutrophilic predominance | 24
thrombocytopenia | 24
platelet count | 24
scrub typhus IgM antibodies | 24
ventilatory support | 24
hemodynamics | 24
inotropic requirement | 24
repeat blood cultures | 120
yeast-like cells | 120
caspofungin | 120
Candida tropicalis | 168
Amphotericin B | 168
fluconazole | 168
voriconazole | 168
micafungin | 168
deranged renal parameters | 168
liver function test | 168
coagulation profile | 168
anuric | 168
metabolic acidosis | 168
renal replacement therapy | 168
bradycardia | 168
asystole | 168
death | 168
sepsis | 168
septic shock | 168
multiorgan dysfunction | 168
community-acquired pneumonia | 168
nocardiosis | 168
scrub typhus | 168
candidemia | 168