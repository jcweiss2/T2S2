65 years old | 0
male | 0
admitted to the hospital | 0
hypertension | -4320
benign prostate hyperplasia | -8760
high-grade fever | -240
nausea | -240
vomiting | -240
generalized weakness | -240
intermittent high-grade fever | -720
loss of weight | -720
night-sweats | -720
conscious | 0
well-built | 0
oriented | 0
lethargic | 0
febrile | 0
mild hepatosplenomegaly | 0
conjunctival pallor | 0
hepatosplenomegaly | 0
fatty liver | 0
mild urinary bladder wall thickening | 0
mild cystitis | 0
microcytic hypochromic anemia | 48
leukocytopenia | 48
bicytopenia | 48
raised liver transaminases | 48
total bilirubin | 48
serum triglyceride | 48
plasma fibrinogen | 48
hemoglobin | 48
absolute neutrophil count | 48
total platelet count | 48
serology tests | 48
bone marrow and trephine biopsies | 192
erythroid hyperplasia | 192
megaloblastic erythropoiesis | 192
erythroid and lymphophagocytosis | 192
lactate dehydrogenase | 192
hyperferritinemia | 192
hyponatremia | 192
decreased total protein | 192
MTB | 192
Rifampicin | 192
CECT thorax and abdomen | 192
mild hepatomegaly | 192
prostatomegaly | 192
PET Scan | 192
hepatomegaly | 192
external iliac lymphadenopathy | 192
disseminated tuberculosis | 192
fever | 360
hypertriglyceridemia | 360
pancytopenia | 360
hemophagocytosis | 360
hyperferritinemia | 360
supportive measures | 360
broad-spectrum intravenous antibiotics | 360
transfused with PRBC | 360
modified Anti-Tubercular Treatment | 360
methylprednisolone | 360
Intravenous Immunoglobulin | 360
breathlessness | 384
SpO2 | 384
intensive care unit | 384
hemoglobin | 384
leukocytopenia | 384
total platelet count | 384
Urea | 384
LDH | 384
AST | 384
creatinine | 384
ALT | 384
status epilepticus | 384
poor Glasgow Coma Scale | 384
intubated | 384
declared dead | 480