35 years old | 0
female | 0
morbidly obese | 0
alcohol use disorder | 0
admitted to the hospital | 0
decreased urine output | 0
anasarca | 0
alcoholic cirrhosis | 0
acute kidney injury | 0
liver dysfunction | 0
MELD score of 32 | 0
shock | 0
transfer to the medical intensive care unit | 0
initiation of hemodialysis | 0
initiation of vasopressors | 0
initiation of broad-spectrum antibiotics | 0
weaned off vasopressors | 504
purpuric plaques on the bilateral lower extremities | 504
retiform purpuric plaques with central necrotic eschar | 504
indurated stellate red-brown plaques | 504
peau d'orange on the abdomen | 504
normal calcium | 504
hypoalbuminemia | 504
low phosphorus | 504
excisional biopsy | 504
calcification within small vessels | 504
fat necrosis | 504
calciphylaxis | 504
treatment with intravenous sodium thiosulfate | 504
treatment with vitamin K | 504
treatment with pentoxifylline | 504
treatment with zoledronic acid | 504
medical maggot therapy | 504
application of pathogen-free maggot larvae | 504
maggot therapy for wound debridement | 504
debridement of necrotic tissue | 528
serosanguinous oozing | 528
removal of maggots | 528
debridement including a 3-cm-deep concavity | 528
palpably hollowed eschar | 528
massive hemorrhage from a site of debridement | 552
hemorrhagic shock | 552
transfusion of 8 units of blood | 552
discontinuation of subcutaneous heparin | 552
intermittent bleeding from deep wounds | 552
control of bleeding with pressure dressings | 552
improvement of skin | 1008
no new lesions | 1008
softening of indurated plaques | 1008
recovery of renal function | 1008
discontinuation of hemodialysis | 1008
placement of a percutaneous gastrostomy tube | 1344
pneumoperitoneum | 1344
septic shock | 1344
death | 1344