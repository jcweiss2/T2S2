28 years old|0
male|0
African American|0
multiple sclerosis|-4320
admitted to medical telemetry|0
elevated white blood cell count|0
elevated creatinine kinase|0
lactate|0
no evidence of acute infiltrate or consolidation|0
scattered hypodensities|0
started on broad spectrum antibiotics|0
vancomycin|0
piperacillin/tazobactam|0
levetiracetum|0
acetaminophen|0
gram positive cocci in clusters|48
Staphylococcus pettenkoferi|72
no evidence of valvular vegetations or regurgitation|48
multiple nonconvulsive focal seizures|48
levetiracetum 500 mg twice a day|48
vancomycin|48
ceftriaxone|48
continued to spike fevers|96
no growth|48
no growth|72
transoesophageal echocardiogram|96
no evidence of valvular vegetations|96
micro-perforations|96
trace to mild aortic regurgitation|96
no surgical intervention|96
magnetic resonance imaging|120
numerous white matter lesions|120
clinically monitor off antibiotics|120
levetiracetum 1500 mg BID|120
lacosamide 100 mg BID|120
septic shock|-4320
CoNS bacteremia|-4320
treated empirically with broad spectrum antibiotics|-4320
negative TTE|-4320
lumbar puncture|-4320
no infectious etiology|-4320
discharged|-4320
steroids|-4320
multiple sclerosis flare|-4320
demyelinating lesions|-4320
discontinued antibiotics|-4320
negative blood cultures|-4320
discharged|0
primary care follow up|0
neurology follow up|0
fevers|0
CoNS bacteremia|0
new valvular regurgitation|96
perforations|96
possible endocarditis|96
no risk factors|0
no intravenous drug abuse|0
no poor dental health|0
no long term intravenous indwelling catheters|0
mild aortic regurgitation|96
no signs of CHF|96
no symptoms of CHF|96
same CoNS species|-4320
no prolonged antibiotic course|-4320
negative culture data|-4320
no valvular hardware|0
extremely rare|0
limited TTE|-4320
treated for CoNS bacteremia|-4320
TEE|96
aortic valve perforations|96
regurgitation|96
endocarditis|96
emerging organisms|0
clinical suspicion|0
recognizing CoNS|0
possible causative bacterium|0
TEE as sensitive imaging modality|0
