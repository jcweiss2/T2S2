17 days old | 0
female | 0
premature | 0
admitted to the NICU | 0
failure to thrive | 0
severe metabolic derangements | 0
severe diarrhea | 0
intractable diarrhea | 0
African American | 0
34 5/7 weeks gestation | 0
vaginal delivery | 0
Penta screen abnormal | -672
meconium-stained amniotic fluid | -672
rupture of membranes for 5 hours | -672
Apgar scores 8 and 9 | -672
birthweight 2.445 kg | -672
length 47 cm | -672
head circumference 34 cm | -672
intubated for surfactant administration | -672
extubated to nasal continuous positive airway pressure | -672
treated with ampicillin and gentamicin | -672
diagnosis of clinical sepsis | -672
started on feeds of breastmilk via orogastric tube | -672
developed extensive watery diarrhea | -240
down 25% from birthweight | -240
metabolic acidosis | -240
acute kidney injury | -240
electrolyte derangements | -240
hypernatremia | -240
hyperkalemia | -240
hyperchloremia | -240
hyperglycemia | -240
unconjugated hyperbilirubinemia | -240
started on phototherapy | -240
leukocytosis | -240
I:T ratio of 0.10 | -240
made NPO | -240
electrolyte abnormalities corrected | -240
stool studies sent | -240
campylobacter antigen positive | -240
treated with azithromycin | -240
mother's breastmilk sent for microbial studies | -240
coagulase negative staph positive | -240
E. coli positive | -240
blood cultures negative | -240
started on various feeding regimens | -168
relapse of profuse diarrhea | -168
electrolyte derangements | -168
cessation of enteral feeds | -168
transferred to our institution | 0
receiving TPN with SMOFlipid | 0
signs of moderate dehydration | 0
sunken eyes | 0
dry skin | 0
capillary refill about 4 s | 0
loose stools | 0
infectious disease and gastrointestinal consults | 0
stool studies negative | 0
full sepsis work-up negative | 0
maternal HIV testing negative | 0
GI pathogen PCR panel negative | 0
stool positive for abundant leukocytes and occult blood | 0
stool and blood cultures negative | 0
stool osmotic gap 30 mOsm/kg | 0
newborn screen results positive for glucose-6-phosphate dehydrogenase deficiency | 0
worsening unconjugated hyperbilirubinemia | 24
TPN-induced cholestasis | 24
diarrhea despite strict NPO | 24
secretory diarrhea suspected | 24
EGD and flexible sigmoidoscopy visually normal | 48
duodenal biopsy showed well-preserved enterocytes | 48
electrolyte abnormalities | 48
hyponatremia | 48
hypochloremia | 48
stool sodium and chloride significantly increased | 48
urine sodium and chloride decreased | 48
started on trophic feeds with Enfalyte | 72
advanced to amino acid-based formula | 72
relapse of severe diarrhea | 120
congenital secretory diarrhea genetic panel positive | 120
homozygous mutation for MYO5B c.1462del | 120
diagnosed with MVID | 120
treatment with IV nutritional support | 120
correction of electrolyte imbalance | 120
transferred to a bowel transplant center | 168
transferred back to our institution | 240
maintained on intravenous TPN | 240
awaiting bowel transplant | 240
nephrocalcinosis developed | 240
attributed to dehydration | 240
managed with fluids | 240