63 years old | 0
woman | 0
admitted to the Emergency Department | 0
fever (T 39°C) lasting for 10 days | -240
diarrhea | -240
wet | 0
confused | 0
febrile (T 40°C) | 0
heart rate 121 bpm | 0
blood pressure 85/50 mmHg | 0
SpO2 95% | 0
fluid challenge with normal saline | 0
leukopenia (2190/mm3) | 0
low neutrophil count (1690/mm3) | 0
low lymphocyte count (440/mm3) | 0
thrombocytopenia (33000/mm3) | 0
high C-reactive protein (157 mg/L) | 0
high D-dimers (65.588 FEUng/mL) | 0
high lactic dehydrogenase (1098 mmol/l) | 0
mild renal insufficiency (1.41 mg/dl) | 0
unremarkable arterial gas analysis | 0
positive serology testing (IgG+, IgM-) for SARS-CoV-2 | 0
negative nasopharyngeal swab test | 0
diffuse pulmonary basal lobe opacifications on CT scan | 0
blood cultures obtained | 0
urine cultures obtained | 0
empiric antibiotic therapy with meropenem | 0
empiric antibiotic therapy with gentamycin | 0
admitted to COVID-19 ICU | 0
no subsequent repeated nasopharyngeal swabs confirmed active COVID-19 | 0
no gastric tube samples confirmed active COVID-19 | 0
further decrease in leukocytes during ICU stay | 24
further decrease in platelets during ICU stay | 24
diffuse intravascular coagulation (DIC) | 24
blood transfusions required | 24
fresh frozen plasma transfusions required | 24
negative microbiological cultures | 24
no septic foci found | 24
bone marrow aspirate excluded acute leukemia | 24
sedated after two days from ICU admission | 48
intubated after two days from ICU admission | 48
mechanical ventilation after two days from ICU admission | 48
worsening clinical conditions | 48
incoming multiorgan failure | 48
extubated three days later | 96
mental confusion after extubation | 96
unresponsiveness to external stimuli after extubation | 96
EEG showing non-convulsive status epilepticus (NCSE) | 96
diffuse slow background activity on EEG | 96
epileptiform discharges on EEG | 96
status epilepticus severity scale (STESS) rating 3 | 96
ineffective benzodiazepine I.V. bolus | 96
started I.V. levetiracetam (3000 mg daily) | 96
SE resolution after two days | 168
normal cerebral spinal fluid (CSF) examination | 96
negative CSF for neurotropic viruses | 96
unremarkable brain MRI | 96
remained in ICU for 11 days | 264
transferred to Internal Medicine Unit | 264
discharged home after 20 days | 480
no neurological sequelae at discharge | 480
referred to ED 11 days later | 504
worsening mental slowing | 504
aphasia | 504
afebrile | 504
no other symptoms | 504
motor seizure during ED stay | 504
right upper limb jerks | 504
bilateral tonic-clonic seizure | 504
confused | 504
partially oriented | 504
hypertonic left lower limb | 504
hyposthenic left lower limb | 504
unremarkable laboratory tests | 504
unremarkable brain CT scan | 504
EEG showing sub-continuous epileptiform discharges | 504
focal convulsive SE diagnosis | 504
STESS rating 5 | 504
admitted to Neurology Unit | 504
new brain MRI showing DWI signal alterations | 504
right occipitoparietal signal alterations | 504
bilateral frontoparietal paramedian signal alterations | 504
cortical distribution | 504
no gadolinium enhancement | 504
second CSF examination normal | 504
negative PCR for SARS-CoV-2 | 504
negative PCR for neurotropic viruses | 504
negative autoimmune panel for encephalitis | 504
persistent positive serology (IgG+, IgM-) | 504
negative nasopharyngeal swab | 504
mildly increased IL-6 | 504
mildly increased IL-8 | 504
negative whole-body PET-CT scan | 504
lacosamide 200 mg bid started | 504
motor signs ceased | 504
persistent confusion | 504
psychiatric symptoms appeared | 504
behavioral disturbances | 504
persecutory ideation | 504
aggressiveness | 504
levetiracetam withdrawn | 504
valproic acid (30 mg/kg/day) started | 504
dexamethasone (16 mg/day) started | 504
clinical improvement after six days | 600
SE resolution on EEG | 600
control brain MRI negative | 816
discharged home after 34 days | 816
alert | 816
oriented | 816
able to follow commands | 816
compliant | 816
no focal neurological deficits | 816
repetitive | 816
fatuous | 816
lacosamide 200 mg bid continued | 816
valproic acid 1250 mg daily continued | 816
slightly improved after 45 days | 1296
no further seizures | 1296
EEG showing mild diffuse slowing | 1296
no epileptiform activity | 1296
