39 years old | 0
female | 0
admitted for elective cardiac surgery | -24
cadaveric renal transplant | -8760
renal transplant failed | -6720
chronic vesicoureteral reflux | 0
chronic end-stage renal disease | 0
on chronic renal dialysis | 0
secondary hyperparathyroidism | 0
secondary arterial hypertension | 0
chronic anaemia | 0
iron supplements | 0
atorvastatin | 0
aspirin | 0
amlodipine | 0
erythropoietin | 0
vitamin D supplements | 0
worsening dyspnoea | -432
malnourished and cachectic | 0
diastolic murmur | 0
bibasal lung crepitations | 0
severe mitral stenosis | 0
severely calcified mitral annulus | 0
sub-valvular apparatus | 0
mean gradient of 10 mmHg | 0
mitral valve area of 0.8 cm2 | 0
severe tricuspid regurgitation | 0
preserved biventricular ejection fraction | 0
coronary angiography | 0
no flow-limiting coronary lesions | 0
urea 111 | 0
creatinine 4.7 | 0
phosphorus 10 | 0
calcium 8.6 | 0
parathormone hormone 725 | 0
mitral valve replacement | 0
mechanical prosthesis | 0
tricuspid valve repair | 0
annuloplasty ring | 0
transfusion of multiple blood products | 0
coagulopathy | 0
bleeding | 0
cardiopulmonary bypass | 0
intensive care unit | 0
renal replacement therapy | 0
extubated | 48
warfarin therapy | 72
transferred to the floor | 96
develop skin lesions | 168
necrotic ulcers | 168
fingertips | 168
thigh | 168
calciphylaxis | 168
tissue biopsies | 168
abundant deposition of calcium | 168
necrotic changes | 168
histopathological diagnosis | 168
conservative treatment | 168
enzymatic debridement | 168
collagenase-based ointment | 168
frequent dressings | 168
empirical prophylactic antibiotics | 168
transferred to local district hospital | 456
worsening wound infection | 1080
sepsis | 1080
deceased | 1080