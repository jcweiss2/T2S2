7-day-old | 0
female | 0
newborn | 0
admitted to the Department of Neonatology | 0
poor feeding | -24
bloody stools | -24
loss of consciousness | -24
cesarean section | -168
antenatal period uncomplicated | -168
no history suggestive of infections in the mother | -168
birth weight 3300g | -168
temperature 35.6°C | 0
heart rate 170 beats per minute | 0
respiratory rate 65 times per minute | 0
capillary refill time >3 seconds | 0
blood pressure 35/23mmHg | 0
unresponsive | 0
dry mucous membranes | 0
diminished pulses | 0
mottled cold extremities | 0
decreased urine output | 0
abdominal distention | 0
no abdominal wall cellulitis | 0
white blood cell count 38.51×10^9/L | 0
polymorphonuclear cells 49% | 0
lymphocytes 38.8% | 0
monocytes 12.2% | 0
hemoglobin 14.6g/dL | 0
platelet count 279×10^9/L | 0
C-reactive protein 37mg/L | 0
prothrombin time 16.2 sec | 0
activated partial thromboplastin time 34 sec | 0
necrotizing enterocolitis confirmed | 0
pneumatosis intestinalis | 0
portal venous gas | 0
ascitic fluid examination | 6
WBC count 2815×10^6/L | 6
polymorphonuclear cells 56% | 6
lymphocytes 15% | 6
monocytes/macrophages 29% | 6
red blood cell count 55×10^6/L | 6
blood culture collected | 0
fecal culture collected | 0
no bacterial growth | 0
normal saline administered | 0
dopamine administered | 0
empiric antibiotic therapy started | 0
ceftazidime administered | 0
penicillin G sodium administered | 0
abdominal distension increased | 2
soy sauce-colored urine | 2
jaundice | 2
hemoglobin concentration decreased | 2
direct antiglobulin test negative | 2
acid elution results negative | 2
red blood cells transfused | 2
blood potassium 8.7mmol/L | 2
premature ventricular contractions | 2
continuous renal replacement therapy initiated | 2
vancomycin administered | 2
meropenem administered | 2
antibiotics for meningitis administered | 2
coagulation tests abnormal | 13
fibrin degradation products increased | 13
D-Dimer increased | 13
disseminated intravascular coagulation | 13
clinical metagenomic next-generation sequencing positive for C. perfringens | 13
explorative laparotomy not performed | 13
patient died | 48
C. perfringens infection | 0
massive intravascular hemolysis | 0
septic shock | 0
organ failure | 0
renal failure | 0
acute kidney failure | 0
hyperkalemia | 0
multiple organ failure | 48