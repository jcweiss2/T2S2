43 years old|0
male|0
admitted to the Emergency Department|0
fever|-48
sneezing|-48
fatigue|-48
sore throat|-48
dry cough|-48
no dyspnea|-48
mild cognitive impairment since birth|0
arterial hypertension|0
systemic lupus erythematosus|0
lupus nephritis|0
mycophenolate|0
prednisone|0
family history negative for cancer|0
family history negative for endocrinopathy|0
family history negative for inflammatory diseases|0
parents dead|0
no children|0
fever (38 °C)|0
oxygen saturation 94% in room air|0
respiratory rate 18 breaths/min|0
chest auscultation decreased breath sounds|0
chest auscultation coarse crackles in both lung bases|0
white blood cell count 7110/μL|0
mild lymphocytopenia 650/μL|0
D-dimer 0.73 μg/ml|0
C-reactive protein 62 mg/L|0
PCT 94 ng/mL|0
hemoglobin within normal limits|0
platelets within normal limits|0
serum electrolytes within normal limits|0
creatinine within normal limits|0
liver function test results within normal limits|0
arterial blood gas analysis pH 7.44|0
arterial blood gas analysis pO2 75 mm Hg|0
arterial blood gas analysis pCO2 37 mm Hg|0
SARS-CoV-2 RNA positivity|0
chest computed tomography bilateral ground-glass opacities|0
hyperdense and irregular foci in thoracic vertebral bodies|0
diagnosis of SARS-CoV-2 pneumonia|0
empirical antibiotic therapy with piperacillin/tazobactam|0
oxygen support|0
hospital day 12 general condition improved|288
C-reactive protein normalized 3.5 mg/L|288
blood culture tests negative|288
urine culture tests negative|288
serum PCT remained elevated 84 ng/mL|288
serum CTN 2120 pg/mL|288
carcinoembryonic antigen 108 ng/mL|288
total calcium 9.3 mg/dL|288
ionized calcium 1.21 mmol/L|288
thyrotropin 1.29 μU/mL|288
thyroxine 13.2 pg/mL|288
right laterocervical swelling|288
neck ultrasound inhomogeneously echogenic lymph nodes|288
neck ultrasound small punctate calcifications|288
neck ultrasound nonhomogeneous thyroid with multiple nodules|288
largest thyroid nodule diameter 30 mm|288
fine-needle aspiration|288
diagnosis of MTC|288
CTN in aspiration needle washout fluid >2000 pg/mL|288
PCT:CTN ratio 3.96|288
neck computed tomography scan negative for lesions|288
lung computed tomography scan negative for lesions|288
abdomen computed tomography scan negative for lesions|288
multiple sclerotic lesions dorsal spine level|288
multiple sclerotic lesions hip bone level|288
fluorine-18 fluorodeoxyglucose PET/CT increased tracer uptake right laterocervical lymph nodes|288
fluorine-18 fluorodeoxyglucose PET/CT slight tracer uptake thyroid|288
fluorine-18 fluorodeoxyglucose PET/CT slight tracer uptake dorsal vertebral bodies|288
total thyroidectomy|288
bilateral cervical lymph node dissection|288
histologic examination confirmed MTC|288
neoplastic cells positive for CTN|288
neoplastic cells positive for carcinoembryonic antigen|288
neoplastic cells positive for synaptophysin|288
neoplastic cells positive for chromogranin A|288
neoplastic cells positive for thyroglobulin|288
MTC metastases in 3 of 12 lymph nodes|288
largest lymph node metastasis 30 mm|288
MTC classified as T1b-N1a, stage III|288
blood tests 48 hours post-surgery CTN 986 pg/mL|336
blood tests 48 hours post-surgery PCT 16 ng/mL|336
hospital day 22 SARS-CoV-2 swabs negative|528
discharged|528
prednisone 5 mg/die|528
ramipril 10 mg/die|528
levothyroxine 50 μg/die|528
cholecalciferol 800 IU/die|528
calcium carbonate 1 g/die|528
6-month follow-up scheduled|Approx. 4320 (6 months)
(18)F-fluorodihydro-xyphenylalanine PET no thyroid lodge fixation|Approx. 4320
(18)F4 fluorodihydro-xyphenylalanine PET no cervical lymph node fixation|Approx. 4320
multiple osteoblastic foci dorsal vertebral metameres|Approx. 4320
multiple osteoblastic foci sternum|Approx. 4320
multiple osteoblastic foci right scapula|Approx. 4320
CTN 921 pg/mL|Approx. 4320
PCT 16 ng/mL|Approx. 4320
RET gene analysis planned|Approx. 4320
