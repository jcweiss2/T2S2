18 years old | 0
male | 0
admitted to the hospital | 0
fever | 0
cough | 0
fatigue | 0
dyspnea | 0
anorexia | 0
diarrhea | 0
vomiting | 0
abdominal pain | 0
GI symptoms | 0
abdominal CT performed | 0
ultrasonography performed | 0
ground-glass opacities at the base of the lungs | 0
GI abnormalities on CT | 0
sepsis | 0
abdominal distention | 0
GI bleeding | 0
ischemic bowel disease | 0
hypercoagulable state | 0
contrast-enhanced abdominopelvic CT | 0
abnormal liver function tests | 0
contrast-enhanced ultrasonography | 0
capillary perfusion of abdominal organs | 0
imminent kidney failure | 0
contrast-enhanced fluid-filled colon | 0
luminal distention | 0
bowel wall thickening | 0
mucosal hyperenhancement | 0
peri enteric fat stranding | 0
mesenteric inflammation | 0
vascular engorgement | 0
pneumatosis | 0
portal venous gas | 0
acute pan colitis | 0
subpleural patchy air space opacity | 0
diffuse concentric mural thickening | 0
submucosal edema of the colon | 0
adjacent pericolic fat stranding | 0
mild free fluid in the peritoneal cavity | 0
pneumoperitoneum | 0
acute diverticulitis | 0
ileus | 0
GI perforation | 0
notable ascites | 0
intramural bowel gas | 0
mesenteric ischemia | 0
periportal edema | 0
hematomas at retroperitoneum | 0
abdominal wall hematoma | 0
rectosigmoid hematoma | 0
small bowel obstruction | 0
cecal wall thickening | 0
ileocolonic intussusception | 0
ileocolic intussusception | 0
acute appendicitis | 0
multisystem inflammatory syndrome in children | 0
Kawasaki-like presentations | 0
mucocutaneous symptoms | 0
non-compressible appendix | 0
dilated appendix | 0
mural hyperemia | 0
periappendiceal mesenteric fat stranding | 0
periappendiceal edema | 0
ascites | 0
thickened terminal ileum | 0
luminal dilatation | 0
wall thickening of the appendix | 0
wall thickening of the colon | 0
calcified deposit within the appendix | 0
pelvic free fluid | 0
enlarged lymph nodes | 0
appendiceal perforation | 0
small rim-enhancing fluid collections | 0
thromboembolic complications | 0
endothelial damage | 0
hypercoagulation | 0
microvascular involvement | 0
end-organ ischemia | 0
bowel loops ischemia | 0
spleen infarction | 0
kidneys infarction | 0
liver infarction | 0
superior mesenteric artery thrombotic occlusion | 0
intestinal gangrene | 0
dilated ileal loops | 0
non-enhancing bowel walls | 0
deep venous thrombosis | 0
acute pulmonary thromboembolism | 0
acute myocardial infarction | 0
CT angiography performed | 0
non-occlusive AMI | 0
thrombosis of distal SMA branches | 0
thromboembolic occlusion of SMA | 0
decreased peristalsis | 0
interloop fluid | 0
increased intraluminal contents | 0
stasis | 0
SMV thrombosis | 0
filling defect in the SMV | 0
diffuse small bowel wall thickening | 0
mesenteric fat stranding | 0
mesenteric venous congestion | 0
intra-abdominal hemorrhage | 0
extraperitoneal hematoma | 0
intramuscular hematoma | 0
iliopsoas hematoma | 0
rectus sheath hematoma | 0
active bleeding | 0
hyperdense fresh hematoma | 0
fluid-fluid level formation | 0
pelvic extraperitoneal hemorrhage | 0
centers of active bleeding | 0
massive right iliopsoas muscle hematoma | 0
extravasation extending to the retroperitoneal area | 0
small low-density area in the left iliopsoas muscle | 0
spontaneous iliopsoas muscle hematoma | 0
