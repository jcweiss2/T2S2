48 years old | 0 | 0 
male | 0 | 0 
admitted to the hospital | 0 | 0 
toothache | -96 | 0 
dyspnea | -96 | 0 
chest pain | -96 | 0 
sweating | -96 | 0 
tachyarrhythmia | -96 | 0 
sore throat | -96 | 0 
fever | -96 | 0 
gross swelling of the lower right cheek | 0 | 0 
submandibular and mental regions were erythematous and warm on palpation | 0 | 0 
difficulties in opening the jaw | 0 | 0 
inflammatory changes of the mucous membrane of his oral cavity | 0 | 0 
treated at home with ceftriaxone-steroids-based | -96 | 0 
ineffective treatment | -48 | 0 
worsened condition | -48 | 0 
dyspnea | -48 | 0 
chest pain | -48 | 0 
increase in the amount of white blood cells | 0 | 0 
neutrophils | 0 | 0 
C-reactive protein | 0 | 0 
orotracheal intubation | 0 | 0 
left pleural effusion | 0 | 0 
mediastinitis | 0 | 0 
right parapharyngeal abscess | 0 | 0 
drainage of the right neck | 0 | 0 
left chest drain | 0 | 0 
intravenous antibiotic therapy | 0 | 0 
piperacillin sodium plus tazobactam sodium | 0 | 48 
worsened clinical condition | 48 | 48 
transferred to an Intensive Care Unit | 48 | 48 
air collection in the right submandibular | 48 | 48 
air collection in the left carotid | 48 | 48 
air collection in the retroesophageal and pretracheal spaces | 48 | 48 
cervical necrotizing fasciitis with DNM | 48 | 48 
bilateral pleural effusions | 48 | 48 
additive pleural drain | 72 | 72 
abscesses in the cervical spaces | 72 | 72 
extensive mediastinal empyema | 72 | 72 
left pleural effusion | 72 | 72 
right hydropneumothorax | 72 | 72 
aggressive mediastinal debridement | 72 | 72 
VATS | 72 | 72 
incision and drainage of the neck abscesses | 72 | 72 
oral tooth extraction | 72 | 72 
purulent fluid in the cavity below was drained and packed | 72 | 72 
Streptococcus anginosus | 72 | 72 
Gemella morbillorum | 72 | 72 
Staphylococcus lugdunensis | 72 | 72 
antibiotic therapy | 72 | 168 
Amoxicillin | 72 | 168 
Metronidazole | 72 | 168 
dismissed in better health conditions | 168 | 168