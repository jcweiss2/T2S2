38 years old | 0
female | 0
admitted to the hospital | 0
septic shock | 0
streptococcal necrotising fasciitis | 0
thoracic trauma | -48
amoxicilline | 0
clindamycine | 0
linezolid | 0
infection spread | 0
pneumothorax | 0
Stenotrophomonas maltophilia | 0
Citrobacter spp. | 0
Aspergillus spp. | 0
Mucor spp. | 0
liposomal amphotericin B | 9
HBOT therapy | 9
Enterococcus faecium | 9
Enterobacter gallinarum | 9
Pseudomonas aeruginosa | 9
Citrobacter sedlakii | 9
Stenotrophomonas maltophilia | 9
Candida albicans | 9
Aspergilus fumigatus | 9
Aspergilus terreus | 9
mucormycosis | 11
Lichtheimia ramosa | 11
Rhizopus arrhizus | 11
cefepime | 11
ciprofloxacine | 11
sulfamethoxazole-trimethoprime | 11
metronidazole | 11
pozaconazole | 11
isavuconazole | 11
monocyte deactivation | 11
IFN-γ | 11
nivolumab | 27
PD-1 expression | 27
T lymphocyte PD-1 expression | 27
tissue culture negative | 28
PCR negative | 34
RRT weaning | 39
extubation | 43
reconstructive surgery | 52
skin grafting | 52
discharged | 1320