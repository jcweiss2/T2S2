76 years old | 0
    woman | 0
    subjective fevers | 0
    nonproductive cough | 0
    dyspnea | 0
    admitted to the intensive care unit | 0
    acute hypoxic respiratory failure | 0
    COVID-19 infection | 0
    blood pressure 110/53 mm Hg | 0
    pulse rate 124 beats/min | 0
    respiratory rate 31 breaths/min | 0
    oxygen saturation 79% | 0
    temperature 102.3°F | 0
    severe respiratory distress | 0
    tachycardia | 0
    diffusely decreased breath sounds | 0
    crackles | 0
    hypertension | 0
    hyperlipidemia | 0
    hypothyroidism | 0
    acute dyspnea | 0
    hypoxia | 0
    COVID-19-induced acute respiratory distress syndrome | 0
    acute pulmonary embolism | 0
    acute heart failure | 0
    septic shock | 0
    cardiac tamponade | 0
    acute coronary syndrome | 0
    viral pneumonia | 0
    bacterial pneumonia | 0
    viral cardiomyopathy | 0
    potassium 2.2 mEQ/L | 0
    creatinine 1.79 mg/dL | 0
    C-reactive protein 23.10 mg/L | 0
    interleukin-6 781.46 mg/L | 0
    lactate dehydrogenase 334 U/L | 0
    ferritin 457 ng/mL | 0
    procalcitonin 15.20 ng/mL | 0
    prothrombin time 18.9 seconds | 0
    fibrinogen >600 mg/dL | 0
    white blood cell count 16.1 cells/L | 0
    92.7% neutrophils | 0
    IgG 1622 mg/dL | 0
    SARS-CoV-2 positive | 0
    troponin 0.03 ng/dL | 0
    high-sensitivity troponin peaked at 503 ng/L | 0
    proBNP 35,000 pg/mL | 0
    diffuse bilateral pulmonary edema vs infiltrates | 0
    worsening diffuse bilateral pulmonary opacities/infiltrates vs edema | 0
    electrocardiogram no signs of ischemia | 0
    normal sinus rhythm | 0
    short PR interval 72 ms | 0
    left ventricular hypertrophy | 0
    QTc interval 680 ms | 0
    previous echocardiograms normal LV ejection fraction | 0
    no wall motion abnormalities | 0
    transthoracic echocardiogram severely decreased LV systolic function | 0
    segmental wall motion abnormalities | 0
    akinesis of the distal segments of the left ventricle | 0
    preserved function at the base | 0
    akinesis of the mid and distal portions of the right ventricle | 0
    preserved function at the base of the free wall | 0
    ejection fraction 25%-30% | 0
    intubated | 0
    limited bedside TTE normal cardiac EF 55% | 0
    shock state | 0
    vasopressor support with norepinephrine | 0
    ARDSnet protocol | 0
    treated with tocilizumab 480 mg | 0
    treated with tocilizumab 240 mg | 0
    intravenous immunoglobulin 25 g for 5 days | 0
    ceftriaxone | 0
    cefdinir | 0
    cefepime | 0
    cytokine storm | 0
    leukocytosis | 0
    not treated with hydroxychloroquine | 0
    not treated with azithromycin | 0
    prolonged QTc interval | 0
    worsening bilateral airspace opacities vs vascular congestion | 0
    treated with intravenous furosemide 40 mg | 0
    cardiac enzymes elevated | 0
    repeat bedside TTE LVEF 20%-25% | 0
    severe viral myocarditis | 0
    transferred to a tertiary center | 0
    LVEF 25%-30% | 0
    wall motion abnormalities | 0
    non-ST-elevation myocardial infarction | 0
    viral cardiomyopathy | 0
    treated with therapeutic enoxaparin | 0
    LVEF recovered to 50% | 48
    mildly reduced LV systolic function | 48
    mid-septal and apical hypokinesis | 48
    mildly reduced right ventricular function | 48
    blood cultures negative | 48
    respiratory cultures negative | 48
    inflammatory markers improved | 48
    inflammatory markers worsened again | 48
    IL-6 downtrend from 781.46 mg/L to 171.82 mg/L | 48
    high-sensitivity troponin decreased from 503 ng/L to 418 ng/L | 48
    not candidate for extracorporeal membrane oxygenation | 48
    transferred back to intensive care unit | 48
    SARS-CoV-2-induced myocardial injury | 0
    cytokine storm | 0
    acute myocardial injury | 0
    hemodynamic instability | 0
    shock state | 0
    viral myocarditis | 0
    Takotsubo cardiomyopathy | 0
    therapeutic enoxaparin | 0
    early cardiac biomarkers | 0
    noninvasive imaging | 0
    cardiology involvement | 0
    cardiac complications | 0

    76 years old | 0
    woman | 0
    subjective fevers | 0
    nonproductive cough | 0
    dyspnea |$|$0
    admitted to the intensive care unit | 0
    acute hypoxic respiratory failure | 0
    COVID-19 infection | 0
    blood pressure 110/53 mm Hg | 0
    pulse rate 124 beats/min | 0
    respiratory rate 31 breaths/min | 0
    oxygen saturation 79% | 0
    temperature 102.3°F | 0
    severe respiratory distress | 0
    tachycardia | 0
    diffusely decreased breath sounds | 0
    crackles | 0
    hypertension | 0
    hyperlipidemia | 0
    hypothyroidism | 0
    acute dyspnea | 0
    hypoxia | 0
    COVID-19-induced acute respiratory distress syndrome | 0
    acute pulmonary embolism | 0
    acute heart failure | 0
    septic shock | 0
    cardiac tamponade | 0
    acute coronary syndrome | 0
    viral pneumonia | 0
    bacterial pneumonia | 0
    viral cardiomyopathy | 0
    potassium 2.2 mEQ/L | 0
    creatinine 1.79 mg/dL | 0
    C-reactive protein 23.10 mg/L | 0
    interleukin-6 781.46 mg/L | 0
    lactate dehydrogenase 334 U/L | 0
    ferritin 457 ng/mL | 0
    procalcitonin 15.20 ng/mL | 0
    prothrombin time 18.9 seconds | 0
    fibrinogen >600 mg/dL | 0
    white blood cell count 16.1 cells/L | 0
    92.7% neutrophils | 0
    IgG 1622 mg/dL | 0
    SARS-CoV-2 positive | 0
    troponin 0.03 ng/dL | 0
    high-sensitivity troponin peaked at 503 ng/L | 0
    proBNP 35,000 pg/mL | 0
    diffuse bilateral pulmonary edema vs infiltrates | 0
    worsening diffuse bilateral pulmonary opacities/infiltrates vs edema | 0
    electrocardiogram no signs of ischemia | 0
    normal sinus rhythm | 0
    short PR interval 72 ms | 0
    left ventricular hypertrophy | 0
    QTc interval 680 ms | 0
    previous echocardiograms normal LV ejection fraction | 0
    no wall motion abnormalities | 0
    transthoracic echocardiogram severely decreased LV systolic function | 0
    segmental wall motion abnormalities | 0
    akinesis of the distal segments of the left ventricle | 0
    preserved function at the base | 0
    akinesis of the mid and distal portions of the right ventricle | 0
    preserved function at the base of the free wall | 0
    ejection fraction 25%-30% | 0
    intubated | 0
    limited bedside TTE normal cardiac EF 55% | 0
    shock state | 0
    vasopressor support with norepinephrine | 0
    ARDSnet protocol | 0
    treated with tocilizumab 480 mg | 0
    treated with tocilizumab 240 mg | 0
    intravenous immunoglobulin 25 g for 5 days | 0
    ceftriaxone | 0
    cefdinir | 0
    cefepime | 0
    cytokine storm | 0
    leukocytosis | 0
    not treated with hydroxychloroquine | 0
    not treated with azithromycin | 0
    prolonged QTc interval | 0
    worsening bilateral airspace opacities vs vascular congestion | 0
    treated with intravenous furosemide 40 mg | 0
    cardiac enzymes elevated | 0
    repeat bedside TTE LVEF 20%-25% | 0
    severe viral myocarditis | 0
    transferred to a tertiary center | 0
    LVEF 25%-30% | 0
    wall motion abnormalities | 0
    non-ST-elevation myocardial infarction | 0
    viral cardiomyopathy | 0
    treated with therapeutic enoxaparin | 0
    LVEF recovered to 50% | 48
    mildly reduced LV systolic function | 48
    mid-septal and apical hypokinesis | 48
    mildly reduced right ventricular function | 48
    blood cultures negative | 48
    respiratory cultures negative | 48
    inflammatory markers improved | 48
    inflammatory markers worsened again | 48
    IL-6 downtrend from 781.46 mg/L to 171.82 mg/L | 48
    high-sensitivity troponin decreased from 503 ng/L to 418 ng/L | 48
    not candidate for extracorporeal membrane oxygenation | 48
    transferred back to intensive care unit | 48
    SARS-CoV-2-induced myocardial injury | 0
    cytokine storm | 0
    acute myocardial injury | 0
    hemodynamic instability | 0
    shock state | 0
    viral myocarditis | 0
    Takotsubo cardiomyopathy | 0
    therapeutic enoxaparin | 0
    early cardiac biomarkers | 0
    noninvasive imaging | 0
    cardiology involvement | 0
    cardiac complications | 0