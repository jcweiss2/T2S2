22 years old | 0
female | 0
distant history of alcohol use | -20160
distant history of cocaine use | -20160
presented to the emergency room | 0
one week history of nausea | -168
one week history of vomiting | -168
subjective fevers | -168
myalgias | -168
fatigue | -168
denied chest pain | 0
denied dyspnea | 0
denied cough | 0
no recent illicit substance use | 0
sinus tachycardia of 130 beats/min | 0
temperature of 36.9 degrees Celsius | 0
blood pressure of 75/40 mmHg | 0
oxygen saturations of 90% on room air | 0
elevated jugular venous pressure of 9 cm | 0
heart sounds difficult to hear on auscultation | 0
elevated white blood cell count of 14.4 × 109/L | 0
neutrophil count of 13.0 × 109/L | 0
normal cardiac troponin I | 0
normal creatinine | 0
normal electrolytes | 0
normal beta-HCG | 0
urine toxicology negative for illicit drugs | 0
electrocardiogram showed sinus tachycardia | 0
small voltages in the limb leads | 0
chest X-ray showed generous sized cardiac silhouette | 0
clear lung fields | 0
admitted into the intensive care unit | 0
given fluids | 0
ionotropic support with norepherine | 0
pipericillin-tazobactam started | 0
vancomycin started | 0
blood cultures drawn | 0
nasopharyngeal swab conducted | 0
positive for Influenza A H1N1 | 0
oseltamivir initiated | 0
remained hypotensive | 0
echocardiogram performed | 24
moderate sized pericardial effusion | 24
maximal diameter of 1.5 cm | 24
right ventricular diastolic collapse | 24
significant respiratory variation on mitral valve annular doppler velocity | 24
urgent pericardiocentesis conducted | 24
improvement of hemodynamic status | 24
withdrawl of all ionotropic support | 24
pericardial drain inserted | 24
repeat echocardiogram two days later | 72
resolution of pericardial effusion | 72
absence of echocardiographic findings of tamponade | 72
pericardial effusion negative for bacterial cultures | 72
pericardial effusion negative for acid fast bacilli | 72
pericardial effusion negative for malignancy | 72
serologic testing for HIV negative | 72
serologic testing for Hepatitis B negative | 72
serologic testing for Hepatitis C negative | 72
high dose ibuprofen initiated | 72
colchicine initiated | 72
pericardial drain removed | 336
repeat echocardiogram within two weeks | 336
no return of pericardial effusion | 336
discharged from the hospital | 336
