31 years old | 0
female | 0
previous cesarean section | -720
second cesarean section | -17
suprapubic abdominal pain | -72
bilateral flank pain | -72
dysuria | -72
nauria | -72
vomiting | -72
diarrhea | -72
afebrile | -72
subjective rigors | -72
chills | -72
hypotension | -72
leukocytosis | -72
elevated serum lactate | -72
intravenous fluid volume resuscitation | 0
empiric broad spectrum intravenous antibiotic therapy | 0
admitted to ICU | 0
sepsis without established source | 0
urologic examination | 0
radiologic examinations | 0
urinalysis | 0
urosepsis | 0
postpartum sepsis | 0
suction dilation & curettage (D&C) | 0
laparoscopic examination | 0
intra-abdominal viscera examination | 0
white blood cell count rose | 24
septic shock worsened | 24
leukemoid reaction | 24
disseminated intravascular coagulation (DIC) | 24
potential infection with Clostridium species | 24
supra-cervical hysterectomy | 48
bilateral salpingectomy | 48
abdominal compartment syndrome | 48
grossly enlarged uterus | 48
acute and chronic endo-myometritis | 48
necrotic features | 48
acute salpingitis | 48
necrotic gynecologic tissue | 48
puerperal septic source | 48
intravenous immunoglobulin (IVIg) | 48
exploratory laparotomy | 120
abdominal washout | 120
vacuum-assisted closure (VAC) device | 120
abdominal washout | 168
Wittmann temporary abdominal fascia Velcro prosthetic patch | 168
wound VAC | 168
exploratory laparotomy | 288
abdominal washout | 288
tightening of Wittmann abdominal fascia patch | 288
wound VAC | 288
abdominal washout | 336
closure of abdominal fascia | 336
white blood cell count normalized | 360
discharged from ICU | 408
discharged from hospital | 600
follow-up in clinic | 720
doing well | 720
toxic shock syndrome | 0
endometritis | 0
sepsis secondary to C. sordellii | 0
tissue samples sent to CDC | 0
microscopic examination of uterine tissue | 504
extensive endometrial necrosis | 504
hemorrhage | 504
fibrin deposition | 504
neutrophilic infiltration | 504
edematous changes | 504
focal granulation tissue | 504
lymphoplasmacytic infiltrate | 504
thrombosed vessels | 504
uterine contents positive for C. sordellii | 504
IHC staining | 504
PCR testing | 504