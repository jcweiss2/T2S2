65 years old | 0
male | 0
hypertension | 0
subarachnoid hemorrhage | 0
external ventricular drain | 0
coiling | 0
admitted to the medical intensive care unit | 0
septic shock | 192
Clostridioides difficile infection | 192
leukocytosis up to 39.5 K/uL | 192
creatinine level of 1.86 mg/dL | 192
vancomycin liquid 125 mg every 6 hours through a nasogastric tube | 192
IV metronidazole 500 mg every 8 hours | 192
worsening sepsis | 288
no improvement in diarrhea | 288
fidaxomicin 200 mg per NG tube twice daily | 288
worsening abdominal pain | 336
distension | 336
acute hypoxemic respiratory failure | 336
mechanical ventilation | 336
computed tomography scan of the abdomen and pelvis with IV and oral contrast | 336
diffuse severe bowel wall thickening in the sigmoid colon and rectum | 336
colonic distension up to 6 cm | 336
toxic megacolon | 336
flexible sigmoidoscopy | 336
extensive pseudomembranes up to 50 cm from the anal verge | 336
laparoscopic loop ileostomy with colonic lavage | 336
IV metronidazole | 336
vancomycin irrigation through Foley catheter in the efferent limb of the loop ileostomy | 336
weaned off vasopressors | 336
persistent diarrhea | 336
fever | 336
leukocytosis | 336
consultation by gastroenterology team | 336
antibiotics held for 24 hours | 360
polyethylene glycol preparation through Foley catheter | 360
donor stool administration through Foley catheter | 384
resolution of leukocytosis | 456
resolution of diarrhea | 456
transferred to general medical floor | 456
discharged to rehabilitation facility | 456
repeat colonoscopy in 6 months | 4320
resolution of CDI | 4320
successful reversal of ileostomy | 4320
