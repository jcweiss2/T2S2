74 years old | 0
female | 0
Japanese | 0
schizophrenia | -720
high-grade fever | -24
unaware of febrile status | -24
no chest pain | -24
no cough | -24
no dyspnea | -24
no palpitation | -24
no urinary complaints | -24
no bowel complaints | -24
no history of tuberculosis | -24
no history of malignancy | -24
no previous hospital admissions | -24
no smoking | -24
no alcohol | -24
no illicit drugs | -24
no recent travel history | -24
admitted to the hospital | 0
fever 39.1°C | 0
pulse rate 110 beats/min | 0
blood pressure 100/60 mmHg | 0
respiratory rate 24 times/min | 0
99% oxygen saturation | 0
level of consciousness E4V4M6 | 0
non-tender mass in the lower right back | -720
mass awareness for 1 month | -720
leukocytosis 23 300 cells/mm3 | 0
polymorphic neutrophil predominance | 0
hemoglobin 8.6 g/dL | 0
platelet count 339 000/mm3 | 0
CPK 125 IU/L | 0
blood urea nitrogen 23.3 mg/dl | 0
creatinine 0.97 mg/dl | 0
C-reactive protein 15.26 mg/dl | 0
blood sugar 116 mg/dl | 0
HbA1c 5.4% | 0
HIV test negative | 0
urinalysis +/− protein | 0
urinalysis 1+ nitrite | 0
urinalysis 2+ leukocyte | 0
urine glucose negative | 0
urine occult blood negative | 0
urine ketones negative | 0
subcutaneous abscess suspected | 0
ultrasound examination | 12
low echoic mass | 12
CT detected large mass | 12
surgical drainage | 24
post-procedural septic shock | 24
M. morganii detected in fluid | 24
M. morganii detected in urine culture | 24
blood cultures negative | 24
repeat CT with intravenous contrast | 48
right renal abscess | 48
staghorn calculus | 48
retroperitoneum abscess improvement | 48
iliopsoas abscess | 48
urinary tract infection | -24
M. morganii infection | -24
meropenem administered | 24
salvage nephrectomy | 72
post-operative recovery | 96
intravenous meropenem | 96
oral levofloxacin | 168
discharged to nursing home | 336