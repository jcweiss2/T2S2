65 years old | 0
male | 0
admitted to the hospital | 0
abdominal pain | -168
abdominal distension | -168
obstipation | -168
discoloration of abdominal skin | -168
liposuction of the abdomen | -168
gastric bypass | -7224
morbid obesity | -7224
tachycardia | 0
tachypnoea | 0
normal blood pressure | 0
subcutaneous emphysema of abdominal skin | 0
blackish discoloration of the abdominal skin | 0
erythema | 0
diffuse tenderness | 0
no rebound tenderness | 0
contrast CT scan of the abdomen | 0
hold up of the contrast in the small intestine | 0
jejunum dilation | 0
proximal ileal loops dilation | 0
no free fluid in the abdomen | 0
specks of air in the abdomen | 0
exploratory laparotomy | 24
dead necrotic abdominal skin excision | 24
subcutaneous tissue excision | 24
anterior rectus sheath healthy | 24
copious seropurulent fluid in the perifascial planes | 24
mid ileal loop kinked | 24
adhered to the duodenojejunal junction | 24
obstruction | 24
obstruction relieved | 24
mid jejunum perforation | 24
perforation repaired | 24
linea alba closed | 24
IV fluids | 24
nasogastric aspiration | 24
total parenteral nutrition | 24
altered sensorium | 288
hyponatremia | 288
sepsis secondary to pneumonia | 288
IV antibiotics | 288
E. Coli growth | 288
Enterococcus growth | 288
Acticoat dressings | 288
wound improved | 336
granulations appeared | 336
soakage reduced | 336
high risk for skin grafting | 336
intermittent fever | 336
persistent tachycardia | 336
allograft application | 336
exudate reduced | 336
dressing changed once daily | 336
autologous skin grafting | 672
graft took up well | 672
uneventful recovery | 672
incisional hernia | 8760
incisional hernia repair | 8760
back to regular activities | 17544
