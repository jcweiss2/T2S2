53 years old | 0
male | 0
admitted to the hospital | 0
altered mental status | 0
hypotension | 0
fever | 0
respiratory distress |,0
diabetic nephropathy | 0
requirement of renal replacement therapy | 0
diabetic retinopathy | 0
bilateral amaurosis | 0
cardiac arrest | 0
acute respiratory failure | 0
cardiopulmonary resuscitation | 0
return to spontaneous blood circulation | 0
orotracheal intubation | 0
normocytic normochromic anemia | 0
mixed hyperbilirubinemia | 0
conserved renal function | 0
no electrolyte disorders | 0
CT angiography negative for pulmonary embolism | 0
positive polymerase chain reaction assay for SARS-CoV-2 | 0
respiratory distress | 0
no vaccination | 0
unknown COVID-19 variant | 0
neurological examination | 0
somnolent | 0
alertable | 0
obeying simple orders | 0
intact brainstem reflexes | 0
normal motor function | 0
normal sensitive function | 0
brain CT showing supratentorial bilateral frontal leukoencephalopathy | 0
calcified atheromatous plaques | 0
deterioration of mental status | 0
stupor | 0
severe hypoglycemia | 0
glucose level of 18 mg/dl | 0
MRI showing symmetric focal high intensity signals | 0
glucose normalization | 0
mental status improvement | 0
multiple comorbidities | 0
worsen respiratory status | 0
end-of-life symptom management order | 0
ESMO protocol implemented | 0
