33 years old | 0
female | 0
African American | 0
admitted to the hospital | 0
history of recurrent progressive metastatic squamous cell carcinoma | -4032
cervical cancer | -4032
initial definitive external pelvic chemoradiation | -4032
chemotherapy weekly with cisplatin | -4032
intracavitary high-dose rate brachytherapy | -4032
recurrent disease in upper abdomen | -672
recurrent disease in iliac bone | -672
sepsis | -672
pancreatitis | -672
small bowel resection | -672
permanent ostomy formation | -672
treated with pembrolizumab | -96
painful hyperpigmented maculopapular rash | -72
blister-like lesions | -72
maculopapular rash on lower back | -72
maculopapular rash on feet | -72
maculopapular rash on forehead | -48
maculopapular rash on trunk | -48
maculopapular rash on thighs | -48
painful blistering of lips | -48
ocular involvement | -48
biopsy | -24
diagnosis of SJS/TEN | -24
apoptotic keratinocytes | -24
lymphocytic infiltration | -24
transfer to local University Burn Intensive Care Unit | 0
moderate distress | 0
desquamative rash | 0
odynophagia | 0
worsening mouth ulcers | 0
Staphylococcus epidermidis sepsis | 0
treated with IV vancomycin | 0
started on solumedrol | 0
improvement in cutaneous symptoms | 24
dermatology consultation | 24
ophthalmology consultation | 24
burn consultation | 24
gynecologic oncology consultation | 24
topical antibiotic ointment | 24
cyclosporine | 24
artificial tears | 24
erythromycin ointment | 24
silverlon dressing | 24
dampened 10-ply gauze | 24
burn net | 24
aggressive nutritional supplementation | 24
protein supplementation | 24
micronutrient supplementation | 24
vitamin C supplementation | 24
weekly nutrition labs | 24
intravaginal betamethasone therapy | 24
estrogen therapy | 24
discontinuation of cyclosporine | 48
initiation of prednisone | 48
improvement of symptoms | 72
tapering of corticosteroid | 72
episode of fever | 120
episode of hypotension | 120
empiric meropenem | 120
empiric vancomycin | 120
blood cultures grew Klebsiella | 120
treated with ciprofloxacin | 120
discharge to home | 168