18 years old | 0
female | 0
history of intravenous drug use | -720
extraction of all maxillary teeth | -600
mandibular dental infection | -480
treated with oral amoxicillin | -480
low grade fevers | -120
sudden deterioration in mental status | -120
admitted to the hospital | 0
altered mental status | 0
fever | 0
chills | 0
chest pain | 0
dyspnea | 0
nausea | 0
vomiting | 0
diarrhea | 0
skin lesions | 0
numbness | 0
tingling | 0
weakness of the lower extremities | 0
prominent holosystolic murmur at the apex | 0
petechial rash | 0
encephalopathy | 0
facial droop | 0
slurred speech | 0
intubated for airway protection | 24
leukocytosis | 24
87.6% neutrophils | 24
platelet count of 17 × 10^9/L | 24
liver and kidney functions were within normal | 24
declined a HIV test | 24
innumerable acute to subacute embolic infarcts in both cerebral and cerebellar hemispheres | 24
proximal right internal carotid artery T-shaped acute thrombus | 24
occlusion of the right middle cerebral artery | 24
subarachnoid hemorrhage in the right parietal region and around the posterior aspect of the midbrain | 24
echo densities on the tricuspid, aortic, and mitral valves | 24
vegetations on the tricuspid, aortic, and mitral valves | 24
blood culture grew S. marcescens | 24
S. marcescens isolate was pansensitive susceptible to ceftriaxone, cefepime, ceftazidime, meropenem, gentamicin, tobramycin, amikacin, ciprofloxacin, and levofloxacin | 24
antibiotic was changed to cefepime | 72
cardiothoracic surgery consulted | 72
poor candidate for surgery due to deterioration in neurological status | 72
neurological status continued to deteriorate | 120
no cough or gag reflex | 120
pupils were fixed and mid-dilated | 120
family decided to withdraw care | 120
discharged to hospice care | 120