59 years old | 0
man | 0
admitted to the hospital | 0
large symptomatic anterior mediastinal mass | 0
progressively more short of breath | -8760
significantly decreased exercise tolerance | -8760
intermittent fevers | -8760
leukocytosis | -8760
evaluated in Pakistan by a cardiologist | -8760
echocardiogram | -8760
stress test | -8760
mediastinal and right pleural base mass | -8760
additional radiological imaging | -8760
chest X-ray | -8760
large mass in the right pleural space | -8760
CT scan of the chest | -8760
large inhomogeneous mass | -8760
near total compression of the right atrium | -8760
total compression of the lung | -8760
significant compression atelectasis | -8760
biopsy of the mass | -8760
thymoma | -8760
traveled to the United States | 0
persistent right pleural based mass | 0
compression of the right atrium | 0
compression of the right lung | 0
pathology slides reviewed by two separate institutions | 0
diagnosis confirmed to be thymoma | 0
discussion regarding treatment options | 0
elected to undergo surgical resection | 0
pre-operative evaluation | 0
febrile to 103° | 0
significant leukocytosis of 30,000 | 0
admitted to the thoracic surgery service | 0
chest X-ray | 0
large right pleural mass | 0
repeat transthoracic echocardiogram | 0
normal ventricular function | 0
no vegetations | 0
continued compression of the right atrium | 0
Duplex ultrasound of the lower extremities | 0
no deep venous thromboses | 0
blood cultures | 0
urine cultures | 0
negative cultures | 0
hematology/oncology service consulted | 0
bone marrow biopsy | 0
peripheral smear | 0
negative bone marrow biopsy | 0
negative peripheral smear | 0
Infectious Disease service consulted | 0
started on intravenous antibiotics | 0
intermittent fevers | 0
leukocytosis | 0
compression atelectasis of the right lung | 0
massive tumor necrosis | 0
surgical resection on hospital day 2 | 48
endotracheally intubated | 48
double-lumen endotracheal tube | 48
transesophageal echocardiography | 48
left lateral decubitus position | 48
extended right posterolateral thoracotomy incision | 48
right pleural cavity explored | 48
enormous mass | 48
involved all three lobes of the right lung | 48
mass opened | 48
purulent fluid | 48
necrotic tumor mass | 48
culture sent | 48
frozen section | 48
suspicious for lymphoma | 48
deferred definitive diagnosis | 48
discussion with oncologist | 48
deferred resection | 48
chest tubes placed | 48
wound closed | 48
transferred to cardiothoracic ICU | 48
postoperative day 1 | 72
septic | 72
vasopressor support | 72
aggressive fluid resuscitation | 72
weaned off vasopressors | 96
weaned off ventilator | 48
extubated | 48
transferred to medical/surgical unit | 48
chest tubes | 48
minimal drainage | 48
daily chest X-rays | 48
noticeable improvement in right lung | 48
final pathology | 48
T cells | 48
neoplastic epithelial cells | 48
type B1 thymoma | 48
Salmonella species | 48
non-typhoidal | 48
intravenous antibiotic coverage changed to cefepime | 48
transitioned to oral antibiotics | 240
discharged home on post-operative day 10 | 240
antibiotic therapy | 240
follow-up plan | 240
repeat CT four weeks later | 672
presence of the mass | 672
no significant change in size | 672
doing well | 672
effort-induced shortness of breath | 672
decision for surgical resection | 672
readmitted on March 14, 2013 | 672
right thoracotomy | 672
complete resection of tumor mass | 672
partial right lower lobectomy | 672
echocardiogram intraoperatively | 672
large mass compressing right atrium | 672
specimen completely resected | 672
marked improvement in compression | 672
tolerated procedure well | 672
postoperative course uneventful | 672
intensive care unit for 1 day | 672
transferred to surgical floor | 672
postoperative day 2 | 672
shortness of breath resolved | 672
significant improvement on chest X-ray | 672
chest tube discontinued | 672
sent home on postoperative day 5 | 672
complete 1 week of antibiotic therapy | 672
