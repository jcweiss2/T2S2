49 years old | 0
female | 0
esophageal squamous cell carcinoma | 0
neoadjuvant chemotherapy | 0
minimally invasive Ivor-Lewis esophagectomy | 0
postoperative day 3 | 72
increased inflammatory indexes | 72
CRP 178.2 ng/mL | 72
postoperative day 4 | 96
endoscopy | 96
CT scan | 96
large anastomotic leak | 96
giant wound cavity in the pleural space | 96
fibrosis | 96
abundant necrotic tissue | 96
acute respiratory distress syndrome | 96
sepsis | 96
intensive care | 96
ventilatory support | 96
antibiotic therapy | 96
anastomotic dehiscence | 96
EVAC therapy | 96
Esosponge placement | 96
14 treatment sessions | 96
over 35 days | 96
leak improvement | 96
cavity size improvement | 96
healthy-appearing granulation tissue | 96
inflammatory indexes improvement | 96
clinical conditions improvement | 96
endoscopic findings confirmed by CT scans | 96
no complications observed | 96
after 14th session | 96
endoscopic evaluation | 96
cleaner cavity | 96
smaller cavity (1 cm) | 96
placement of fully covered SEMS | 96
liquid diet | 96
leak healing | 96
stents kept for 3 weeks each | 96
endoscopy after SEMS removal | 96
esophagram after SEMS removal | 96
leak resolution | 96
tiny persistent depression | 96
no symptoms of recurrent fistula formation | 96
over 6 months | 96
