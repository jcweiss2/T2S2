41 years old | 0
female | 0
severe mitral regurgitation | -6 years
mitral valve replacement | -6 years
high profile bioprosthesis size 31 | -6 years
abnormal position of the bio-prosthesis strut | 0
narrowing of the left ventricular outflow tract | 0
mean systolic gradient of 35 mmHg | 0
left ventricular outflow tract obstruction | 0
smallish left ventricular cavity | 0
redo MVR | 0
mechanical valve size 29 Carbomedics | 0
posterior MV leaflet resected | 0
severe calcification | 0
significant bleeding from the chest tubes | 10
hemodinamic instability | 10
surgical re-exploration for bleeding | 10
cardiopulmonary bypass | 10
aortic cross clamp | 10
cardioplegia | 10
left atrium opened | 10
no problem with the new mechanical mitral valve | 10
no tears identified | 10
tear in the posterior wall of the LVOT | 10
repair of the tear | 10
transfer to intensive care unit | 10
stable condition | 10
died | 192
sepsis | 192
disseminated intravascular coagulopathy | 192