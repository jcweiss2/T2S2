43 years old | 0
male | 0
schizophrenia | 0
asthma | 0
polysubstance use disorder | 0
IVDU | 0
admitted to the hospital | 0
fever | 0
chills | 0
left-sided pleuritic chest pain | 0
methicillin-sensitive Staphylococcus aureus TV endocarditis | -2628
paraspinal abscess | -2628
percutaneous drainage | -2628
6 weeks of intravenous antibiotic therapy | -2628
febrile | 0
tachycardic | 0
normotensive | 0
adequate oxygen saturation | 0
intravenous antimicrobial therapy | 0
transthoracic echocardiography | 0
30-mm mobile mass on the TV | 0
vegetation | 0
evaluated by a multidisciplinary heart valve team | 0
care provided by a multispecialty team | 0
psychiatry | 0
specialized social work | 0
7 days of appropriate antimicrobial therapy | 168
continued to be febrile | 168
positive blood cultures | 168
septic pulmonary emboli | 168
tricuspid valve replacement | 168
refused an open surgical procedure | 168
debulk the TV vegetation | 168
percutaneous vacuum-assisted device | 168
consent obtained | 168
general anesthesia | 168
endotracheal tube | 168
left-sided central venous catheter | 168
TEE guidance | 168
vegetation measuring 32 × 26 mm | 168
mild tricuspid regurgitation | 168
right ventricle not dilated | 168
normal systolic function | 168
TV annulus measured at 37 mm | 168
no vegetations on other cardiac valves | 168
AngioVac vacuum-assisted thrombectomy system | 168
extracorporeal circuit | 168
in-line filter | 168
debulking TV vegetations | 168
reducing bacterial load | 168
inflow cannula advanced | 168
extracorporeal circulation initiated | 168
real-time debulking | 168
TEE guidance | 168
additional manipulations | 168
satisfactory debulking | 168
flow stopped | 168
largest components removed | 168
small residual components | 168
moderate TR | 168
no structural damage | 168
components retrieved | 168
visual inspection | 168
culture | 168
hemodynamically stable | 168
vegetation cultures positive | 168
methicillin-sensitive Staphylococcus aureus | 168
6 weeks of antibiotic therapy | 168
suboxone | 168
manage opioid use disorder | 168
discharged | 720
represented with methicillin-resistant Staphylococcus aureus bacteremia | 2160
transesophageal echocardiography | 2160
no abscess | 2160
no worsening vegetation | 2160
6 weeks of antimicrobial therapy | 2160
discharged home | 2592