48 years old | 0
    male | 0
    admitted with altered mental status | 0
    found covered in urine and feces | -24
    confused | -24
    bed ridden | -672
    cough | -672
    diarrhea | -672
    body temperature 35.8°C | 0
    tachycardic (118 beats/minute) | 0
    tachypneic (28 breaths/minute) | 0
    minimal accessory muscle use | 0
    oxygen saturation 100% | 0
    diminished breath sounds on lung bases | 0
    soft abdomen | 0
    distended abdomen | 0
    non-tender abdomen | 0
    bilateral pitting edema in feet | 0
    acute hypoxemic respiratory failure | 0
    tachypnea up to 40 breaths/min | 0
    oxygen saturation 85% on room air | 0
    intubated | 0
    transferred to intensive care | 0
    bilateral pleural effusions | 0
    small pericardial effusion | 0
    large heterogeneous splenomegaly | 0
    ascites | 0
    mesenteric anasarca | 0
    soft-tissue anasarca | 0
    diffuse cerebral atrophy | 0
    severe hyperferritinemia | 0
    blood culture negative | 0
    sputum culture negative | 0
    urine culture negative | 0
    HBsAg negative | 0
    HBsAb negative | 0
    hepatitis C antibody negative | 0
    EBV PCR negative | 0
    SARS-CoV-2 RNA PCR negative | 0
    HIV 1,2 antigen/antibody test negative | 0
    HTLV-1/2 antibodies negative | 0
    CMV DNA PCR ordered | 0
    antinuclear antibodies negative | 0
    anti-double stranded DNA negative | 0
    Beta-2 Glycoprotein 1 antibody negative | 0
    C3 complement negative | 0
    C4 complement negative | 0
    paracentesis performed | 48
    thoracentesis performed | 48
    pleural fluid exudative | 48
    pleural fluid lymphocytic | 48
    cytology negative for malignant cells | 48
    flow cytometry T cell predominance | 48
    T cell rearrangement study positive | 48
    repeat chest CT suggestive of bilateral pneumonia | 48
    bone marrow biopsy hemophagocytic activity | 48
    no evidence of leukemia | 48
    no evidence of lymphoma | 48
    no evidence of plasma cell carcinoma | 48
    no evidence of metastatic carcinoma | 48
    elevated Interleukin 2 Receptor CD25 Soluble | 48
    HLH diagnosis confirmed | 48
    treated with fluids | 0
    treated with vasopressors | 0
    treated with broad-spectrum antibiotics | 0
    worsening renal function | 120
    anasarca | 120
    renal replacement therapy initiated | 120
    HLH-94 protocol initiated | 288
    dexamethasone 20 mg daily | 288
    etoposide 75 mg/m2 | 288
    cardiac arrest | 298
    pulseless electrical activity | 298
    ROSC after 7 min | 298
    refractory shock | 312
    died | 312
    severe hyperkalemia 7.0 meq/L | 298
    hyperphosphatemia 16.1 mg/dL | 298
    hypocalcemia 6.3 mg/dL | 298
    hyperuricemia 11.0 mg/dL | 298
    elevated BUN 66 mg/dL | 298
    elevated creatinine 5.78 mg/dL | 298
    suspicion of TLS | 298
    CMV PCR positive | 298
    TLS diagnosed | 298
    