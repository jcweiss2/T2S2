male | 0
premature birth | 0
emergency cesarean delivery | 0
abruptio placenta | 0
birth weight 1090g | 0
Apgar 4 and 8 | 0
respiratory distress | 0
respiration rate 65 breaths per min | 0
chest retraction | 0
CPAP machine | 0
positive end expiratory pressures 6 | 0
inspired oxygen 30% | 0
cloudy eyes | 0
ectropion | 0
dry ichthyotic skin | 0
typical male genitalia | 0
bilateral undescended testicles | 0
height 75th percentile | 0
weight 25th percentile | 0
head circumference 25th percentile | 0
temperature 36.2°C | 0
heart rate 167 beats per min | 0
normal neurological examination | 0
normal breath sounds | 0
no organomegaly | 0
normal blood count | 0
normal electrolytes | 0
normal liver function | 0
respiratory distress syndrome | 0
ground-glass opacity on X-ray | 0
minor respiratory acidosis | 0
surfactant dosage | 0
continued CPAP assistance | 12
bowel movement | 12
trophic feeding | 72
breast milk | 72
abdominal distension | 144
tachycardia | 144
tachypnea | 144
thrombocytopenia | 144
neutropenia | 144
raised C-reactive protein | 144
meropenem | 144
vancomycin | 144
stopped tropic feeding | 216
antibiotics discontinued | 216
feeding restarted | 216
high-flow oxygen treatment | 336
relapses of unexplained apnea | 504
septic examination negative | 504
brain MRI normal | 504
nasogastric tube | 504
conjugated hyperbilirubinemia | 504
neonatal cholestasis workup | 504
persistent conjugated hyperbilirubinemia | 504
total bilirubin 69.8 umol/L | 504
total parenteral nutrition | 504
genetic studies | 504
X-ray of spine normal | 504
echocardiogram normal | 504
eye test normal | 504
skull X-ray showed craniosynostosis | 504
hepatosplenomegaly not seen | 504
normal-appearing gallbladder | 504
no signs of biliary atresia | 504
albumin level decline | 504
bilirubin rise | 504
AST rise | 504
ALT rise | 504
multiple albumin infusions | 504
infectious etiology investigation | 504
TSH normal | 504
T3 normal | 504
T4 normal | 504
cortisol normal | 504
metabolic disorders negative | 504
galactosemia negative | 504
tyrosinemia type 1 negative | 504
whole-exome sequencing | 672
NOTCH2 gene mutation | 672
heterozygous variant c.1076c>T | 672
p. (Ser359Phe) | 672
chr1: 120512166 | 672
severe cyanosis | 936
apnea | 936
bradycardia | 936
cardio-respiratory resuscitation | 936
intubation | 936
mechanical breathing | 936
epinephrine | 936
septic shock | 936
multiorgan failure | 936
disseminated intravascular coagulation | 936
acute renal damage | 936
capillary leak syndrome | 936
death | 2400
NOTCH2 gene | -2400
ALGS2 | -2400
pathogenic variant | -2400
c.1076c>T | -2400
p. (Ser359Phe) | -2400
chr1: 120512166 | -2400
heterozygous | -2400
autosomal dominant | -2400
neonatal cholestasis | -2400
cholestasis | -2400
liver disease | -2400
genetic disorder | -2400
NOTCH2 mutation | -2400
ALGS | -2400
JAG1 | -2400
NOTCH2 | -2400
craniosynostosis | -2400
ichthyosis | -2400
respiratory distress syndrome | -2400
sepsis | -2400
biliary atresia | -2400
TPN-associated cholestasis | -2400
Hajdu-Cheney syndrome | -2400
Serpentine fibula polycystic renal syndrome | -2400
cancer | -2400
genetic counseling | -2400
familial screening | -2400
neonatal intensive care unit | -2400
pediatric gastroenterology | -2400
clinical nutrition | -2400
liver transplantation | -2400
whole-exome sequencing | -2400
next-generation sequencing | -2400
NOTCH2 gene sequencing | -2400
 Twist Family BHLH Transcription Factor 1 | -2400
TWIST1 | -2400
JAG1/NOTCH | -2400
NOTCH2 signaling | -2400
NOTCH2 mutation | -2400
ALGS2 diagnosis | -2400
cholestasis gene panel | -2400
neonatal cholestasis | -2400
genetic testing | -2400
molecular diagnosis | -2400
genetic counseling | -2400
familial screening | -2400
NOTCH2 gene mutation | -2400
heterozygous variant | -2400
c.1076c>T | -2400
p. (Ser359Phe) | -2400
chr1: 120512166 | -2400
autosomal dominant | -2400
ALGS2 | -2400
neonatal cholestasis | -2400
liver disease | -2400
genetic disorder | -2400
NOTCH2 mutation | -2400
ALGS | -2400
JAG1 | -2400
NOTCH2 | -2400
craniosynostosis | -2400
ichthyosis | -2400
respiratory distress syndrome | -2400
sepsis | -2400
biliary atresia | -2400
TPN-associated cholestasis | -2400
Hajdu-Cheney syndrome | -2400
Serpentine fibula polycystic renal syndrome | -2400
cancer | -2400
genetic counseling | -2400
familial screening | -2400
neonatal intensive care unit | -2400
pediatric gastroenterology | -2400
clinical nutrition | -2400
liver transplantation | -2400
whole-exome sequencing | -2400
next-generation sequencing | -2400
NOTCH2 gene sequencing | -2400
 Twist Family BHLH Transcription Factor 1 | -2400
TWIST1 | -2400
JAG1/NOTCH | -2400
NOTCH2 signaling | -2400
NOTCH2 mutation | -2400
ALGS2 diagnosis | -2400
cholestasis gene panel | -2400
neonatal cholestasis | -2400
genetic testing | -2400
molecular diagnosis | -2400
genetic counseling | -2400
familial screening | -2400
NOTCH2 gene mutation | -2400
heterozygous variant | -2400
c.1076c>T | -2400
p. (Ser359Phe) | -2400
chr1: 120512166 | -2400
autosomal dominant | -2400
ALGS2 | -2400
neonatal cholestasis | -2400
liver disease | -2400
genetic disorder | -2400
NOTCH2 mutation | -2400
ALGS | -2400
JAG1 | -2400
NOTCH2 | -2400
craniosynostosis | -2400
ichthyosis | -2400
respiratory distress syndrome | -2400
sepsis | -2400
biliary atresia | -2400
TPN-associated cholestasis | -2400
Hajdu-Cheney syndrome | -2400
Serpentine fibula polycystic renal syndrome | -2400
cancer | -2400
genetic counseling | -2400
familial screening | -2400
neonatal intensive care unit | -2400
pediatric gastroenterology | -2400
clinical nutrition | -2400
liver transplantation | -2400
whole-exome sequencing | -2400
next-generation sequencing | -2400
NOTCH2 gene sequencing | -2400
 Twist Family BHLH Transcription Factor 1 | -2400
TWIST1 | -2400
JAG1/NOTCH | -2400
NOTCH2 signaling | -2400
NOTCH2 mutation | -2400
ALGS2 diagnosis | -2400
cholestasis gene panel | -2400
neonatal cholestasis | -2400
genetic testing | -2400
molecular diagnosis | -2400
genetic counseling | -2400
familial screening | -2400
NOTCH2 gene mutation | -2400
heterozygous variant | -2400
c.1076c>T | -2400
p. (Ser359Phe) | -2400
chr1: 120512166 | -2400
autosomal dominant | -2400
ALGS2 | -2400
neonatal cholestasis | -2400
liver disease | -2400
genetic disorder | -2400
NOTCH2 mutation | -2400
ALGS | -2400
JAG1 | -2400
NOTCH2 | -2400
craniosynostosis | -2400
ichthyosis | -2400
respiratory distress syndrome | -2400
sepsis | -2400
biliary atresia | -2400
TPN-associated cholestasis | -2400
Hajdu-Cheney syndrome | -2400
Serpentine fibula polycystic renal syndrome | -2400
cancer | -2400
genetic counseling | -2400
familial screening | -2400
neonatal intensive care unit | -2400
pediatric gastroenterology | -2400
clinical nutrition | -2400
liver transplantation | -2400
whole-exome sequencing | -2400
next-generation sequencing | -2400
NOTCH2 gene sequencing | -2400
 Twist Family BHLH Transcription Factor 1 | -2400
TWIST1 | -2400
JAG1/NOTCH | -2400
NOTCH2 signaling | -2400
NOTCH2 mutation | -2400
ALGS2 diagnosis | -2400
cholestasis gene panel | -2400
neonatal cholestasis | -2400
genetic testing | -2400
molecular diagnosis | -2400
genetic counseling | -2400
familial screening | -2400
NOTCH2 gene mutation | -2400
heterozygous variant | -2400
c.1076c>T | -2400
p. (Ser359Phe) | -2400
chr1: 120512166 | -2400
autosomal dominant | -2400
ALGS2 | -2400
neonatal cholestasis | -2400
liver disease | -2400
genetic disorder | -2400
NOTCH2 mutation | -2400
ALGS | -2400
JAG1 | -2400
NOTCH2 | -2400
craniosynostosis | -2400
ichthyosis | -2400
respiratory distress syndrome | -2400
sepsis | -2400
biliary atresia | -2400
TPN-associated cholestasis | -2400
Hajdu-Cheney syndrome | -2400
Serpentine fibula polycystic renal syndrome | -2400
cancer | -2400
genetic counseling | -2400
familial screening | -2400
neonatal intensive care unit | -2400
pediatric gastroenterology | -2400
clinical nutrition | -2400
liver transplantation | -2400
whole-exome sequencing | -2400
next-generation sequencing | -2400
NOTCH2 gene sequencing | -2400
 Twist Family BHLH Transcription Factor 1 | -2400
TWIST1 | -2400
JAG1/NOTCH | -2400
NOTCH2 signaling | -2400
NOTCH2 mutation | -2400
ALGS2 diagnosis | -2400
cholestasis gene panel | -2400
neonatal cholestasis | -2400
genetic testing | -2400
molecular diagnosis | -2400
genetic counseling | -2400
familial screening | -2400
NOTCH2 gene mutation | -2400
heterozygous variant | -2400
c.1076c>T | -2400
p. (Ser359Phe) | -2400
chr1: 120512166 | -2400
autosomal dominant | -2400
ALGS2 | -2400
neonatal cholestasis | -2400
liver disease | -2400
genetic disorder | -2400
NOTCH2 mutation | -2400
ALGS | -2400
JAG1 | -2400
NOTCH2 | -2400
craniosynostosis | -2400
ichthyosis | -2400
respiratory distress syndrome | -2400
sepsis | -2400
biliary atresia | -2400
TPN-associated cholestasis | -2400
Hajdu-Cheney syndrome | -2400
Serpentine fibula polycystic renal syndrome | -2400
cancer | -2400
genetic counseling | -2400
familial screening | -2400
neonatal intensive care unit | -2400
pediatric gastroenterology | -2400
clinical nutrition | -2400
liver transplantation | -2400
whole-exome sequencing | -2400
next-generation sequencing | -2400
NOTCH2 gene sequencing | -2400
 Twist Family BHLH Transcription Factor 1 | -2400
TWIST1 | -2400
JAG1/NOTCH | -2400
NOTCH2 signaling | -2400
NOTCH2 mutation | -2400
ALGS2 diagnosis | -2400
cholestasis gene panel | -2400
neonatal cholestasis | -2400
genetic testing | -2400
molecular diagnosis | -2400
genetic counseling | -2400
familial screening | -2400
NOTCH2 gene mutation | -2400
heterozygous variant | -2400
c.1076c>T | -2400
p. (Ser359Phe) | -2400
chr1: 120512166 | -2400
autosomal dominant | -2400
ALGS2 | -2400
neonatal cholestasis | -2400
liver disease | -2400
genetic disorder | -2400
NOTCH2 mutation | -2400
ALGS | -2400
JAG1 | -2400
NOTCH2 | -2400
craniosynostosis | -2400
ichthyosis | -2400
respiratory distress syndrome | -2400
sepsis | -2400
biliary atresia | -2400
TPN-associated cholestasis | -2400
Hajdu-Cheney syndrome | -2400
Serpentine fibula polycystic renal syndrome | -2400
cancer | -2400
genetic counseling | -2400
familial screening | -2400
neonatal intensive care unit | -2400
pediatric gastroenterology | -2400
clinical nutrition | -2400
liver transplantation | -2400
whole-exome sequencing | -2400
next-generation sequencing | -2400
NOTCH2 gene sequencing | -2400
 Twist Family BHLH Transcription Factor 1 | -2400
TWIST1 | -2400
JAG1/NOTCH | -2400
NOTCH2 signaling | -2400
NOTCH2 mutation | -2400
ALGS2 diagnosis | -2400
cholestasis gene panel | -2400
neonatal cholestasis | -2400
genetic testing | -2400
molecular diagnosis | -2400
genetic counseling | -2400
familial screening | -2400
NOTCH2 gene mutation | -2400
heterozygous variant | -2400
c.1076c>T | -2400
p. (Ser359Phe) | -2400
chr1: 120512166 | -2400
autosomal dominant | -2400
ALGS2 | -2400
neonatal cholestasis | -2400
liver disease | -2400
genetic disorder | -2400
NOTCH2 mutation | -2400
ALGS | -2400
JAG1 | -2400
NOTCH2 | -2400
craniosynostosis | -2400
ichthyosis | -2400
respiratory distress syndrome | -2400
sepsis | -2400
biliary atresia | -2400
TPN-associated cholestasis | -2400
Hajdu-Cheney syndrome | -2400
Serpentine fibula polycystic renal syndrome | -2400
cancer | -2400
genetic counseling | -2400
familial screening | -2400
neonatal intensive care unit | -2400
pediatric gastroenterology | -2400
clinical nutrition | -2400
liver transplantation | -2400
whole-exome sequencing | -2400
next-generation sequencing | -2400
NOTCH2 gene sequencing | -2400
 Twist Family BHLH Transcription Factor 1 | -2400
TWIST1 | -2400
JAG1/NOTCH | -2400
NOTCH2 signaling | -2400
NOTCH2 mutation | -2400
ALGS2 diagnosis | -2400
cholestasis gene panel | -2400
neonatal cholestasis | -2400
genetic testing | -2400
molecular diagnosis | -2400
genetic counseling | -2400
familial screening | -2400
NOTCH2 gene mutation | -2400
heterozygous variant | -2400
c.1076c>T | -2400
p. (Ser359Phe) | -2400
chr1: 120512166 | -2400
autosomal dominant | -2400
ALGS2 | -2400
neonatal cholestasis | -2400
liver disease | -2400
genetic disorder | -2400
NOTCH2 mutation | -2400
ALGS | -2400
JAG1 | -2400
NOTCH2 | -2400
craniosynostosis | -2400
ichthyosis | -2400
respiratory distress syndrome | -2400
sepsis | -2400
biliary atresia | -2400
TPN-associated cholestasis | -2400
Hajdu-Cheney syndrome | -2400
Serpentine fibula polycystic renal syndrome | -2400
cancer | -2400
genetic counseling | -2400
familial screening | -2400
neonatal intensive care unit | -2400
pediatric gastroenterology | -2400
clinical nutrition | -2400
liver transplantation | -2400
whole-exome sequencing | -2400
next-generation sequencing | -2400
NOTCH2 gene sequencing | -2400
 Twist Family BHLH Transcription Factor 1 | -2400
TWIST1 | -2400
JAG1/NOTCH | -2400
NOTCH2 signaling | -2400
NOTCH2 mutation | -2400
ALGS2 diagnosis | -2400
cholestasis gene panel | -2400
neonatal cholestasis | -2400
genetic testing | -2400
molecular diagnosis | -2400
genetic counseling | -2400
familial screening | -2400
NOTCH2 gene mutation | -2400
heterozygous variant | -2400
c.1076c>T | -2400
p. (Ser359Phe) | -2400
chr1: 120512166 | -2400
autosomal dominant | -2400
ALGS2 | -2400
neonatal cholestasis | -2400
liver disease | -2400
genetic disorder | -2400
NOTCH2 mutation | -2400
ALGS | -2400
JAG1 | -2400
NOTCH2 | -2400
craniosynostosis | -2400
ichthyosis | -2400
respiratory distress syndrome | -2400
sepsis | -2400
biliary atresia | -2400
TPN-associated cholestasis | -2400
Hajdu-Cheney syndrome | -2400
Serpentine fibula polycystic renal syndrome | -2400
cancer | -2400
genetic counseling | -2400
familial screening | -2400
neonatal intensive care unit | -2400
pediatric gastroenterology | -2400
clinical nutrition | -2400
liver transplantation | -2400
whole-exome sequencing | -2400
next-generation sequencing | -2400
NOTCH2 gene sequencing | -2400
 Twist Family BHLH Transcription Factor 1 | -2400
TWIST1 | -2400
JAG1/NOTCH | -2400
NOTCH2 signaling | -2400
NOTCH2 mutation | -2400
ALGS2 diagnosis | -2400
cholestasis gene panel | -2400
neonatal cholestasis | -2400
genetic testing | -2400
molecular diagnosis | -2400
genetic counseling | -2400
familial screening | -2400
NOTCH2 gene mutation | -2400
heterozygous variant | -2400
c.1076c>T | -2400
p. (Ser359Phe) | -2400
chr1: 120512166 | -2400
autosomal dominant | -2400
ALGS2 | -2400
neonatal cholestasis | -2400
liver disease | -2400
genetic disorder | -2400
NOTCH2 mutation | -2400
ALGS | -2400
JAG1 | -2400
NOTCH2 | -2400
craniosynostosis | -2400
ichthyosis | -2400
respiratory distress syndrome | -2400
sepsis | -2400
biliary atresia | -2400
TPN-associated cholestasis | -2400
Hajdu-Cheney syndrome | -2400
Serpentine fibula polycystic renal syndrome | -2400
cancer | -2400
genetic counseling | -2400
familial screening | -2400
neonatal intensive care unit | -2400
pediatric gastroenterology | -2400
clinical nutrition | -2400
liver transplantation | -2400
whole-exome sequencing | -2400
next-generation sequencing | -2400
NOTCH2 gene sequencing | -2400
 Twist Family BHLH Transcription Factor 1 | -2400
TWIST1 | -2400
JAG1/NOTCH | -2400
NOTCH2 signaling | -2400
NOTCH2 mutation | -2400
ALGS2 diagnosis | -2400
cholestasis gene panel | -2400
neonatal cholestasis | -2400
genetic testing | -2400
molecular diagnosis | -2400
genetic counseling | -2400
familial screening | -2400
NOTCH2 gene mutation | -2400
heterozygous variant | -2400
c.1076c>T | -2400
p. (Ser359Phe) | -2400
chr1: 120512166 | -2400
autosomal dominant | -2400
ALGS2 | -2400
neonatal cholestasis | -2400
liver disease | -2400
genetic disorder | -2400
NOTCH2 mutation | -2400
ALGS | -2400
JAG1 | -2400
NOTCH2 | -2400
craniosynostosis | -2400
ichthyosis | -2400
respiratory distress syndrome | -2400
sepsis | -2400
biliary atresia | -2400
TPN-associated cholestasis | -2400
Hajdu-Cheney syndrome | -2400
Serpentine fibula polycystic renal syndrome | -2400
cancer | -2400
genetic counseling | -2400
familial screening | -2400
neonatal intensive care unit | -2400
pediatric gastroenterology | -2400
clinical nutrition | -2400
liver transplantation | -2400
whole-exome sequencing | -2400
next-generation sequencing | -2400
NOTCH2 gene sequencing | -2400
 Twist Family BHLH Transcription Factor 1 | -2400
TWIST1 | -2400
JAG1/NOTCH | -2400
NOTCH2 signaling | -2400
NOTCH2 mutation | -2400
ALGS2 diagnosis | -2400
cholestasis gene panel | -2400
neonatal cholestasis | -2400
genetic testing | -2400
molecular diagnosis | -2400
genetic counseling | -2400
familial screening | -2400
NOTCH2 gene mutation | -2400
heterozygous variant | -2400
c.1076c>T | -2400
p. (Ser359Phe) | -2400
chr1: 120512166 | -2400
autosomal dominant | -2400
ALGS2 | -2400
neonatal cholestasis | -2400
liver disease | -2400
genetic disorder | -2400
NOTCH2 mutation | -2400
ALGS | -2400
JAG1 | -2400
NOTCH2 | -2400
craniosynostosis | -2400
ichthyosis | -2400
respiratory distress syndrome | -2400
sepsis | -2400
biliary atresia | -2400
TPN-associated cholestasis | -2400
Hajdu-Cheney syndrome | -2400
Serpentine fibula polycystic renal syndrome | -2400
cancer | -2400
genetic counseling | -2400
familial screening | -2400
neonatal intensive care unit | -2400
pediatric gastroenterology | -2400
clinical nutrition | -2400
liver transplantation | -2400
whole-exome sequencing | -2400
next-generation sequencing | -2400
NOTCH2 gene sequencing | -2400
 Twist Family BHLH Transcription Factor 1 | -2400
TWIST1 | -2400
JAG1/NOTCH | -2400
NOTCH2 signaling | -2400
NOTCH2 mutation | -2400
ALGS2 diagnosis | -2400
cholestasis gene panel | -2400
neonatal cholestasis | -2400
genetic testing | -2400
molecular diagnosis | -2400
genetic counseling | -2400
familial screening | -2400
NOTCH2 gene mutation | -2400
heterozygous variant | -2400
c.1076c>T | -2400
p. (Ser359Phe) | -2400
chr1: 120512166 | -2400
autosomal dominant | -2400
ALGS2 | -2400
neonatal cholestasis | -2400
liver disease | -2400
genetic disorder | -2400
NOTCH2 mutation | -2400
ALGS | -2400
JAG1 | -2400
NOTCH2 | -2400
craniosynostosis | -2400
ichthyosis | -2400
respiratory distress syndrome | -2400
sepsis | -2400
biliary atresia | -2400
TPN-associated cholestasis | -2400
Hajdu-Cheney syndrome | -2400
Serpentine fibula polycystic renal syndrome | -2400
cancer | -2400
genetic counseling | -2400
familial screening | -2400
neonatal intensive care unit | -2400
pediatric gastroenterology | -2400
clinical nutrition | -2400
liver transplantation | -2400
whole-exome sequencing | -2400
next-generation sequencing | -2400
NOTCH2 gene sequencing | -2400
 Twist Family BHLH Transcription Factor 1 | -2400
TWIST1 | -2400
JAG1/NOTCH | -2400
NOTCH2 signaling | -2400
NOTCH2 mutation | -2400
ALGS2 diagnosis | -2400
cholestasis gene panel | -2400
neonatal cholestasis | -2400
genetic testing | -2400
molecular diagnosis | -2400
genetic counseling | -2400
familial screening | -2400
NOTCH2 gene mutation | -2400
heterozygous variant | -2400
c.1076c>T | -2400
p. (Ser359Phe) | -2400
chr1: 120512166 | -2400
autosomal dominant | -2400
ALGS2 | -2400
neonatal cholestasis | -2400
liver disease | -2400
genetic disorder | -2400
NOTCH2 mutation | -2400
ALGS | -2400
JAG1 | -2400
NOTCH2 | -2400
craniosynostosis | -2400
ichthyosis | -2400
respiratory distress syndrome | -2400
sepsis | -2400
biliary atresia | -2400
TPN-associated cholestasis | -2400
Hajdu-Cheney syndrome | -2400
Serpentine fibula polycystic renal syndrome | -2400
cancer | -2400
genetic counseling | -2400
familial screening | -2400
neonatal intensive care unit | -2400
pediatric gastroenterology | -2400
clinical nutrition | -2400
liver transplantation | -2400
whole-exome sequencing | -2400
next-generation sequencing | -2400
NOTCH2 gene sequencing | -2400
 Twist Family BHLH Transcription Factor 1 | -2400
TWIST1 | -2400
JAG1/NOTCH | -2400
NOTCH2 signaling | -2400
NOTCH2 mutation | -2400
ALGS2 diagnosis | -2400
cholestasis gene panel | -2400
neonatal cholestasis | -2400
genetic testing | -2400
molecular diagnosis | -2400
genetic counseling | -2400
familial screening | -2400
NOTCH2 gene mutation | -2400
heterozygous variant | -2400
c.1076c>T | -2400
p. (Ser359Phe) | -2400
chr1: 120512166 | -2400
autosomal dominant | -2400
ALGS2 | -2400
neonatal cholestasis | -2400
liver disease | -2400
genetic disorder | -2400
NOTCH2 mutation | -2400
ALGS | -2400
JAG1 | -2400
NOTCH2 | -2400
craniosynostosis | -2400
ichthyosis | -2400
respiratory distress syndrome | -2400
sepsis | -2400
biliary atresia | -2400
TPN-associated cholestasis | -2400
Hajdu-Cheney syndrome | -2400
Serpentine fibula polycystic renal syndrome | -2400
cancer | -2400
genetic counseling | -2400
familial screening | -2400
neonatal intensive care unit | -2400
pediatric gastroenterology | -2400
clinical nutrition | -2400
liver transplantation | -2400
whole-exome sequencing | -2400
next-generation sequencing | -2400
NOTCH2 gene sequencing | -2400
 Twist Family BHLH Transcription Factor 1 | -2400
TWIST1 | -2400
JAG1/NOTCH | -2400
NOTCH2 signaling | -2400
NOTCH2 mutation | -2400
ALGS2 diagnosis | -2400
cholestasis gene panel | -2400
neonatal cholestasis | -2400
genetic testing | -2400
molecular diagnosis | -2400
genetic counseling | -2400
familial screening | -2400
NOTCH2 gene mutation | -2400
heterozygous variant | -2400
c.1076c>T | -2400
p. (Ser359Phe) | -2400
chr1: 120512166 | -2400
autosomal dominant | -2400
ALGS2 | -2400
neonatal cholestasis | -2400
liver disease | -2400
genetic disorder | -2400
NOTCH2 mutation | -2400
ALGS | -2400
JAG1 | -2400
NOTCH2 | -2400
craniosynostosis | -2400
ichthyosis | -2400
respiratory distress syndrome | -2400
sepsis | -2400
biliary atresia | -2400
TPN-associated cholestasis | -2400
Hajdu-Cheney syndrome | -2400
Serpentine fibula polycystic renal syndrome | -2400
cancer | -2400
genetic counseling | -2400
familial screening | -2400
neonatal intensive care unit | -2400
pediatric gastroenterology | -2400
clinical nutrition | -2400
liver transplantation | -2400
whole-exome sequencing | -2400
next-generation sequencing | -2400
NOTCH2 gene sequencing | -2400
 Twist Family BHLH Transcription Factor 1 | -2400
TWIST1 | -2400
JAG1/NOTCH | -2400
NOTCH2 signaling | -2400
NOTCH2 mutation | -2400
ALGS2 diagnosis | -2400
cholestasis gene panel | -2400
neonatal cholestasis | -2400
genetic testing | -2400
molecular diagnosis | -2400
genetic counseling | -2400
familial screening | -2400
NOTCH2 gene mutation | -2400
heterozygous variant | -2400
c.1076c>T | -2400
p. (Ser359Phe) | -2400
chr1: 120512166 | -2400
autosomal dominant | -2400
ALGS2 | -2400
neonatal cholestasis | -2400
liver disease | -2400
genetic disorder | -2400
NOTCH2 mutation |