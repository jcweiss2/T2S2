30 years old | 0  
    female | 0  
    polysubstance abuse | -72  
    anxiety | -72  
    depression | -72  
    admitted to the Emergency Department | 0  
    unresponsive | 0  
    found in bathtub | -24  
    injected intravenous heroin | -24  
    administered NARCAN 4 mg intranasally | -24  
    no improvement of respiratory status | -24  
    no improvement of level of consciousness | -24  
    arrived at ED | 0  
    unresponsive to verbal stimuli | 0  
    unresponsive to painful stimuli | 0  
    intermittently moaning | 0  
    administered NARCAN 4 mg intravenously | 0  
    no significant improvement in mental status | 0  
    intubated | 0  
    airway protection | 0  
    administered etomidate 20 mg | 0  
    administered succinylcholine 100 mg | 0  
    axillary temperature 25.8°C | 0  
    pulse rate 55 | 0  
    respiratory rate 16 | 0  
    blood pressure 94/40 | 0  
    wet clothes removed | 0  
    warm blankets applied | 0  
    temperature-sensing Foley inserted | 0  
    clear yellow urine 35 ml | 0  
    topical warming with Bair Hugger system | 0  
    warm saline bags placed in axillae | 0  
    warm saline bags placed on groins | 0  
    administered 2 L warmed IV normal saline | 0  
    hyperkalemia 5.6 mmol/L | 0  
    creatinine 1.16 mg/dL | 0  
    hyperglycemia 385 mg/dL | 0  
    hypocalcemia 7.2 mmol/L | 0  
    leukocytosis 16,000 | 0  
    EKG atrial fibrillation | 0  
    EKG Osborne waves | 0  
    central venous access obtained | 0  
    transferred to intensive care unit | 0  
    continued warming with IV fluids | 0  
    bladder irrigation | 0  
    administered regular insulin 10 units | 0  
    administered calcium gluconate | 0  
    became normotensive | 24  
    became normothermic | 24  
    repeat EKG normal rate | 24  
    repeat EKG normal rhythm | 24  
    repeat EKG normal QRS complex | 24  
    Osborne waves resolved | 24  
    extubated | 48  
    following commands | 48  
    answering questions appropriately | 48  
    addiction medicine consulted | 72  
    discharged home | 72  
    friends heard medical stories | -48  
    induced cooling | -48  
    placed in bathtub | -24  
    filled tub with ice | -24  
    inserted ice cubes rectally | -24  
    hypothermia | 0  
    hyperkalemia | 0  
    hypocalcemia | 0  
    hypothermia therapy | -48  
    neurological protection | -48  
    cardiac protection | -48  
    cerebral metabolism reduced | -48  
    decreased intracellular acidosis | -48  
    decreased free radical oxygen production | -48  
    decreased cerebral edema | -48  
    minimized risk of thrombosis | -48  
    decreased infarct size | -48  
    reduced myocardial injury | -48  
    preserved adenosine triphosphate | -48  
    improved blood flow | -48  
    bradycardia risk | -48  
    reduced cardiac output | -48  
    hypotension risk | -48  
    infection risk | -48  
    bleeding risk | -48  
    insulin resistance | -48  
    decreased gastrointestinal mobility | -48  
    reduced cytochrome P450 activity | -48  
    decreased medication clearance | -48  
    electrolyte abnormalities | -48  
    rewarmed 0.2-0.5°C per hour | 24  
    passive rewarming | 0  
    active rewarming | 0  
    removed wet clothes | 0  
    warm blankets | 0  
    Bair Hugger | 0  
    warmed IV fluids | 0  
    heating packs groin | 0  
    heating packs axilla | 0  
    IV fluids irrigation orogastric tube | 0  
    IV fluids irrigation Foley catheter | 0  
    Osborne waves resolved | 24  
    EKG normalized | 24  
    free of arrhythmias | 24  
    no conflicts of interest | 0  
    