90 years old | 0
male | 0
admitted to the hospital | 0
impaired consciousness | 0
respiratory failure | 0
unconscious in a bathtub | -1
chronic cerebral infarct | -8760
Glasgow Coma Scale component scores: E1 V1 M3 | 0
body temperature was 36.1 °C | 0
blood pressure was 154/110 mmHg | 0
pulse rate was 113/min | 0
respiratory rate was 24 breaths/min | 0
SpO2 was 60% | 0
poor inflation of the right chest | 0
diminished respiratory sounds in the right lower lung | 0
intubated with SLT | 0
blood pressure dropped | 0
septic shock | 0
piperacillin/tazobactam | 0
azithromycin | 0
noradrenalin (NAD) 0.3 μg/kg/min | 0
vasopressin (AVP) 1 unit/hour | 0
hydrocortisone 100 mg | 0
dobutamine (DOB) | 0
chest radiography | 1
computed tomography | 1
right middle and lower lung infiltrates | 1
no abnormality in the left lung | 1
arterial blood gas analysis | 1
PaO2 64 mmHg | 1
PaCO2 53 mmHg | 1
pH 7.10 | 1
unilateral distension of left thorax | 1
right thorax did not fully elevate | 1
SLT replaced with DLT | 6
ILV started | 6
arterial blood gas analysis | 6
PaO2 103 mmHg | 6
FiO2: right 1.0, left 0.6 | 6
mean arterial blood pressure (MAP) increased | 6
NAD reduced | 6
DOB reduced | 6
continuous hemodiafiltration | 6
arterial blood gas analysis | 25
PaO2 75 mmHg | 25
FiO2: right 0.5, left 0.5 | 25
arterial blood gas analysis | 45
PaO2 94 mmHg | 45
FiO2: right 0.5, left 0.4 | 45
ILV discontinued | 45
conventional two-lung ventilation | 45
arterial blood gas analysis | 55
PaO2 87 mmHg | 55
PaCO2 41 mmHg | 55
pH 7.33 | 55
vasopressors discontinued | 55
continuous hemodiafiltration discontinued | 55
DLT replaced with SLT | 81
ventilator set to pressure support mode | 81
FiO2 0.3 | 81
PEEP 8 cmH2O | 81
inspiratory pressure 8 cmH2O | 81
extubated | 147