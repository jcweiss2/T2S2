2 years old | 0
castrated male domestic shorthair cat | 0
weighing 4.7 kg | 0
presented to a university teaching hospital | 0
chronic kidney disease | -unknown
diagnosed with chronic kidney disease | -unknown
bloodwork | -unknown
acute and progressively ataxic | -2
vomiting | -2
leukocytosis | -2
neutrophilia | -2
lymphocytosis | -2
mild azotemia | -2
blood urea nitrogen 45 mg/dl | -2
creatinine 2.2 mg/dl | -2
progressive tetraparesis | 0
concerns for respiratory depression | 0
referred for further evaluation | 0
bradycardic | 0
heart rate 120 bpm | 0
tachypneic | 0
48 breaths/min | 0
stuporous mentation | 0
tetraplegia | 0
absent withdrawals | 0
absent peripheral reflexes | 0
weak gag reflex | 0
absent menace response | 0
short shallow breaths | 0
mild hypercapnia | 0
mild azotemia | 0
urinalysis | 0
urine specific gravity 1.018 | 0
moderate bacteriuria | 0
rare presence of white blood cells | 0
minimal red blood cells | 0
accidental ingestion of baclofen | -4
baclofen 10 mg | -4
ingested dose 2.1 mg/kg | -4
hemodialysis recommended | 0
IV fluid therapy | 0
lactated Ringer’s solution | 0
10 ml/h | 0
hemodialysis catheter placement | 0
hemodialysis initiated | 1.5
neonatal extracorporeal circuit | 1.5
blood flow 90 ml/min | 1.5
ultrafiltration flow rate 100 ml/h | 1.5
5 h hemodialysis | 1.5
sodium profiling 150 mmol/l | 1.5
sodium phosphate supplementation | 1.5
lactated Ringer’s solution increased to 150 ml/h | 1.5
anticoagulation with heparin | 1.5
target activated clotting time 180-220 s | 1.5
progressive hypercapnia | 2.5
respiratory acidosis | 2.5
propofol administered | 2.5
endotracheal intubation | 2.5
propofol CRI | 2.5
manual ventilation | 2.5
worsening hypercapnia | 3.5
mechanical ventilation initiated | 3.5
FiO2 100% | 3.5
positive end-expiratory pressure 1 cmH2O | 3.5
respiratory rate 18 breaths/min | 3.5
target tidal volume 10.5 ml/kg | 3.5
peak flow rate 7.1 l/min | 3.5
severe hemorrhage |(note: The assistant message seems cut off or incomplete. You can choose to ignore it. However, if you want me to proceed to answer the user's message, please provide the complete case description.)
