42 years old | 0
    female | 0
    underwent DALK in the left eye with big bubble technique | 0
    recipient stromal flap partially dissected | 0
    air injected into remaining stroma | 0
    donor button cut 8.25 mm | 0
    donor DM peeled off | 0
    donor button placed over recipient DM | 0
    sutured with recipient rim | 0
    donor cornea age 36 years | 0
    donor cornea in situ cornea excision | 0
    surgery had gone well | 0
    postoperative day 1 | 24
    whitish infiltrates along graft-host junction | 24
    severe anterior chamber reaction | 24
    postoperative keratitis | 24
    graft removed | 24
    replaced by another stromal graft | 24
    removed graft sent for microbiology | 24
    corneal scrapings from recipient rim sent for microbiology | 24
    host DM clear and intact | 24
    residual infiltrates in host rim | 24
    repeat-deep anterior lamellar keratoplasty (reDALK) | 24
    clinical picture worse | 48
    infiltrates along entire graft host junction | 48
    hypopyon | 48
    topical vancomycin started | 27
    topical ceftazidime started | 27
    Gram-negative Bacilli identified | 48
    topical antibiotics increased to half hourly | 48
    Klebsiella pneumoniae resistant to multiple antibiotics identified | 72
    imipenem drops started | 72
    gatifloxacin drops added | 72
    infiltrates extended toward center of graft | 96
    hypopyon persisted | 96
    therapeutic penetrating keratoplasty (TPK) | 168
    infiltrates observed in host DM | 168
    graft clear without infiltrates | 192
    hypopyon resolved | 192
    imipenem continued | 192
    gatifloxacin continued | 192
    prednisolone drops added | 264
    unaided vision 6/60 | 1008
    vision improved to 6/18 with pin hole | 1008
    graft clear | 1008
    anterior segment quiet | 1008
    normal intraocular pressure | 1008
    pathogen eradicated | 1008
    <|eot_id|>
    42 years old | 0
    female | 0
    underwent DALK in the left eye with big bubble technique | 0
    recipient stromal flap partially dissected | 0
    air injected into remaining stroma | 0
    donor button cut 8.25 mm | 0
    donor DM peeled off | 0
    donor button placed over recipient DM | 0
    sutured with recipient rim | 0
    donor cornea age 36 years |5
    donor cornea in situ cornea excision |5
    surgery had gone well |0
    postoperative day 1 |24
    whitish infiltrates along graft-host junction |24
    severe anterior chamber reaction |24
    postoperative keratitis |24
    graft removed |24
    replaced by another stromal graft |24
    removed graft sent for microbiology |24
    corneal scrapings from recipient rim sent for microbiology |24
    host DM clear and intact |24
    residual infiltrates in host rim |24
    repeat-deep anterior lamellar keratoplasty (reDALK) |24
    clinical picture worse |48
    infiltrates along entire graft host junction |48
    hypopyon |48
    topical vancomycin started |27
    topical ceftazidime started |27
    Gram-negative Bacilli identified |48
    topical antibiotics increased to half hourly |48
    Klebsiella pneumoniae resistant to multiple antibiotics identified |72
    imipenem drops started |72
    gatifloxacin drops added |72
    infiltrates extended toward center of graft |96
    hypopyon persisted |96
    therapeutic penetrating keratoplasty (TPK) |168
    infiltrates observed in host DM |168
    graft clear without infiltrates |192
    hypopyon resolved |192
    imipenem continued |192
    gatifloxacin continued |192
    prednisolone drops added |264
    unaided vision 6/60 |1008
    vision improved to 6/18 with pin hole |1008
    graft clear |1008
    anterior segment quiet |1008
    normal intraocular pressure |1008
    pathogen eradicated |1008