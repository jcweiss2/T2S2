64 years old | 0
male | 0
polysubstance abuse | -672
hypertension | -672
ischaemic heart disease | -672
admitted to the hospital | 0
COVID-19 positive | 0
asymptomatic | 0
asymptomatic bradycardia | 0
sinus bradycardia | 0
electrocardiogram | 0
right heart axis | 0
incomplete right bundle branch block | 0
downsloping depression of the ST-segment | 0
T inversion | 0
normotensive | 0
good pulse volume | 0
good oxygen saturation | 0
pansystolic murmur | 0
moderate aortic regurgitation | 0
thickened aortic valve | 0
dilated left ventricular chamber | 0
ejection fraction of 70% | 0
no pericardial effusion | 0
pulmonary artery systolic pressure | 0
no foot oedema | 0
trial of bolus intravenous atropine | 0
intravenous infusion of dopamine | 0
transcutaneous cardiac pacing | 12
intravenous infusion of noradrenaline | 12
heart rate improved | 12
blood pressure decreased | 24
transvenous pacing | 24
shortness of breath | 24
chest pain | 24
sweating | 24
re-implantation of transvenous pacing | 24
abdominal pain | 96
no bowel movements | 96
vomiting | 96
streaks of blood on diapers | 96
severe metabolic acidosis | 96
high anion gap | 96
free-flow gastric decompression | 96
computed tomography examination of the abdomen | 96
inflammatory or infective changes | 96
right inguinal hernia | 96
small bowel and mesenteric content | 96
proximal bowel dilatation | 96
obstruction | 96
clinical deterioration | 120
multiorgan failure | 120
persistent hyperglycaemia | 120
cardiorenal syndrome | 120
anuria | 120
worsening metabolic acidosis | 120
fulminant hepatic failure | 120
worsening transaminitis | 120
hyperbilirubinemia | 120
thrombocytopaenia | 120
coagulopathy | 120
N-acetylcysteine regime | 120
third space loss | 120
global pericardial effusion | 120
right ventricular wall thickness | 120
double strengths of triple inotropic support | 120
haemodialysis | 120
sustained slow-efficiency dialysis | 120
continuous veno-venous hemofiltration | 120
repeated cycles of fresh-frozen plasma | 120
packed cells | 120
platelet concentrate | 120
empirical antibiotics | 120
meropenem | 120
death | 144