36 years old | 0
pregnant woman | 0
gravida 2 para 1 | 0
38–39 weeks of gestation | 0
admitted to the hospital | 0
severe pre-eclampsia | 0
obesity class 3 | 0
body mass index: 41.84 kg/m² | 0
oligohydramnios | 0
amniotic fluid index=3 | 0
suspicion of intrauterine growth restriction | 0
COVID-19 | 0
estimated fetal weight of 2200 g | 0
10 regular antenatal visits | -672
blood pressure normal | -672
systolic: 90–110 mm Hg | -672
diastolic: 60–80 mm Hg | -672
at 38 weeks BP 170/110 mm Hg | -24
urinary protein of +2 | -24
diagnosis of severe PE | -24
treated with MgSO4 intravenously | 0
COVID-19 screening | 0
IgG antibody reactive | 0
chest radiograph normal | 0
RT-PCR test performed | 0
abnormal non-stress test | 0
low variability | 0
late deceleration | 0
suspected IUGR | 0
caesarean section performed | 0
sterilization | 0
meconium-stained amniotic fluid | 0
birth weight 2190 g | 0
height 38 cm | 0
1 min Apgar score 7 | 0
5 min Apgar score 8 | 0
maternal COVID-19 molecular test negative | 24
BP decreased | 48
urine output decreased | 48
BP: 100/60 mm Hg | 48
urine output: 160 mL/13 hours | 48
fluid resuscitation | 48
BP still low | 72
BP: 96/54 mm Hg | 72
severe anaemia | 72
haemoglobin: 3.8 g/dL | 72
ultrasound revealed free fluid | 72
internal bleeding | 72
exploratory laparotomy performed | 72
uterus enlarged | 72
atonic | 72
Couvelaire uterus | 72
haematoma in left adnexa | 72
modified B-lynch procedure attempted | 72
supracervical hysterectomy performed | 72
blood loss 1200 mL | 72
fluid input 2300 mL | 72
3 units of whole blood transfusion before surgery | 72
2 units of whole blood during surgery | 72
ICU treatment | 72
ventilator mode PSIMV | 72
positive end expiratory pressure 6 cm H₂O | 72
fraction of inspired oxygen 100% | 72
GCS E4VxM6 | 72
oxygen saturation 97–100% | 72
ventilator support continued | 72
transfusion-related acute lung injury risk | 72
anaemia | 72
hypoalbuminaemia | 72
thrombocytopenia | 72
hyponatraemia | 72
hypokalaemia | 72
non-steroidal anti-inflammatory drugs administered | 72
ceftriaxone administered | 72
albumin administered | 72
packed red cell transfusion | 72
serum electrolyte correction | 72
rhonchi detected | 96
pulmonary oedema suspected | 96
pneumonia differential diagnosis | 96
furosemide administered | 96
meropenem administered | 96
blood culture performed | 96
SARS-CoV-2 molecular tests repeated | 96
RT-PCR positive | 168
COVID:19 with bacterial pneumonia | 168
remdesivir commenced | 168
blood culture no growth | 168
BP consistently elevated | 168
BP >150/90 mm Hg | 168
isosorbide dinitrate administered | 168
nicardipine administered | 168
ventilator maintained for a week | 168
ventilator removed | 192
NRBM maintained | 192
oxygen saturation 97–98% | 192
D-dimer increased | 216
heparin administered | 216
fever | 216
temperature 37.8°C | 216
antipyretics administered | 216
incisional wound bleeding | 264
vital signs normal | 264
fever resolving | 264
wound care performed | 264
convalescent plasma transfusion | 264
ultrasound performed | 264
haematoma superficial to fascia | 264
heparin stopped | 312
no incisional bleeding | 312
RT-PCR negative | 360
RT-PCR negative | 456
Enterococcus gallinarum detected | 432
antibiotics changed | 432
levofloxacin commenced | 432
ciprofloxacin commenced | 432
stable vital signs | 576
BP 126/73 mm Hg | 576
oxygen saturation 95–96% | 576
incisional wound healed | 576
discharged | 600
38–39 weeks of gestation |/home/bruno/chatgpt-assistant/events_processing
