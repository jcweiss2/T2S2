47 years old | 0
female | 0
dysuria | -168
vomiting | -168
right lower back pain | -168
altered level of consciousness | -168
abdominal pain | -168
urinary disorders | -168
fever | -168
loss of appetite | -168
admitted to hospital | 0
treated with antibiotics | -168
nitrofurantoin | -168
dehydration | 0
blood pressure 122/97 mmHg | 0
axillary temperature 35 °C | 0
heart rate 90 beats per minute | 0
respiratory rate 24 breaths per minute | 0
oxygen saturation 92% | 0
soft and painless abdomen | 0
bilateral lung crackles | 0
normal heart auscultation | 0
increased urea level | 0
increased creatinine level | 0
Proteus mirabilis | 0
resistant to nitrofurantoin | 0
treated with cephalothin | 0
acute pyelonephritis | 0
acute renal failure | 0
mechanical ventilation | 48
vasopressor for septic shock | 48
transferred to ICU | 48
piperacillin–tazobactam | 48
anti-HIV test | 48
dialysis | 48
leukopenia | 48
lymphopenia | 48
anemia | 48
urea level increased to 194 mg/dL | 48
creatinine level increased to 6.28 mg/dL | 48
erythroblasts detected | 48
multiple organ dysfunction | 72
coagulopathy | 72
renal failure | 72
circulatory failure | 72
pulmonary failure | 72
petechiae on chest and abdomen | 72
diffuse bleeding in oral cavity | 72
lesions in oral mucosa | 72
severe anemia | 72
received packed red blood cells | 72
structures suspected to be bacteria or fungi | 72
blood culture negative for bacteria | 72
presence of yeasts | 72
anuria | 96
cyanotic extremities | 96
refractory shock | 96
yeast-like structures suspected to be yeasts | 96
phagocytized by monocytes | 96
micafungin initiated | 96
died | 96
H. capsulatum confirmed | 96
anti-HIV test result positive | 96