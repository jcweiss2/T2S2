42 years old | 0
male | 0
admitted to the hospital | 0
severe abdominal pain | 0
fever | -72
body temperature 39°C | 0
jaundice | 0
severe weakness | 0
ill | 0
adynamic | 0
yellowness of the skin and sclera | 0
hot skin | 0
body temperature 38.9°C | 0
heart rate 100 beats per 1 minute | 0
blood pressure 110/70 mm Hg | 0
abdominal pain | -72
pain in the right hypochondrium | -72
radiating to the lower back | -72
chills | -72
subfebrile temperature | -72
rise in body temperature to 38.5°C | -72
diagnosed with acute pyelonephritis | -240
antibiotic therapy | -240
oral ciprofloxacin | -240
analgesics | -240
ketoprophen | -240
nimesulide | -240
abdominal pain sharply increased | 0
spread to the entire right half of the abdomen | 0
rebound tenderness | 0
yellowness of the skin and sclera | 0
darkening of the urine | 0
viral hepatitis | -6840
cholecystostomy | -6840
tumor of the pancreatic head | -6840
suspected | -6840
pancreatoduodenectomy | -6840
cholecystectomy | -6840
external drainage of the pancreatic remnant duct | -6840
pancreatic drainage spontaneously migrated | -6840
no further complications | -6840
formation of a spontaneous internal fistula | -6840
discharged | -6720
diagnosed with DM | -5760
insulin therapy | -5760
smoked | -0
consumed alcohol | -0
worked as a driver | 0
free gas under the right hemidiaphragm | 0
heterogeneity of the liver shadow | 0
small gas-fluid levels in its tissue | 0
signs of bowel paresis | 0
hemoglobin 113 g/l | 0
erythrocytes 4.0×10^12/l | 0
leukocytes 13.9×10^9/l | 0
neutrophils 90% | 0
platelets 279×10^9/l | 0
ALT 810 U/l | 0
AST greater than 913 U/l | 0
amylase 5 U/l | 0
total bilirubin 277 μmol/l | 0
glucose 28.0 mmol/l | 0
creatinine 49 μmol/l | 0
prothrombin index 65% | 0
INR 1.28 | 0
rupture of the liver abscess | 0
peritonitis | 0
emergency surgery | 0
midline laparotomy | 0
brownish muddy fluid | 0
organs of the upper abdomen fixed | 0
purulent-hemorrhagic fluid | 0
liver tissue debris | 0
abscess cavity | 0
intraoperative endoscopy | 0
no ulcer in the gastric stump | 0
anastomosed jejunal loop | 0
efferent jejunal loop freed | 0
abscess cavity flushed | 0
abdominal cavity flushed | 0
drained | 0
prolonged mechanical ventilation | 24
inotropic support with epinephrine | 24
sepsis | 24
blood procalcitonin 5.1 ng/ml | 24
Staphylococcus haemolyticus | 24
Klebsiella pneumoniae | 24
Escherichia coli | 24
vancomycin | 24
meropenem | 24
vancomycin and amikacin | 48
right-sided pneumonia | 240
bilateral pleural effusions | 240
pleural cavities drained | 240
transferred from intensive care unit | 336
surgical ward | 336
gradual improvement | 336
echography | 336
CT | 336
reduction of the liver lesion | 336
discharged | 960
subphrenic drains | 960
draining fluid | 960
serous-purulent | 960
bile staining | 960
drains removed | 1200
outpatient visit | 1200
satisfactory condition | 1936
works occasionally as a driver | 1936
insulin | 1936
enzyme replacement therapy | 1936
echography | 1936
liver tissue healed | 1936
no signs of biliary hypertension | 1936
magnetic resonance imaging | 1936
non-dilated bile ducts | 1936
pancreatic remnant | 1936
non-dilated Wirsung duct | 1936
mild hyperglycemia | 1936
low serum amylase | 1936
normal ranges | 1936