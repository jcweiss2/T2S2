25 years old | 0
female | 0
obesity | 0
body mass index (BMI) 40.1 kg/m2 | 0
polycystic ovary syndrome | 0
iodine allergy | 0
gastritis | 0
admitted to receive LAGB procedure | 0
LAGB procedure | 0
band placed laparoscopically | 0
pars flaccida technique | 0
discharged on the third day | 72
uneventful post-operative course | 0
weight dropped to 95 kg | -1248
occasional malaise | -1248
feverishness | -1248
recurrent upper respiratory tract infections | -1248
readmitted to the surgery department | -1560
fever | -1560
signs of port site infection | -1560
port removed | -1560
discharged after a day | -1559
occasional malaise | -1248
feverishness | -1248
gastroscopy | -936
no signs of a functioning band or its erosion | -936
readmitted to another surgical department | -744
suspicion of band infection | -744
laparoscopy with conversion to laparotomy | -744
band removed | -744
bacterial culture revealed E. coli band infection | -744
targeted antibiotics administered | -744
minimal surgical wound infection | -736
discharged | -736
returned with hectic fever | -728
elevated levels of white blood cell counts (WBC) | -728
elevated levels of C-reactive protein (CRP) | -728
abdominal computed tomography (CT) scan | -728
peritoneal adhesions | -728
abdominal and mediastinal lymphadenopathy | -728
left pleural effusion | -728
broad-spectrum antibiotics administered | -728
chest CT scan | -728
increased parenchymal density | -728
referred to the pulmonology department | -728
elevated levels of Ca-125 antigen | -728
elevated levels of CRP | -728
elevated levels of WBC | -728
elevated levels of γ-glutamyltransferase (GGTP) | -728
elevated levels of D-dimer | -728
elevated levels of procalcitonin | -728
hypoalbuminemia | -728
IgA deficiency | -728
bone marrow biopsy | -728
reactive changes due to infection | -728
no parasite infection | -728
broad-spectrum antibiotics and antifungal agents continued | -728
immunoglobulin therapy administered | -728
sudden abdominal pain | -720
signs of septic shock | -720
urgent laparotomy | -720
massive peritoneal adhesions | -720
moderate ascites | -720
swabbed for culture | -720
liver, omental and peritoneal surgical biopsy | -720
suspecting malignant neoplasm | -720
histopathological examination | -720
chronic granulomatous inflammation | -720
Ziehl-Neelsen stain negative | -720
transferred to the intensive care unit | -720
bronchial lavage and peritoneal effusion tested for Mycobacterium tuberculosis DNA | -720
negative result | -720
suspecting atypical mycobacteriosis | -720
ethambutol, clarithromycin and amikacin introduced | -720
antifungal and antiparasitic agents introduced | -720
total parenteral nutrition introduced | -720
patient’s status stabilized | -720
CRP and WBC levels decreased | -720
persisting fever lowered | -720
corticosteroids administered | -720
enteral nutrition introduced | -720
good effect | -720
discharged | -696
postoperative specimen (omentum fragment) tested further genetically | -696
M. tuberculosis DNA revealed | -696
corticosteroids discontinued | -696
isoniazid, rifampicin, pyrazinamide and streptomycin administered | -696
therapy completed | -480
abdominal CT scan | -480
no pathological findings | -480
fever and malaise withdrew | -480
no symptoms | 0