62 years old | 0
male | 0
diabetes mellitus | 0
hypertension | 0
abdominal pain | 0
palpable pulsatile epigastric mass | 0
bilateral total hip replacements | -672
infection of hip replacements | -672
treated with levofloxacin | -672
treated with teicoplanin | -672
treated with vancomycin | -672
implants removed | -672
joint spacers implanted | -672
blood cultures demonstrated MRSA | -672
blood cultures demonstrated proteus mirabilis | -672
fever | -672
CT demonstrated septic spleen | -336
splenectomy | -336
recurrent sepsis | -120
white blood count of 12,000/mm3 | -120
CT angiography revealed paravisceral aortic pseudoaneurysm | -120
paravisceral aortic pseudoaneurysm | -120
placement of covered stent into CA attempted | 0
placement of covered stent into CA unsuccessful | 0
midline laparotomy | 0
exposure of paravisceral aorta | 0
exposure of infrarenal aorta | 0
division of crura of diaphragm | 0
aortic clamping | 0
opening of pseudoaneurysm | 0
removal of infected tissues and necrotic aortic wall | 0
reconstruction of CA not feasible | 0
ligation of distal CA | 0
excision of pseudoaneurysm | 0
repair of aorta with cryopreserved human aortic allograft patch | 0
aortic cross clamp time 34 min | 0
postoperative stay in intensive care unit | 24
blood cultures confirmed MRSA infection | 24
tissue culture from aortic wall free from bacteria | 24
dismissed from hospital | 168
meropenem treatment | 168
1-year follow-up | 8760
control CTA showed patent SMA and renal arteries | 8760
no pseudoaneurysm or symptom of infection | 8760