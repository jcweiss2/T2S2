male | 0
neonate | 0
born at 37 weeks of gestation | -168
caesarean section | -168
breech presentation | -168
Apgar scores were 8 and 9 | -168
admitted to NICU | 0
7 days of life | 0
chest retractions | 0
fever | 0
38.5°C | 0
pale | 0
moderate tachypnoea | 0
dyspnoea | 0
bilateral fine gasps | 0
chest X-ray showed accentuated bronchovascular markings | 0
WBC count was 11.9 × 10^9/L | 0
polymorphonuclear cells, 59.4% | 0
C-reactive protein level was within a normal range | 0
blood culture was sterile | 0
RSV type A was identified | 0
nasopharyngeal samples were negative for bacteria | 0
empirical antibiotic therapy | 0
penicillin 150,000 IU/kg/die | 0
gentamicin 5 mg/kg/die | 0
nCPAP was started | 2
increasing fraction of oxygen | 2
i.v. systemic corticosteroids | 2
chest X-ray scan showed opacities | 24
upper right and hilar-perihilar left lung regions | 24
antibiotics were discontinued | 96
clinical improvement | 96
sterile blood culture | 96
RSV detection in the nasopharyngeal samples | 96
normal procalcitonin levels | 96
nCPAP was replaced with high-flow nasal cannula | 96
clinical conditions of the baby worsened | 120
severe hypotension | 120
i.v. fluids | 120
catecholamine support | 120
septic shock | 120
chest X-ray displayed massive opacification | 120
right upper and left lower lobes of the lungs | 120
heart ultrasound revealed a moderately hypertrophic interventricular septum | 120
wide-spectrum antibiotics | 120
ampicillin 150 mg/kg/die | 120
gentamicin 5 mg/kg/die | 120
cefotaxime 100 mg/kg/die | 120
nasal-CPAP was re-started | 120
WBC count was 23.2 × 10^9/L | 120
polymorphonuclear cells, 77.7% | 120
C-reactive protein level increased to 15.2 mg/dL | 120
blood culture yielded S. pneumoniae serotype 3 | 120
CSF culture was sterile | 120
i.v. cefotaxime was administered | 120
nCPAP was discontinued | 312
baby was discharged home | 312
clinical course was uneventful | 312
neurodevelopmental outcome was within the normal range | 936
at 18 months of age | 936