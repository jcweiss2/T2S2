28 years old | 0 | 0 
male | 0 | 0 
farmer | 0 | 0 
admitted to the hospital | 0 | 0 
ingestion of two fresh tablets of Celphos | -4 | -4 
vomiting | -4 | 0 
abdominal pain | -4 | 0 
agitated | 0 | 0 
anxious | 0 | 0 
irritable | 0 | 0 
pulse rate not palpable | 0 | 0 
blood pressure not recordable | 0 | 0 
heart rate 110/min | 0 | 0 
respiratory rate 28/min | 0 | 0 
oxygen saturation 95% | 0 | 0 
sinus tachycardia | 0 | 0 
T wave inversion in lead 3 | 0 | 0 
intravenous crystalloids | 0 | 24 
IV magnesium sulphate | 0 | 24 
IV calcium gluconate | 0 | 24 
IV hydrocortisone | 0 | 24 
IV dopamine | 0 | 24 
IV noradrenaline | 0 | 24 
gastric lavage with potassium permanganate | 0 | 0 
activated charcoal | 0 | 24 
arterial blood gas analysis | 0 | 0 
metabolic acidosis | 0 | 0 
pH 7.2 | 0 | 0 
HCO3 8 mmol/L | 0 | 0 
PCO2 33 mmol/L | 0 | 0 
intubated | 0 | 0 
shifted to ICU | 0 | 0 
BP 60-80 mmHg | 6 | 6 
PR 120/min | 6 | 6 
RR 20/min | 6 | 6 
input/output 3L/300 ml | 6 | 24 
monomorphic ventricular tachycardia | 48 | 48 
DC cardio-version | 48 | 48 
IV amiodarone | 48 | 96 
cardiac bio-markers raised | 48 | 336 
normal sinus rhythm | 48 | 336 
ABG pH 7.4 | 96 | 96 
HCO3 18 mmol/L | 96 | 96 
CO2 42 mmol/L | 96 | 96 
BP 70/50-90/60 mmHg | 96 | 96 
blood urea 100 mg/dl | 96 | 96 
serum creatinine 4.5 mg/dl | 96 | 96 
urine output 400 ml/24 hours | 96 | 96 
AST/ALT 80/90 IU/L | 96 | 96 
ALP 200 U/L | 96 | 96 
S bilirubin 2.5 mg/dl | 96 | 96 
kidney failure | 96 | 168 
liver failure | 96 | 168 
BP 100/70 mmHg | 120 | 120 
PR 110/min | 120 | 120 
RR 22/min | 120 | 120 
TLC 14000/mm3 | 120 | 120 
Urea 200 mg/dl | 120 | 120 
S. creatinine 7.5 mg/dl | 120 | 120 
urine output 400 ml/24 hours | 120 | 120 
ABG pH 7.1 | 120 | 120 
HCO3 10 mmol/L | 120 | 120 
haemodialysis | 120 | 120 
haemodialysis | 168 | 168 
blood urea 70 mg/dl | 168 | 168 
creatinine 4.0 mg/dl | 168 | 168 
urine output 1200 ml/24 hours | 168 | 168 
extubated | 144 | 144 
shifted to SDU | 192 | 192 
vitals normal | 192 | 336 
liver and kidney functions improving | 192 | 336 
discharged | 336 | 336