Mayer-Rokitansky-Küster-Hauser syndrome | 0 | 0 
27 years old | 0 | 0 
female | 0 | 0 
admitted to the clinic | 0 | 0 
lower abdominal pain | -336 | 0 
bilateral pelvic pain | -336 | 0 
denied routinely irrigating or dilating her neovagina | -672 | 0 
penetrative sexual intercourse every couple of weeks | -672 | 0 
had not had intercourse in a few months | -720 | 0 
CT imaging of the abdomen | 0 | 0 
tubular, heterogenous, fluid-filled structure | 0 | 0 
outpatient referral to the gynecologist | 0 | 24 
abdominal pain acutely worsened | 24 | 24 
presented to the local Emergency Department | 24 | 24 
diaphoresis | 24 | 24 
significant distress due to pain | 24 | 24 
vitals were unremarkable on presentation | 24 | 24 
leukocytosis | 24 | 24 
absolute neutrophils | 24 | 24 
repeat abdominal CT | 24 | 24 
increasing inflammatory process | 24 | 24 
received empiric intravenous piperacillin-tazobactam | 24 | 24 
transferred emergently to the hospital | 24 | 48 
notably hypotensive | 48 | 48 
tachycardic | 48 | 48 
afebrile | 48 | 48 
tachypneic | 48 | 48 
oxygen saturation of 95 % | 48 | 48 
received four IV fluid boluses | 48 | 48 
antimicrobials were empirically changed | 48 | 48 
taken emergently to the operative room | 48 | 72 
exploratory laparotomy | 72 | 72 
cystoscopy | 72 | 72 
vaginoscopy | 72 | 72 
normal bladder and urethra | 72 | 72 
entirely obliterated introitus | 72 | 72 
diffuse intra-abdominal spillage of the mucus | 72 | 72 
perforated sigmoid neovagina | 72 | 72 
about one liter of purulent fluid was drained | 72 | 72 
three intrabdominal drains were placed | 72 | 72 
post-operatively, the patient remained intubated | 72 | 192 
requiring mechanical ventilation | 72 | 192 
septic shock requiring three vasopressor agents | 72 | 192 
antimicrobials were transitioned | 120 | 120 
peritoneal culture growing gram-negative rods | 120 | 120 
blood cultures remained negative | 120 | 192 
peritoneal cultures finalized to Bacterioides thetaioaomicron | 168 | 168 
Bacterioides caccae | 168 | 168 
Actinomyces species | 168 | 168 
antimicrobials were changed | 168 | 168 
weaned off vasopressors | 192 | 192 
extubated | 192 | 192 
transferred to the general floor | 288 | 288 
Infectious Diseases team was consulted | 288 | 288 
additional susceptibilities for the Bacteroides species were requested | 288 | 288 
discharged home | 360 | 360 
abdominal wound vacuum | 360 | 360 
IV piperacillin-tazobactam for four weeks | 360 | 504 
experienced generalized malaise | 504 | 504 
diffuse abdominal pain | 504 | 504 
readmitted with sepsis | 504 | 504 
laboratory data revealed white blood count | 504 | 504 
absolute neutrophil count | 504 | 504 
d-dimer | 504 | 504 
lactate | 504 | 504 
CT of the chest, abdomen and pelvis | 504 | 504 
bilateral pleural effusions | 504 | 504 
loculated left pleural effusion | 504 | 504 
multiple new abdominal abscesses | 504 | 504 
transcutaneous drainage catheter in pelvis | 504 | 504 
open anterior midline wound with wound vacuum | 504 | 504 
hypoxemia | 504 | 504 
transferred to the intensive care unit | 504 | 504 
IV piperacillin-tazobactam was continued | 504 | 504 
underwent placement of a right perihepatic drain | 504 | 528 
aspiration of 20 mL of purulence | 528 | 528 
unsuccessful drainage of peri-splenic collection | 528 | 528 
blood cultures remained negative | 528 | 528 
interventional radiology was reconsulted | 528 | 528 
drained 350 mL of pus from the right perinephric abscess | 528 | 528 
drained 90 mL of pus from her perisplenic abscess | 528 | 528 
broad-spectrum PCR was sent on the drained fluid | 528 | 528 
improved clinically | 528 | 768 
antimicrobials were narrowed | 768 | 768 
discharged based on the susceptibilities | 768 | 768 
broad spectrum PCR from the fluid was positive | 768 | 768 
followed up at the adult infectious diseases clinic | 864 | 864 
continued on ampicillin-sulbactam | 864 | 864 
plans to reimage | 864 | 864 
clinically improved | 864 | 864 
repeat CT abdomen demonstrated decreased in the size of right and left sub-phrenic abscesses | 1008 | 1008 
transitioned from IV ampicillin-sulbactam to oral amoxicillin-clavulanate | 1008 | 1008 
complete resolution of the abscesses | 1008 | 1008