70 years old | 0
male | 0
emergency esophageal diversion | -720
injury to the cervical esophagus | -720
spinal surgery | -720
gastric pull-up procedure | -168
anastomotic leakage | -168
endoscopy | -168
esophageal stent | -168
local cervical infection | -504
sepsis | -504
arterial hypertonus | 0
non-active smoking status | 0
ischemic stroke | 0
incomplete senso-motoric hemiparesis | 0
thyroidectomy | 0
open prostatectomy | 0
prostate cancer | 0
malnutrition | 0
systemic inflammation | 0
jugular phlegmon | 0
cervical phlegmon | 0
hemoglobin level of 6.7 g/dL | 0
white blood cell count of 6400 cells/μL | 0
platelet count of 210 × 103/μL | 0
creatinine level of 0.76 mg/dL | 0
unremarkable liver and cholestasis parameters | 0
albumin level of 2.8 g/dL | 0
dislodged esophageal stent | 0
extraesophageal air and fluid-filled cavity | 0
esophageal perforation | 0
infected cavity | 0
esophageal stenosis | 0
stent removal | 0
endoscopic vacuum therapy | 168
EsoSponge system | 168
jugular and cervical phlegmon resolved | 336
repeated endoscopic balloon dilatation | 336
subtotal esophageal resection | 504
reconstruction using a free-jejunal graft interposition | 504
CT angiography | 504
partial sternotomy | 504
laparotomy | 504
jejunal segment harvested | 504
left carotid artery and the left jugular vein used as recipient vessels | 504
graft implanted in an isoperistaltic position | 504
cervical anastomosis performed in an end-to-end fashion | 504
upper mediastinal gastro-jejunostomy in a side-to-side fashion | 504
upper sternum resected | 504
soft tissue defect covered with a sternocleidomastoid muscle flap | 504
abdominal reconstruction achieved by an end-to-end jejunojejunostomy | 504
oral alimentation reestablished | 720
daily speech therapy | 720
anastomotic healing confirmed radiologically and endoscopically | 720
patient transferred to a rehabilitation clinic | 720