45 years old | 0
    male | 0
    admitted to the ICU | 0
    fever | -168
    cough | -168
    generalized weakness | -168
    loose motions | -168
    altered sensorium | -48
    herpetiform rash on the back | -168
    rash becoming generalized | -168
    petechiae | -168
    ecchymotic patch | -168
    disoriented | 0
    irritable | 0
    not obeying verbal commands | 0
    moving all limbs | 0
    no lymphadenopathy | 0
    no eschar | 0
    chronic alcoholism | 0
    heavy smoking | 0
    severe thrombocytopenia | 0
    raised urea | 0
    raised creatinine | 0
    raised liver enzymes | 0
    increased serum bilirubin | 0
    increased lactate | 0
    increased ammonia | 0
    normal coagulation parameters | 0
    normal fibrinogen | 0
    oropharyngeal bleeding | 0
    platelet transfusion | 0
    severe metabolic acidosis | 0
    fluid resuscitation | 0
    improved urine output | 0
    started on broad spectrum antibiotics | 0
    intubated | 0
    mechanical ventilator support | 0
    neurologic deterioration | 0
    hemodynamic deterioration | 0
    respiratory deterioration | 0
    normal MRI brain | 0
    generalized retiform purpuric rash | 0
    high grade fever | 0
    hypotension | 0
    blood negative for malaria parasite | 0
    negative dengue serology | 0
    negative Leptospira serology | 0
    presumptive diagnosis of meningococcemia | 0
    awaiting blood culture report | 0
    negative Gram stains of skin biopsy | 0
    negative serum Neisseria meningitidis Ag detection | 0
    negative urine Neisseria meningitidis Ag detection | 0
    lumbar puncture not performed | 0
    negative venereal disease research laboratory | 0
    negative CARBOGEN | 0
    negative rapid plasma reagin card test |:0
    negative acute hepatitis profile | 0
    negative vasculitis workup | 0
    sterile blood cultures | 0
    sterile urine culture | 0
    Weil-Felix test OX-2 titer 1:320 | 0
    Weil-Felix test OX-19 titer 1:40 | 0
    Weil-Felix test OX-K titer 1:40 | 0
    negative Orientia tsutsugamushi serology | 0
    started on doxycycline | 0
    no increase in titers after 1 week | 168
    developed bullous eruptions | 24
    skin biopsy findings | 24
    negative direct immunofluorescence study | 24
    prominent vasculitis | 24
    improved neurologically | 48
    improved hemodynamically | 48
    extubated | 48
    shifted out of ICU | 48
    improved serum creatinine | 48
    elevated liver enzymes | 48
    decreased serum bilirubin | 48
    retiform rash fading | 48
    clinical improvement | 48
    discharged | 336
