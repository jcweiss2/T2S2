2 years old | 0
male | 0
admitted to pediatric polyclinic | 0
fever | -168
upper respiratory tract infection | -168
treated for upper respiratory tract infection | -168
fever again | -168
delivery by cesarean section | -17520
birth weight 3450 g | -17520
length 50 cm | -17520
head circumference 35 cm | -17520
hospitalized at newborn intensive care unit | -17520
hyperbilirubinemia | -17520
neonatal sepsis | -17520
no reproduction in blood culture | -17520
no reproduction in urinary culture | -17520
no frequent admissions to hospital | -17520
no hospitalization | -17520
no known disease in family history | 0
body weight 12.5 kg | 0
height 87 cm | 0
physical examination normal | 0
body temperature 37.2 oC | 0
WBC 19.2x103/µL | 0
Hb 10.7 g/dL | 0
HTC 31.9% | 0
MCV 74 fL | 0
RDW 16.8 | 0
Plt 332000x103/µL | 0
C-reactive protein 3.04 mg/dL | 0
biochemical parameters normal | 0
urine dipstick positive for leukocytes | 0
urine dipstick negative for blood/hemoglobin | 0
urine dipstick negative for nitrite | 0
12-14 leukocytes in urinary sediment | 0
abundant amorphous crystals in urinary sediment | 0
urinary system ultrasound revealed 7.5-mm stone | 0
grade 2 hydronephrosis | 0
urinary culture detected R. ornithinolytica | 0
sensitive to trimethoprim/sulfamethoxazole | 0
sensitive to amoxicillin/clavulanic acid | 0
sensitive to gentamicin | 0
sensitive to cefuroxime axetil | 0
resistant to ampicillin | 0
urine sample obtained with catheter | 0
culture obtained with catheter | 0
tests for stone etiology ordered | 0
oral cefuroxime axetil started | 0
urinary culture taken with catheter | 24
R. ornithinolytica reproduced | 24
antibiotic sensitivity report same as former | 24
urine cultured on EMB | 24
urine cultured on blood agar | 24
colonies proliferated | 24
gram-negative bacilli isolated | 24
bacterial identification using VITEK-2 | 24
immunoglobulins normal | 24
calcium/creatinine normal | 24
oxalate normal | 24
citrate normal | 24
magnesium normal | 24
uric acid normal | 24
grade 2 hydronephrosis | 24
endoscopic stone removal | 24
double J catheter introduced | 24
remission of hydronephrosis | 24
follow-up at nephrology clinic | 24
follow-up at pediatric urology clinic | 24
urinary stone ultrasound image | 0
R. ornithinolytica confirmed | 24
cefuroxime therapy for 10 days | 24
follow-up urine culture negative | 240
