18 years old | 0
male | 0
admitted to the hospital | 0
fever | -72
rash | -72
acne | -672
minocycline | -672
increased WBC count | 0
eosinophilia | 0
systemic involvement | 0
diffuse erythematous or maculopapular eruption | 0
pruritis | 0
DRESS syndrome |;0
fever persisted | 0
rash persisted | 0
discharged | 24
