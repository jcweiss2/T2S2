46 years old | 0
male | 0
motorcyclist | 0
admitted to the emergency department | 0
road traffic collision | -1
erythematous changes over the trunk | 0
severe abnormalities of the extremities | 0
bilateral lung contusions | 0
mild hemothorax | 0
fractures of the right third to fifth ribs | 0
liver laceration | 0
minor active bleed | 0
empiric trans-arterial embolization | 0
Gelfoam | 0
sinus tachycardia | 0
ventricular premature complex (VPC) | 0
elevated troponin-I | 0
echocardiogram | 0
no cardiac wall abnormality | 0
no pericardial effusion | 0
10 French pigtail chest catheter | 96
left pleural effusion | 96
chest radiography (CXR) | 96
hemithorax white-out | 96
fluid amount | 96
pigtail catheter size not revised | 120
transferred to a regular hospital ward | 240
stable condition | 240
chest pigtail catheter removed | 240
shortness of breath | 264
recurrent massive left pleural effusion | 264
echo-guided pigtail insertion | 264
minimal turbid fluid drained | 264
culture of drainage fluid positive for Staphylococcus aureus (S. aureus) | 264
symptoms temporarily improved | 264
severe chest pain | 288
worsening shortness of breath | 288
frequent VPC | 288
cardiomegaly | 288
severe purulent pericardial effusion | 288
purulent pericarditis | 288
cardiac tamponade | 288
pericardiectomy | 288
debridement | 288
purulent exudate removed | 288
right atrium/superior vena cava (RA/SVC) junction tear | 288
RA/SVC junction tear repaired | 288
oxacillin administered | 288
gentamycin administered | 288
dyspnea with desaturation | 504
bilateral lung pleural effusion | 504
empyema | 504
decortication surgery | 504
multiple bilateral loculated effusions and exudates removed | 504
intravenous administration of antibiotics | 504
recovered | 720
discharged | 720