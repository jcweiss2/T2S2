11 years old | 0
male | 0
admitted to the hospital | 0
fever | -96
nausea | -96
abdominal pain | -96
pneumonia | -6048
hospitalized | 0
vital signs stable | 0
clear breathing sound | 0
direct tenderness on the right side of abdomen | 0
elevated C-reactive protein | 0
elevated procalcitonin | 0
normal whole blood cell count | 0
bowel wall thickening in the terminal ileum | 0
enlarged lymph nodes along the ileocolic artery | 0
administration of intravenous antibiotics | 0
diarrhea | 24
hypotension | 72
inotropic agents | 72
transferred to intensive care unit | 72
elevated white blood cell count | 72
elevated platelet count | 72
elevated serum CRP | 72
elevated procalcitonin | 72
elevated serum aspartate aminotransferase | 72
elevated serum alanine aminotransferase | 72
elevated pro-brain natriuretic peptide | 72
elevated prothrombin time | 72
elevated activated partial thromboplastin time | 72
elevated fibrinogen level | 72
elevated D-dimer level | 72
cardiomegaly on chest X-ray | 96
hypoalbuminemia | 96
intravenous immunoglobulin | 96
conjunctival injection | 144
cracked lips | 144
strawberry tongue | 144
KDSS | 144
high-dose aspirin | 144
fever subsided | 192
erythematous papular rash | 192
finger desquamation | 192
transferred to general ward | 192
aspirin dose reduced | 192
desquamation of the left wrist | 312
desquamation of the perianal area | 312
elevated inflammation markers normalized | 312
coagulopathy normalized | 312
cardiomegaly not detected | 312
pleural effusion not detected | 312
enlarged lymph nodes reduced | 312
coronary artery dilatation reduced | 312
discharged | 312
SARS-CoV-2 antibody test positive | 0
SARS-CoV-2 PCR test negative | 0
SARS-CoV-2 IgM test negative | 0
SARS-CoV-2 IgG test positive | 0
lung parenchymal consolidation | 144
MIS-C | 0