72 years old | 0
    woman | 0
    presented with cough | -168
    presented with shortness of breath | -168
    presented with weakness | -168
    hypoxia | 0
    oxygen saturation of 80% | 0
    admitted for COVID-19 pneumonia | 0
    superimposed with bacterial pneumonia | 0
    sepsis | 0
    hypertension | 0
    hypothyroidism | 0
    obesity | 0
    treatment with dexamethasone | 0
    treatment with albuterol | 0
    nasal cannula oxygen | 0
    prophylactic therapeutic dosing of enoxaparin | 0
    blood cultures grew gram-positive cocci in clusters | 0
    vancomycin | 0
    meropenem | 0
    doxycycline | 0
    intravenous piggyback set to gravity infiltrated | -384
    infiltration caused mild swelling | -384
    infiltration caused pain | -384
    worsening respiratory failure | -384
    endotracheal intubation | -384
    transfer to intensive care unit | -384
    started on norepinephrine | -384
    proned periodically | -384
    gradual improvement of respiratory status | -384
    medication administration via triple lumen central catheter | -384
    blood draws via triple lumen central catheter | -384
    no peripheral intravenous catheters in left hand or arm | -384
    poor peripheral venous access | -384
    left hand displayed worsened swelling | 0
    large dorsal purplish bulla | 0
    responsive to yes or no questions | 0
    reported pain in hand | 0
    reported pain in distal forearm | 0
    unable to flex fingers | 0
    denied numbness | 0
    vascular surgery consultation | 0
    no signs of arterial insufficiency | 0
    arterial duplex ultrasound | 0
    Doppler examination | 0
    computed tomography demonstrated hematoma of dorsal wrist | 0
    venous duplex ultrasound | 0
    no evidence of venous thrombosis | 0
    nonsurgical management | 0
    local wound care | 0
    hand surgery consultation | 72
    symptoms continued to worsen | 72
    examination found faint ulnar and radial Doppler signals | 72
    cool fingers | 72
    considerable blistering | 72
    mottling | 72
    intrinsic minus posturing | 72
    worsened pain with passive extension of IP and MCP joints | 72
    limited active range of motion | 72
    compartment pressures of 52 and 54 mm Hg in hypothenar eminence | 72
    compartment pressures of 40 and 42 mm Hg in thenar eminence | 72
    delta pressures ranged between -2 and 30 mm Hg | 72
    compartment syndrome diagnosis | 72
    decompressive fasciotomy | 72
    thenar and hypothenar muscle groups severely edematous | 72
    dorsal incisions over second and fourth metacarpals | 72
    release interosseous and adductor compartments | 72
    evacuate dorsal hematoma | 72
    all compartments released | 72
    dorsal fasciotomies closed loosely | 72
    improved pain | 168
    range of motion limited | 168
    improved flexion and extension to <10° | 168
    improved swelling | 168
    improved flexion and extension to >10° | 216
    oppose thumb to middle finger | 216
    dorsal wound with superficial necrosis | 216
    dorsal wound with eschar ulnarly | 216
    discharged | 744
    physical therapy | 744
    composite fist formed | 744
    fully extend fingers | 744
    necrotic eschar debrided serially | 2016
    wound fully healed | 4872
    mild scar contracture | 4872
    wrist flexion limited to 60° | 4872
    full wrist extension | 4872
    full range of motion in digit IP and MCP joints | 4872
    forearm supination | 4872
    forearm pronation | 4872
    wrist radial deviation | 4872
    wrist ulnar deviation | 4872
    Disabilities of the Arm, Shoulder, and Hand score 60 of 100 | 4872
    very satisfied with outcome | 4872
    resolution of neuropathic pain symptoms | 4872
    written informed consent obtained | 4872
    no benefits related to subject | 4872
    <|eot_id|>
    72 years old | 0
    woman | 0
    presented with cough | -168
    presented with shortness of breath | -168
    presented with weakness | -168
    hypoxia | 0
    oxygen saturation of 80% | 0
    admitted for COVID-19 pneumonia | 0
    superimposed with bacterial pneumonia |3
    sepsis | 0
    hypertension | 0
    hypothyroidism | 0
    obesity | 0
    treatment with dexamethasone | 0
    treatment with albuterol | 0
    nasal cannula oxygen | 0
    prophylactic therapeutic dosing of enoxaparin | 0
    blood cultures grew gram-positive cocci in clusters | 0
    vancomycin | 0
    meropenem | 0
    doxycycline | 0
    intravenous piggyback set to gravity infiltrated | -384
    infiltration caused mild swelling | -384
    infiltration caused pain | -384
    worsening respiratory failure | -384
    endotracheal intubation | -384
    transfer to intensive care unit | -384
    started on norepinephrine | -384
    proned periodically | -384
    gradual improvement of respiratory status | -384
    medication administration via triple lumen central catheter | -384
    blood draws via triple lumen central catheter | -384
    no peripheral intravenous catheters in left hand or arm | -384
    poor peripheral venous access | -384
    left hand displayed worsened swelling | 0
    large dorsal purplish bulla | 0
    responsive to yes or no questions | 0
    reported pain in hand | 0
    reported pain in distal forearm | 0
    unable to flex fingers | 0
    denied numbness | 0
    vascular surgery consultation | 0
    no signs of arterial insufficiency | 0
    arterial duplex ultrasound | 0
    Doppler examination | 0
    computed tomography demonstrated hematoma of dorsal wrist | 0
    venous duplex ultrasound | 0
    no evidence of venous thrombosis | 0
    nonsurgical management | 0
    local wound care | 0
    hand surgery consultation | 72
    symptoms continued to worsen | 72
    examination found faint ulnar and radial Doppler signals | 72
    cool fingers | 72
    considerable blistering | 72
    mottling | 72
    intrinsic minus posturing | 72
    worsened pain with passive extension of IP and MCP joints | 72
    limited active range of motion | 72
    compartment pressures of 52 and 54 mm Hg in hypothenar eminence | 72
    compartment pressures of 40 and 42 mm Hg in thenar eminence | 72
    delta pressures ranged between -2 and 30 mm Hg | 72
    compartment syndrome diagnosis | 72
    decompressive fasciotomy | 72
    thenar and hypothenar muscle groups severely edematous | 72
    dorsal incisions over second and fourth metacarpals | 72
    release interosseous and adductor compartments | 72
    evacuate dorsal hematoma | 72
    all compartments released | 72
    dorsal fasciotomies closed loosely | 72
    improved pain | 168
    range of motion limited | 168
    improved flexion and extension to <10° | 168
    improved swelling | 168
    improved flexion and extension to >10° | 216
    oppose thumb to middle finger | 216
    dorsal wound with superficial necrosis | 216
    dorsal wound with eschar ulnarly | 216
    discharged | 744
    physical therapy | 744
    composite fist formed | 744
    fully extend fingers | 744
    necrotic eschar debrided serially | 2016
    wound fully healed | 4872
    mild scar contracture | 4872
    wrist flexion limited to 60° | 4872
    full wrist extension | 4872
    full range of motion in digit IP and MCP joints | 4872
    forearm supination | 4872
    forearm pronation | 4872
    wrist radial deviation | 4872
    wrist ulnar deviation | 4872
    Disabilities of the Arm, Shoulder, and Hand score 60 of 100 | 4872
    very satisfied with outcome | 4872
    resolution of neuropathic pain symptoms | 4872
    written informed consent obtained | 4872
    no benefits related to subject | 4872

    