54 years old|0  
    female|0  
    admitted to the hospital|0  
    progressively worsening altered mental status|0  
    weakness|0  
    symptoms ongoing for several months| -4320  
    alert|0  
    oriented to self|0  
    oriented to time|0  
    oriented to place|0  
    oriented to situation|0  
    mild decline in baseline cognitive function|0  
    elevated blood pressure|0  
    moon facies|0  
    weakness in bilateral lower extremities|0  
    reduced strength in bilateral hip flexors|0  
    inability to ambulate independently|0  
    sensation intact|0  
    reflexes intact|0  
    diabetes mellitus| -4320  
    recently uncontrolled diabetes mellitus| -4320  
    recent diagnosis of hypertension| -4320  
    requiring anti-hypertensive therapy| -4320  
    past medical history of remote early-stage breast cancer| -4320  
    underwent bilateral total mastectomy| -4320  
    received adjuvant hormonal therapy| -4320  
    non-smoker|0  
    rare alcohol use|0  
    profound hypokalemia|0  
    alkalemia|0  
    aldosterone normal|0  
    aldosterone/renin ratio normal|0  
    direct renin decreased|0  
    serum random cortisol elevated|0  
    serum ACTH elevated|0  
    dexamethasone suppression testing abnormal|0  
    8 mg dexamethasone did not suppress AM cortisol|0  
    AM cortisol 84.6 mcg/dL|0  
    serum chromogranin level elevated|0  
    CT imaging of the chest|0  
    CT imaging of the abdomen|0  
    CT imaging of the pelvis|0  
    bilateral pulmonary lesions|0  
    intraabdominal lymphadenopathy|0  
    bilateral diffuse adrenal gland thickening|0  
    multiple hepatic metastases|0  
    2.5 cm lesion at the pancreatic tail|0  
    pancreatic lesion visualized on MRI abdomen|0  
    bone scan negative for metastatic lesions|0  
    pituitary MRI negative for a pituitary mass|0  
    underwent electromyogram of bilateral lower extremities|0  
    electromyogram abnormal|0  
    suggestive of severe proximal myopathy|0  
    underwent muscle biopsy|0  
    muscle biopsy reported as severe generalized myofiber atrophy|0  
    biopsy of liver lesion|0  
    metastatic NET, G1|0  
    well differentiated NET, grade-1|0  
    Ki-67 proliferative index <3%|0  
    mitotic rate not reported|0  
    neoplastic cells positive for synaptophysin|0  
    neoplastic cells positive for chromogranin|0  
    neoplastic cells positive for caudal-type homeobox 2 (CDX2)|0  
    neoplastic cells negative for calretinin|0  
    neoplastic cells negative for inhibin|0  
    neoplastic cells negative for S100|0  
    neoplastic cells negative for cytokeratin-7 (CK7)|0  
    neoplastic cells negative for GATA binding protein 3 (GATA-3)|0  
    neoplastic cells negative for thyroid transcription factor-1 (TTF-1)|0  
    germline genetic testing not completed|0  
    clinical presentation concerning for recurrent and metastatic breast cancer|0  
    differential diagnosis ruled out|0  
    Guillain-Barre syndrome considered|0  
    electromyography findings ruled out Guillain-Barre syndrome|0  
    muscle biopsy ruled out Guillain-Barre syndrome|0  
    muscle biopsy negative for evidence of inflammation|0  
    muscle biopsy negative for vasculitis|0  
    other autoimmune myositis conditions ruled out|0  
    negative serum markers|0  
    negative muscle biopsy findings|0  
    hypercortisolemia|0  
    liver tissue biopsy findings of NET|0  
    muscle biopsy findings|0  
    elevated serum cortisol|0  
    elevated serum ACTH|0  
    weakness secondary to glucocorticoid-induced myopathy|0  
    diagnosed with metastatic ACTH-producing NET|0  
    primary tumor suspected in pancreas|0  
    tumor burden not high|0  
    malignant hypercortisolism difficult to control|0  
    poor prognostic feature|0  
    invasive diagnostic procedures avoided|0  
    started on octreotide acetate 100 mg twice daily|0  
    minimal improvement|0  
    started on ketoconazole 400 mg twice daily|0  
    titrated up to 600 mg three times daily|0  
    received 38 days of oral ketoconazole|0  
    slight decrease in ACTH and cortisol levels|0  
    no meaningful change in motor strength appreciated|0  
    started abiraterone acetate 500 mg twice daily|0  
    serum cortisol reduction immediate|0  
    serum cortisol started downtrend by day 3|72  
    cortisol levels completely normalized with 10 days of starting AA|240  
    complete resolution of hypercortisolemia|240  
    cortisol-induced myopathy remained stable|240  
    concern for durability of response|240  
    underwent bilateral adrenal artery embolization|240  
    AA discontinued after 14 days of treatment|336  
    discharged to rehabilitation facility|336  
    admitted to medical intensive care unit one week after discharge|432  
    management of septic shock secondary to pneumonia|432  
    ultimately succumbed|432  

<|eot_id|>
