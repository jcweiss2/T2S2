male | 0
34 weeks of gestation | 0
caesarean section | 0
central placenta previa with hemorrhage | 0
hyperthyroidism | -672
dexamethasone | -24
admitted to the neonatal intensive care unit | 0
intubated | 0
respiratory distress | 0
pulmonary hemorrhage | 0
high-frequency oscillatory ventilation (HFOV) | 0
inhalational nitric oxide | 72
PPHN | 72
surfactant | 0
umbilical venous catheter (UVC) | 0
umbilical artery catheter (UAC) | 0
hydrocortisone (HC) | 0
circulatory failure | 0
hypotension | 0
intensive inotropic support | 0
epinephrine | 0
dopamine | 0
weaned HC | 120
mean arterial pressure (MAP) raised | 168
blood exchange | 0
albumin | 0
hyperbilirubinemia | 0
acute hypokalemia | 336
potassium replacement | 336
oral repletion | 336
fetal echocardiography | -672
structurally normal heart | -672
pediatric cardiology consultation | 24
transthoracic echocardiogram (TTE) | 24
right-to-left shunting of blood | 24
patent ductal arteriosus (PDA) | 24
bidirectional shunting | 24
mean pulmonary artery pressure (PAP) | 72
LVEF | 72
atrial left-right shunt | 72
patent ductal shunt | 72
PPHN ameliorated | 264
mean PAP decreased | 264
echocardiography repeated | 720
profound cardiomegaly | 720
harsh systolic ejection murmur | 720
severe thickening of the IVS | 720
mild thickening of the posterior left ventricular wall (LVPW) | 720
hypertrophic cardiomyopathy (HCM) | 720
propranolol | 720
captopril | 720
24-hour Holter electrocardiographic monitoring | 720
arrhythmia | 720
serial transesophageal echocardiograms | 720
thickness of the IVS decreased | 1440
supplemental oxygen discontinued | 720
tandem mass spectroscopy analysis | 720
exome sequencing | 720
discharged from hospital | 1080
post-discharge follow-up | 1440
MAP | 1440
cardiologic evaluation | 1440