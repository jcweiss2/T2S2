51 years old | 0
female | 0
admitted to the hospital | 0
osteoarthritis | -672
acetabular dysplasia | -672
total hip arthroplasty | 0
famotidine | -2
glycopyrrolate | -2
spinal block | -2
bupivacaine | -2
midazolam | -2
oxygen | -2
anesthesia | -2
blood loss | -2
fluid administered | -2
urine output | -2
arterial blood gas analysis | -2
pH 7.386 | -2
PaCO2 42.5 mmHg | -2
PaO2 164.7 mmHg | -2
HCO3 24.6 mM/L | -2
SaO2 99.8% | -2
Hb 10.1 g/dl | -2
recovery room | 0
blood pressure 110/60 mmHg | 0
heart rate 65 beats/min | 0
pulse oximetry 99% | 0
complained of being cold | 0
shivered | 0
covered with a warm blanket | 0
dizziness | 3
slight cyanosis | 3
blood test | 3
chemical test | 3
coagulation | 3
hemoglobin 7.9 g/dl | 3
hematocrit 24.3% | 3
hypovolemia | 3
central venous catheter | 3
lidocaine | 3
local anesthesia | 3
venipuncture | 3
J-inducing wire | 3
catheter insertion | 3
blood absorption | 3
packed red blood cells | 3
emergency blood test | 3
Hemovac | 3
computed tomography | 6
iopromide | 6
contrast medium | 6
heaviness in chest | 6
oxygen | 6
arterial blood gas analysis | 6
pH 7.406 | 6
PaCO2 36.8 mmHg | 6
PaO2 109.6 mmHg | 6
HCO3-11.5 mM/L | 6
SaO 299.3% | 6
electrocardiogram | 6
echo cardiogram | 6
cardiac enzyme test | 6
chest X-ray | 6
hydrothorax | 6
sono guide | 6
Chiba needle | 6
pleural effusion | 6
pig tail catheter | 6
contrast medium drainage | 6
catheter replacement | 6
catheter fixation | 9
vital signs monitoring | 9
anaphylaxis | 9
cardiopulmonary side-effects | 9
chest X-ray | 12
hydrothorax disappearance | 12
catheter removal | 168
discharged | 336