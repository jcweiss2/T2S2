22 years old | 0
woman | 0
presented to the emergency with dyspnea | -72
denied cough | 0
denied sputum | 0
denied chest pain | 0
denied other respiratory symptoms | 0
denied symptoms of upper extremity weakness | 0
denied symptoms of lower extremity weakness | 0
denied blurred vision | 0
denied swallowing difficulty | 0
speech problem (nasal speech) | -4320
treated by ENT surgeons | -4320
treated by speech therapist | -4320
history of substance abuse | absent | 0
recent drug intake | absent | 0
labored breathing | 0
respiratory rate of 40 breaths/minute | 0
confused | 0
SaO2 85% | 0
blood pressure 146/98 mm Hg | 0
pulse 104/minute and regular | 0
body temperature 36.7°C | 0
pedal edema absent | 0
neck vein engorgement absent | 0
mild crackles at both lung fields | 0
arterial blood gas analysis pH7.314 | 0
arterial blood gas analysis PaCO2 56.7 mm Hg | 0
arterial blood gas analysis PaO2 92.2 mmHg | 0
arterial blood gas analysis oxygen saturation 90% | 0
chest X-ray no definite infiltration | 0
chest X-ray reduced lung volume | 0
white blood cell count 6980 μL | 0
hemoglobin 12.5 g/dL | 0
platelet count 345000 μL | 0
blood glucose 94 mg/dL | 0
BUN/Cr 12/0.8 mg/dL | 0
AST/ALT 24/25 units/L | 0
chest CT scan no pulmonary thromboembolism | 0
ECG sinus tachycardia | 0
echocardiography normal systolic function | 0
echocardiography normal diastolic function | 0
respiratory failure imminent | 0
supplemental oxygen | 0
transferred to intensive care unit | 0
mechanically ventilated | 0
rapid sequence induction | 0
IV midazolam 3 mg | 0
succinylcholine 70 mg | 0
SaO2 improved to 100% | 0
unable to breathe without mechanical support | 0
muscle relaxant effect worn off | 0
ENT surgeon assessment | 0
upper airway obstruction absent | 0
considered neuromuscular disorders | 0
considered Guillain–Barre syndrome | 0
considered MG | 0
physical examination normal | 0
neurological examination normal | 0
cerebrospinal fluid analysis normal | 0
diagnosis of MG | 0
electromyography decremental response | 0
pharmacological Jolly test incremental responses | 0
acetylcholine receptor antibody titer 12.4 nmol/L | 0
condition improved | 0
pyridostigmine bromide 720 mg/day | 0
prednisolone 30 mg/day | 0
intravenous gamma-globulin 400 mg/kg/day | 0
weaning from ventilator failed | 336
tracheostomy performed | 336
successfully weaned from ventilator | 1344
discharged | 1344
advised thymectomy | 1344
developed respiratory distress | 1344
respiratory arrest | 1344
signs and symptoms of sepsis | 1344
successfully intubated | 1344
resuscitated | 1344
prednisolone stepped up | 1344
pyridostigmine stepped up | 1344
antibiotics | 1344
fluid | 1344
intravenous gamma-globulin 400 mg/kg/day | 1344
finally discharged | 576
thymus follicular hyperplasia | 576
currently followed up | 576
responded well with maintenance steroid | 576
responded well with pyridostigmine | 576
