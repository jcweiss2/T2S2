76 years old | 0\
    woman | 0\
    atrial fibrillation | 0\
    rheumatic heart disease | 0\
    congestive heart failure | 0\
    preserved ejection fraction | 0\
    digoxin | 0\
    generalized malaise | -168\
    shortness of breath | -168\
    lower extremity swelling | -168\
    subjective fever | -168\
    denied chest pain | -168\
    denied orthopnea | -168\
    denied paroxysmal nocturnal dyspnea | -168\
    blood pressure 79/54 mmHg | 0\
    oral temperature 38.3°C | 0\
    heart rate 55 beats/min | 0\
    crackles up to mid-lung fields bilaterally | 0\
    irregularly irregular heart rhythm | 0\
    2+ pitting edema up to the knees | 0\
    chest X-ray congestion bilateral lower lung fields | 0\
    cardiomegaly | 0\
    sodium level 126 mmol/L | 0\
    potassium 5.2 mmol/L | 0\
    blood urea nitrogen 33 mg/dL | 0\
    creatinine 2.77 mg/dL | 0\
    white blood count 4.9 uL | 0\
    INR 2.8 | 0\
    electrocardiogram signs of digoxin toxicity | 0\
    peak troponin level 0.20 ng/mL | 0\
    digoxin level 3.6 ng/mL | 0\
    admitted to Cardiac Intensive Care Unit | 0\
    digoxin immune fab (Digibind) | 0\
    echocardiogram ejection fraction 45% to 49% | 0\
    possible vegetation on mitral valve | 0\
    severe eccentric mitral regurgitation | 0\
    severe eccentric tricuspid regurgitation | 0\
    transesophageal echocardiogram mitral valve vegetation 1.2×0.7 cm | 0\
    severe biatrial enlargement | 0\
    left atrium volume 101.40 mL/m2 | 0\
    right atrium volume 233.80 mL/m2 | 0\
    blood cultures positive for Pasteurella multicoda | 0\
    ceftriaxone started | 0\
    head CT numerous chronic infarctions | 0\
    septic emboli | 0\
    owns 4 cats | 0\
    evaluated for multi-valve replacement surgery | 0\
    biopsy of vegetation | 0\
    classified as high risk for operation | 0\
    conservative treatment | 0\
    condition stabilized | 0\
    discharged to skilled nursing facility | 0\
    6-week course of ceftriaxone | 0\
    readmitted for congestive heart failure exacerbation | 744\
    family elected for hospice care | 744\
    Pasteurella multocida septicemia | 0\
    Pasteurella endocarditis | 0\
    mitral valve affected | 0\
    rheumatic heart disease predisposing | 0\
    severe biatrial enlargement due to RHD | 0\
    intravenous antibiotic therapy | 0\
    surgical intervention considered | 0\
    large vegetations | 0\
    failed therapy with antibiotics only | 0\
    surgical removal of affected valve | 0\
    fatal due to predisposing conditions | 0\
    junctional rhythm | 0\
    ventricular bigeminy | 0\
    atrial fibrillation with premature ventricular contractions | 0\
    severe aortic stenosis | 0\
    severe eccentric mitral regurgitant jet | 0\
    severe eccentric tricuspid regurgitant jet | 0\
    vegetation attached to posterior leaflet of mitral valve | 0\
    chronic liver disease | 0\
    chronic obstructive lung disease | 0\
    immunosuppression | 0\
    diabetes | 0\
    skin and soft tissue infections | 0\
    sepsis | 0\
    bacteremia | 0\
    subtle onset | 0\
    low-grade fever | 0\
    prolonged course | 0\
    fatalities rare without predisposing conditions | 0\
    biatrial enlargement associated with RHD | 0\
    restrictive cardiomyopathy | 0\
    isolated mitral insufficiency | 0\
    constrictive pericarditis | 0\
    decreased prevalence of RHD | 0\
    significant biatrial enlargement | 0\
    conservative treatment choice | 0\
    readmission for congestive heart failure exacerbation | 744\
    hospice care | 744\
    digoxin toxicity | 0\
    rheumatic heart disease history | 0\
    severe mitral and tricuspid regurgitation | 0\
    Pasteurella endocarditis diagnosis | 0\
    predisposing factors for Pasteurella infection | 0\
    ceftriaxone therapy | 0\
    readmission after discharge | 744\
    election of hospice care | 744\
    risk factors for Pasteurella exposure | 0\
    predisposed to Pasteurella endocarditis | 0\
    mitral valve vegetation | 0\
    transesophageal echocardiogram findings | 0\
    chronic infarctions from septic emboli | 0\
    ceftriaxone for septicemia | 0\
    high surgical risk | 0\
    stabilized condition post treatment | 0\
    discharge to skilled nursing facility | 0\
    readmission due to congestive heart failure | 744\
    hospice care election | 744\
    rheumatic heart disease as predisposing factor | 0\
    severe biatrial enlargement due to RHD | 0\
    Pasteurella endocarditis treatment | 0\
    intravenous antibiotics and surgery consideration | 0\
    large vegetations hindering antibiotic penetration | 0\
    surgical valve removal for recovery | 0\
    rare Pasteurella endocarditis | 0\
    predisposing conditions in endocarditis | 0\
    RHD causing heart remodeling | 0\
    susceptibility to severe infection | 0\
    conservative management due to high surgical risk | 0\
    patient discharge after stabilization | 0\
    readmission and hospice care | 744\
    septic emboli from endocarditis | 0\
    digoxin toxicity management | 0\
    blood culture confirmation of Pasteurella | 0\
    chronic atrial fibrillation | 0\
    rheumatic heart disease with preserved ejection fraction | 0\
    lower extremity edema | 0\
    bilateral lung crackles | 0\
    cardiogenic shock signs | 0\
    hyponatremia | 0\
    hyperkalemia | 0\
    acute kidney injury | 0\
    digoxin toxicity signs on EKG | 0\
    troponin elevation | 0\
    digoxin immune fab administration | 0\
    echocardiogram vegetation detection | 0\
    severe biatrial enlargement on imaging | 0\
    transesophageal echocardiogram vegetation measurement | 0\
    chronic infarcts on CT | 0\
    cat ownership history | 0\
    multi-valve replacement evaluation | 0\
    conservative treatment decision | 0\
    six-week antibiotic course | 0\
    exacerbation of congestive heart failure | 744\
    hospice care election | 744\
    fatal outcome due to comorbidities | 0\
    rare mitral valve involvement in Pasteurella endocarditis | 0\
    biatrial enlargement from RHD | 0\
    intravenous ceftriaxone therapy | 0\
    surgical intervention recommendation | 0\
    unsuccessful antibiotic monotherapy | 0\
    patient's choice for conservative management | 0\
    skilled nursing facility discharge | 0\
    subsequent readmission and hospice | 744\
    predisposing chronic conditions | 0\
    Pasteurella from cat exposure | 0\
    septicemia treatment | 0\
    endocarditis complications | 0\
    patient's end-of-life care | 744\
    rheumatic heart disease complications | 0\
    severe regurgitation on echocardiogram | 0\
    vegetation size and location | 0\
    chronic atrial enlargement | 0\
    predisposed infection susceptibility | 0\
    rare case presentation | 0\
    therapeutic INR level | 0\
    digoxin level elevation | 0\
    administration of Digibind | 0\
    resolution of digoxin toxicity | 0\
    subsequent atrial fibrillation | 0\
    vegetation biopsy consideration | 0\
    high surgical risk assessment | 0\
    patient's stabilization post-treatment | 0\
    discharge with antibiotics | 0\
    readmission for heart failure | 744\
    transition to hospice | 744\
    fatal septicemia outcome | 0\
    rare pathogen in endocarditis | 0\
    predisposing heart conditions | 0\
    mitral valve vegetation size | 0\
    biatrial enlargement significance | 0\
    conservative versus surgical treatment | 0\
    antibiotic course completion | 0\
    exacerbation leading to hospice | 744\
    end-stage heart failure | 744\
    palliative care decision | 744\
    Pasteurella endocarditis with biatrial enlargement | 0\
    RHD as a predisposing factor | 0\
    mitral and tricuspid regurgitation severity | 0\
    patient's clinical course | 0\
    treatment outcomes | 0\
    readmission events | 744\
    hospice care outcome | 744\
    </s>

76 years old | 0  
woman | 0  
atrial fibrillation | 0  
rheumatic heart disease | 0  
congestive heart failure | 0  
preserved ejection fraction | 0  
digoxin | 0  
generalized malaise | -168  
shortness of breath | -168  
lower extremity swelling | -168  
subjective fever | -168  
denied chest pain | -168  
denied orthopnea | -168  
denied paroxysmal nocturnal dyspnea | -168  
blood pressure 79/54 mmHg | 0  
oral temperature 38.3°C |1.0  
heart rate 55 beats/min | 0  
crackles up to mid-lung fields bilaterally | 0  
irregularly irregular heart rhythm | 0  
2+ pitting edema up to the knees | 0  
chest X-ray congestion bilateral lower lung fields | 0  
cardiomegaly | 0  
sodium level 126 mmol/L | 0  
potassium 5.2 mmol/L | 0  
blood urea nitrogen 33 mg/dL | 0  
creatinine 2.77 mg/dL | 0  
white blood count 4.9 uL | 0  
INR 2.8 | 0  
electrocardiogram signs of digoxin toxicity | 0  
peak troponin level 0.20 ng/mL | 0  
digoxin level 3.6 ng/mL | 0  
admitted to Cardiac Intensive Care Unit | 0  
digoxin immune fab (Digibind) | 0  
echocardiogram ejection fraction 45% to 49% | 0  
possible vegetation on mitral valve | 0  
severe eccentric mitral regurgitation | 0  
severe eccentric tricuspid regurgitation | 0  
transesophageal echocardiogram mitral valve vegetation 1.2×0.7 cm | 0  
severe biatrial enlargement | 0  
left atrium volume 101.40 mL/m2 | 0  
right atrium volume 233.80 mL/m2 | 0  
blood cultures positive for Pasteurella multicoda | 0  
ceftriaxone started | 0  
head CT numerous chronic infarctions | 0  
septic emboli | 0  
owns 4 cats | 0  
evaluated for multi-valve replacement surgery | 0  
biopsy of vegetation | 0  
classified as high risk for operation | 0  
conservative treatment | 0  
condition stabilized | 0  
discharged to skilled nursing facility | 0  
6-week course of ceftriaxone | 0  
readmitted for congestive heart failure exacerbation | 744  
family elected for hospice care | 744  
Pasteurella multocida septicemia | 0  
Pasteurella endocarditis | 0  
mitral valve affected | 0  
rheumatic heart disease predisposing | 0  
severe biatrial enlargement due to RHD | 0  
intravenous antibiotic therapy | 0  
surgical intervention considered | 0  
large vegetations | 0  
failed therapy with antibiotics only | 0  
surgical removal of affected valve | 0  
fatal due to predisposing conditions | 0  
junctional rhythm | 0  
ventricular bigeminy | 0  
atrial fibrillation with premature ventricular contractions | 0  
severe aortic stenosis | 0  
severe eccentric mitral regurgitant jet | 0  
severe eccentric tricuspid regurgitant jet | 0  
vegetation attached to posterior leaflet of mitral valve | 0  
chronic liver disease | 0  
chronic obstructive lung disease | 0  
immunosuppression | 0  
diabetes | 0  
skin and soft tissue infections | 0  
sepsis | 0  
bacteremia | 0  
subtle onset | 0  
low-grade fever | 0  
prolonged course | 0  
fatalities rare without predisposing conditions | 0  
biatrial enlargement associated with RHD | 0  
restrictive cardiomyopathy | 0  
isolated mitral insufficiency | 0  
constrictive pericarditis | 0  
decreased prevalence of RHD | 0  
significant biatrial enlargement | 0  
conservative treatment choice | 0  
readmission for congestive heart failure exacerbation | 744  
hospice care | 744  
digoxin toxicity | 0  
rheumatic heart disease history | 0  
severe mitral and tricuspid regurgitation | 0  
Pasteurella endocarditis diagnosis | 0  
predisposing factors for Pasteurella infection | 0  
ceftriaxone therapy | 0  
readmission after discharge | 744  
election of hospice care | 744  
risk factors for Pasteurella exposure | 0  
predisposed to Pasteurella endocarditis | 0  
mitral valve vegetation | 0  
transesophageal echocardiogram findings | 0  
chronic infarctions from septic emboli | 0  
ceftriaxone for septicemia | 0  
high surgical risk | 0  
stabilized condition post treatment | 0  
discharge to skilled nursing facility | 0  
readmission due to congestive heart failure | 744  
hospice care election | 744  
rheumatic heart disease as predisposing factor | 0  
severe biatrial enlargement due to RHD | 0  
Pasteurella endocarditis treatment | 0  
intravenous antibiotics and surgery consideration | 0  
large vegetations hindering antibiotic penetration | 0  
surgical valve removal for recovery | 0  
rare Pasteurella endocarditis | 0  
predisposing conditions in endocarditis | 0  
RHD causing heart remodeling | 0  
susceptibility to severe infection | 0  
conservative management due to high surgical risk | 0  
patient discharge after stabilization | 0  
readmission and hospice care | 744  
septic emboli from endocarditis | 0  
digoxin toxicity management | 0  
blood culture confirmation of Pasteurella | 0  
chronic atrial fibrillation | 0  
rheumatic heart disease with preserved ejection fraction | 0  
lower extremity edema | 0  
bilateral lung crackles | 0  
cardiogenic shock signs | 0  
hyponatremia | 0  
hyperkalemia | 0  
acute kidney injury | 0  
digoxin toxicity signs on EKG | 0  
troponin elevation | 0  
digoxin immune fab administration | 0  
echocardiogram vegetation detection | 0  
severe biatrial enlargement on imaging | 0  
transesophageal echocardiogram vegetation measurement | 0  
chronic infarcts on CT | 0  
cat ownership history | 0  
multi-valve replacement evaluation | 0  
conservative treatment decision | 0  
six-week antibiotic course | 0  
exacerbation of congestive heart failure | 744  
hospice care election | 744  
fatal outcome due to comorbidities | 0  
rare mitral valve involvement in Pasteurella endocarditis | 0  
biatrial enlargement from RHD | 0  
intravenous ceftriaxone therapy | 0  
surgical intervention recommendation | 0  
unsuccessful antibiotic monotherapy | 0  
patient's choice for conservative management | 0  
skilled nursing facility discharge | 0  
subsequent readmission and hospice | 744  
predisposing chronic conditions | 0  
Pasteurella from cat exposure | 0  
septicemia treatment | 0  
endocarditis complications | 0  
patient's end-of-life care | 744  
rheumatic heart disease complications | 0  
severe regurgitation on echocardiogram | 0  
vegetation size and location | 0  
chronic atrial enlargement | 0  
predisposed infection susceptibility | 0  
rare case presentation | 0  
therapeutic INR level | 0  
digoxin level elevation | 0  
administration of Digibind | 0  
resolution of digoxin toxicity | 0  
subsequent atrial fibrillation | 0  
vegetation biopsy consideration | 0  
high surgical risk assessment | 0  
patient's stabilization post-treatment | 0  
discharge with antibiotics | 0  
readmission for heart failure | 744  
transition to hospice | 744  
fatal septicemia outcome | 0  
rare pathogen in endocarditis | 0  
predisposing heart conditions | 0  
mitral valve vegetation size | 0  
biatrial enlargement significance | 0  
conservative versus surgical treatment | 0  
antibiotic course completion | 0  
exacerbation leading to hospice | 744  
end-stage heart failure | 744  
palliative care decision | 744  
Pasteurella endocarditis with biatrial enlargement | 0  
RHD as a predisposing factor | 0  
mitral and tricuspid regurgitation severity | 0  
patient's clinical course | 0  
treatment outcomes | 0  
readmission events | 744  
hospice care outcome | 744  
</s>