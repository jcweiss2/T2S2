58 years old|0
female|0
brought to the emergency room|0
complaints of lethargy|0
fever|0
watery, non-bloody diarrhea|0
diarrhea for 2 days|0
confused|-48
progressively became lethargic|-48
fever (maximum temperature of 39.4 °C at home)|-48
no history of loss of consciousness|0
no history of shortness of breath|0
no history of cough|0
no recent travel|0
no exposure to sick contacts|0
hypertension|0
losartan|0
rheumatoid arthritis|0
tofacitinib 11 mg once daily|0
CKD stage 3A|0
COPD|0
current smoker|0
smoking history of 20 pack-year|0
no alcohol use|0
no illicit drug use|0
temperature of 39.4 °C|0
heart rate of 112 bpm|0
respiratory rate of 20 per minute|0
blood pressure 127/75 mmHg|0
oxygen saturation 85% on room air|0
oxygen saturation improved to 100% on 3 L nasal cannula|0
drowsy|0
intermittently follow commands|0
clear breath sounds bilaterally|0
normal heart sounds|0
non-distended abdomen|0
non-tender abdomen|0
normal bowel sounds|0
oriented to place and person|0
not oriented to time|0
no focal neurological deficits|0
no neck rigidity|0
negative meningeal signs|0
no rashes|0
WBC 17,400 cells/μL|0
87% neutrophils|0
hemoglobin 10.7 g/dL|0
platelet count 235,000/μL|0
sodium 126 mEq/L|0
potassium 3.0 mEq/L|0
bicarbonate 19.3 mEq/L|0
BUN 32 mg/dL|0
creatinine 2 mg/dL (baseline 1.3 mg/dL)|0
AST 260 U/L|0
ALT 40 U/L|0
CK 347,700 U/L|0
negative Hepatitis A IgM antibody|0
negative Hepatitis B surface antigen|0
negative Hepatitis B core IgM antibody|0
negative Hepatitis C antibodies|0
stool studies: no WBC|0
normal stool osmolality|0
normal calprotectin|0
negative urine culture|0
negative blood culture|0
negative stool culture|0
positive urine Legionella pneumophila serogroup 1 antigen|0
urinalysis: 51-100/hpf WBC|0
urinalysis: 6-10/hpf RBC|0
urinalysis: 3+ occult blood|0
chest X-ray bibasilar densities|0
right pleural effusion|0
CT head: no acute intracranial abnormality|0
CT chest/abdomen/pelvis: patchy right basilar opacities|0
colonic diverticulosis|0
no diverticulitis|0
started on broad-spectrum antibiotics|0
sepsis of unknown source|0
antibiotics changed to azithromycin|0
improvement in mental status|24
improvement in diarrhea|24
worsening renal function|24
worsening CK|24
anuria|24
signs of volume overload|24
started on hemodialysis|24
transferred to ICU|24
vasopressor requirements|24
remained in ICU for 7 days|168
received 14-day azithromycin course|168
tofacitinib discontinued|0
weaned off pressors|168
supplementary oxygen requirement reduced|168
started on midodrine|168
rhabdomyolysis resolved|168
discharged after 17 days|408
complete renal recovery in 2 months|1344
