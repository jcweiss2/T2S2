80 years old | 0
male | 0
admitted to the hospital | 0
history of cardiovascular risk factors | -672
history of hypertension | -672
history of type 2 diabetes | -672
history of tabagism | -672
vague and diffuse abdominal pain | 0
physical examination | 0
no signs of peritonitis | 0
normal vital signs | 0
no free fluid in the abdomen | 0
emergency ultrasound | 0
leucocytosis | 0
elevated PCR | 0
increased LDH | 0
contrast-enhanced CT scan | 0
extensive thrombosis affecting SMA | 0
thrombosis affecting SMV | 0
no involvement of the portal vein | 0
marked thinning of the small bowel wall | 0
lack of contrast-enhancement | 0
no luminal dilatation | 0
no air-fluid levels | 0
intramural gas | 0
pneumatosis intestinalis | 0
gas in the SMA | 0
gas in the branches of the SMA | 0
no gas in the SMV | 0
no gas in the portal vein | 0
emergency surgery | 12
excision of multiple necrotic bowel loops | 12
transferred to the intensive care unit | 12
died the next day | 24
multiple organ dysfunction syndrome | 24
ischemia-reperfusion events | 24
systemic inflammatory response syndrome | 24