29 years old | 0
woman | 0
referred to intensive care unit | 0
chronic ulcerative pancolitis | -35040
autoimmune hepatitis | -35040
cirrhosis (Child-Pugh C) | -35040
treated with azathioprine | -35040
treated with corticosteroids | -35040
prednisone 30 mg per day | -35040
consulted emergency department | -96
fever | -96
left leg pain | -96
diarrhoea | -96
septic shock | -10
temperature 39.4°C | 0
heart rate 120 beats per minute | 0
blood pressure 70/50 mm Hg | 0
oxygen saturation 50% | 0
acute respiratory distress | 0
Glasgow Coma Score 8 | 0
no stiff neck | 0
purpuric erythema 10 cm posterior left thigh | 0
mechanical ventilation | 0
large-volume expansion | 0
catecholaminergic support by adrenaline | 0
cardiac arrest | 0
low-flow time 5 minutes | 0
acute renal failure (creatinemia 204 μmol/L) | 0
increased creatinine kinase level (930 IU/L) | 0
disseminated intravascular coagulation | 0
platelets 40 × 10^9/L | 0
D-dimer >10 000 ng/L | 0
prothrombin time 17% | 0
leucopenia (3800 cells/mm³) | 0
hepatocellular failure (factor V 30%, bilirubin 99 μ/L) | 0
lactate level 16 mmol/L | 0
C-reactive protein 13.4 mg/L | 0
broad-spectrum antibiotic therapy (piperacillin–tazobactam, vancomycin, amikacin) | 0
clindamycin added | 2
bullae | 0
superficial excoriations | 0
erythema | 0
subcutaneous fat infiltration in legs | 0
diagnosis of necrotizing soft tissue infection | 0
surgery | 4
extensive debridement of tissues | 4
tissues not necrotizing | 4
E. coli growth in samples | 0
antibiotic therapy changed to cefotaxime | 0
continuous renal replacement therapy | 0
anuric renal failure | 0
continuous bleeding of surgical wound | 0
haemorrhagic shock | 0
massive transfusions | 0
disseminated intravascular coagulation worsened | 0
skin lesions extensive | 24
subcutaneous crackles | 24
second surgery debridement | 24
extension of soft tissue cellulitis | 24
lake of bleeding | 24
necrotizing fascia | 24
patient died | 24
E. coli strain phylogenetic group C | 0
virulence factors (yersiniabactin, aerobactin, salmochelin, hemolysin, cytotoxic necrotizing factor 1, Hra, P fimbriae pilin) | 0
genes associated with virulence plasmidic region (hlyF, ompTp, etsC, iss) | 0
immunocompromised | 0
liver cirrhosis (Child-Pugh C) | 0
azathioprine | 0
corticosteroids | 0
fatal necrotizing soft tissue infection | 24
septic shock before death | 24
failure of immune system | 0
deficient bactericidal activity of IgM | 0
soft tissue infections prevalence 2-11% | 0
Staphylococcus aureus | 0
Streptococcus pyogenes | 0
bullae present in 15% of necrotizing soft tissue infections | 0
virulence factors (PAI IIJ96, conserved virulence plasmidic region) | 0
cnf1 toxin | 0
activation of RhoGTPases | 0
aware E. coli responsible for necrotizing soft tissue infections | 0
conflict of interest none declared | 0
