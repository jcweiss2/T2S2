36 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
pregnant | 0 | 0 | Factual
admitted to hospital | 0 | 0 | Factual
recurrent vomiting | -72 | 0 | Factual
epigastric pain | -72 | 0 | Factual
uterine fibroid | -672 | 0 | Factual
weight loss | -672 | 0 | Factual
no change in bowel habits | 0 | 0 | Negated
no hematemesis | 0 | 0 | Negated
no rectal bleeding | 0 | 0 | Negated
no hematuria | 0 | 0 | Negated
no passing stones | 0 | 0 | Negated
using iron tablets | -672 | 0 | Factual
markedly dehydrated | 0 | 0 | Factual
drowsy | 0 | 0 | Factual
blood pressure 126/76 mmHg | 0 | 0 | Factual
pulse rate 94 min–1 | 0 | 0 | Factual
respiratory rate 30 min–1 | 0 | 0 | Factual
temperature 36.6°C | 0 | 0 | Factual
no lymphadenopathy | 0 | 0 | Negated
no thyromegaly | 0 | 0 | Negated
no edema | 0 | 0 | Negated
uterus size of 40 weeks | 0 | 0 | Factual
tender epigastric area | 0 | 0 | Factual
drowsy and hypotonic | 0 | 0 | Factual
brisk deep tendon reflexes | 0 | 0 | Factual
no obvious focal neurological sign | 0 | 0 | Negated
planter reflexes were down-going | 0 | 0 | Factual
chest and cardiovascular systems were unremarkable | 0 | 0 | Factual
hemoglobin 8.7 g/dl | 0 | 0 | Factual
WBCs 7000 μl–1 | 0 | 0 | Factual
platelets 445 000 μl–1 | 0 | 0 | Factual
ESR 109 mm/h | 0 | 0 | Factual
toxic granulation of WBCs | 0 | 0 | Factual
BUN 4.4 mmol/l | 0 | 0 | Factual
creatinine 59 μmol/l | 0 | 0 | Factual
HCO3 22 mmol/l | 0 | 0 | Factual
Na 138 mmol/l | 0 | 0 | Factual
Ca 4.8 mmol/l | 0 | 0 | Factual
uric acid 508 μmol/l | 0 | 0 | Factual
lactic acid 1.2 mmol/l | 0 | 0 | Factual
phosphorous 0.8 mmol/l | 0 | 0 | Factual
HIV serology was negative | 0 | 0 | Factual
calcium at 14 weeks’ gestation was 2.43 mmol/l | -504 | -504 | Factual
ALT 4 u/l | 0 | 0 | Factual
AST 11 u/l | 0 | 0 | Factual
ALP 150 u/l | 0 | 0 | Factual
total protein 72 g/l | 0 | 0 | Factual
albumen 30 g/l | 0 | 0 | Factual
cholesterol 4.05 mmol/l | 0 | 0 | Factual
triglyceride 3.59 mmol/l | 0 | 0 | Factual
PTH 3 pg/ml | 0 | 0 | Factual
TSH 0.68 mIU/l | 0 | 0 | Factual
free thyroxin 16.6 pmol/l | 0 | 0 | Factual
cortisol 1849 nmol/l | 0 | 0 | Factual
vitamin D 15 ng/ml | 0 | 0 | Factual
normal saline infusion | 0 | 24 | Factual
intramuscular calcitonin | 0 | 24 | Factual
transferred to medical intensive care unit | 0 | 24 | Factual
rupture membrane | 24 | 24 | Factual
urgent cesarean section | 24 | 24 | Factual
hemodialysis | 24 | 24 | Factual
bleeding | 24 | 24 | Factual
hypotension | 24 | 24 | Factual
blood transfusion | 24 | 24 | Factual
delivery of a baby girl | 24 | 24 | Factual
removal of uterine masses | 24 | 24 | Factual
histopathology report was consistent with leiomyoma | 24 | 24 | Factual
septicemia | 48 | 72 | Factual
septic shock | 48 | 72 | Factual
vasopressors | 48 | 72 | Factual
broad-spectrum antibiotics | 48 | 72 | Factual
postoperative laboratory test results | 72 | 72 | Factual
CT scan of the chest and pelvis showed no evidence of mass lesion | 72 | 72 | Factual
MRI of the brain showed evidence of infarcts | 72 | 72 | Factual
MRA revealed evidence of vasospasm | 72 | 72 | Factual
diffuse ischemic changes secondary to hypoxic insult | 72 | 72 | Factual
condition began to improve | 96 | 120 | Factual
discharged home | 168 | 168 | Factual
final diagnosis of humoral hypercalcemia associated with a uterine fibroid | 168 | 168 | Factual
serum calcium remained within the normal range | 168 | 744 | Factual