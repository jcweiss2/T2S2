19 years old | 0 | 0 
male | 0 | 0 
army officer | 0 | 0 
admitted to the hospital | 0 | 0 
fever | -120 | 0 
arthralgia | -120 | 0 
myalgia | -120 | 0 
headache | -120 | 0 
productive cough | -120 | 0 
yellowish sputum | -120 | 0 
chest heaviness | -120 | 0 
dyspnea | -120 | 0 
diarrhea | -120 | 0 
reduced oral intake | -120 | 0 
conscious | 0 | 0 
dehydrated | 0 | 0 
cold peripheries | 0 | 0 
febrile | 0 | 0 
temperature of 38.5°C | 0 | 0 
hypotensive | 0 | 0 
blood pressure of 81/53 mmHg | 0 | 0 
tachycardic | 0 | 0 
146 beats per minute | 0 | 0 
tachypnoeic | 0 | 0 
30 breaths per minute | 0 | 0 
oxygen saturation of 75-80% | 0 | 0 
coarse crepitation | 0 | 0 
tenderness at epigastric region | 0 | 0 
palpable liver | 0 | 0 
no cervical lymph nodes | 0 | 0 
no inguinal lymph nodes | 0 | 0 
no axillary lymph nodes | 0 | 0 
haemoglobin of 11.3 g/dL | 0 | 0 
low white blood cell count | 0 | 0 
0.5 × 10^6/L | 0 | 0 
neutrophil predominance | 0 | 0 
86.1% | 0 | 0 
platelet count of 80 × 10^6/L | 0 | 0 
C-reactive protein of 28.28 mg/dL | 0 | 0 
acute kidney injury | 0 | 0 
serum sodium of 137 mmol/L | 0 | 0 
serum potassium of 3.7 mmol/L | 0 | 0 
serum urea of 14 mmol/L | 0 | 0 
serum creatinine of 206 μmol/L | 0 | 0 
liver function tests normal | 0 | 0 
serum albumin of 22 g/dL | 0 | 0 
creatinine kinase of 351 IU/L | 0 | 0 
arterial blood gases on room air | 0 | 0 
pH of 7.378 | 0 | 0 
pCO2 of 37 mmHg | 0 | 0 
pO2 of 52.7 mmHg | 0 | 0 
O2 saturation of 89% | 0 | 0 
HCO3 of 21.7 mmol/L | 0 | 0 
Dengue NS-1 Antigen negative | 0 | 0 
IgG and IgM antibody negative | 0 | 0 
chest radiograph showed consolidation | 0 | 0 
right upper lobe consolidation | 0 | 0 
left lower lobe consolidation | 0 | 0 
diagnosis of severe community acquired pneumonia | 0 | 0 
acute kidney injury | 0 | 0 
resuscitation with normal saline | 0 | 12 
non-invasive ventilation | 0 | 12 
inotropic support | 12 | 72 
intravenous ceftriaxone | 0 | 48 
intravenous azithromycin | 0 | 48 
intubation | 12 | 12 
mechanical ventilation | 12 | 72 
bronchoscopy | 48 | 48 
haemoserous and greenish secretion | 48 | 48 
repeated chest radiograph | 48 | 48 
worsening consolidation | 48 | 48 
abscess formation | 48 | 48 
intravenous meropenem | 48 | 72 
intravenous cloxacillin | 48 | 72 
antiviral oseltamivir | 48 | 72 
continuous venous-venous haemofiltration | 48 | 72 
severe metabolic acidosis | 48 | 72 
oliguric acute kidney injury | 48 | 72 
persistent spiking of temperature | 48 | 72 
worsening of septic parameters | 48 | 72 
refractory hypotension | 48 | 72 
death | 72 | 72 
blood cultures negative | 0 | 72 
atypical bacterial serologies negative | 0 | 72 
Leptospiral serologies negative | 0 | 72 
Hepatitis B/C serologies negative | 0 | 72 
HIV serologies negative | 0 | 72 
respiratory viruses screening negative | 0 | 72 
tracheal aspiration positive for MDR Acinetobacter baumannii | 48 | 72 
bronchoalveolar lavage positive for MDR Acinetobacter baumannii | 48 | 72 
MDR Acinetobacter baumannii susceptible to polymyxin B | 48 | 72 
minimum inhibitory concentration of 0.5 μg/ml | 48 | 72 
MDR Acinetobacter baumannii resistant to penicillin group | 48 | 72 
MDR Acinetobacter baumannii resistant to ampicillin/sulbactam | 48 | 72 
MDR Acinetobacter baumannii resistant to third generation cephalosporins | 48 | 72 
MDR Acinetobacter baumannii resistant to fluoroquinolone | 48 | 72 
MDR Acinetobacter baumannii resistant to carbapenem group | 48 | 72 
PCR for carbapenemases genes NDM, OXA-23, OXA 24 or OXA-58 not performed | 0 | 72