54 years old | 0
male | 0
Korean | 0
admitted to the hospital | 0
jaundice | -168
body temperature 39.2℃ | 0
resting heart rate 90 beats per minute | 0
respiratory rate 16 breaths per minute | 0
blood pressure 125/80 mm Hg | 0
generalized erythematous maculopapular rash | 0
moist erosions on the patient's lips | 0
moist erosions on the buccal mucosa | 0
moist erosions on the oropharynx | 0
bilateral conjunctival injection | 0
hemoglobin 13.5 g/dL | 0
white blood cell count 8,630/mm3 | 0
eosinophils 0.11 | 0
C-reactive protein 4.1 mg/dL | 0
erythrocyte sedimentation rate 4.0 mm/hr | 0
aspartate aminotransferase (AST) 318 IU/L | 0
alanine transaminase (ALT) 650 IU/L | 0
prothrombin time (PT) 57% | 0
total bilirubin 8.4 mg/dL | 0
albumin 3.1 g/dL | 0
creatinine 0.8 mg/dL | 0
laboratory tests negative for hepatitis A | 0
laboratory tests negative for hepatitis B | 0
laboratory tests negative for hepatitis C | 0
subepidermal clefting | 0
bulla formation | 0
necrotic keratinocytes | 0
vacuolar degeneration | 0
infiltration of lymphocytes | 0
blood culture negative | 0
occupational exposure to TCE | -672
worked at a factory producing spoons | -672
urinary trichloroacetic acid level 22 mg/L | -336
diagnosis of hypersensitivity syndrome caused by TCE | 0
initiating intravenous methylprednisolone | 0
fever 40.2℃ | 0
regained strength | 12
AST 67 IU/L | 408
ALT 167 IU/L | 408
total bilirubin 4.2 mg/dL | 408
discharged | 408
prescribed prednisolone 60 mg once daily | 408
visited emergency department | 408 + 120
dyspnea | 408 + 120
left pneumonic infiltration | 408 + 120
pleural effusion | 408 + 120
hemoglobin 9.0 g/d | 408 + 120
white blood cell count 2,470/mm3 | 408 + 120
platelet count 135,000/mm3 | 408 + 120
AST 36 IU/L | 408 + 120
ALT 38 IU/L | 408 + 120
PT 34% | 408 + 120
total bilirubin 3.1 mg/dL | 408 + 120
blood culture yielded methicillin-sensitive Staphylococcus aureus | 408 + 120
transferred to the medical intensive care unit | 408 + 120
bradycardia | 408 + 126
asystole | 408 + 126
death | 408 + 126