72 years old | 0
male | 0
admitted to the hospital | 0
mechanical fall | -72
lying on the floor at home | -72
history of Stage IVA squamous cell carcinoma | -2176
completed concurrent chemoradiotherapy | -2176
weakness | 0
pain in right wrist | 0
pain in left hip | 0
epiphora | 0
pain in left eye | 0
limited range of motion of both hips | 0
minimal erythema | 0
palpable trace effusion | 0
tenderness to palpation | 0
matted eyelashes | 0
mucopurulent conjunctival secretions | 0
corneal edema | 0
hypopyon | 0
fibrinous membrane in pupil | 0
pupil fixed and non-reactive | 0
white blood cell count 6.6 K/cmm | 0
thrombocytopenia | 0
renal impairment | 0
procalcitonin 5.13 ng/mL | 0
blood cultures exhibited growth of Gram-positive cocci | 0
Group C Streptococcus dysgalactiae subsp. equisimilis identified | 0
ophthalmology consultation | 0
B scan ultrasound of the left eye | 0
vitreous debris | 0
aqueous and vitreous tap of left eye | 0
intravitreal injection of vancomycin and ceftazidime | 0
vitreous culture yielded growth of Streptococcus dysgalactiae subsp. equisimilis | 0
transthoracic echocardiography | 72
bicuspid aortic valve | 72
mild to moderate aortic regurgitation | 72
normal left ventricular function | 72
mild to moderate dilatation | 72
normal right ventricular size and function | 72
aortic valve vegetation | 144
anterior mitral valve leaflet vegetation | 144
transesophageal echocardiography | 216
small mobile vegetation on the non-coronary cusp of the aortic valve | 216
thickened aortic root | 216
echodensity in the posterior aspect of the aortic root | 216
moderate aortic valve vegetation | 216
mitral valve thickening | 216
mobile echodensity on the posterior mitral valve | 216
mild-moderate mitral valve regurgitation | 216
treated with vancomycin | 0
treated with penicillin G | 48
infective endocarditis | 0
left eye vision worsened | 48
intravitreal injection in left eye | 48
treated with topical trimethoprim/sulfamethoxazole | 48
treated with prednisolone acetate | 48
treated with atropine | 48
scheduled for vitrectomy | 120
no light perception in left eye | 120
vitrectomy cancelled | 120
orthopedic service examination | 0
no septic arthritis | 0
no fracture or dislocation | 0
no soft tissue swelling | 0
magnetic resonance imaging of thoracic and lumbar spine | 0
no evidence of infection | 0
otolaryngologists examination | 0
no infection or new lesions | 0
all blood cultures negative | 0
transferred to another facility | 240
aortic valve replacement | 288
acute heart failure | 288
hypoxic respiratory distress | 288
pulmonary edema | 288
BiPAP | 288
dobutamine | 288
prosthetic valve replacement | 312
aortic root abscess debrided | 312
transferred to general medicine floor | 336