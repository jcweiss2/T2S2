40 years old | 0
male | 0
admitted to a local hospital | 0
fever (39 °C) | 0
diarrhea | 0
oxygen saturation of 60% | 0
gradual onset of dyspnea | 0
confusion | 0
shock | 0
bleeding spots on the chest and abdomen | 0
florid spots on the lower limbs | 0
platelet count (PLT) of 26 × 109/L | 0
blood urea nitrogen (BUN) level of 13.9 mmol/L | 0
creatinine (CRE) level of 330 μmol/L | 0
urine protein level of 3+ | 0
positivity for the HFRS anti-IgM antibody | 0
history of hypertension | 0
usual blood pressure 160/100 mmHg | -8760
fatty liver | 0
diagnosed with HFRS | 0
treated with ventilator-assisted ventilation | 0
fluid replacement | 0
norepinephrine to increase the blood pressure | 0
admitted to the Department of Intensive Care | 0
septic shock | 0
decompensated metabolic acidosis | 0
AKI | 0
multiple organ failure | 0
continuous renal replacement therapy (CRRT) | 0
sedation and analgesia | 0
plasma transfusions | 0
platelet transfusions | 0
left nasal cavity filled with an expanded sponge | -24
left nasal cavity bleeding | -24
left nasal alar became purple and swollen | -12
massive nasal necrotic lesions | 0
microbial cultures from the lesion samples revealed growth of mucormycetes | 0
identified as Rhizopus oryzae complex | 0
bronchoalveolar lavage fluid culture confirmed Aspergillus growth | 0
PCR strains identified Aspergillus fumigatus | 0
bronchoalveolar lavage fluid galactomannan (GM) 1.29 | 0
serum GM 4.99 | 0
diagnosed with rhinomucormycosis | 0
pulmonary aspergillosis | 0
systemic caspofungin | 0
voriconazole | 0
caspofungin: loading dose: 70 mg/d | 0
caspofungin: post-35 mg/d | 0
voriconazole: loading dose: 400 mg/12 h | 0
voriconazole: post-100 mg/12 h | 0
nasal cavity rinsed with 10 mL saline | 0
kept dry for 1 h | 0
filled with sterile dressing containing 2.5 mg/mL amphotericin B for 4 h | 0
filled with sterile dressing containing 5% sodium bicarbonate for 1 h | 0
left nasal scab fell off | 288
large tissue defect remained | 288
computed tomography revealed no orbitocerebral involvement | 288
bronchoalveolar lavage fluid culture revealed no fungal growth | 288
lung imaging findings gradually returned to normal | 288
urine output recovered | 288
renal function recovered | 288
weaning from the ventilator | 264
discontinuation of caspofungin | 312
discontinuation of voriconazole | 336
recovered | 672
discharged | 672
