22 years old | 0
female | 0
admitted to the intensive care unit | 0
general malaise | -168
myalgia | -168
dyspnea | -168
subjective fevers | -168
anorexia | -168
nasal discharge | -168
congestion | -168
abdominal pain | -168
increased vaginal pain | -168
dysuria | -168
unprotected sex | -720
afebrile | 0
tachycardic | 0
hypotensive | 0
white blood cell count 6200/µL | 0
white blood cell count 19,500/µL | 0
platelet count 23,000/µL | 0
creatinine 1.33 mg/dL | 0
creatinine 0.5 mg/dL | 0
alanine transaminase 36 U/L | 0
aspartate transaminase 59 U/L | 0
alkaline phosphatase 466 U/L | 0
total bilirubin 2.9 mg/dL | 0
serum lactic acid level 4.9 mmol/L | 0
chest radiography bilateral pleural effusions | 0
CT abdomen and pelvis hepatic abscesses | 0
bile duct dilatation | 0
mild splenomegaly | 0
right sided Bartholin gland cyst | 0
ultrasound hepatic abscesses | 0
reactive gall bladder thickening | 0
Fusobacterium necrophorum growth | 0
meropenem started | 0
transferred to our hospital | 72
febrile (102.4°F) | 72
tachycardic | 72
tachypneic | 72
blood pressure 157/97 | 72
oxygen saturation 100% | 72
high flow nasal cannula | 72
lung crackles | 72
right upper quadrant abdominal tenderness | 72
labial erythema | 72
edema | 72
white blood cell count 14,700/µL | 72
hemoglobin 11 g/dL | 72
platelet count 16,000/µL | 72
erythrocyte sedimentation rate 31 mm/h | 72
serum lactate dehydrogenase 323 U/L | 72
alkaline phosphatase 129 U/L | 72
c-reactive protein 17.05 mg/dL | 72
fibrinogen 349 mg/dL | 72
haptoglobin 59 mg/dL | 72
COVID-19 PCR negative | 72
HIV negative | 72
urine gonorrhea and chlamydia PCR negative | 72
CT neck no abscess | 72
CT chest septic emboli | 72
multifocal pneumonia | 72
bilateral pleural effusion | 72
hepatic abscess worsening | 72
meropenem transitioned to piperacillin-tazobactam | 72
respiratory status improved | 72
transferred to general medicine ward | 144
nasal cannula | 144
thoracentesis | 192
pleural fluid removed 800 mL | 192
exudative pleural fluid | 192
fungal smear negative | 192
acid-fast stain negative | 192
gram stain 4+ granulocytes | 192
bacterial culture no growth | 192
CT chest abdomen pelvis multifocal pneumonia | 216
pleural effusions | 216
necrotizing pneumonia | 216
pulmonary abscess | 216
hepatic abscesses | 216
right perineal fluid collection | 216
VATS washout | 240
decortication | 240
pleural rind acid fast negative | 240
fibrinous pleuritis | 240
empyema | 240
cultures 1+ granulocytes | 240
pelvic examination | 240
right labial abscess | 240
incision and drainage | 240
clear serous fluid | 240
thick white caseous material | 240
gram stain 3+ granulocytes | 240
Candida albicans growth | 240
CT abdomen pelvis right iliac vein thrombus | 360
echocardiography no vegetations | 360
diagnosis of Lemierre syndrome | 360
ceftriaxone | 360
metronidazole | 360
discharged | 408
symptoms improved | 408
amoxicillin-clavulanate | 408
