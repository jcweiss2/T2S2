70 years old | 0
    male | 0
    admitted to the hospital | 0
    sudden headache | -48
    deteriorating consciousness | -48
    pancreatic tumor resection | -17520
    prostatic cancer resection | -17520
    body temperature 36.0°C | 0
    heart rate 79/min irregular | 0
    blood pressure 123/70 mmHg | 0
    oxygen saturation 100% (O2 10 l/min) | 0
    respiratory rate 12/min | 0
    Japan Coma Scale III-100 | 0
    Glasgow Coma Scale E1V2M5 | 0
    pupils 2 mm/4 mm | 0
    light reflex ±/± | 0
    left concomitant deviation | 0
    right paresis | 0
    white blood cell count 7800/µl | 0
    C-reactive protein 0.23 mg/dl | 0
    atrial fibrillation rhythm | 0
    multiple brain infarctions | 0
    no thrombus detected by transthoracic echocardiography | 0
    left atrial thrombus identified by transesophageal echocardiography | 0
    carotid echography not performed | 0
    cardiogenic cerebral infarction | 0
    conscious disturbance worsened | 0
    intubated | 0
    unfractionated heparin 15,000 U | 0
    edaravone 30 mg × 2 | 0
    fever 38.5°C | 24
    rapid drop of blood pressure | 28
    septic shock | 28
    white blood cell count 28,300/µL | 28
    hemoglobin 14.3 g/dL | 28
    platelet count 25.6 × 104/µL | 28
    total protein 6.2 g/dL | 28
    albumin 3.4 g/dL | 28
    total bilirubin 0.7 mg/dL | 28
    aspartate aminotransferase 22 U/L | 28
    alanine aminotransferase 16 U/L | 28
    lactase dehydrogenase 194 U/L | 28
    alkaline phosphatase 189 U/L | 28
    creatine kinase 114 U/L | 28
    blood urea nitrogen 11.0 mg/dL | 28
    creatinine 0.99 mg/dL | 28
    C-reactive protein 1.38 mg/dL | 28
    prothrombin time 79.0% | 28
    activated partial thromboplastin time 66.0 s | 28
    fibrinogen 686 mg/dL | 28
    S. pneumoniae detected in blood | 28
    S. pneumoniae detected in sputum | 28
    slight infiltration in lower right lung field | 28
    no spleen observed | 28
    spinal fluid test normal | 28
    community-acquired pneumonia | 28
    OPSI | 28
    ceftriaxone 2 g × 2 | 28
    IVIG 5 g × 3 days | 28
    fluid resuscitation | 28
    0.5 γ noradrenaline | 28
    mechanical ventilation | 28
    edaravone discontinued due to severe infection | 28
    condition improved | 28
    catecholamines reduced | 72
    extubated | 96
    free from mechanical ventilation | 96
    catecholamine-dependent condition prolonged | 96
    noradrenaline discontinued | 192
    unfractionated heparin 15,000 U/day continued | 192
    switched to warfarin | 192
    moved to different hospital for rehabilitation | 216
<|eot_id|>