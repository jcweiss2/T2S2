35 years old | 0
    female | 0
    history of Crohn’s disease | 0
    sepsis-like syndrome | 0
    cholestasis | 0
    noncaseating granulomatous hepatitis | 0
    low-grade fever | 0
    chills | 0
    nonspecific abdominal pain | 0
    nonbilious emesis | 0
    no cough | 0
    no dysuria | 0
    no skin rashes | 0
    CD status postright hemicolectomy in 2013 | -87600
    adhesion-related small bowel obstruction status postadhesiolysis in 2020 | -35040
    off disease-modifying therapy for last 5 years | -43800
    generalized anxiety disorders | 0
    bipolar disorders | 0
    ill appearance | 0
    toxic appearance | 0
    tachycardia (126 beats per minute) | 0
    hypotension (80/50 mmHg) | 0
    fever (38.8°C) | 0
    diffuse abdominal tenderness | 0
    no focal guarding | 0
    no rigidity | 0
    low hemoglobin (8.2 g/dl) | 0
    leukopenia (WCC 2.5 X 109/L) | 0
    thrombocytopenia (76 X 109/L) | 0
    elevated serum lactate (4.3 mmol/L) | 0
    elevated C-reactive protein (60.6 mg/l) | 0
    acute kidney injury | 0
    elevated serum creatinine (2.15 mg/dl) | 0
    high serum calcium (11.0 mg/dl) | 0
    normal total bilirubin (0.7 mg/dl) | 0
    elevated ALT (66 U/l) | 0
    elevated alkaline phosphatase (175 U/l) | 0
    negative urinalysis | 0
    unremarkable chest X-rays | 0
    admitted to intensive care unit | 0
    presumed intra-abdominal sepsis | 0
    acute cholecystitis | 0
    cholangitis | 0
    treated with fluid resuscitation | 0
    empiric antibiotics (vancomycin and piperacillin/tazobactam) | 0
    CT abdomen (mild gallbladder wall thickening, pericholecystic fluid) | 0
    no gallstones | 0
    no active Crohn’s flare-up | 0
    MRI (mild cholecystitis, no stones, normal biliary ducts) | 0
    continued fever despite antibiotics | 0
    cholecystectomy | 0
    acalculous cholecystitis | 0
    normal intraoperative cholangiogram | 0
    gallbladder histology (mild nonspecific acalculous cholecystitis) | 0
    worsening liver biochemistry postcholecystectomy | 96
    ALT increase (240 U/L) | 96
    ALP increase (200 U/L) | 96
    total bilirubin increase (6.2 mg/dl) | 96
    direct bilirubin (5.0 mg/dl) | 96
    CT and MRI (normal postoperative changes, no collections, normal biliary ducts) | 96
    ERCP (clear biliary ducts) | 96
    negative viral serologies | 96
    negative autoimmune screening | 96
    normal IgG, IgM, IgA | 96
    normal transferrin saturation | 96
    normal ferritin | 96
    normal ceruloplasmin | 96
    no hepatotoxic medications | 96
    hepatology consultation | 96
    liver biopsy (acute hepatitis, noncaseating granulomas, giant cells) | 96
    no primary biliary cirrhosis | 96
    no primary sclerosing cholangitis | 96
    no autoimmune hepatitis | 96
    negative infectious workup | 96
    negative AAFP stain | 96
    negative Giemsa stain | 96
    negative QuantiFERON gold assay | 96
    negative Coccidiosis serology | 96
    negative Brucella serology | 96
    negative Bartonella serology | 96
    negative Coxiella serology | 96
    negative Histoplasma urine antigen | 96
    hypercalcemia resolved | 96
    normalized renal function | 96
    low PTH | 96
    normal PTH-related peptide | 96
    normal Vitamin D3 1,25-OH | 96
    normal ACE levels | 96
    Chest CT (small ground-glass pulmonary nodules, no lymphadenopathy) | 96
    antibiotics discontinued on Day 14 | 336
    interdisciplinary discussions | 336
    oral steroids instituted | 336
    prednisone taper | 336
    discharged | 336
    clinical improvement | 432
    ALT normalization (70 U/l) | 432
    ALP normalization (69 U/l) | 432
    <|eot_id|>
    