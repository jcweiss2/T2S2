11 years old | 0
female | 0
febrile illness | -48
abdominal pain | -48
vomiting | -48
seizures | -48
repetitive focal to bilateral tonic-clonic seizures | -48
normal neurodevelopment | 0
unremarkable personal and family medical history | 0
admitted to ICU | 0
sedated | 0
intubated | 0
mechanically ventilated | 0
EEG showed slow background with extreme delta brushes | 48
extensive diagnostic work-up | 0
hyperproteinorrachy | 0
rhinovirus DNA in PCR panel on nasal exudate | 0
continuous convulsive seizures | 552
focal clonic jerks of the right hemibody | 552
bilateral clonic jerking | 552
seizure burden peaked | 624
abundant epileptiform EEG activity | 624
focal to bilateral tonic-clonic seizures | 624
brain MRI negative | 0
T2-FLAIR bilateral hyperintensity of the claustra | 168
T2-FLAIR hyperintensity of the left cuneus | 816
failure of anesthetics | 0
failure of antiseizure medications | 0
failure of immunotherapy | 0
ketogenic diet started | 768
anakinra started | 816
seizures reduced by 50% | 840
seizures stopped | 864
discharged from ICU | 1152
anakinra stopped | 1344
candida albicans sepsis | 1344
focal seizures persisted | 1344
IV midazolam | 1152
focal seizures became less frequent | 3264
transferred to rehabilitation | 3264
relapse of seizures | 5232
seizures controlled with IV midazolam | 5232
discharged home | 6480
lacosamide | 6480
phenobarbital | 6480
clobazam | 6480
weaned ketogenic diet | 6480
low carbohydrate diet | 6480
no clinical seizures | 15552
moderate intellectual disability | 15552
milder impact on verbal functioning | 15552
able to go back to school | 15552
support teacher | 15552