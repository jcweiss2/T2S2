history of coronary artery disease | -2160
history of myocardial infarction | -2160
history of ischemic dilated cardiomyopathy | -2160
pocket infection of cardiac resynchronization therapy defibrillator | 0
erythema and discomfort around left upper chest implant site | -720
edema and serosanguinous drainage | -720
oral amoxicillin treatment | -720
nonbacteremic | 0
afebrile | 0
severely reduced left ventricular systolic function | 0
ejection fraction of 20%–25% | 0
global hypokinesis of the left ventricle | 0
no evidence of vegetations | 0
leads scarred to lateral wall of superior vena cava | 0
transvenous lead extraction | 0
cardiac resynchronization therapy defibrillator pocket capsule dissected out | 0
device removed | 0
coronary sinus and right atrial leads extracted | 0
right ventricular lead extraction | 0
hypotensive | 0
large pericardial effusion | 0
emergency midsternotomy | 0
bleeding manually controlled with pressure | 0
cardiopulmonary bypass instituted | 0
5-mm tear in superior cavoatrial junction | 0
perforation in right atrium | 0
oozing hematoma at level of innominate vein | 0
lesions repaired with multiple 4-0 polypropylene sutures | 0
right ventricular lead capped and abandoned | 0
intra-aortic balloon pump placed | 0
multiple blood transfusions | 0
coagulopathy | 0
transfusions of cryoprecipitate, platelets, fresh frozen plasma, and factor VII | 0
chest closed | 0
severe cardiogenic shock | 24
multiorgan failure | 24
hypotensive | 24
vasopressin, epinephrine, and norepinephrine administration | 24
hypoxic respiratory failure | 24
mechanical ventilation | 24
liver failure | 24
albumin and multiple blood products | 24
broad-spectrum antibiotics | 24
oliguric | 24
continuous venovenous hemodialysis | 48
bilateral, symmetrical cyanotic changes | 72
vasopressor administration stopped | 72
upper- and lower-digit ischemia | 216
dry gangrene | 216
dull pain | 216
no ability to move fingers and toes | 216
bilateral stiffness | 216
2+ pitting edema | 216
nonexistent capillary refill time | 216
palpable 2+ peripheral pulses | 216
Doppler study showed flat waveforms | 216
intra-aortic balloon pump removed | 168
endotracheal tube removed | 168
albumin discontinued | 264
liver enzymes returned to normal limits | 264
kidney function improved | 984
hemodialysis stopped | 984
mental status improved | 984
necrotic lesions treated conservatively | 984
debridement | 648
negative-pressure wound therapy | 648
purulent, foul-smelling material from left infraclavicular operative site | 1296
transferred to facility | 1296
laser extraction of retained lead | 1392
pus drained from subfascial area | 1392
antibiotic regimen | 1392
transvenous implantable cardioverter-defibrillator system implanted | 1536
evaluation of hands and feet | 1536
black skin changes and demarcation lines | 1536
discharged to home health services | 1848
amputation and debridement of necrotic feet | 2556
amputation of fingers scheduled | 2556