3 years old | 0
    female | 0
    admitted to the hospital | 0
    fever | -168
    cough | -168
    respiratory distress | -168
    decreased mental status | -168
    positive rapid antigen test result | -120
    oseltamivir | -120
    condition deteriorated | -120
    difficult breathing | -120
    sleepiness | -120
    impending respiratory failure | 0
    decreased mental status | 0
    blood pressure 117/67 mmHg | 0
    heart rate 181 beats/min | 0
    respiratory rate 40/min | 0
    body temperature 37.5℃ | 0
    percutaneous oxygen saturation 91% | 0
    chest wall retraction | 0
    decreased left lung sounds | 0
    drowsy | 0
    intubated | 0
    pH 7.193 | 0
    PaCO2 53.9 mmHg | 0
    PaO2 30.3 mmHg | 0
    bicarbonate 20.3 mmoL/L | 0
    base excess -7.9 | 0
    pancytopenia | 0
    WBC count 710/µL | 0
    absolute neutrophil count 210/µL | 0
    hemoglobin 10.6 g/dL | 0
    platelets 81,000/µL | 0
    C-reactive protein 37.18 mg/dL | 0
    immunoglobulin G 399 mg/dL | 0
    high dose oseltamivir | 0
    intravenous immunoglobulin G | 0
    2009 H1N1 influenza virus detected | 0
    diffuse haziness in left lung | 0
    right upper lung infiltration | 0
    thoracentesis | 0
    turbid chocolate-colored fluid | 0
    chest tube insertion | 72
    increased pleural effusion | 72
    tracheal deviation | 72
    chest computed tomography | 144
    necrotizing pneumonia | 144
    significant left pleural effusion | 144
    persistent high fever 39.1℃ | 144
    leukocytosis | 144
    WBC count 24,250/µL | 144
    absolute neutrophil count 19,640/µL | 144
    broad spectrum antibiotics | 144
    cefotaxime | 144
    vancomycin | 144
    pneumothorax | 168
    chest tube replacement | 168
    waxed-and-waned pneumothorax | 168
    ventilator support | 168
    FiO2 1.0 | 168
    PEEP 5 cmH2O | 168
    TV 90 mL | 168
    percutaneous oxygen saturation near 90% | 168
    peak inspiratory pressure 23-34 cmH2O | 168
    meropenem | 168
    percutaneous oxygen saturation dropped to 77% | 168
    progressive respiratory failure | 168
    persistent purulent pleural effusion | 168
    recurrent massive pneumothorax | 168
    venovenous ECMO support | 168
    multidrug resistant Acinetobacter baumannii | 240
    Stenotrophomonas maltophilia | 240
    blood cultures positive | 240
    tracheal aspirate cultures positive | 240
    pleural fluid cultures positive | 240
    ECMO discontinuation | 240
    blood cultures negative | 432
    tracheal aspirate cultures positive | 432
    pleural fluid cultures positive | 432
    ECMO support duration 6 days | 168
    ventilator weaning | 888
    pH 7.371 | 888
    PaCO2 64.0 mmHg | 888
    PaO2 111.9 mmHg | 888
    bicarbonate 36.3 mmoL/L | 888
    base excess 9.2 | 888
    antibiotics combinations | 888
    isepamicin | 888
    minocyclin | 888
    rifampicin | 888
    ceftazidime | 888
    TMP-SMX | 888
    colistin | 888
    oseltamivir duration 23 days | 552
    mechanical ventilation weaning | 888
    antimicrobials discontinued | 1368
    chest tube removed | 1512
    discharged | 1512
    alert | 1512
    spontaneously breathing | 1512
    no respiratory symptoms | 1512
    chest radiograph improved | 1512
    