70 years old | 0
male | 0
unstable diabetes | 0
arterial hypertension | 0
bilateral bursa with pus discharge from a scrotal fistula | -24
fever | -24
altered general condition | -24
admitted to the hospital | 0
fever of 39° | 0
blood pressure 95/40 cmH2O | 0
heart frequency at 100 beats/minute | 0
testicular examination shows a large, warm, tender bursa | 0
inflammatory signs | 0
presence of an orifice and pus discharge | 0
WBC:1300 | 0
CRP: 340 mg/l | 0
creatinine: 14 mg/l | 0
Procalcitonin 100 ng/ml | 0
abdomino-pelvic scan showed a scrotal collection with air in the perineal and anterior abdominal | 0
received an antibiotic | 0
debridement with drainage of the abscess and resection of areas of necrosis | 2
transferred to the intensive care unit | 2
treated with vasoactive drugs | 2
antiobiotherapy | 2
bourgeoning of the scrotal tissue | 72
ulcerated, bourgeoning lesion on the glans penis | 72
biopsy of the glans | 72
anatomopathological results of the biopsy showed squamous cell carcinoma of the penis | 72
ingual adenopathy not found | 72
MRI of the penis showed the presence of a tumor of the penis extending to the cavernous cavities and the urethra | 72
total penectomy with perineostomy | 96
evolution was favorable | 120
put under surveillance | 120