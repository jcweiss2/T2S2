13 years old | 0
male | 0
admitted to the hospital | 0
fever | -24
limping | -24
left-sided knee pain | -24
knee without visible changes | -24
pain and tenderness at the infrapatellar ligament | -24
elevated leucocytes | -24
elevated C-reactive protein (CRP) | -24
radiography of the knee and leg was normal | -24
sent home | -24
continued to be febrile | -24
admitted to the pediatric department | 0
suspicion of soft tissue infection surrounding the knee | 0
ultrasound of the knee was normal | 24
staphylococci were cultured from blood | 72
IV vancomycin treatment was initiated | 72
knee was red and swollen | 72
cutaneous micro-ulcerations | 72
MRI showed synovitis with knee joint effusion | 72
signs of medullary osteomyelitis in the proximal tibia | 72
subperiostal fluid accumulation | 72
elevated CRP | 72
elevated sedimentation rate (SR) | 72
acute arthroscopy with synovectomy and lavage of the knee joint | 72
cultures from the medullary canal grew MRSA | 72
cultures from blood grew MRSA | 72
cultures from nasal swaps grew MRSA | 72
biopsy materials from the knee grew MRSA | 72
MRSA strain was positive for PVL | 72
wounds were debrided every other day | 120
pain increased | 120
CRP and leucocytes continued to rise | 120
MRI showed progression of the infection | 168
renewed surgical debridement | 168
patient became septic | 168
developed multiple bilateral pulmonary infiltrates | 168
admitted to the ICU | 168
oral linezolid was added to the antimicrobial treatment | 168
patient’s general condition improved | 192
returned to the orthopedic ward | 192
clinical and biochemical improvement continued | 240
CRP rose again | 360
MRI showed a new subperiostal abscess | 360
progression of the osteomyelitis | 360
renewed surgery | 360
patient’s condition improved | 360
discharged | 1176
followed in the outpatient clinic | 1176
frequent clinical, biochemical, and radiological controls | 1176
osteomyelitis progressed radiologically | 1176
follow-up MRI | 1260
supplemented by computer tomography (CT) | 1260
bone and leukocyte scintigraphy | 1260
no active infection | 1260
radiological signs eventually subsided | 1512
plain radiography showed a normal tibia | 2112
fever persisted for 51 days | 0
CRP and SR were elevated for 23 weeks | 0