23-year-old pregnant Caucasian woman | 0
referred for fetal echocardiogram at 20 weeks gestation | -1680
congenital heart disease | 0
DORV with normally related great arteries | 0
remote VSD | 0
moderate to severe hypoplastic mitral valve | 0
hypoplastic left ventricle | 0
APV syndrome | 0
to-and-fro flow across dysplastic and rudimentary pulmonary valve tissue | 0
moderate degree of stenosis | 0
peak velocity of 3.0 m/s across rudimentary pulmonary valve tissue | 0
severely dilated main and branch pulmonary arteries | 0
below normal right ventricular systolic function | 0
no evidence of ductus arteriosus | 0
polyhydramnios | 0
amnioreduction | 0
22q11.2 deletion | 0
DiGeorge syndrome | 0
delivered at 36 weeks gestation | -576
cesarean section | -576
breech position | -576
premature rupture of membranes | -576
severe polyhydramnios | -576
birth weight 2300 grams | 0
cyanotic at birth | 0
apneic at birth | 0
intubation | 0
initial blood gas pH 7.17 | 0
pCO2 69 | 0
pO2 21 | 0
oxygen saturations 70% | 0
admission to cardiovascular intensive care unit | 0
hypoxic on 100% fractional inspired oxygen | 0
inhaled nitric oxide | 0
prone positioning | 0
profoundly hypoxic | 0
cyanotic female neonate | 0
dysmorphic features consistent with 22q.11 deletion | 0
to-and-fro murmur along left sternal border | 0
postnatal transthoracic echocardiogram | 0
DORV with sub-aortic VSD | 0
side-by-side great arteries | 0
aortic-mitral fibrous discontinuity | 0
severely hypoplastic mitral valve | 0
z-score −5.1 | 0
minimal antegrade flow | 0
non-apex forming left ventricle | 0
thickened and dysplastic aortic valve leaflets | 0
normal annular measurements | 0
aortic valve annulus 0.9 cm | 0
z-score +3.2 | 0
aortic sinuses 1.22 cm | 0
z-score +3 | 0
no evidence of coarctation of aorta | 0
aortic isthmus 0.4 cm | 0
z-score −1.2 | 0
dysplastic and rudimentary pulmonary valve leaflets | 0
mild valvar stenosis | 0
severe/free insufficiency | 0
to-and-fro flow on color Doppler | 0
severely dilated main pulmonary artery | 0
13 mm | 0
z-score +5.42 | 0
severely dilated branch pulmonary arteries | 0
LPA 7.5 mm | 0
z-score +3.99 | 0
RPA 8 mm | 0
z-score +4.21 | 0
dilated right ventricle | 0
hypertrophied right ventricle | 0
severely depressed systolic function | 0
fractional shortening 19% | 0
partially restrictive atrial septum | 0
left to right shunting | 0
refractory cardiogenic shock | 0
severe hypoxemia | 0
surgical intervention within first 12 hours of life | 12
atrial septectomy | 12
branch pulmonary artery plication | 12
over sewing of main pulmonary artery | 12
placement of right 3.5 mm modified Blalock-Taussig"Thomas shunt | 12
failed to separate from cardiopulmonary bypass | 12
ongoing severe ventricular dysfunction | 12
transitioned to ECMO support | 12
hemothorax | 12
acute kidney injury | 12
required continuous renal replacement therapy | 12
profoundly immunocompromised | 12
severe lymphopenia | 12
hypogammaglobinemia | 12
developed septic shock | 24
Serratia marcescens septicemia | 24
abdominal compartment syndrome | 24
requiring abdominal decompression | 24
washout | 24
continued to deteriorate hemodynamically | 24
multi-organ failure | 24
profound neurological impairment | 24
decision of comfort care | 24
died on post-operative day 31 | 744
