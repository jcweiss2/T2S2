48 years old | 0
male | 0
chronic pancreatitis | 0
alcohol dependency | 0
septic shock | 0
cellulitic, oedematous and mottled discoloration of genitalia and perineum | 0
Fournier’s Gangrene | 0
radical debridement | 0
urology | 0
plastic surgery | 0
general surgery | 0
copious amounts of pus | 0
left inguinal canal | 0
large left-sided retroperitoneal collection | 0
two large drains placed | 0
peritoneal cavity examination | 0
no intra-peritoneal collection | 0
computed tomography scan | 0
acute-on-chronic pancreatitis | 0
focal necrosis at head of pancreas | 0
fluid tracking from pancreas into retroperitoneum | 0
subcutaneous emphysema in left flank | 0
inotropic support | 0
intravenous antibiotic therapy | 0
further debridement | 24
medial thigh pouches created | 24
testes | 24
wounds dressed with vacuum-assisted closure device | 24
polymicrobial growths isolated | 24
piperacillin/tazobactam | 24
histology confirmed necrotizing fasciitis | 24
3-week course of intravenous therapy | 48
switched to oral antibiotics | 168
acute pancreatitis managed conservatively | 0
nasogastric feeding | 0
diabetes mellitus type 2 | 0
oral treatment | 0
multiple debridements | 72
VAC changes | 72
abdomino/perineal skin defect ready for resurfacing | 168
split-skin grafting | 168
100% graft uptake | 192
discharged | 192
follow-up review | 384
excellent recovery | 384