76 years old | 0
male | 0
Caucasian | 0
admitted to the hospital | 0
bloody diarrhea | -96
intermittent abdominal pain | -96
vomiting | -96
dizziness | -96
generalized weakness | -96
watery foul-smelling diarrhea | -216
weight loss | -216
celiac disease | -4380
gluten-free diet | -4380
non-compliant with gluten-free diet | -672
afebrile | 0
tachycardic | 0
severely hypotensive | 0
cachectic | 0
severely dehydrated | 0
hyperactive bowel sounds | 0
diffuse abdominal tenderness | 0
microcytic hypochromic anemia | 0
metabolic acidosis | 0
hypoalbuminemia | 0
hypokalemia | 0
acute renal failure | 0
severe coagulopathy | 0
septic shock | 0
gastrointestinal infection | 0
hemolytic uremic syndrome | 0
gastrointestinal malignancy | 0
ischemic colitis | 0
intravenous fluids | 0
antibiotics | 0
sodium bicarbonate drip | 0
fresh frozen plasma | 0
electrolyte supplementation | 0
emergent hemodialysis | 0
hypotension improved | 24
anion-gap metabolic acidosis improved | 24
ARF improved | 24
severe coagulopathy improved | 24
ferritin level | 24
low serum iron | 24
normal total iron-binding capacity | 24
low iron saturation | 24
thyrotropin | 24
vitamin B12 | 24
folate | 24
total bilirubin | 24
lactate dehydrogenase | 24
peripheral blood smear | 24
blood cultures | 24
urine cultures | 24
stool cultures | 24
fecal leukocytes | 24
Clostridium difficile toxin PCR assay | 24
ova and parasites | 24
intravenous antibiotics discontinued | 48
colonoscopy | 48
esophagogastroduodenoscopy | 48
normal colonic and rectal mucosa | 48
flattened mucosa | 48
mucosal nodularity | 48
duodenal biopsies | 48
active chronic inflammation | 48
intraepithelial lymphocytosis | 48
subtotal villous blunting | 48
celiac crisis | 48
intravenous vitamin K | 48
parenteral nutrition | 48
methylprednisolone | 48
transferred to general medicine floor | 120
gluten-free diet | 120
oral budesonide | 120
oral steroid discontinued | 240
discharged | 240
follow-up | 8760
substantial improvement | 8760
asymptomatic | 8760