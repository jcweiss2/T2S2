38 years old | 0
female | 0
13th week of pregnancy | 0
abdominal discomfort | -24
nausea | -24
vomiting | -24
no fever | -24
no vaginal discharge | -24
admitted to the emergency room | 0
evaluated in the Obstetric Emergency Department | 0
discharged home | 0
returned to the ER | 144
persistent abdominal pain | 144
nausea | 144
vomiting | 144
tachycardic | 144
diffuse abdominal pain | 144
guarding on the right quadrants | 144
neutrophilia | 144
low prothrombinemia | 144
acute renal failure | 144
high procalcitonin | 144
high c-reactive protein | 144
abdominal ultrasound | 144
moderate fluid in all quadrants | 144
good foetal vitality | 144
surgical consultation | 144
hypotension | 144
general abdominal guarding | 144
hyperlacticaemia | 144
hypokalaemia | 144
hyperglycaemia | 144
septic shock with an abdominal source | 144
emergency exploratory laparotomy | 144
generalised purulent peritonitis | 144
perforated acute appendicitis | 144
appendicectomy | 144
abdominal washing | 144
laparostomy | 144
admitted to the Intensive Care Unit | 144
septic shock | 144
need for vasopressor therapy | 144
need for dialysis | 144
intravenous piperacillin-tazobactam antibiotherapy | 144
laparostomy revision | 192
marked bowel oedema | 192
bowel distention | 192
mild intraabdominal soiling | 192
further peritoneal lavage | 192
new laparostomy with progressive closure technique | 192
surgical revision | 240
abdominal cavity primary closed | 240
antibiotherapy adjusted | 288
piperacillin-tazobactam suspended | 288
amoxicillin with clavulanic acid started | 288
transferred to the obstetrics ward | 432
discharged home | 336
elective caesarean section | 1008
gave birth to a healthy child | 1008
post-partum follow-up consultation | 1344
ventral hernia | 1344
child thriving without neurological or other impairments | 1344