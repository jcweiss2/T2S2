54 years old | 0
man | 0
presented to the hospital with melena | 0
hemoglobin of 6.7 g/dL | 0
history of transhiatal esophagectomy | -78840
left neck anastomosis | -78840
esophageal adenocarcinoma | -78840
esophagogastroduodenoscopy | 0
5-cm clean-based ulcer on the anterior surface of the gastric conduit above the diaphragmatic impression | 0
suspected ischemic etiology | 0
biopsies taken of the ulcer edge | 0
reactive foveolar mucosa | 0
intraepithelial lymphocytosis | 0
fibrinopurulent exudate | 0
no dysplasia | 0
size of the ulceration | 0
suspicion of post-esophagectomy complication | 0
outpatient surgical referral | 0
discharged on proton pump inhibitors | 0
presented with hematemesis | 720
hemoglobin nadir of 4.8 g/dL | 720
esophagogastroduodenoscopy in the intensive care unit | 720
deeper, hematin-stained ulcer base | 720
rhythmic pulsations corresponding to cardiac contractions | 720
pulsations suggested ulcer may be abutting a cardiac ventricle | 720
chest computed tomography | 720
suspicion of ulcer erosion to the heart | 720
urgent thoracic surgery consult | 720
gastrocardiac fistula confirmed | 720
intraoperative visualization of a large defect in the ventricular wall arising from the gastric conduit | 720
repaired using a bovine pericardial patch | 720
multiple short-term complications after esophagectomy | -78840
failure to wean from mechanical ventilation | -78840
pneumonia | -78840
reintubation | -78840
sepsis | -78840
pulmonary edema | -78840
deep wound infection | -78840
gastrocardiac fistula | 720
secondary to ischemia | 720
radiation | 720
peptic ulcer disease | 720
recurrent malignancy | 720
Candida albicans infection | 720
severe peptic ulcer disease | 720
trauma | 720
gastrointestinal bleeding | 720
intermittent bleeding via the fistula | 720
endoscopy reveals a gastric ulcer on the cardiac surface | 720
clot within a pulsatile ulcer base | 720
acute-onset and rapidly progressive deterioration due to exsanguination through the fistula | 720
surgical repair techniques | 720
closing the defect using sutures | 720
pericardial patches | 720
endoscopic findings can be variable | 720
appropriate radiologic studies | 720
surgical exploration | 720
timely diagnosis | 720
surgical management crucial to good outcomes | 720
biopsies taken of the ulcer edge |2 0
