40 years old | 0
female | 0
admitted to the emergency department | 0
fever | -72
minor headache | -72
abdominal pain | -72
postpartum care | -504
cesarean section | -504
neck swelling | -264
needle aspiration | -264
thyroid gland examination | -264
no specific findings in thyroid gland | -264
vital signs measured | 0
body temperature 40.6 ℃ | 0
blood pressure 100/48 mmHg | 0
heart rate 100 bpm | 0
respiratory rate 18 breaths/min | 0
no specific findings in thyroid gland | 0
no neck stiffness | 0
no tonsil hypertrophy | 0
no abdominal tenderness | 0
no abnormal breath sounds | 0
no costal spine angle tenderness | 0
no signs of infection at cesarean section site | 0
no signs of infection at thyroid fine-needle aspiration site | 0
colposcopy performed | 0
no specific findings in colposcopy | 0
bicytopenia | 0
hemoglobin 14.0 g/dL | 0
platelets 133000/μL | 0
absolute neutrophil count 2512/μL | 0
total bilirubin level 0.3 mg/dL | 0
liver enzyme level measurement | 0
aspartate transaminase 65 U/L | 0
alanine transaminase 35 U/L | 0
thyroid function test | 0
T3 65.1 ng/dL | 0
free T4 0.88 ng/dL | 0
urinalysis | 0
one white blood cell/high-powered field | 0
C-reactive protein level 4.46 mg/dL | 0
chest radiograph normal | 0
abdominal computed tomography | 0
no prominent infectious focus | 0
antipyretic drug administered | 0
fever subsided | 0
vital signs remained stable | 0
discharged | 96
broad-spectrum antibiotics prescribed | 96
referral to infectious disease outpatient department | 96
returned to emergency department | 120
fever 38 ℃ | 120
decreased blood pressure 60/30 mmHg | 120
thrombocytopenia | 120
platelets 94000/μL | 120
total bilirubin level 3.1 mg/dL | 120
liver enzyme levels | 120
aspartate transaminase 202 U/L | 120
alanine transaminase 444 U/L | 120
renal function indicators | 120
blood urea nitrogen 42.1 mg/dL | 120
creatinine 3.35 mg/dL | 120
multiorgan failure | 120
ferritin level 3429.0 μg/L | 120
triglyceride level 957 mg/dL | 120
admitted to intensive care unit | 120
broad-spectrum antibiotics administered | 120
steroids administered | 120
high-dose steroid regimen not administered | 120
bone marrow biopsy performed | 120
hemophagocytic lymphohistiocytosis diagnosed | 120
thrombocytopenia worsened | 120
serum ferritin levels increased | 120
condition rapidly deteriorated | 120
died | 144
hematochezia | 144
disseminated intravascular coagulation | 144