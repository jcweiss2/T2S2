43 years old | 0
African American | 0
male | 0
admitted to the hospital | 0
uncontrolled HIV | -6720
nonadherence to antiretroviral therapy | -6720
chronic hepatitis B infection | -6720
progressive confusion | -168
fevers | -168
upper respiratory symptoms | -168
rhinorrhea | -168
denies cough | -168
denies shortness of breath | -168
denies chest pain | -168
denies headache | -168
denies abdominal pain | -168
HIV diagnosed | -5040
lost to follow-up | -5040
HIVAN | -3360
pneumocystis pneumonia | -3360
positive M184V mutation | -3360
ART treatment | -3360
abacavir | -1680
dolutegravir | -1680
lamivudine | -1680
poor adherence | -1680
inconsistent follow-up | -1680
last known CD4 count | -720
febrile | 0
tachycardic | 0
cachexia | 0
oral thrush | 0
non-blanching maculopapular rashes | 0
confusion | 0
somnolence | 0
pancytopenia | 0
WBC | 0
neutrophils | 0
lymphocytes | 0
monocytes | 0
hemoglobin | 0
platelets | 0
acute kidney injury | 0
serum creatinine | 0
lactate | 0
liver function tests | 0
AST | 0
ALT | 0
HIV viral load | 0
CD4 count | 0
reactivated chronic HBV | 0
HBcAb IgM | 0
HBcAb IgG | 0
HBsAg | 0
HBsAb | 0
HBV viral load | 0
empiric treatment for meningitis | 0
vancomycin | 0
ceftriaxone | 0
acyclovir | 0
ampicillin | 0
fluconazole | 0
LP | 24
cryptococcal meningitis | 24
seizures | 96
intubation | 96
transfer to the intensive care unit | 96
elevated ferritin | 96
elevated triglycerides | 96
elevated fibrinogen | 96
elevated soluble IL-2 receptor alpha | 96
HLH considered | 96
dexamethasone | 192
dolutegravir | 192
emtricitabine-tenofovir | 192
improved progressively | 192
discharged | 504
HIV viral load | 1008
HBV viral load | 1008
outpatient follow-up | 1008