Event | Time
found to have a segment-V space-occupying lesion in the liver | -8760
transarterial embolization | -8760
began taking sorafenib | -4320
stopped sorafenib due to dizziness, skin ulcers, and other symptoms | -3024
CT scan found enlarged lesions in liver segment V | -2592
radiation therapy performed | -2592
history of hepatitis B | -8760
serological tests for various viruses | -8760
donor suffered brain death from a car accident | -8760
HLA matching of donor and recipient | -8760
transplantation process smooth | 0
59 years old | 0
female | 0
Piggyback LT performed | 0
developed acute renal failure and a hematoma around the liver | 0
received intravenous administration of hepatitis B immunoglobulin | 24
received immunosuppressive drugs | 24
continuous hemodialysis and intermittent infusion of blood products | 24
active bleeding in the abdominal cavity ceased | 24
renal function gradually recovered | 24
pathological analyses confirmed diagnosis of HCC | 24
massive tumor necrosis observed | 24
liver function began to improve | 240
developed regular and repeated fevers | 240
serum PCT levels began to rise | 240
serum PCT levels dropped | 312
blood cultures were negative | 312
cytomegalovirus, Epstein–Barr virus were negative | 312
rash advanced into erythematous macules and papules | 432
sputum culture suggested presence of infections | 456
changed tacrolimus administration to sirolimus | 480
added mycophenolate mofetil | 480
abdominal incision split and was sutured again | 744
performed bone marrow aspiration | 800
bone marrow pathology report revealed no special lesions | 800
FISH analysis of peripheral blood detected donor lymphocytes | 800
skin biopsy specimens exhibited acute lt-GVHD | 800
assembled multidisciplinary team (MDT) | 800
continued to use steroids, tacrolimus, G-CSF, and anti-infective therapy | 800
rash significantly reduced | 800
general condition continued to deteriorate | 800
serum ferritin levels increased | 800
esophageal and oral ulcers worsened | 800
temperature rose to 39.4°C, experienced hallucinations | 944
succumbed to septic shock and MODS | 1320