1½ year-old male child | 0
admitted to the Pediatric Intensive Care Unit | 0
fever | -360
loose motions | -360
cough | -240
cold | -240
productive cough | -240
post-tussive vomiting | -240
breathlessness | -240
measles at 8½ months old | -4320
incomplete immunization | -4320
OPV vaccine | -4320
BCG vaccine | -4320
lethargic | 0
pale | 0
dusky | 0
shallow respiration | 0
pulse rate 130/minute | 0
bounding pulse | 0
blood pressure 100/65 mm Hg | 0
depressed anterior fontanel | 0
dry tongue | 0
pallor | 0
no icterus | 0
no edema | 0
no cyanosis | 0
no clubbing | 0
no lymphadenopathy | 0
no skin rashes | 0
altered sensorium | 0
generalized hypotonia | 0
sluggish reflexes | 0
flexed plantar | 0
lost skin turgor | 0
malnourished | 0
protein energy malnutrition (PEM) | 0
diagnosed with diarrhea | 0
severe dehydration | 0
respiratory infection | 0
hemoglobin 11g% | 0
leukocytosis | 0
thrombocytopenia | 0
negative peripheral smear for malarial parasite | 0
normal liver function tests | 0
normal renal function tests | 0
negative Widal test | 0
normal chest X-ray | 0
blood culture | 0
stool culture | 0
greenish yellow liquid stool | 0
mucus in stool | 0
no blood in stool | 0
no parasitic elements in stool | 0
25–30 pus cells/high power field | 0
no red blood cells in stool | 0
no ova in stool | 0
no cysts of parasites in stool | 0
IV fluids | 0
Inj. Cefotaxime | 0
Inj. Amikacin | 0
Inj. Calcium gluconate | 0
IV IgG | 0
ventilator on admission | 0
Inj. Metronidazole added after 4 days | 96
respiratory symptoms subsided after 2 weeks | 336
ventilator taken off after 2 weeks | 336
total protein 5.1g% after 3 weeks | 504
albumin 2.6g% after 3 weeks | 504
hemoglobin reduced to 8.7g% after 3 weeks | 504
leukocytosis persisted after 3 weeks | 504
stool sample sent after 7 days | 168
Gram stain for Campylobacter negative | 168
Campylobacter Charcoal Differential Agar culture | 168
MacConkey agar culture | 168
V. vulnificus identified | 168
lactose-fermenting colonies | 168
oxidase-positive colonies | 168
halophilic vibrio | 168
sensitive to amikacin | 168
resistant to amoxicillin-clavulanic acid | 168
resistant to cefotaxime | 168
resistant to nalidixic acid | 168
resistant to co-trimoxazole | 168
resistant to tetracycline | 168
resistant to norfloxacin | 168
another stool culture after 4 days | 96
Klebsiella pneumoniae in ET secretions | 168
Acinetobacter species in ET secretions | 168
sensitive to imipenem | 168
sensitive to netilmycin | 168
Inj. Imipenem started | 168
Inj. Ciprofloxacin started | 168
Inj. Promethazine every 6 hours | 168
nebulization with ipratropium bromide | 168
transferred to ward after 1 month | 672
Inj. Amikacin in ward for 13 days | 672
discharged | 672
no complaints at discharge | 672
stable condition at discharge | 672
