65 years old | 0
African American | 0
female | 0
BMI 26.5 | 0
daily smoker | 0
history of peptic ulcer disease | 0
treated with omeprazole | 0
surgical history of hysterectomy | 0
admitted to the hospital | 0
complaints of worsening left sided abdominal pain | -336
nausea | -336
emesis | -336
hematochezia | -336
anorexia | -336
10-pound weight loss | -336
focalized peritoneal signs | 0
elevated white blood count | 0
potassium of 3.0 mmol/L | 0
albumin of 2.3 g/dL | 0
sigmoid diverticulitis | 0
pericolonic abscess | 0
treated with intravenous levofloxacin | 0
treated with metronidazole | 0
drain placement | 0
purulent fluid drained | 0
streptococcus viridans | 0
gram negative rods | 0
proteus species | 0
open Hartmann’s operation | 72
perforated diverticulitis | 72
serositis | 72
abscess formation | 72
fibrous adhesions | 72
fat necrosis | 72
granulation tissue | 72
negative for malignancy | 72
peri-operative antibiotics | 72
IV cefepime | 72
IV metronidazole | 72
mild hypotension | 24
tachycardia | 24
fluid resuscitation | 24
epidural infusion suspended | 24
clear liquid diet | 24
minimal intake | 24
no evidence of bowel function | 24
epidural analgesic catheter removed | 96
total parenteral nutrition | 120
hyponatremia | 168
hypochloremia | 168
bilateral adrenal enlargement | 192
bilateral adrenal gland hemorrhage/infarction | 192
low cortisol level | 192
random serum cortisol level | 192
hydrocortisone sodium succinate | 192
clinical status improved | 216
blood pressure stabilized | 216
heart rate stabilized | 216
return of bowel function | 216
discharged to a rehabilitation facility | 336
steroids tapered down | 336
prednisone | 336
follow up | 744
steroid dependence | 1056
no signs of adrenal recovery | 1056
hydrocortisone | 1056
continued on hydrocortisone | 1056