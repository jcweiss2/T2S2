64 years old | 0
    male | 0
    human immunodeficiency virus (HIV)/AIDS | 0
    CD4 count on admission <10 cells/mm3 | 0
    antiretroviral therapy | 0
    Kaposi Sarcoma | 0
    treated with radiation | 0
    pancytopenia | 0
    managed with thrice weekly filgrastim | 0
    left orbital apex syndrome | 0
    Aspergillus fumigatus sinusitis | 0
    managed initially on isavuconazonium sulfate | 0
    admitted to our facility for acute management of a suspected invasive mold infection | 0
    isavuconazonium sulfate discontinued | 0
    liposomal amphotericin-b started | 0
    voriconazole started | 0
    Aspergillus fumigatus recovered from surgical cultures | 0
    liposomal amphotericin-b discontinued | 0
    voriconazole changed to posaconazole 300 mg daily | 312
    hospital day 13 | 312
    hospital day 20 | 480
    fever of 39.9°C | 480
    elevated lactate of 2.6 mmol/L | 480
    absolute neutrophil count greater than 1000 cells/mm3 | 480
    blood cultures obtained | 480
    urinalysis | 480
    chest x-ray | 480
    increasing drainage from KS lesions on the thigh | 480
    considered as a potential infection source | 480
    broad empiric antibiotic therapy initiated with IV vancomycin 1250 mg IV every 12 hours | 480
    broad empiric antibiotic therapy initiated with cefepime 2000 mg IV every 8 hours | 480
    encephalopathy | 480
    rigors | 480
    persistent fever | 480
    hypotension | 480
    tachypnea | 480
    cefepime changed to piperacillin/tazobactam 4.5 g extended IV infusion every 8 hours | 480
    IV fluid bolus given | 480
    concern for cefepime related encephalopathy | 480
    Wound Care Team consulted | 480
    right thigh KS lesion with increased sloughing and drainage | 480
    musty odor | 480
    hospital day 22 | 528
    blood culture sets positive for P. mendocina | 528
    PICC line removed | 504
    catheter tip culture | 504
    repeat blood cultures | 504
    bacterial growth not detected | 504
    antibiotic susceptibilities requested for cefepime | 528
    antibiotic susceptibilities requested for ceftazidime | 528
    antibiotic susceptibilities requested for levofloxacin | 528
    antibiotic susceptibilities requested for meropenem | 528
    piperacillin-tazobactam Etest strips unavailable | 528
    antibiotic therapy adjusted to ceftazidime | 528
    total 10-day course from first negative blood culture | 528
    ultimate source of infection unclear | 528
    open wound (no cultures obtained from this site) | 528
    blood cultures cleared quickly | 528
    infection successfully treated | 528
    concern for cefepime related encephalopathy | 528
    inability to document in vitro susceptibility of piperacillin-tazobactam | 528
    unnecessary anaerobic coverage | 528
    patient received all treatment for infection during 44-day total hospital stay | 1056
    successfully discharged | 1056

    