Here is the table of events and timestamps:

18 years old | 0
male | 0
hepatitis C-related cirrhosis | 0
recurrent hepatic encephalopathies | 0
chronic portal vein thrombosis | 0
underwent LT | 0
construction of an end-to-side anastomosis of the donor portal vein to the superior mesenteric vein | 0
construction of an end-to-end bile duct anastomosis | 0
construction of an iliac conduit | 0
massive venous bleeding from local varices | -24
recovered well after surgery | -24
normal liver graft function | -24
five months after LT, stenosis of the bile duct anastomosis | -120
biliary leakage | -120
elevated liver enzymes in a cholestatic pattern | -120
treated with a pigtail | -120
six weeks later, a FCSCEMS was inserted | -84
persisting leakage | -84
no further signs of leakage after stent extraction | -84
hepatitis C reinfection | -84
recurrent stenosis of the biliary anastomosis | -84
treated with ERCP | -84
balloon dilatations | -84
placements of a total of 7 pigtails | -84
stent placements | -84
biopsy-proven significant fibrosis | -12
treated with pegylated interferon and ribavirin | -12
thirty-four months after LT | -12
scheduled for an elective ERCP | -12
elective ERCP | -12
biliary pigtail exchange | -12
large portobiliary fistula at the site of the anastomosis | -12
slight hemobilia from the papilla | -12
placed a FCSEMS inside the bile duct | -12
septic shock | 48
admitted to the intensive care unit | 48
hemodynamic support and empiric broad-spectrum antibiotic treatment | 48
computed tomography and subsequent angiography | 48
no evidence of persistent fistula | 48
chronic obliteration of the iliac conduit | 48
partial perfusion of the hepatic artery by gastroduodenal collaterals | 48
anuric kidney failure | 48
continuous venovenous hemofiltration | 48
intermittent hemodialysis | 48
four months later, the patient was scheduled for FCSEMS replacement | 0
FCSEMS replacement | 0
no evidence of persisting leakage on cholangiogram | 0
no relevant stenosis | 0
fifty-month follow-up | 0
no evidence of recurrent stenosis or portobiliary fistula | 0