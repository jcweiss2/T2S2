54 years old | 0
male | 0
presented to the hospital | 0
fever | -168
cough | -168
progressive dyspnea | -168
syncope | -168
healthy state before onset of symptoms | -168
co-workers tested positive for SARS-CoV-2 | -168
nausea | 0
intermittent vomiting | 0
mild diarrhea | 0
denied previous medical history | 0
not taking any medications | 0
social history: 8 pack-years cigarette smoking 20 years ago | 0
temperature 38.3°C | 0
blood pressure 117/75 mmHg | 0
pulse 83 beats per minute | 0
respiratory rate 22 breaths per minute | 0
oxygen saturation 80% on room air | 0
bilateral rales | 0
negative influenza A and B tests | 0
high pretest probability of COVID-19 | 0
nasopharyngeal swab positive for SARS-CoV-2 | 0
mild lymphopenia | 0
elevated lactate dehydrogenase (315 U/L) | 0
elevated ferritin (3626 ng/mL) | 0
elevated D-dimer (1.34 mg/L) | 0
elevated inter-leukin-6 (13 pg/mL) | 0
elevated troponin-I (0.37 ng/mL) | 0
bilateral alveolar infiltrates on chest X-ray | 0
S1Q3T3 pattern on electrocardiogram | 0
acute respiratory distress syndrome (ARDS) | 0
septic shock | 0
intubated | 0
mechanical ventilation initiated | 0
norepinephrine initiated (0.01 μg/kg/min) | 0
bedside transthoracic echocardiogram performed | 0
large right-heart thrombus-in-transit through TV into RV | 0
preserved RV systolic function | 0
low-molecular-weight heparin (enoxaparin) started | 0
admitted to isolation unit | 0
hydroxychloroquine started | 0
azithromycin started | 0
cytokine release storm | 0
tocilizumab given | 0
limited transthoracic echocardiogram after 1 week | 168
preserved RV systolic function | 168
no evidence of thrombus | 168
LMWH continued | 0
minimal ventilator support required | 168
tracheostomy performed | 336
percutaneous endoscopic gastrostomy tube placed | 336
oxygen requirements decreased to 3–4 L | 336
continuous positive airway pressure support at night | 336
discharged to long-term acute care facility | 624
apixaban 5 mg twice a day started | 624
elevated D-dimer followed | 0
thrombocytopenia not observed | 0
elevated inflammatory markers | 0
cardiac injury | 0
hemostatic disturbances | 0
ARDS | 0
hypotension | 0
hypoxia | 0
vasovagal mechanism suspected | 0
preserved RV size | 0
minor myocardial damage | 0
peak troponin-I 0.37 ng/mL | 0
no clinical deterioration concerning PE | 0
intermediate low-risk PE category | 0
LMWH selected over unfractionated heparin | 0
elevated white cell count (5.41×103/µL) | 0
elevated neutrophils (4.56×103/µL) | 0
decreased lymphocytes (0.59×103/µL) | 0
elevated glucose (132 mg/dL) | 0
elevated blood urea nitrogen (22 mg/dL) | 0
elevated serum creatinine (1.08 mg/dL) | 0
decreased sodium (128 mmol/L) | 0
normal potassium (3.7 mmol/L) | 0
decreased chloride (88 mmol/L) | 0
normal carbon dioxide (26 mmol/L) | 0
normal pH arterial (7.41) | 0
normal pCO2 arterial (38.3 mmHg) | 0
normal pO2 arterial (104.3 mmHg) | 0
normal bicarbonate arterial (23.8 mmol/L) | 0
decreased total protein (6.6 g/dL) | 0
decreased albumin (3.4 g/dL) | 0
normal total bilirubin (0.5 mg/dL) | 0
elevated alanine aminotransferase (37 U/L) | 0
elevated aspartate aminotransferase (43 U/L) | 0
normal alkaline phosphatase (46 U/L) | 0
elevated total creatine kinase (147 U/L) | 0
elevated venous lactic acid (1.5 mmol/L) | 0
elevated procalcitonin (0.36 ng/mL) | 0
elevated interleukin-6 (13 pg/mL) | 0
