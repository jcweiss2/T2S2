18 years old | 0
male | 0
admitted to the hospital | 0
ulcerative colitis (UC) | 0
chronic inflammatory bowel disorder (IBD) | 0
megacolon | 0
failing systemic therapy | 0
infection | 0
hospitalization | 0
institutional review board approval | 0
ethics committee approval | 0
study protocol approval | 0
publication of data approval | 0
informed written consent | 0
transferred from another hospital | -24
intensive care unit (ICU) admission | 0
acute respiratory deterioration | 0
UC diagnosis | -672
infliximab administration | -216
infliximab administration | -528
intensive supportive therapy | 0
septic shock | 0
moderate acute respiratory distress syndrome | 0
acute kidney failure | 0
invasive ventilation | 0
renal replacement therapy | 0
hemodynamically unstable | 0
septic cardiomyopathy (SCM) | 0
reduced systolic left ventricular function | 0
reduced systolic right ventricular function | 0
left ventricular ejection fraction <15% | 0
positive inotropic therapy | 0
