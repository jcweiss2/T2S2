Here is the table of events and timestamps:

| Event | Timestamp |
| --- | --- |
| 59-year-old female | 0 |
| blood type: O, Rh positive | 0 |
| segment-V space-occupying lesion in the liver | -672 |
| suspected of being liver cancer | -672 |
| transarterial embolization | -672 |
| sorafenib | -336 |
| stopped due to dizziness, skin ulcers, and other symptoms | -224 |
| radiation therapy | -224 |
| prescribed dose: PTV5400cGy/18f, and a dose rate of 0.6–1 Gy/min | -224 |
| total of seven radiotherapy treatments | -224 |
| Piggyback LT | 0 |
| acute renal failure | 0 |
| hematoma around the liver | 0 |
| hepatitis B immunoglobulin | 1 |
| intravenous administration | 1 |
| immunosuppressive drugs, including steroids and tacrolimus | 1 |
| initial goal was to maintain the tacrolimus blood level at ~10 ng/mL | 1 |
| continuous hemodialysis and intermittent infusion of fresh frozen plasma, leukocyte-depleted red blood cells, and other blood products | 1 |
| active bleeding in the abdominal cavity ceased and renal function gradually recovered | 1 |
| pathological analyses confirmed the diagnosis of HCC | 10 |
| massive tumor necrosis was observed (necrosis accounted for ~90%, while the surviving tumor accounted for ~10%) | 10 |
| liver function began to improve | 10 |
| aspartate aminotransferase (AST), alanine aminotransferase (ALT), gamma-glutamyl transpeptidase (GGT), and alkaline phosphatase (ALP) levels all returned to normal | 10 |
| regular and repeated fevers of 37–39°C, peaking at 23:00 h daily | 10 |
| procalcitonin (PCT) levels began to rise to 10.3 ng/mL | 10 |
| blood cultures were negative, and cytomegalovirus, Epstein–Barr virus (EBV) were negative | 13 |
| fever did not subside, and obscure red spots were also observed on the patient’s chest | 13 |
| no symptoms such as itching, and the Nikolsky sign was negative | 13 |
| changed the tacrolimus administration to sirolimus and added mycophenolate mofetil to maintain immune suppression | 17 |
| sputum culture suggested the presence of Acinetobacter baumannii and methicillin-resistant Staphylococcus aureus (MRSA) infections | 18 |
| the patient’s rash advanced into erythematous macules and papules, and spread to the limbs, palms, neck, and face | 19 |
| oral examination revealed white ulcers on both sides of the buccal mucosa and lips | 19 |
| severe bone marrow suppression was observed, as well as a white blood cell (WBC) count of 0.86 × 10^9/L, a platelet (PLT) count of 35 × 10^9/L, and a hemoglobin (HGB) level of 70 g/L | 19 |
| transferred to the intensive care unit | 19 |
| a dermatologist hypothesized that the rash may be a drug-related adverse reaction and recommended gamma globulin administration (2500 mg, 3 days) | 19 |
| skin biopsy on the patient’s left chest and performed fluorescence in situ hybridization (FISH) of the peripheral blood | 19 |
| abdominal incision split and was sutured again | 29 |
| bone marrow aspiration to determine the cause of the bone marrow suppression | 32 |
| bone marrow pathology report revealed no special lesions in the morphology of granulocytes, red blood cells, or megakaryocytes | 32 |
| FISH analysis of the peripheral blood followed by flow cytometry detected 3% donor lymphocytes | 33 |
| skin biopsy specimens exhibited epidermal dyskeratosis, basic vacuolization, and lymphocytic infiltrates, which were consistent with grade-1 acute lt-GVHD | 33 |
| differential diagnoses include bacterial, fungal, and viral infections, drug reactions, toxic epidermal necrolysis, and hemophagocytic syndrome | 33 |
| collective findings, together with the clinical course, were consistent with the diagnosis of lt-GVHD | 33 |
| analysis of serum T-lymphocyte subsets revealed that the ratio of CD4:CD8 was reversed (1:13.3 instead of 2:1) | 33 |
| serum immunoglobin M was reduced to 0.3 g/L | 33 |
| despite continuous platelet transfusion and the use of thrombopoietin (TPO), the patient’s PLT count dropped to 3.2 × 10^9/L | 33 |
| the patient’s serum immunoglobin M level was reduced to 0 g/L | 55 |
| succumbed to septic shock and multiple organ dysfunction syndrome (MODS) | 55 |