64 years old | 0
male | 0
hepatitis C virus infection | 0
alcohol-related cirrhosis | 0
hepatocellular carcinoma | 0
liver transplant | 0
ABO-identical liver transplant | 0
cytomegalovirus-seronegative donor | 0
toxoplasma-seropositive donor | 0
cytomegalovirus-seropositive recipient | 0
toxoplasma-seropositive recipient | 0
body mass index 24.5 kg/m2 | 0
Child–Pugh score A6 | 0
model end-stage liver disease score 10 | 0
transfusion of 2 units of concentrated red cells | 0
transfusion of 4 units of fresh frozen plasma | 0
tacrolimus | 0
Corticosteroid | 0
methylprednisolone | 0
increase in hepatic enzymes | -216
aspartate aminotransferase increase | -216
alanine aminotransferase increase | -216
hepatic biopsy | -216
acute cellular rejection | -216
steroid pulse therapy | -216
methylprednisolone | -216
recovery | -160
discharge | -160
readmission | 216
fever | 216
skin rash | 216
diarrhea | 216
leukopenia | 216
anemia | 216
low hemoglobin | 216
low blood pressure | 216
skin biopsy | 216
spongiosis | 216
basal cell hydropic changes | 216
apoptotic keratinocytes | 216
lymphocytic exocytosis | 216
satellite-cell necrosis | 216
subepidermal cleft formation | 216
grade III of acute GVHD | 216
myelogram | 240
hypoplastic bone marrow | 240
aplasia | 240
single-cell necrosis | 240
gastrointestinal symptoms | 240
gland abscesses | 240
mucosal denudation | 240
macrochimerism | 240
donor T-lymphocyte macrochimerism | 240
methylprednisolone | 216
antithymocyte globulin | 216
pulmonary insufficiency | 288
renal insufficiency | 288
agranulocytosis | 288
multi-organ failure | 288
death | 288