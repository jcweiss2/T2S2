33 years old | 0 | 0 
female | 0 | 0 
admitted to the hospital | 0 | 0 
nausea | -24 | 0 
vomiting | -24 | 0 
abdominal pain | -24 | 0 
discharged | -36 | -36 
hospitalized for recurrent pericarditis | -36 | -36 
treated with colchicine | -36 | -12 
febrile | 0 | 0 
hypotensive | 0 | 0 
leukocytosis | 0 | 0 
elevated serum lactate | 0 | 0 
acute kidney injury | 0 | 0 
acute transaminitis | 0 | 0 
severe coagulopathy | 0 | 0 
normal serum troponin | 0 | 0 
negative comprehensive toxicology screen | 0 | 0 
normal sinus rhythm | 0 | 0 
normal biventricular function | 0 | 0 
no valvular disease | 0 | 0 
no pericardial effusion | 0 | 0 
sepsis suspected | 0 | 0 
fluid resuscitated | 0 | 24 
broad-spectrum antibiotics | 0 | 24 
vasopressor therapy | 0 | 24 
severe multisystem organ failure | 24 | 24 
intubated | 24 | 24 
paralyzed | 24 | 24 
intravascular volume repletion | 24 | 48 
intravenous vasopressors | 24 | 48 
stress-dose steroids | 24 | 48 
high-dose vitamin B12 | 24 | 48 
Swan-Ganz catheter placed | 24 | 24 
distributive shock | 24 | 24 
cardiac output 7.4 l/min | 24 | 24 
pulmonary artery diastolic pressure 8 mm Hg | 24 | 24 
systemic vascular resistance indexed 1572 dynes/s/cm5/m2 | 24 | 24 
cardiogenic shock | 48 | 48 
high filling pressures | 48 | 48 
low CO | 48 | 48 
high systemic vascular resistance | 48 | 48 
elevated troponin | 48 | 48 
severe biventricular failure | 48 | 48 
left ventricular ejection fraction 15% | 48 | 48 
intravenous milrinone | 48 | 72 
continuous renal replacement therapy | 48 | 120 
PRBC transfusion | 48 | 48 
CO normalized | 72 | 72 
troponin decreased | 72 | 72 
multisystem organ failure improved | 72 | 72 
neutropenic | 96 | 96 
recovery of LVEF to 50-55% | 144 | 144 
weaned from vasopressors | 240 | 240 
taken off CRRT | 240 | 240 
extubated | 312 | 312 
hair loss | 576 | 576 
admitted to taking 60 tablets of 0.6 mg of colchicine | 0 | 0 
elevated serum colchicine level | 30 | 30 
elevated whole blood colchicine level | 14 | 14 
hypertension | -36 | 0 
pulmonary emboli | -36 | 0 
polysubstance abuse | -36 | 0 
discharged from hospital | 432 | 432 
outpatient rehabilitation | 432 | 432 
complete renal recovery | 432 | 432 
complete hepatic recovery | 432 | 432 
complete cardiac recovery | 432 | 432