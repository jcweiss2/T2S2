67 years old | 0
male | 0
coronary heart disease | 0
atrial fibrillation | 0
heart failure | 0
admitted to the hospital | 0
dyspnea | 0
rapid AF | 0
treated with diuretics | 0
treated with milrinone | 0
treated with nitrate | 0
RFCA of AF | -72
discharged from the hospital | 72
chest discomfort | -432
fever | -432
confusion | -432
gazing upwards | -432
mild limb seizures | -432
vomiting | -432
temperature 41°C | -432
WBC 5.2 × 10^9/L | -432
hsCRP 18.56 mg/L | -432
supraventricular tachycardia | -432
hypothermia therapy | -432
admitted to emergency department | -432
temperature 37.9°C | 0
blood pressure 99/73 mm Hg | 0
pulse rate 78 beats/min | 0
ECG showed AF | 0
NT-proBNP 1550.00 pg/mL | 0
alanine aminotransferase 21 U/L | 0
cardiac troponin I 3.95 μg/L | 0
WBC 10.58 × 10^9/L | 0
neutrophil 97.2% | 0
hsCRP 26.0 mg/L | 0
fecal occult blood 3+ | 0
cerebral CT did not reveal any abnormal findings | 0
pulmonary CT did not reveal any abnormal findings | 0
CECT showed suspicious thrombus in left atrial appendage | 0
fasting | 0
GI decompression | 0
antibiotic treatment | 0
imipenem/cilastatin | 0
linezolid | 0
regained consciousness | 24
repeated epileptic seizures | 24
cerebral MRI showed lacuna infarctions | 48
emergency EGD | 48
small and deep ulcer at 30 cm from incisors | 48
esophageal stenting | 48
self-expanding, polyester-covered, length 100 mm, width 18 mm | 48
WBC counts decreased | 72
hsCRP level decreased | 72
epileptic seizures went away | 72
acid reflux | 120
temperature increased | 168
WBC counts increased | 168
cardiac CECT showed esophageal-mediastinum fistula | 168
encapsulated effusion | 168
pneumatosis behind left atrium | 168
post wall of LA depression | 168
mediastinal abscess | 168
AEF | 168
surgical repair planned | 168
right thoracotomy incision | 192
membranaceous and funicular adhesions | 192
tight adhesion between esophagus and pericardium | 192
6 mm diameter fistula in the anterior wall of esophagus | 192
tight adhesion between LA and pericardium | 192
bleeding at the posterior wall of LA | 192
Rid-muscle flap pedicled with vessels | 192
repair LA posterior wall and fistula between esophagus and LA | 192
pleuroclysis using povidone iodine and nature saline | 192
transferred to intensive care unit | 216
out-of-control sepsis | 216
infectious shock | 216
repeated fever | 216
chills | 216
metabolic acidosis | 216
hypotension | 216
tachycardia | 216
oliguria | 216
death | 240