57 years old | 0
    woman | 0
    fever | -72
    diarrhea | -72
    tetracycline | -72
    fatigue | -72
    admitted to a local general hospital | -72
    elevated transaminase levels | -72
    bicytopenia | -72
    reduced prothrombin time activity | -72
    HAV-IgM negative | -72
    HBs antigen negative | -72
    HCV antibody negative | -72
    VCM-IgM negative | -72
    CMV antigenemia negative | -72
    AMA negative | -72
    ASMA negative | -72
    HTLV-1 antibody negative | -72
    HIV antibody negative | -72
    encephalopathy | -72
    confusion | -72
    slow movement | -72
    bone marrow biopsy | -72
    increased numbers of mature histiocytes | -72
    hemophagocytosis | -72
    FH | -72
    HPS | -72
    steroid pulse therapy | -72
    CHDF | -72
    transferred to our hospital | 0
    liver transplantation | 0
    severe respiratory failure | 72
    tracheal intubation | 72
    mechanical ventilation | 72
    CT chest bronchial wall thickening | 72
    bilateral diffuse infiltration shadow of lungs | 72
    bronchoscopic pseudomembranous formation | 72
    β-D-glucan level increased | 72
    Aspergillus galactomannan antigen level >5.0 | 72
    CRP 2.52 mg/dl | 72
    PCT 0.4 ng/mL | 72
    pH 7.32 | 72
    PaO2 89.4 mmHg | 72
    PaCO2 53.9 mmHg | 72
    HCO3− 19.3 mmol/L | 72
    PaO2/FiO2 149 | 72
    endobronchial biopsy | 72
    active inflammation | 72
    necrotic tissue | 72
    filamentous fungal hyphae infiltration | 72
    Aspergillus fumigatus isolated | 72
    Burkholderia cepacia isolated | 72
    pseudomembranous ITBA | 72
    ARDS | 72
    bacterial pneumonia | 72
    IPA | 72
    pulmonary edema | 72
    unable to perform BAL | 72
    broad-spectrum antibiotics | 72
    imipenem | 72
    voriconazole | 72
    caspofungin | 72
    β-D-glucan level decreased | 72
    tracheobronchial pseudomembrane scarring | 72
    septic shock | 72
    Burkholderia cepacia | 72
    ARDS | 72
    died | 1368
    
