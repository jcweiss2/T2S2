31 years old | 0
female | 0
non-smoking | 0
Caucasian | 0
no past medical history | 0
admitted to the hospital | 0
sudden-onset severe headache | -840
left arm numbness | -840
cranial computed tomography (CT) scan | -840
grade 2 SAH | -840
ruptured right middle cerebral artery aneurysm | -840
percutaneous endovascular coil embolization | -840
fever | -672
chills | -672
constant abdominal pain | -672
purulent uterine discharge | -672
empiric antibacterial therapy | -672
sepsis | -672
septic shock | -672
transferred to the intensive care unit | -672
body temperature 38.3 °C | -672
invasive blood pressure 90/65 mmHg | -672
heart rate 135/min | -672
arterial oxygen saturation 82 % | -672
mild disorientation | -672
slower capillary refill | -672
coarse rales | -672
sequential organ failure assessment (SOFA) score 4 | -672
hemoglobin 6.8 g/dL | -672
d-dimers 4.58 μg/mL | -672
C-reactive protein 322 mg/L | -672
fibrinogen concentration 6.4 mL | -672
blood culture showed E. coli | -672
chest radiography | -672
pulmonary nodules | -672
transvaginal ultrasound | -672
enlarged uterus | -672
complete loss of zonal anatomy | -672
abdominal magnetic resonance imaging (MRI) | -672
enlarged heterogenous myometrial mass | -672
splenic metastatic lesion | -672
serum β-human chorionic gonadotrophin (β-hCG) 232,085 mUI/mL | -672
suction evacuation and curettage | -672
pathology report confirmed choriocarcinoma diagnosis | -672
International Federation of Gynecology and Obstetrics (FIGO) modified WHO prognostic scoring system | -672
total score of 12 | -672
high risk of developing resistance to single-drug chemotherapy | -672
initiation of multiagent chemotherapy regimen | -672
low-dose etoposide | -672
cisplatin | -672
EMA/CO regimen | -24
etoposide | -24
methotrexate | -24
actinomycin D | -24
cyclophosphamide | -24
vincristine | -24
six cycles of EMA/CO | 0
β-hCG levels plateaued above normal | 0
restaging with MRI of the brain | 24
18F-fluorodeoxyglucose (FDG) positron emission tomography (PET)/CT scan | 24
decreased pulmonary nodules | 24
decreased uterine mass | 24
low standardized uptake value (SUV) of <3.8 | 24
revised FIGO score 7 | 24
therapeutic regimen changed to EP/EMA | 24
etoposide plus cisplatin | 24
etoposide, methotrexate, and actinomycin D | 24
normalization of β-hCG | 168
completion of three cycles | 168
grade 3 neutropenia | 48
incorporation of granulocyte colony stimulating factor (G-SCF) | 48
dose reduction of both etoposide and actinomycin D | 48
grade 2 alopecia | 48
grade 2 nausea | 48
dexamethasone | 48
ondansetron | 48
grade 2 fatigue | 168
use of male condoms | 0
follow-up | 1680
disease-free for almost two years | 1680