66 years old | 0
male | 0
Caucasian | 0
admitted to the hospital | 0
pain during defecation | -144
hematochezia | -48
coronary artery bypass surgery | -6720
percutaneous coronary intervention | -6720
chronic obstructive pulmonary disease | -6720
diabetes | -6720
myelo-dysplastic syndrome | -6720
75-pack years of smoking | -6720
Plavix | -6720
ASA | -6720
antihypertensive drugs | -6720
colonoscopy | 0
unstable bleeding | 0
hypotensive | 0
normal heart rate | 0
fever | 0
tenderness in the lower left quadrant | 0
anaemic | 0
infected | 0
intravenous fluid | 0
blood cultures | 0
intravenous antibiotics | 0
acute contrast-enhanced computer tomography | 0
retroperitoneal bleeding | 0
left external iliac artery | 0
emergency damage control endo-grafting | 0
Fluency covered stentgraft | 0
temperature fluctuating | 72
intermittent left-sided abdominal pain | 72
septic | 72
CT-scan | 72
hematoma | 72
air near the covered stent | 72
sigmoidal colon | 72
Clostridium tertium bacterium | 72
white blood count decreasing | 72
C-reactive-protein concentration decreasing | 72
control CT-scan | 216
infected hematoma regression | 216
thickening of the sigmoid colon | 216
exploratory laparotomy | 216
fistula | 216
Hartmann’s procedure | 216
infected stent removal | 216
femoro-femoral bypass operation | 216
intensive care unit | 216
hypotension | 216
pain | 216
slow recovery | 216
histological examination | 216
diverticulitis | 216
abscess | 216
inflammation | 216
perforation | 216
infection in the left groin | 504
CT-scan | 504
intravenous antibiotics | 504
re-incision | 504
drainage | 504
rinsing of the abscess cavity | 504
discharged | 720
oral antibiotics | 720
control appointment | 1008
no signs of vascular prosthesis infection | 1008
antibiotics discontinued | 1008
stress | 1008
colostomy | 1008
gratefulness | 1008