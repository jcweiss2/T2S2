68 years old | 0
male | 0
admitted to the Emergency Department | 0
fever | -72
wheezing | -72
arterial hypertension | 0
dyslipidemia | 0
Atorvastatin 80 mg once daily | 0
Candesartan 32 mg OD | 0
SARS-CoV-2 positive | 0
bilateral interstitial pneumonia | 0
HRCT severity score 15/20 | 0
BP 117/74 mmHg | 0
HR 83 bpm | 0
SpO2 79% | 0
sinus rhythm at 85 bpm | 0
narrow QRS complex | 0
normal atrioventricular conduction | 0
normal intraventricular conduction | 0
no ST-T segment abnormalities | 0
Azithromycin 500 mg OD | 0
Methylprednisolone 20 mg BID | 0
Remdesivir 200 mg OD | 0
Enoxaparin 6000 UI BID | 0
Insulin Lispro 6/8/8 UI TID | 0
High Flow Nasal Cannula FiO2 45% | 0
antihypertensive therapy discontinued | 0
statin therapy discontinued | 0
clinical status improved | 672
HRCT severity score 5/20 | 600
sudden worsening of dyspnea | 672
increased heart rate | 672
ST-T segment morphological alterations | 672
BP 154/75 mmHg | 672
HR 85 bpm | 672
SpO2 97% | 672
sinus rhythm at 78 bpm | 672
ST-elevation ≥ 2 mm in DI, aVL, V1-V4 | 672
STEMI diagnosis | 672
Acetylsalicylic acid 300 mg | 672
Ticagrelor 180 mg | 672
Bisoprolol 2.5 mg | 672
Atorvastatin 80 mg | 672
hypokinesis in mid-apical anterior segment | 672
no intra-cardiac thrombi | 672
PCI performed | 672
critical stenosis of LAD | 672
PTCA with DES | 672
transfer delay 3 hours 23 minutes | 672
left hemiplegia | 696
NIHSS score 7 | 696
acute right frontal ischemic lesion | 696
no fibrinolysis | 696
discharge | 1176
no residual neurologic deficit | 1344
