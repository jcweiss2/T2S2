65 years old | 0
female | 0
ovarian cancer | 0
relapsed ovarian cancer | 0
carboplatin treatment | 0
dyspnea | -0.33
wheezing | -0.33
hypotension | -0.33
confusion | -0.33
infusion stopped | -0.33
transferred to ICU | -0.33
intubated | -0.33
adrenaline infused | -0.33
fluids infused | -0.33
corticosteroids infused | -0.33
cardiac ultrasound performed | -0.33
acute coronary syndrome excluded | -0.33
ECG performed | -0.33
troponin I measured | -0.33
pulmonary embolism ruled out | -0.33
spiral CT scan of lungs performed | -0.33
Swan-Ganz catheter inserted | -0.33
pulmonary capillary wedge pressure measured | -0.33
central venous pressure measured | -0.33
ventilated | -0.33
blood cultures drawn | -0.33
urine cultures drawn | -0.33
abdomen ultrasound performed | -0.33
brain CT scan performed | -0.33
fever | 144
ventilator-associated pneumonia diagnosed | 144
bronchoalveolar lavage drawn | 144
antibiotics administered | 144
septic | 144
died | 144