59 years old | 0
male | 0
Pakistani | 0
admitted to the hospital | 0
short of breath | -8760
decreased exercise tolerance | -8760
intermittent fevers | -8760
leukocytosis | -8760
evaluated by cardiologist | -8760
echocardiogram | -8760
stress test | -8760
mediastinal and right pleural base mass | -8760
chest X-ray | -8760
large mass in the right pleural space | -8760
computed tomography scan | -8760
large inhomogeneous mass | -8760
compression of the right atrium | -8760
compression of the lung | -8760
compression atelectasis | -8760
biopsy of the mass | -8760
diagnosis of thymoma | -8760
traveled to the United States | -720
CT scan of the chest | -720
persistent right pleural based mass | -720
compression of the right atrium | -720
compression of the right lung | -720
pathology slides reviewed | -720
diagnosis confirmed to be thymoma | -720
discussion with patient and family | -24
elected to undergo surgical resection | -24
febrile | -24
leukocytosis | -24
admitted to thoracic surgery service | -24
chest X-ray | -24
large right pleural mass | -24
transthoracic echocardiogram | -24
normal ventricular function | -24
no vegetations | -24
compression of the right atrium | -24
Duplex ultrasound | -24
no deep venous thromboses | -24
blood and urine cultures | -24
negative cultures | -24
hematology/oncology service consulted | -24
bone marrow biopsy | -24
peripheral smear | -24
negative results | -24
Infectious Disease service consulted | -24
started on intravenous antibiotics | -24
surgical resection of mass | 48
endotracheally intubated | 48
transesophageal echocardiography | 48
extended right posterolateral thoracotomy incision | 48
exploration of right pleural cavity | 48
enormous mass | 48
purulent fluid and necrotic tumor mass | 48
frozen section | 48
suspicious for lymphoma | 48
deferred resection of mass | 48
chest tubes placed | 48
wound closed | 48
transferred to cardiothoracic intensive care unit | 48
septic | 72
vasopressor support | 72
aggressive fluid resuscitation | 72
weaned off vasopressors | 96
weaned off ventilator | 96
extubated | 96
transferred to medical/surgical unit | 96
chest tubes remained in place | 96
daily chest X-rays | 96
noticeable improvement in right lung | 96
final pathology | 120
thymoma | 120
Salmonella species | 120
non-typhoidal | 120
intravenous antibiotic coverage changed | 120
transitioned to oral antibiotics | 240
discharged home | 240
follow-up plan | 240
repeat CT scan | 672
mass without significant change | 672
effort-induced shortness of breath | 672
decision to undergo surgical resection | 672
readmitted to hospital | 720
right thoracotomy | 744
complete resection of tumor mass | 744
partial right lower lobectomy | 744
echocardiogram | 744
large mass compressing right atrium | 744
specimen resected | 744
marked improvement in compression of right atrium | 744
tolerated procedure well | 744
transferred to surgical floor | 768
shortness of breath resolved | 768
significant improvement on chest X-ray | 768
chest tube discontinued | 768
sent home | 840
completed antibiotic therapy | 1008