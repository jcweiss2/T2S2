39 years old | 0
male | 0
admitted to the hospital | 0
malaise | -168
encephalopathy | -168
septic shock | 0
blood cultures grew MSSA | 0
fluid cultures from left elbow olecranon bursa grew MSSA | 0
fluid cultures from right foot abscess grew MSSA | 0
concern for endocarditis with systemic emboli | 0
retained foreign objects on chest radiograph | 0
retained foreign objects on abdominal radiograph | 0
transesophageal echocardiography (TEE) was negative for vegetation | 0
MSSA pulmonary septic emboli | 0
retained foreign body in the right upper pulmonary artery sub-segmental branch | 0
retained guide wire extending from the inferior vena cava (IVC) to the left iliac and left common femoral vein | 0
motor vehicle accident | -3840
femoral central venous access placement | -3840
guide wire presence | -3840
plan for re-imaging and retrieval | -3840
lost to follow up | -3840
interventional radiology removed the IVC portion of the wire | 24
unable to retrieve the right pulmonary artery portion of the wire | 24
started on antibiotic regimen | 24
clearance of bacteremia | 168
resolution of symptoms | 168
no chronic lifelong suppression therapy | 168
discharged | 168