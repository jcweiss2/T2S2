23 years old | 0
woman | 0
referred to medical high-dependency unit | 0
hypogastric pain | -168
vomiting | -168
suicide attempt 7 years ago | -1344
expressive aphasia | 0
vertigo | 0
unsteady gait | 0
severe metabolic acidosis | 0
hyperlactataemia | 0
brain computed tomography | 0
lumbar puncture | 0
treated with 680 mmol i.v. bicarbonate | 0
infusions | 0
antipyretics | 0
pyrexia | 0
toxicology screening showed ethylene glycol traces | 0
glycolic acid in urine | 0
immediate therapy with i.v. ethanol | 0
lost consciousness | 16
developed convulsions | 16
intubated | 16
admitted to intensive care unit | 16
aspiration pneumonia | 16
sepsis | 16
renal failure | 16
ethylene glycol poisoning confirmed | 16
treatment included antibiotics for pneumonia | 16
continuous haemodiafiltration | 16
CRRT with bicarbonate-buffered solutions | 16
citrate-calcium module | 16
estimated citrate level 4.0–4.7 mmol/L | 16
improvement of consciousness | 168
extubation attempt on day 7 | 168
failed extubation on day 8 due to sputum retention | 192
reintubation | 192
dilatation tracheostomy on day 12 | 288
required two revisions due to bleeding | 288
referred to tertiary hospital on day 16 | 384
intractable metabolic alkalosis | 384
two organ failures | 384
bleeding from tracheostomy | 384
initial bronchoscopy | 384
eliminated atelectasis | 384
secured open bronchial tree | 384
microbiology specimens | 384
ceasing antibiotics after 5 days (day 21) | 504
echocardiography showed reduced ejection fraction | 504
thrombus in right internal jugular vein | 504
chest X-ray showed infiltration of right lower lobe | 504
metabolic alkalosis on admission to tertiary centre | 384
hypernatraemia | 384
urea 37 mmol/L | 384
serum creatinine 422 μmol/L | 384
total to ionised calcium ratio 2.42 | 384
total plasma protein 107.7 g/L | 384
electrophoresis performed | 384
immunoassay on free light chains on day 21 | 504
free kappa 170 mg/L | 504
free lambda 106 mg/L | 504
kappa/lambda ratio 1.61 | 504
treated with CRRT | 384
RCA | 384
trisodium citrate | 384
calcium chloride replacement | 384
calcium-free lactate-buffered solution | 384
dialysate flow 1.5 L/h | 384
plasmatic natrium lowered by 10 mmol/L | 408
dialysate flow increment to 2.2 L/h | 408
normal acid-base parameters reached on day 20 | 480
restored consciousness | 480
weaning of respiratory support | 480
decannulated on day 22 | 528
CRRT ceased on day 23 | 552
diuresis restored | 552
transferred back to regional hospital | 552
improving slowly | 552
discharged home on day 48 | 1152
no need for renal replacement therapy | 1152
healed tracheostomy | 1152
normal renal functions | 1152
taking care of child | 1152
hyperlactataemia |7.0
brain computed tomography |0
lumbar puncture |0
treated with 680 mmol i.v. bicarbonate |0
infusions |0
antipyretics |0
pyrexia |0
toxicology screening showed ethylene glycol traces |0
glycolic acid in urine |0
immediate therapy with i.v. ethanol |0
lost consciousness |16
developed convulsions |16
intubated |16
admitted to intensive care unit |16
aspiration pneumonia |16
sepsis |16
renal failure |16
ethylene glycol poisoning confirmed |16
treatment included antibiotics for pneumonia |16
continuous haemodiafiltration |16
CRRT with bicarbonate-buffered solutions |16
citrate-calcium module |16
estimated citrate level 4.0–4.7 mmol/L |16
improvement of consciousness |168
extubation attempt on day 7 |168
failed extubation on day 8 due to sputum retention |192
reintubation |192
dilatation tracheostomy on day 12 |288
required two revisions due to bleeding |288
referred to tertiary hospital on day 16 |384
intractable metabolic alkalosis |384
two organ failures |384
bleeding from tracheostomy |384
initial bronchoscopy |384
eliminated atelectasis |384
secured open bronchial tree |384
microbiology specimens |384
ceasing antibiotics after 5 days (day 21) |504
echocardiography showed reduced ejection fraction |504
thrombus in right internal jugular vein |504
chest X-ray showed infiltration of right lower lobe |504
metabolic alkalosis on admission to tertiary centre |384
hypernatraemia |384
urea 37 mmol/L |384
serum creatinine 422 μmol/L |384
total to ionised calcium ratio 2.42 |384
total plasma protein 107.7 g/L |384
electrophoresis performed |384
immunoassay on free light chains on day 21 |504
free kappa 170 mg/L |504
free lambda 106 mg/L |504
kappa/lambda ratio 1.61 |504
treated with CRRT |384
RCA |384
trisodium citrate |384
calcium chloride replacement |384
calcium-free lactate-buffered solution |384
dialysate flow 1.5 L/h |384
plasmatic natrium lowered by 10 mmol/L |408
dialysate flow increment to 2.2 L/h |408
normal acid-base parameters reached on day 20 |480
restored consciousness |480
weaning of respiratory support |480
decannulated on day 22 |528
CRRT ceased on day 23 |552
diuresis restored |552
transferred back to regional hospital |552
improving slowly |552
discharged home on day 48 |1152
no need for renal replacement therapy |1152
healed tracheostomy |1152
normal renal functions |1152
taking care of child |1152
