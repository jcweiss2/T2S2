48 years old | 0
male | 0
Spanish-speaking | 0
admitted to the hospital | 0
shortness of breath | -168
cough | -168
central chest pain | -168
feeling of warmth | -168
hypertension | -6720
hyperlipidemia | -6720
chronic back pain | -6720
lisinopril | -6720
atorvastatin | -6720
over-the-counter analgesics | -6720
temperature 36.4 Celsius | 0
heart rate 87/minute | 0
blood pressure 126/73 mm of Hg | 0
respiratory rate 22/minute | 0
oxygen saturation 95% | 0
white blood cell count 9,000/cumm | 0
neutrophil count 76.6% | 0
lymphocyte count 15.4% | 0
absolute lymphocyte count 1.40 K/mm | 0
lactic acid level 1.3 mmol/L | 0
erythrocyte sedimentation rate (ESR) 62 mm/hr | 0
c-reactive protein (CRP) 8.66 mg/dl | 0
troponin <0.03 ng/ml | 0
procalcitonin 0.19 ng/ml | 0
normal sinus rhythm | 0
no ST or T wave changes | 0
hypo inflation | 0
perihilar air space opacities | 0
atelectasis | 0
bilateral ground glass opacities | 0
ceftriaxone | 0
azithromycin | 0
tachycardic | 12
hypoxic | 12
fevers | 12
SARS CoV-2 positive | 12
hydroxychloroquine | 12
non-invasive ventilation | 72
endotracheal intubation | 120
transfer to the intensive care unit | 120
prone position | 120
ST elevations | 192
troponin level peaked at 0.10 ng/ml | 192
clopidogrel | 192
allergy to aspirin | 192
evaluated by Cardiology | 192
acute coronary syndrome | 192
serial ECGs | 216
ST changes resolved | 216
coronary catheterization deferred | 216
focal pericarditis | 216
elevated ESR 122 mm/hr | 240
elevated CRP 17.86 mg/dl | 240
cytokine storm | 240
methylprednisolone | 240
dexamethasone | 240
deep vein thrombosis | 240
prophylactic dose of anticoagulation | 240
therapeutic anticoagulation | 240
intravenous plasma | 240
critical respiratory status | 240
normal left ventricular function | 336
no regional wall motion abnormalities | 336
discharged | -1