34 years old | 0
male | 0
admitted to the hospital | 0
fatigue | -168
back pain | -168
abdominal pain | -168
nausea | -168
vomiting | -168
dyspnea | -24
hemoptysis | -24
temperature 35.9 °C | -24
systolic blood pressure 70 mmHg | -24
heart rate 100 beats per minute | -24
respiratory rate 19 breaths per minute | -24
oxygen saturation 60% | -24
jaundice | -24
abdominal pain over the right upper quadrant | -24
ubiquitous coarse crackles | -24
bilateral patchy infiltrates | -24
mild normochromic, normocytic anemia | -24
bilirubin 8.45 mg/dL | -24
severe thrombocytopenia | -24
acute renal failure | -24
leukocytosis | -24
elevated C-reactive protein | -24
elevated procalcitonin | -24
community acquired pneumonia with sepsis | -24
piperacillin/tazobactam | -24
ciprofloxacin | -24
endotracheal intubation | -16
extracorporeal membrane oxygenation (ECMO) therapy | -16
combined metabolic and respiratory acidosis | 0
hypoxemia | 0
extended confluent infiltrates | 0
severe adult respiratory distress syndrome (ARDS) | 0
diffuse alveolar hemorrhage | 0
intravascular hemolysis | 0
drop of hemoglobin | 0
reduced haptoglobin | 0
increased lactate dehydrogenase | 0
coagulation compromised | 0
fibrinogen levels below detection limit | 0
packed red blood cells transfused | 0
fibrinogen transfused | 0
muddy-brown casts | 0
acanthocytes | 0
hyperkalemia | 0
continuous venovenous renal replacement therapy | 0
plasmapheresis | 0
volume therapy | 0
sodium bicarbonate | 0
extracorporeal cytokine absorbent filter | 0
prednisolone | 0
fulminant multi-organ failure | 17
death | 17
fibrin monomers negative | 17
anti-glomerular basement antibodies negative | 17
anti-nuclear antibodies negative | 17
anti-neutrophil cytoplasmic antibodies negative | 17
schistocytes detected | 17
ADAMTS-13 activity reduced | 17
LipL32-PCR detecting Leptospira interrogans DNA positive | 24
Leptospira interrogans serovar icterohaemorrhagiae strain 17 detected | 24
pet rat identified as transmitting vector | -672