26 years old | 0
female | 0
thin built | 0
57 kg | 0
body mass index 20.2 | 0
admitted to the emergency department | 0
lump in the right upper quadrant of her abdomen | 0
malaena | 0
pale | 0
anicteric | 0
pulse rate of 120/min | 0
blood pressure of 90/60 mm of Hg | 0
respiratory rate of 25/min | 0
tender lump in the right upper quadrant | 0
probable suspicion of an infected bilioma | 0
no symptoms suggestive of hepatic failure | 0
aggressive resuscitation | 0
progressive pallor | 8
hypotension | 8
further episodes of malena | 8
high index of suspicion for an iatrogenic vasculobiliary pathology | 8
emergency ultrasound | 8
free fluid in lower abdomen | 8
encysted collection around liver | 8
bidirectional flow pattern on Doppler signal | 8
emergency computed tomography (CT) abdomen | 8
vascular reconstruction | 8
haemoglobin of 5.6 g/dl | 8
slightly elevated hepatic enzymes | 8
normal coagulation profile | 8
resuscitated with IV fluids | 8
packed red blood cells transfused | 8
contrast-enhanced computer-aided tomography | 8
perihepatic collection | 8
contrast spillage in the gallbladder fossa | 8
HAPA | 8
involving the right hepatic artery | 8
reconstructed image | 8
deteriorated | 16
urgent unavailability of angio-embolisation | 16
urgent exploratory laparotomy | 16
abdomen accessed with a right subcostal incision | 16
subphrenic and supracolic compartments containing altered clotted blood evacuated | 16
right hepatic artery isolated | 16
controlled proximally | 16
ruptured pseudoaneurysmal sac opened | 16
minimal back bleeding | 16
excised | 16
pseudoanerysm sac identified | 16
metal clip eroding in the right hepatic artery | 16
rent in the wall of the right hepatic artery repaired | 16
refashioning of the edges | 16
no other associated visceral injuries | 16
arterial anatomy showed the most common prevalent pattern | 16
single right hepatic artery arising from trunk of common hepatic | 16
5 cm after gastroduodenal artery branch | 16
pathology of the site did not allow to comment of 'Moynihan hump/Caterpillar hump' | 16
no active bile leak from cystic duct stump | 16
ligated again | 16
liver bed | 16
peritoneal lavage given | 16
wide bore drain kept in the Morrison's pouch | 16
haemostasis achieved | 16
wound closed in two layers | 16
received 3 units of packed red blood cells postoperatively | 24
post-operative course uneventful | 24
superficial surgical site infection | 24
wound dressings | 24
discharged on day 12 | 288
follow-up as outpatient at 6 months | 4320
no signs of delayed biliary stricture or liver dysfunction | 4320
ultrasound and Doppler assessment at hepatic hilum | 4320
bidirectional flow | 4320
plan to follow-up the patient for at least 2 years | 4320
laparoscopic cholecystectomy | -672
metal clip | -672
cystic artery stump | -672
pseudoaneurysm | 8
HAPA | 8
right hepatic artery | 8
erosion of metal clip | 8
haemobilia | 0
gastrointestinal haemorrhage | 0
melena | 0
jaundice | 0
abdominal pain | 0
anemia | 0
upper gastrointestinal endoscopy | 8
CT scan | 8
angiographic reconstruction | 8
hyperdense areas | 8
transarterial embolisation | 16
coiling | 16
exploratory laparotomy | 16
excise the aneurysm | 16
repair the artery | 16