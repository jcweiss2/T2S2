55 years old | 0
    male | 0
    admitted to the intensive care unit | 0
    motorcycle accident | 0
    sternal lesions | 0
    humeral lesions | 0
    D4 vertebral fracture | 0
    D9 vertebral fracture | 0
    hypertensive pneumothorax | 0
    Glasgow Coma Score 14/15 | 0
    intracapsular spleen haematoma | 0
    multiple fractures of the pelvis | 0
    empirical therapy with ceftazidime | 120
    empirical therapy with gentamicin | 120
    abrupt onset of fever | 168
    temperature >38.5°C | 168
    clinical features of septic shock | 168
    severe leucocytosis | 168
    low platelet count | 168
    vasoactive amines | 168
    mechanical ventilation | 168
    no hemodialytic treatment | 168
    monolateral purulent pleural suffusion | 168
    thoracic drainage | 168
    copious purulent leakage | 168
    two sets of blood samples taken for culture | 168
    growth of pleomorphic Gram-positive microorganisms | 250
    identification by MALDI-TOF failed | 250
    identification achieved by 16S rRNA PCR amplification and sequencing | 250
    metabolic profile evaluated by API20A | 250
    antimicrobial susceptibility testing performed by Etest | 250
    empirical treatment with vancomycin | 336
    empirical treatment with meropenem | 336
    discontinued vancomycin | 336
    discontinued meropenem | 336
    recovered from sepsis | 336
    <|eot_id|>
    