58 years old | 0
    man | 0
    visited a local hospital | 0
    sore throat | 0
    diagnosed with moderate pneumonia | -408
    COVID-19 | -408
    managed with oxygen | -408
    glucocorticoids | -408
    increased oxygen requirements | -408
    worsened pneumonia | -408
    developed severe respiratory fatigue | -391
    diagnosed with ARDS | -391
    hypertension | 0
    intubated | 0
    mechanical ventilation | 0
    tocilizumab | 0
    transferred to intensive care unit | 0
    venovenous ECMO | 0
    computed tomography showed bilateral and peripheral ground-glass and consolidative pulmonary opacities | 0
    developed hypotension | 9
    intra-abdominal bleed | 9
    right hemicolectomy | 9
    hemostasis confirmed | 9
    ileostoma created | 9
    histopathological examination revealed absence of morphological abnormalities | 9
    absence of aneurysms | 9
    absence of stenosis | 9
    absence of thrombi | 9
    absence of bacteria | 9
    absence of fungi | 9
    ileostoma exhibited ischemic changes | 27
    stomal reconstruction | 27
    ischemic changes adjacent to stoma | 27
    surgical wound necrosis | 27
    repeated debridement | 27
    no fungi in culture | 27
    thrombi | 27
    Mucorales | 27
    Grocott staining showed Mucorales invasion | 27
    respiratory improvement | 0
    SARS-CoV-2 antigen negative | 29
    SARS-CoV-2 antigen negative | 31
    multiple organ failure | 46
    death | 46
    autopsy revealed necrosis | 46
    thrombus in common iliac vein | 46
    necrosis of small intestine | 46
    necrosis of liver | 46
    necrosis of gall bladder | 46
    necrosis of right kidney | 46
    necrosis of spleen | 46
    Mucorales in thrombi | 46
    Mucorales in necrotic organs | 46
    Mucorales in stomach | 46
    Mucorales in urinary bladder | 46
    Rhizopus oryzae identified | 46
    absence of Mucorales in nasal cavity | 46
    absence of Mucorales in pharyngeal mucosa | 46
    absence of Mucorales in trachea | 46
    absence of Mucorales in lungs | 46
    absence of SARS-CoV-2 S proteins | 46
    myofibroblast proliferation | 46
    lymphocyte proliferation | 46
    diffuse alveolar damage | 46
    cytomegalovirus infection | 46
    no significant inflammation in heart | 46
    sepsis | 46
    multi-organ failure | 46
    mucormycosis | 46
    death | 46
    
    <|eot_id|>
    58 years old | 0
    man | 0
    visited a local hospital | 0
    sore throat | 0
    diagnosed with moderate pneumonia | -408
    COVID-19 | -408
    managed with oxygen | -408
    glucocorticoids | -408
    increased oxygen requirements | -408
    worsened pneumonia | -408
    developed severe respiratory fatigue | -391
    diagnosed with ARDS | -391
    hypertension | 0
    intubated | 0
    mechanical ventilation | 0
    tocilizumab | 0
    transferred to intensive care unit | 0
    venovenous ECMO | 0
    computed tomography showed bilateral and peripheral ground-glass and consolidative pulmonary opacities | 0
    developed hypotension | 9
    intra-abdominal bleed | 9
    right hemicolectomy | 9
    hemostasis confirmed | 9
    ileostoma created | 9
    histopathological examination revealed absence of morphological abnormalities | 9
    absence of aneurysms | 9
    absence of stenosis | 9
    absence of thrombi | 9
    absence of bacteria | 9
    absence of fungi | 9
    ileostoma exhibited ischemic changes | 27
    stomal reconstruction | 27
    ischemic changes adjacent to stoma | 27
    surgical wound necrosis | 27
    repeated debridement | 27
    no fungi in culture | 27
    thrombi | 27
    Mucorales | 27
    Grocott staining showed Mucorales invasion | 27
    respiratory improvement | 0
    SARS-CoV-2 antigen negative | 29
    SARS-CoV-2 antigen negative | 31
    multiple organ failure | 46
    death | 46
    autopsy revealed necrosis | 46
    thrombus in common iliac vein | 46
    necrosis of small intestine | 46
    necrosis of liver | 46
    necrosis of gall bladder | 46
    necrosis of right kidney | 46
    necrosis of spleen | 46
    Mucorales in thrombi | 46
    Mucorales in necrotic organs | 46
    Mucorales in stomach | 46
    Mucorales in urinary bladder | 46
    Rhizopus oryzae identified | 46
    absence of Mucorales in nasal cavity | 46
    absence of Mucorales in pharyngeal mucosa | 46
    absence of Mucorales in trachea | 46
    absence of Mucorales in lungs | 46
    absence of SARS-CoV-2 S proteins | 46
    myofibroblast proliferation | 46
    lymphocyte proliferation | 46
    diffuse alveolar damage | 46
    cytomegalovirus infection | 46
    no significant inflammation in heart | 46
    sepsis | 46
    multi-organ failure | 46
    mucormycosis | 46
    death | 46