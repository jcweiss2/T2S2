64 years old | 0
male | 0
admitted to the Intensive Care Unit (ICU) | 0
Escherichia coli Gram-negative septic shock | 0
purulent peritonitis | 0
rectosigmoid junction adenocarcinoma | 0
slightly disoriented | 0
hypotensive | 0
blood pressure of 110/55 mmHg | 0
lactic acidosis | 0
elevated white blood cell count (WBC) of 22680/μL | 0
PCT, 10 ng/mL | 0
renal insufficiency | 0
elevated creatinine, 1.88 mg/dL | 0
hyperglycemia, 263 mg/dL | 0
lactic acidosis (base excess -8.1 mmol/L, lactate 2 mmol/L) | 0
fluids resuscitation (crystalloids and albumin) | 0
broad-spectrum antibiotics | 0
meropenem 3g/24h | 0
metronidazole 1.5g/24h | 0
insulin | 0
invasive monitoring using a Vigileo monitor | 0
emergency surgical intervention | 0
persistence of intestinal subocclusions | 0
sepsis | 0
generalised purulent peritonitis | 0
septic shock | 0
perforation of the rectosigmoid junction adenocarcinoma | 0
rectosigmoid palliative resection | 0
abundant peritoneal lavage | 0
drainage | 0
bacteriological samples from the peritoneal fluid | 0
readmitted to the ICU | 24
intubated | 24
mechanically ventilated | 24
febrile | 24
persistent leukocytosis (WBC of 20090 /μL) | 24
elevated PCT levels (10 ng/mL) | 24
septic encephalopathy (GCS 10 points) | 24
vasoactive support with noradrenaline (0.11 μg/kg/min) | 24
adequate fluid transfusion | 24
minimally invasive haemodynamic monitoring | 24
hyperdynamic state | 24
cardiac output (CO) 7.3 L/min | 24
cardiac index ( CI ) 3.1 L/min/m2 | 24
systemic vascular resistance index (SVRI ) 1897 dyn*s/cm5*m2 | 24
SOFA score was 10 points | 24
APACHE II score was 23 points | 24
blood cultures | 24
urine cultures | 24
vancomycin (2g/24h) | 24
fluconazole (200mg/24h) | 24
adjunctive extracorporeal endotoxin adsorption treatment with an Alteco® LPS Adsorber | 24
double lumen 12Fr catheter introduced into the right femoral vein | 24
adsorber connected to an extracorporeal circuit including an HF 440 blood pump | 24
haemofiltration was not performed | 24
unfractionated heparin used to maintain APTT between 50 and 70 s | 24
blood flow rate set at 150 ml/min | 24
duration of the treatment was 120 minutes | 24
improvement in the hemodynamic status | 48
reduction in the noradrenaline infusion rate from 0.11 μg/kg/min to 0.07 μg/kg/minutes | 48
increase in MAP from 85 mmHg to 99 mmHg | 48
CI pretreatment levels of 3,1 L/min/m2 to 3,7 L/min/m2 | 48
PaO2 reducing from 124 mmHg to 109 mmHg | 48
PaO2/FiO2 from 354 to 311.4 | 48
reduction in PCT levels from 10 ng/mL to 4 ng/mL | 48
decrease in lactate levels from 1.9 mmol/L to 1.37 mmol/L | 48
decrease in the SOFA score from 10 points to 7 points | 48
postoperative complication with a localised peritonitis | 216
ischemic bowel perforation | 216
died | 264
