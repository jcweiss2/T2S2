38 year-old | 0
woman | 0
returned from Bali | -672
no pre travel consultation | -672
no malaria prophylaxis | -672
close contact with people in poor conditions | -672
saw rats around accommodation | -672
recalled mosquito bites | -672
sporadic contact with dogs and cats | -672
no scratching or biting episodes | -672
returned to Portugal asymptomatic | -672
presented to emergency department | -168
fever | -168
chills | -168
malaise | -168
myalgia | -168
conjunctival congestion | -168
unremarkable blood tests | -168
normal chest X-Ray | -168
negative malaria test | -168
negative dengue test | -168
discharged home | -168
acetaminophen treatment | -168
re-evaluated in ambulatory | -144
fever persisted | -144
malaise persisted | -144
myalgia persisted | -144
good general condition | -144
normal physical examination | -144
relative neutrophilia | -144
elevated hepatic aminotransferases | -144
elevated LDH | -144
mildly increased CRP | -144
normal chest X-ray | -144
normal abdominal ultrasonography | -144
blood cultures collected | -144
serologic screen requested | -144
admitted to Infectious Diseases Ward | -144
clinical deterioration | 0
analytical deterioration | 0
shortness of breath | 0
respiratory rate 32/minute | 0
SatO2 90-92% | 0
hypotension | 0
headache | 0
nausea | 0
faint transient macular rash | 0
acutely ill appearance | 0
respiratory alkalosis | 0
pO2/FiO2 ratio 327 | 0
hyperlactacidemia | 0
bilateral interstitial infiltrate | 0
interstitial pneumonia | 0
admitted to ICU | 0
IV fluids | 0
IV ceftriaxone | 0
IV doxycycline | 0
oseltamivir | 0
oxygen support | 0
new microbiological exams requested | 0
condition improved progressively | 24
no invasive ventilation needed | 24
no vasopressive support needed | 24
oliguria reverted | 24
transient hemoglobin decrease | 24
worsening thrombocytopenia | 24
coagulopathy | 24
spontaneous recovery | 24
afebrile by day 4 | 96
discharged from ICU | 120
fully recovered by day 7 | 168
ceftriaxone given for 8 days | 168
doxycycline given for 14 days | 168
discharged from hospital | 312
asymptomatic at discharge | 312
chest X-ray resolution | 312
PCR positive for Rickettsia spp. | 312
negative other microbiological exams | 312
seroconversion confirmed | 624
IgM 1:2048 | 624
IgG 1:4096 | 624
rickettsial DNA detected | 624
R. typhi confirmed | 624
