33 years old | 0
female | 0
fever | -96
cough | -96
dyspnoea | -96
admission | 0
hypoxemia | 0
high-flow nasal cannula therapy | 0
empiric antimicrobial therapy | 0
steroids | 0
methylprednisolone | 0
broad-spectrum antibiotics | 0
pulmonary consolidation | 0
computed tomography scan | 0
percutaneous lung biopsies | 0
histologically | 0
alveolar spaces filled with fibrin balls | 0
fibroblastic tissue | 0
no hyaline membranes | 0
no eosinophils | 0
AFOP diagnosis | 0
transfer to ICU | 0
broad-spectrum antibiotics | 0
high-dose steroids | 0
high-dose immunoglobulins | 0
respiratory failure | 0
orotracheal intubation | 0
mechanical ventilation | 0
invasive ventilation | 0
echocardiography | 0
normal biventricular function | 0
no valve defects | 0
no septal defects | 0
no pulmonary hypertension | 0
venovenous ECMO support | 0
lung rest approach | 0
multidisciplinary team discussion | 336
lung transplantation group | 336
lung transplant emergency waiting list | 336
informed consent | 336
donor lung | 480
bilateral lobar lung transplantation | 480
tacrolimus | 480
methylprednisolone | 480
induction therapy | 480
carbapenem-resistant Pseudomonas aeruginosa pneumonia | 480
exophytic granulation tissue | 480
inflammation | 480
anastomotic stenosis | 480
trachea | 480
bronchopleural fistulae | 512
anastomotic infections | 512
septic shock | 512
bacteraemia | 512
reperfusion syndrome | 512
primary graft dysfunction | 512
severe renal failure | 512
dialysis | 512
critical illness myopathy | 512
prophylactic antifungal therapy | 512
prophylactic antiviral therapy | 512
renal replacement therapy | 512
percutaneous drainage | 512
airway debridement | 512
cryotherapy | 512
electrocautery | 512
laser | 512
bronchoscopic balloon dilatation | 512
immunosuppression | 512
respiratory rehabilitation | 512
weaning ECMO | 672
weaning MV | 1440
tracheostomy | 576
discharge | 720
survival | 8760
no readmissions | 8760
return to normal daily life | 8760
return to social activity | 8760