27 years old | 0
female | 0
sickle cell disease | -8760
autosplenectomy | -8760
Crigler-Najjar syndrome | -8760
cholecystectomy | -8760
hydroxyurea | -8760
discontinued hydroxyurea | -720
right lower extremity ulcer | -720
Voxelotor | -720
Voxelotor 1.5 g oral daily | -720
sickle cell pain crises | -720
fatigue | -720
anemia | -720
admitted to the Emergency Department | 0
bilateral arm pain | 0
back pain | 0
leg pain | 0
dyspnea on exertion | 0
no chest pain | 0
hydromorphone | 0
intravenous fluids | 0
normal saline | 0
supplemental oxygen | 0
hemodynamically stable | 0
anemia | 0
baseline hemoglobin levels | 0
Chest X-ray | 0
no cardiopulmonary infiltrates | 0
admitted to the medical floor | 0
hydromorphone | 0
Oxycontin | 24
maintenance fluids | 24
bedside incentive spirometry | 24
Voxelotor discontinued | 24
bicytopenia | 48
anemia | 48
thrombocytopenia | 48
worsening hemolysis | 48
hyperkalemia | 48
worsening renal function | 48
hypoxia | 48
oxygen saturation 70% | 48
oxygen supplementation | 48
Venturi-Mask | 48
thrombotic thrombocytopenic purpura suspected | 48
LDH 2646 U/L | 48
schistocytes on peripheral blood smear | 48
PLASMIC score 4 | 48
critical care consulted | 48
transferred to the Medical Intensive Care Unit | 48
double-lumen Shiley central venous catheter placed | 48
total plasma exchange therapy | 48
RBCs transfusion | 48
high-dose intravenous methylprednisolone | 48
ADAMTS13 level activity 64.9% | 72
improvement after plasma exchange | 72
platelets improved | 72
creatinine improved | 72
LDH improved | 72
discharged home | 120
Voxelotor restarted | 120
lower dose | 120