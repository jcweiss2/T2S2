21 years old | 0
female | 0
admitted to ICU | 0
high grade fever | -192
chills | -192
respiratory distress | -144
altered sensorium | -48
intubated | -48
mechanical ventilation | -48
shock | 0
vasopressors infusions | 0
edematous peripheries | 0
right upper limb swelling | 0
leukocytopenia | 0
thrombocytopenia | 0
normal prothrombin time | 0
normal activated partial thromboplastin | 0
normal thrombin times | 0
normal fibrinogen levels | 0
right IJV thrombus | 0
absence of venous flow in color Doppler | 0
left IJV and SCV compressible | 0
left IJV and SCV patent | 0
central line insertion in left SCV | 0
radiological confirmation of right IJV thrombus | 0
right IJV thrombus with extension towards right SCV | 0
lower limb Doppler study normal | 0
mild tricuspid regurgitation | 0
ejection fraction <55% | 0
mild dilatation of main pulmonary arteries | 0
left distal pulmonary artery thrombosis | 0
unfractionated heparin started | 0
APC-R | 0
homozygous Factor V Leiden mutation | 0
oral vitamin K anticoagulants started | 24
target INR achieved | 120
heparin stopped | 120
warfarin continued | 120
Dengue IgM positive | 24
hemodynamic status improved | 168
weaned off from ventilator | 168
shock recovered | 168
thrombophilia testing | 168
right upper limb swelling regressed | 168
right IJV and SCV thrombus persisted | 168
partial recanalization | 168
discharged on oral warfarin treatment | 240
father, mother, and younger sister underwent factor 5 Leiden mutation test | 240
factor 5 Leiden mutation test negative | 240