15 years old | 0
female | 0
acute myelogenous leukemia (AML) | 0
standard induction treatment | 0
chemotherapy according to AML-BFM guidelines | 0
second cycle of chemotherapy | -672
pancytopenia | -672
infection with unknown focus | -672
ciprofloxacin | -672
linezolid | -672
meropenem | -672
tobramycin | -672
liposomal amphotericin | -672
after 3 weeks of treatment | -504
tachycardia (140/min) | -504
hypotension (75/41 torr) | -504
lactic acidosis | -504
admitted to the pediatric intensive care unit | 0
transthoracic echocardiography | 0
severely impaired left ventricular ejection fraction (LVEF) of 12% | 0
no dilatation of the left ventricle (LVIDd 38 mm) | 0
electrocardiogram showed sinus tachycardia | 0
incomplete right bundle branch block | 0
NT-proBNP 19 384 pg/ml | 0
high-sensitive troponin T 53.7 pg/ml | 0
fluid therapy | 0
noradrenaline | 0
dobutamine | 0
milrinone | 0
deep sedation | 0
mechanical ventilation | 0
respiratory insufficiency | 0
lactate acidosis worsened (16 mmol/l, pH 6.91) | 0
hypotonic (50/30 torr) | 0
heart rate of 160/min | 0
va-ECMO initiation | 0
cannulation of the left femoral artery and vein | 0
13 Fr/15 cm arterial cannula | 0
21 Fr/55 cm venous cannula | 0
Seldinger technique | 0
sonographic guidance | 0
9 Fr sheath in left superficial femoral artery | 0
ECMO blood flow of 3.3 l/min at 3800 rpm | 0
pre-oxygenator membrane pressure above 350 torr | 0
mean arterial pressure (MAP) 45 torr | 0
noradrenaline (80 µg/min) | 0
vasopressin (2 units/h) | 0
levosimendan (0.5 mg/h) | 0
hydrocortisone (200 mg/d) | 0
residual LVEF 10–15% | 0
CVVHDF | 0
anuric acute kidney injury | 0
continued anti-infective therapy | 0
dose-adjustment of meropenem | 0
ciprofloxacin | 0
metronidazole | 0
cotrimoxazole | 0
liposomal amphotericin B | 0
acyclovir | 0
linezolid replaced by vancomycin | 0
PCT 2.37 ng/ml | 0
CRP 2.98 mg/dl | 0
second day with vaA-ECMO | 24
MAP declined to 40 torr | 24
increased vasopressors | 24
noradrenaline 144 µg/min | 24
vasopressin 4 IE/h | 24
LVEF decreased below 10% | 24
levosimendan infusion stopped | 24
acute ischemic injury of non-cannulated leg | 24
right femoral artery dissection | 24
no embolic event | 24
insufficient blood inflow | 24
low cardiac output | 24
leg ischemia | 24
lactate levels rose to 25 mmol/l | 24
Dacron® conduit on right femoral artery | 24
second arterial cannula (13 Fr/15 cm) | 24
Y-connector connection | 24
ECBF enhanced to 4–5 l/min | 24
pre-oxygenator membrane pressures below 300 torr | 24
MAP maintained at 40–50 torr | 24
ECBF limited by venous drainage pressures below –100 mmHg | 24
sufficient preload verified by echocardiography | 24
inspiratory oxygen fraction increased to 0.55 | 24
prevent harlequin syndrome | 24
impaired lung function | 24
arterial oxygen partial pressure normal | 24
PCT levels rose to 42.5 ng/ml | 24
Hickman catheter explanted | 24
no causal organism identified | 24
broad-complex tachycardia | 24
treated with esmolol | 24
treated with metoprolol | 24
left ventricular function further decreased | 24
aortic valve ceased to open | 24
second venous cannula (21 Fr/55 cm) | 24
right femoral vein into left atrium | 24
percutaneous atrioseptostomy | 24
ECBF 5–6 l/min at 3850–4200 rpm | 24
lactate levels peaked at 29 mmol/l | 24
lactate levels fell instantly | 24
MAP rose from nadir 30 torr | 24
acidosis leveled out | 24
cerebral oximetry showed regional oxygen saturation 60–80% | 24
echocardiography showed left ventricle unloaded | 24
no residual left ventricular function | 24
therapeutic anticoagulation | 24
unfractionated heparin | 24
target partial thrombin time 60–80 s | 24
PCT peaked at 80.4 ng/ml | 72
CRP peaked at 7.23 mg/dl | 72
leukocytes 300/µl | 72
high-sensitive troponin T 343 pg/ml | 72
creatine kinase MB 178 U/l | 72
total creatine kinase 577 U/l | 72
all microbial specimens negative | 72
viral myocarditis excluded | 72
myocardial biopsy | 72
cardiac systolic function gradually recovered | 120
day 5 | 120
ECMO cannulas removed from left femoral vessels | 120
day 7 | 168
ECMO completely removed | 168
LVEF recovered to approximately 30% | 168
mean arterial pressures 60–70 torr | 168
transseptal cannula removal | 168
no relevant atrial communication | 168
CVVHDF stopped | 168
normal renal function | 168
leucocyte count recovered to 1000/µl | 312
day 13 | 312
normal leucocyte values on day 30 | 720
respirator weaning on day 33 | 792
allogenic stem cell transplantation | 1008
discharged after 5 months | 3600
severe critical illness polyneuropathy | 3600
LVEF recovered to approximately 40% | 3600
no ventricular dilatation | 3600
