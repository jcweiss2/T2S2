75 years old | 0
male | 0
admitted to the Department of Urology | 0
diabetes mellitus | -672
hypertension | -672
left flank pain | 0
dysuria | 0
high fever | 0
minimal blood urea nitrogen (BUN) increase | 0
creatinine increase | 0
glycosuria | 0
albuminuria | 0
leukocyturia | 0
urine culture documented an infection from Candida albicans | 0
antimycotic treatment by fluconazole | 0
wide spectrum antibiotic coverage with meropenem | 0
abdominal ultrasound evidenced multiple bilateral kidney stones | 0
left early hydronephrosis | 0
left pyelostomy | 72
septic shock | 72
transferred to the intensive care unit (ICU) | 72
renal function improved | 168
readmitted to the urology department | 168
double J ureteral stent was placed | 168
antimycotic treatment was stopped | 4032
discharged home | 4032
sensory obtundation | 5184
blurred speech | 5184
development of weakness in the right arm and leg | 5184
stuporous but arousable | 5184
right hemiparesis | 5184
sensory-motor aphasia | 5184
erythrocyte sedimentation rate (ESR) increase | 5184
modest monocytosis | 5184
admission computed tomography (CT) scan disclosed a left parietal epidural mass | 5184
magnetic resonance imaging (MRI) disclosed a diffuse ipsilateral hemispheric leptomeningeal enhancement | 5184
emergency surgery at the left fronto-temporal-parietal craniotomy | 5184
durotomy | 5184
en bloc removal of the lesion | 5184
duroplasty was performed by Tutopatch | 5184
bone was repositioned by titanium miniplates | 5184
postoperative course was uneventful | 5188
CT and MRI scans confirming full lesion removal | 5188
antimycotic treatment with amphotericin B | 5188
meropenem | 5188
full midline re-alignment and a small subdural hygroma | 5376
discharged to a rehabilitation facility | 5376
high fever | 7776
impaired consciousness | 7776
aphasia | 7776
fluctuating subcutaneous collection | 7776
subcutaneous and epidural empyema | 7776
re-surgery | 7776
huge, purulent collection was found | 7776
pus was found overlying the rebuilt dural layer | 7776
large spectrum antibiotics were started | 7776
ceftriaxone | 7776
teicoplanin | 7776
no growth of bacteria or fungi was observed from cultures | 8112
therapy was interrupted | 8112
two months post-operative CT scan showed no residual contrast enhancement | 8512
discharged again to a rehabilitation facility | 8512
contrast enhanced MRI was found negative | 10944
premodeled titanium cranioplasty was positioned | 10944
discharged home with no residual deficits | 10944