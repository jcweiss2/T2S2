28 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
attended a health center | -48 | -48 | Factual
fatigue | -48 | 0 | Factual
anosmia | -48 | 0 | Factual
dyspnea | -48 | 0 | Factual
SpO2 levels were 55% | -48 | -48 | Factual
nasal cannula oxygen therapy | -48 | 0 | Factual
SpO2 levels improved to 75% | -48 | 0 | Factual
hospitalized | -48 | -48 | Factual
evaluated at an emergency department | -48 | -48 | Factual
chest radiography | -48 | -48 | Factual
bilateral lung infiltrates | -48 | 0 | Factual
RT-PCR swab tested positive for SARS-CoV-2 infection | -48 | -48 | Factual
admitted in a COVID-19 infirmary unit | -48 | -48 | Factual
non-invasive ventilation support | -48 | -24 | Factual
intubation | -24 | -24 | Factual
invasive mechanical ventilation | -24 | 0 | Factual
ventral decubitus positioning | -24 | 0 | Factual
Escherichia coli detected on sputum culture | -48 | -48 | Factual
methicillin-sensitive Staphylococcus aureus detected on sputum culture | -48 | -48 | Factual
superinfection | -48 | 0 | Factual
amoxicillin | -48 | -40 | Factual
blood culture revealed methicillin-resistant Staphylococcus aureus | -48 | -48 | Factual
methicillin-resistant Staphylococcus aureus dismissed | -48 | -48 | Factual
steady clinical improvement | -24 | 0 | Factual
extubated | 0 | 0 | Factual
discharged | 0 | 0 | Factual
retrosternal thoracalgia | 168 | 168 | Factual
thoracalgia irradiating to the left upper limb | 168 | 168 | Factual
abduction and external rotation limited due to pain | 168 | 168 | Factual
soft tissue swelling of the shoulder and arm | 168 | 168 | Factual
fever | 168 | 168 | Factual
increased levels of C-reactive protein | 168 | 168 | Factual
hemoculture proved negative | 168 | 168 | Factual
urine culture proved negative | 168 | 168 | Factual
chest radiograph | 168 | 168 | Factual
thoracic CT | 168 | 168 | Factual
typical changes compatible with sequelae of Covid-19 pneumonia | 168 | 168 | Factual
admitted for further investigation and treatment planning | 168 | 168 | Factual
gentamicin prescribed | 168 | 216 | Factual
gentamicin administered | 168 | 216 | Factual
thoracic CT with intravenous contrast administration | 216 | 216 | Factual
scapulohumeral synovitis | 216 | 216 | Factual
intra-muscular collections | 216 | 216 | Factual
glenohumeral joint fluid | 216 | 216 | Factual
bilateral shoulder magnetic resonance imaging (MRI) | 240 | 240 | Factual
infraspinatus fossa and subscapular fossa collections | 240 | 240 | Factual
capsular thickening | 240 | 240 | Factual
increased signal intensity post-gadolinium administration | 240 | 240 | Factual
septic arthritis | 240 | 240 | Factual
rotator cuff collections | 240 | 240 | Factual
myonecrosis | 240 | 240 | Factual
aspiration of the infraspinatus fossa collection | 240 | 240 | Factual
seropurulent fluid | 240 | 240 | Factual
drainage catheter | 240 | 240 | Factual
drainage catheter removed | 240 | 240 | Factual
evaluation of the aspirate | 240 | 240 | Factual
direct and culture tests for Mycobacterium tuberculosis | 240 | 240 | Factual
anaerobic and aerobic bacteria | 240 | 240 | Factual
negative results | 240 | 240 | Factual
improvement of left shoulder range of motion | 240 | 288 | Factual
physical rehabilitation exercises | 240 | 288 | Factual
transferred to another hospital | 288 | 288 | Factual
continue physical therapy and rehabilitation exercises | 288 | 288 | Factual