11 years old | 0
female | 0
admitted to the hospital | 0
posterior spinal fusion | -12
propofol | -12
hypotension | -12
blood products | -12
vasopressors | -12
phenylephrine | -12
norepinephrine | -12
extubated | -12
disseminated intravascular coagulation | -24
liver injury | -24
rhabdomyolysis | -24
oliguria | -24
fluid resuscitation | -24
reintubated | -24
high-dose i.v. diuretics | -24
CRRT | 5
selective cytopheretic device | 7
rhabdomyolytic AKI | 0
respiratory failure | 0
severe liver injury | 0
coagulopathy | 0
propofol infusion syndrome | 0
PRIS | 0
cardiac failure | 0
hyperlipidemia | 0
AKI | 0
multiorgan failure | 0
excessive systemic inflammatory response | 0
microvascular dysfunction | 0
capillary leak | 0
tissue ischemia | 0
LE infiltration | 0
toxic byproducts | 0
liver enzymes | 0
pancreatic enzymes | 0
amylase | 0
lipase | 0
triglyceride | 0
white blood count | 0
DIC | 0
protime | 0
partial thromboplastin time | 0
lactate dehydrogenase | 0
d-dimer | 0
haptoglobin | 0
respiratory failure | 0
mechanical ventilation | 0
fraction of inspired oxygen | 0
partial arterial pressure of oxygen | 0
PaO2/fraction of inspired oxygen ratio | 0
broad spectrum antibiotics | 24
procalcitonin | 24
temperature | 24
white blood count | 24
infection | 24
net volume removal | 48
CRRT discontinued | 168
discharged | 480
renal function | 0
urine output | 72
serum creatinine | 0
lactate | 0
bicarbonate | 0
pH | 0
partial pressure of carbon dioxide | 0
ionized calcium | 7
circuit ionized calcium | 7
blood gas analyzer | 7
elution buffer | 24
elution | 24
cytometric analysis | 24
CD11b | 24
mean fluorescent intensity | 24
MFI | 24
sepsis | 120
systemic infection | 120
neutrophils | 0
monocytes | 0
lymphocytes | 0
leukocytes | 0
cell biomarker | 0
systemic inflammation | 0
critically ill patients | 0
device-related adverse events | 0
safety characteristics | 0
efficacy clinical trials | 0
pediatric patients | 0
adult patients | 0
FDA | 0
Investigational Device Exemption | 0
ClinicalTrials.gov | 0
University of Michigan | 0
CytoPherx | 0
Innovative BioTherapies, Inc. | 0
FDA Grant | 0
US FDA | 0