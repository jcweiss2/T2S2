85 years old | 0
female | 0
admitted to the hospital | 0
discomfort | -168
moderate fever | -168
vomiting | -168
referred to the emergency department | -24
CT scan | -24
lower para-oesophageal pleuro-mediastinal collection | -24
thickened wall of the oesophagus | -24
diagnosed with perforated oesophageal cancer | -24
palliation of symptoms | -24
referred to the emergency department of our hospital | -24
conscious | 0
normal breathing | 0
moderately febrile | 0
normal blood pressure | 0
normal heart rate | 0
elevated white blood cell count | 0
elevated C-reactive protein | 0
minimal liver impairment | 0
minimal renal impairment | 0
episode of vomiting | -168
fever | -168
malaise | -168
oral feeding | -168
CT scan | 0
oral contrast | 0
para-oesophageal mediastinal collection | 0
left pleural collection | 0
left thoracotomy | 0
smelly purulent collection | 0
debrided | 0
necrotic tissues removed | 0
distal third of the oesophagus isolated | 0
perforation | 0
necrotic tissues around the perforation removed | 0
mucosal layer exposed | 0
stay sutures placed | 0
mucosal edges grasped with Allis clamp | 0
endoscopic articulating linear cutter used | 0
mucosa sutured | 0
nasogastric tube placed | 0
gastric fundus mobilized | 0
gastric wrap created | 0
chest drainages placed | 0
Escherichia coli cultured | 0
Enterococcus faecalis cultured | 0
postoperative course complicated | 24
left lower lobe pneumonia | 24
systemic infection | 24
multidrug-resistant Klebsiella pneumoniae | 24
CT scan with oral contrast | 216
seal of the repair confirmed | 216
residual collections excluded | 216
resumed creamy diet | 216
chest drains removed | 264
discharged home | 648
normal diet | 648
oesophagogram performed | 744
contrast study of the oesophagus | 744
no transit discomfort | 744