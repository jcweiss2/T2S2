3 years old | 0
male | 0
vaccinated | 0
no significant past medical history | 0
admitted to the pediatric emergency department | 0
chief complaint of cough | 0
cough | -168
nasal congestion | -168
sore throat | -24
no history of fever | -168
no dyspnea | -168
no history of trauma | -168
no recent travel | -168
tolerating solids and liquids well | 0
taking a cough suppressant | -168
taking ibuprofen | -168
symptomatic relief | -168
well appearing | 0
afebrile | 0
hemodynamically stable | 0
temperature 36.7°C | 0
pulse 113 | 0
respiratory rate 23 | 0
pulse oximetry 98% on room air | 0
nasal congestion | 0
erythematous pharynx | 0
able to drink fluids | 0
discharged home | 0
diagnosis of a viral syndrome | 0
presented to another pediatric ED | 72
congestion | 72
sore throat | 72
torticollis | 72
limited range of motion of his neck | 72
drooling | 72
tactile fever | -24
self-resolved | -24
no history of vomiting | 72
temperature 37.5°C | 72
pulse 121 | 72
blood pressure 102/60 | 72
respiratory rate 24 | 72
pulse oximetry 100% on room air | 72
well-appearing and well-hydrated child | 72
diffuse neck tenderness | 72
no associated lymphadenopathy | 72
left-sided torticollis | 72
no significant trismus | 72
no evidence of meningismus | 72
elevated WBC | 72
elevated CRP | 72
mild hypoglycemia | 72
slightly low serum bicarbonate level | 72
concerns for a possible retropharyngeal abscess | 72
soft tissue neck plain film | 72
diffuse paravertebral swelling | 72
2.2 cm linear radiopaque density | 72
possible foreign body | 72
eating fish earlier in the week | -168
given a dose of antibiotics | 72
transferred to another pediatric facility | 72
consultation with a pediatric otolaryngology surgeon | 72
ENT consulted | 72
evaluated the patient | 72
repeat soft tissue neck plain film | 72
2.2 cm linear radiopaque density within the prevertebral soft tissues | 72
taken to the operating room | 72
rigid esophagoscopy | 72
purulent fluid in the cervical esophagus | 72
drained | 72
2 cm fish bone | 72
removed | 72
Penrose drain placed | 72
esophageal perforation | 72
abscess | 72
postoperative computed tomography scan | 72
no residual foreign body | 72
no residual abscess | 72
admitted to the pediatric intensive care unit | 72
broad-spectrum antibiotics | 72
clindamycin | 72
ampicillin/sulbactam | 72
positive wound cultures | 72
Gram stain of gram-positive cocci in pairs | 72
Penrose drain removed | 72
discharged home | 120
tolerating feeds | 120
on oral clindamycin | 120
no evidence of persistent abscess | 120
no esophageal perforation | 120
ENT follow up | 120