64 years old | 0
    male | 0
    alcohol consumption | 0
    liver cirrhosis | 0
    emergency department admission | 0
    two-day history of productive cough | -48
    exertional dyspnea | -48
    temperature 36 °C | 0
    blood pressure 100/60 mmHg | 0
    heart rate 78 bpm | 0
    respiratory rate 19 bpm | 0
    oxygen saturation 96% in ambient air | 0
    round opacity in right upper lobe on chest X-ray | 0
    laboratory tests within normal ranges | 0
    antibiotic therapy started with ceftriaxone and clarithromycin | 0
    sputum culture positive for E. hormaechei | 0
    E. hormaechei sensitive to levofloxacin | 0
    therapy modified to levofloxacin | 0
    systemic respiratory distress syndrome | 48
    intubated | 48
    transferred to ICU | 48
    mechanical ventilation with lung-protective strategy | 48
    hemodynamic instability | 48
    additional blood cultures drawn | 48
    antibiotic therapy escalated to imipenem/cilastatin | 48
    death due to septic shock | 48
