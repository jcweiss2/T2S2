42 years old | 0
Caucasian | 0
female | 0
diagnosed with acetylcholine receptor antibody positive oculo-bulbar myasthenia gravis | -6578
drooping eyelids | -6578
double vision | -6578
difficulty swallowing | -6578
diurnal variation | -6578
characteristic fluctuation of symptoms | -6578
failed bedside swallow evaluation | -6578
aspiration to thin liquids on modified barium swallow | -6578
plasmapheresis | -6578
complete resolution of symptoms | -6578
IVIG | -6578
repetitive nerve stimulation study | -6578
antibody titers confirmed diagnosis of postsynaptic neuromuscular junction disorder | -6578
started pyridostigmine 60 mg 4 times daily | -6578
gradually up-titrated dose of prednisone 30 mg daily | -6578
mycophenolate 1000 milligrams twice daily | -6578
generalized anxiety disorder | 0
allergic rhinitis | 0
recurrence of drooping eyelids | -6578
change in voice | -6578
concerns of impending myasthenia exacerbation | -6578
started regular plasma exchange | -6578
3 exchanges every 4 weeks | -6578
continued prednisone 30 mg daily | -6578
continued mycophenolate 1000 milligrams twice daily | -6578
CT chest showed 6.7 cm lobulated soft tissue mass in anterior mediastinum | -6578
no local invasion | -6578
referred to cardiothoracic surgery for possible thymectomy | -6578
thymectomy put on hold due to patient request | -6578
presented to emergency department with fever | -672
chills | -672
cough with minimal clear sputum production | -672
exertional shortness of breath | -672
decreased sense of taste | -672
decreased sense of smell | -672
decreased appetite | -672
traveled to nearby city two weeks prior to presentation | -1344
no clear history of exposure to sick | 0
no history of similar symptoms in friends or family | 0
chest x-ray showed patchy infiltrates in left lower lobe | 0
elevated white count (12.32×109/L) | 0
lymphopenia (0.78×109/L) | 0
negative respiratory pathogen panel (influenza A/B, Streptococcus pneumonia) | 0
negative urine Legionella | 0
COVID-19 RT-PCR positive | 0
bedside negative inspiratory force (NIF) 65 cm H2O | 0
discharged from emergency department | 0
self-quarantine for fourteen days | 0
follow CDC guidelines | 0
clear instructions to return to emergency department if symptoms worsened | 0
continued immunomodulatory therapy (prednisone, mycophenolate) | 0
plasmapheresis deferred to post quarantine period | 0
recovered from COVID-19 infection | 0
no complications | 0
no symptoms of myasthenic crisis | 0
no myasthenia exacerbation | 0
no changes to immunosuppressive medications | 0
