22 years old | 0
woman | 0
referred by critical care team of district general hospital to regional burns unit | 0
100% TBSA involvement | 0
toxic epidermal necrolysis | 0
GPA (Granulomatosis with polyangiitis) | 0
initially presented to DGH with fever | -240
initially presented to DGH with shortness of breath | -240
initially presented to DGH with feeling generally unwell | -240
chest X-ray demonstrated multiple opacities | -240
CT of chest and abdomen found multiple cavitations | -240
CT of chest and abdomen found pulmonary embolism | -240
CT of chest and abdomen found femoral thrombosis | -240
GPA confirmed | -240
commenced on warfarin | -240
commenced on rituximab | -240
commenced on methylprednisolone | -240
commenced on Immunoglobulins (IgG) | -240
commenced on fluconazole | -240
responded well to treatment | -240
second infusion of rituximab | -168
third infusion of rituximab | -168
prophylactic co-trimoxazole | -168
presented back to DGH with angioedema | -72
developed rash with 90% TBSA | -72
involving oral mucosa | -72
involving ophthalmic mucosa | -72
fluconazole stopped | -72
co-trimoxazole stopped | -72
steroids increased | -72
initial suspicion of Stevens–Johnson syndrome | -72
patient deteriorated | -72
progressed to 100% TBSA | -72
required significant support from critical care team | -72
TEN suspected | -72
TEN confirmed by skin biopsy | -72
initial SCORTEN score of 3 | -72
predicting 35.3% mortality risk | -72
referred to specialist burns centre | -72
transferred to specialist burns centre | -72
piperacillin/tazobactam (Tazocin) commenced | 0
vancomycin commenced | 0
sputum sensitivities | 0
wound swab sensitivities | 0
prednisolone reduced to 40 mg daily | 168
good re-epithelisation of skin | 240
discharged | 504
period of physiotherapy | 504
