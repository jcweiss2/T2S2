54 years old | 0
man | 0
chronic obstructive pulmonary disease | -87600
obstructive sleep apnea | -87600
continuous positive airway pressure | -87600
Fournier’s gangrene | 0
acute renal failure | 0
sepsis | 0
admitted to the emergency department | 0
coronary artery disease | -87600
percutaneous coronary intervention | -87600
stenting | -87600
30 pack-year smoking history | -87600
morbid obesity | 0
respiratory failure | 0
metabolic acidosis | 0
respiratory distress | 0
tachypnea | 0
diffuse bilateral wheezing | 0
mouth opening of three finger-breadths | 0
Mallampati airway classification 3 | 0
thyromental distance of 6 cm | 0
neck circumference of 44 cm | 0
blood oxygen saturation 99% | 0
fraction of inspired oxygen of 0.5 | 0
cyanotic | 0
blood oxygen saturation ~85% | 0
increased intensity during inspiration | 0
coarse, low-pitched wheezing | 0
dyspnea | 0
bronchodilators | 0
elevated prothrombin time of 24 seconds | 0
international normalized ratio, 3.6 | 0
septic shock | 0
awake fiberoptic endotracheal intubation | 0
fiberoptic intubation | 0
semi-Fowler’s position (45°) | 0
bilateral superior laryngeal nerve block | 0
transtracheal instillation of 4% lidocaine | 0
tracheomalacia | 0
endotracheal tube | 0
debridement of Fournier’s gangrene | 0
hypotension | 0
vasoactive agents (phenylephrine) | 0
arterial blood gas pH 7.26 | 0
partial pressure of carbon dioxide 34 mmHg | 0
partial pressure of oxygen 320 mmHg | 0
HCO3− levels of 16.0 | 0
base excess −11 | 0
blood oxygen saturation 100% | 0
remained intubated | 0
transferred to the intensive care unit | 0
antibiotics | 0
inotropic support | 0
pressure-regulated volume control ventilation | 0
fraction of inspired oxygen of 1.0 | 0
respiratory rate of 20 breaths per minute | 0
peak inspiratory pressure of 25 mmHg | 0
positive end-expiratory pressure of 7 mmHg | 0
acute respiratory distress syndrome | 0
computed tomography scan bilateral infiltrates | 0
multiorgan dysfunction | 120
hepatic dysfunction | 120
renal dysfunction | 120
cardiac dysfunction | 120
pulmonary dysfunction | 120
succumbed | 120
respiratory failure |4 0
