40 years old | 0
male | 0
admitted to the hospital | 0
hypertension | -8760
atrial fibrillation | -8760
severe uncontrolled hyperthyroidism | -8760
thyroid storm | -8760
intubation | -8760
central chest pain | -2
palpitation | -2
agitation | -2
nausea | -2
blood pressure 181/112 mmHg | 0
heart rate 140 beats/min | 0
tachypneic | 0
respiratory rate 38/min | 0
temperature 37.6°C | 0
oxygen saturation 85% | 0
anxious | 0
agitated | 0
diffuse goiter | 0
clammy skin | 0
warm skin | 0
bibasilar crackles | 0
fast AF | 0
ST-segment elevation | 0
mild leukocytosis | 0
normal hemoglobin | 0
normal platelets | 0
normal renal function | 0
normal liver function | 0
ProBNP 1100 pg/Ml | 0
thyroid-stimulating hormone undetectable | 0
serum Thyroxin more than 100 pmol/L | 0
Burch-Wartofsky Point Scale 60 | 0
serum troponin T level 1200 ng/L | 0
acute anterior wall MI | 0
thyroid storm | 0
dual antiplatelet therapy | 0
aspirin | 0
clopidogrel | 0
unfractionated heparin infusion | 0
propylthiouracil 200 mg | 0
hydrocortisone 200 mg | 0
cholestyramine 4 mg | 0
Lugol's solution 10 drops | 0
isosorbide dinitrate infusion | 0
furosemide 40 mg | 0
chest pain progression | 2
tachypneic | 2
IV furosemide | 2
isosorbide dinitrate infusion increased | 2
high-risk CAG | 2
coronary angiography | 2
percutaneous coronary intervention | 2
single vessel disease | 2
distal left anterior descending artery 100% embolic occlusion | 2
TIMI 3 | 2
blood flow restored | 2
chest pain settled | 2
ECG changes improved | 2
ejection fraction 35% | 2
anterior wall motion hypokinesia | 2
grade 2 diastolic dysfunction | 2
moderately dilated left atrium | 2
clinical status stabilized | 24
bisoprolol | 24
IV furosemide changed to oral | 24
oxygen saturation improved | 24
ECG exhibited AF with controlled ventricular response | 168
T wave inversion | 168
thyroxin level improved | 168
hydrocortisone tapered down | 168
cholestyramine stopped | 168
Lugol's solution stopped | 168
propylthiouracil switched to carbimazole | 168
discharge | 168
DAPT | 168
rivaroxaban | 168
rosuvastatin | 168
furosemide | 168
bisoprolol | 168
spironolactone | 168
valsartan | 168
clinically stable | 720
compliant with medications | 720
ECG revealed AF with controlled heart rate | 720
T4 level dropped | 720
ejection fraction improved | 1008