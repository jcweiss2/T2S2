66 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
diabetes mellitus | -672 | 0 | Factual
obesity | -672 | 0 | Factual
body mass index 25.3 kg/m2 | -672 | 0 | Factual
consumed rice wine | -672 | 0 | Factual
colonoscopy | 0 | 0 | Factual
colonoscopic polypectomy | 0 | 0 | Factual
endoscopic mucosal resection | 0 | 0 | Factual
hot snare | 0 | 0 | Factual
preventive hemoclips | 0 | 0 | Factual
polyps resected | 0 | 0 | Factual
polyps in right colon | 0 | 0 | Factual
polyps in left colon and rectum | 0 | 0 | Factual
discharged from endoscopy room | 0 | 0 | Factual
right abdominal pain | 24 | 24 | Factual
tenderness | 24 | 24 | Factual
rebound tenderness | 24 | 24 | Factual
severe infection | 24 | 24 | Factual
white blood cell count 21460/mm3 | 24 | 24 | Factual
C-reactive protein level 17.8 mg/dL | 24 | 24 | Factual
blood urea nitrogen level 28 mg/dL | 24 | 24 | Factual
creatinine 2.13 mg/dL | 24 | 24 | Factual
lactic acid 2.4 mmol/L | 24 | 24 | Factual
total bilirubin 1.7 mg/dL | 24 | 24 | Factual
abdominopelvic computed tomography | 24 | 24 | Factual
multiple air bubbles in right lateral abdominal muscles | 24 | 24 | Factual
broad-spectrum antibiotic therapy | 24 | 44 | Factual
piperacillin/tazobactam | 24 | 44 | Factual
emergency exploratory laparotomy | 44 | 44 | Factual
laparoscopic right hemicolectomy | 44 | 44 | Factual
multiple-organ failure | 44 | 44 | Factual
metabolic acidosis | 44 | 44 | Factual
diagnosis of necrotizing fasciitis | 48 | 48 | Factual
surgical debridement and drainage | 48 | 48 | Factual
renal replacement therapy | 48 | 860 | Factual
septic shock | 860 | 860 | Factual
multiple-organ failure | 860 | 860 | Factual
death | 860 | 860 | Factual
imipenem-resistant Acinetobacter baumannii | 72 | 72 | Factual
extended spectrum beta-lactamase negative Escherichia coli | 72 | 72 | Factual
no bacterial growth in blood cultures | 24 | 72 | Factual
no bacterial growth in first surgical wound culture | 48 | 48 | Factual
no pneumoperitoneum | 24 | 24 | Factual
no bowel perforation | 24 | 24 | Factual
no peritonitis | 24 | 24 | Factual
no trauma history | -672 | 0 | Factual
no operation history | -672 | 0 | Factual
no acupuncture | -672 | 0 | Factual
no moxibustion | -672 | 0 | Factual