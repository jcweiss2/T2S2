2 years old | 0
female | 0
chromosomal abnormality of 1p36 deletion syndrome | 0
developmental delay | 0
intellectual disability | 0
seizures | 0
vision problems | 0
hearing problems | 0
distinctive facial features | 0
brain anomalies | 0
orofacial clefting | 0
congenital heart disease | 0
cardiomyopathy | 0
renal anomalies | 0
admitted to the hospital | 0
gastroesophageal reflux | 0
pulmonary arterial banding | -672
ventricular septal defect | -672
Ebstein anomaly | -672
lip alveolus and palate cleft | -672
laryngomalacia | -672
hypothyroidism | -672
psychomotor retardation | -672
home oxygen therapy | -672
tube feeding | -672
upper-gastrointestinal series | 48
fever | 48
diarrhea | 48
high-flow nasal cannula | 48
respiratory distress | 48
stabilized respiration | 72
stabilized circulation | 72
resolved diarrhea | 72
persisted fever | 72
higher fever | 384
tachycardia | 384
mild lactate level elevation | 384
mild decrease of SpO2 | 384
elevated blood urea nitrogen | 384
marginal elevation of C-reactive protein level | 48
negative cultures | 48
abdominal distention | 552
hypotensive shock | 552
thrombocytopenia | 552
renal dysfunction | 552
liver dysfunction | 552
coagulation disorder | 552
mixed acidosis | 552
multiple-organ failure | 552
disseminated intravascular coagulation | 552
mechanical ventilation | 552
inotropes | 552
antibiotics | 552
nasogastric tube | 552
Nélaton’s catheter | 552
skin reddening on the lower extremities and lower abdomen | 566
circulatory failure | 566
no urine production | 566
death | 566
autopsy | 589.5
severe abdominal distention | 589.5
extreme skin reddening | 589.5
intestinal dilation due to gas retention | 589.5
no obvious organic disease | 589.5
congestion in the intestinal wall | 589.5
extensive pneumonia | 589.5
systemic inflammation | 384
septic shock | 552
secondary abdominal compartment syndrome | 552