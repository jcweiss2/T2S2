54 years old | 0
female | 0
non-smoking | 0
underlying stage IV lung adenocarcinoma | 0
brain metastasis | 0
liver metastasis | 0
multiple bone metastasis | 0
ECOG score of 0 | 0
chronic cough | -2160
computed tomography (CT)-guided biopsy | -2160
L858R-positive lung adenocarcinoma | -2160
clinical staging of cT4N3M1b | -2160
erlotinib | -2160
disease progression | -720
osimertinib | -1440
T790M | -1440
chemotherapy | -1080
disease progression | -120
re-biopsy | -120
genomic profiling | -120
ACTDrug next-generation sequencing (NGS)-based assay | -120
L858R/cis-T790M/cis-C797S | -120
brigatinib | 0
afatinib | 0
exertional dyspnea | 48
dry cough | 48
rapid progression | 48
hypercapnic respiratory failure | 48
intubation | 48
leukocytosis | 48
neutrophil predominant | 48
carbon dioxide retention | 48
bilateral interstitial infiltrates | 48
pneumonia | 48
broad-spectrum antibiotics | 48
fever subsided | 96
septic shock improved | 96
oxygenation remained poor | 96
bilateral ground-glass opacities | 96
left lower lung consolidation | 96
intravenous methylprednisolone | 96
oxygenation improved | 144
bilateral infiltrates improved | 144
complete resolution of ground-glass opacities | 336
complete resolution of consolidation | 336
seizure | 504
progressive brain metastasis | 504
brain radiotherapy | 504
progressive septic shock | 576
death | 720