43 years old | 0
male | 0
liver cancer | -672
hepatocellular carcinoma | -672
chronic hepatitis B virus infection | -672
allogeneic liver transplantation | 0
admitted to the hospital | 0
Tacrolimus FK506 | 0
Mycophenolate mofetil | 0
prednisone | 0
low peripheral T cell count | 48
low peripheral B cell count | 48
low peripheral NK cell count | 48
P. sputorum bacteremia | 24
elevated serum procalcitonin | 96
elevated C-reactive protein | 96
elevated peripheral neutrophil granulocyte percentage | 96
imipenem | 96
ceftriaxone/tazobactam | 96
infection controlled | 240
low serum procalcitonin | 240
normal peripheral neutrophil granulocyte percentage | 240
P. sputorum identified by mass spectrometry | 96
P. sputorum identified by 16S rRNA sequencing | 96
P. sputorum identified by pulsed-field gel electrophoresis | 96
antibiotic susceptibility tests | 96
resistant to aztreonam | 96
resistant to cefepime | 96
resistant to ceftazidime | 96
resistant to gentamicin | 96
resistant to meropenem | 96
resistant to tobramycin | 96
susceptible to ceftriaxone | 96
susceptible to ciprofloxacin | 96
susceptible to imipenem | 96
susceptible to levofloxacin | 96
susceptible to minocycline | 96
susceptible to piperacillin | 96
susceptible to piperacillin/tazobactam | 96
susceptible to tetracycline | 96
susceptible to ticarcillin/clavulanic acid | 96
susceptible to tigecycline | 96
susceptible to trimethoprim | 96
intermediate to amikacin | 96
discharged | 240