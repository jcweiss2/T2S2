47 years old | 0
woman | 0
diagnosed with schizophrenia | 0
treated with clozapine | 0
poor adherence to prescribed medication regimen | 0
spouse divorced | -8760
mother passed away | -3600
moved in with son | -72
able to communicate with son | -24
drowsy | -24
incoherent | -24
arrived at emergency department | 0
azotemia | 0
blood urea nitrogen 29 mg/dL | 0
creatinine 2.56 mg/dL | 0
muscle enzyme elevation | 0
creatine kinase 70,758 IU/L | 0
lactate dehydrogenase 933 IU/L | 0
gross hematuria | 0
metabolic acidosis | 0
pH 7.28 | 0
PaCO2 33 mmHg | 0
HCO3- 15.5 mmol/L | 0
anuria | 0
rhabdomyolysis | 0
hemodialysis | 0
mechanical ventilation | 0
respiratory distress | 0
pulmonary edema | 0
leukocytosis | 0
white blood cell count 31,940 cells/μL | 0
high acute phase reactant | 0
C-peptide protein 7.04 mg/dL |)0
sustained fever 38.0oC | 0
sepsis | 0
systemic antibiotics administered | 0
admitted to ICU | 0
continuous renal replacement therapy | 0
low blood pressure | 0
inotropic agents | 0
pulmonary edema improved | 0
extubation | 96
drowsiness persisted | 96
generalized tonic-clonic seizure | 96
no abnormalities on brain MRI | 96
electroencephalogram showed no epileptiform discharge | 96
cerebrospinal fluid analysis | 96
elevated protein levels 61 mg/dL | 96
no evidence of infection in cerebrospinal fluid | 96
organisms not isolated from cerebrospinal fluid | 96
antiepileptic drug prescribed | 96
seizure-like movement subsided | 96
antibiotics administered | 96
extended-spectrum beta-lactamase-resistant Escherichia coli induced urosepsis | 96
leukocytosis did not improve | 96
decreased C-reactive protein levels | 96
fever subsided | 96
prescribed clozapine again | 96
leukocytosis became severe | 102
white blood cell count from 24,970 cells/μL to 72,070 cells/μL over 6 days | 102
fever reappeared 37.8oC | 102
no definite evidence of systemic infection | 102
fever responsive to antipyretic drug | 102
primary hematologic disease unlikely | 102
absence of atypical leukocytes | 102
normal range of white blood cells a month before | -720
severe systemic inflammation | 102
suspicion of underlying myeloproliferative disease | 102
short-term systemic steroids administered | 102
no clinical improvement | 102
serum BCR/ABL1 rearrangement test negative | 102
patient attempted suicide by overdosing on clozapine | 102
clinically suspected NMS caused by clozapine overdose | 102
discontinued clozapine administration | 102
leukocytosis resolved to normal range | 168
white blood cell count 72,070 cells/μL on last dose of clozapine | 102
white blood cell count 7,000 cells/μL 7 days after clozapine withheld | 168
continuous renal replacement therapy switched to intermittent hemodialysis | 168
transferred from ICU to general ward | 168
low-dose clozapine resumed | 168
delusional symptoms | 168
CK elevated 63,046 IU/L | 0
CK decreased to 39 IU/L | 168
discharged alive | 168
no persistent organ failure | 168
