45 years old | 0
male | 0
giant inguinoscrotal hernia | -672
refused surgery | -672
loss of strength | -168
progressive increase of hernia | -168
hernia reached the calves | -168
used a small wagon to transport his hernia | -168
ulcer continuously discharging putrid liquid | -168
systemic inflammatory response syndrome | 0
impairment of coagulation | 0
anemia | 0
severe hyponatremia | 0
complete left-sided pleural effusion | 0
intubation | 1
catecholamine therapy | 1
transferred to the intensive care unit | 1
CT scan | 2
dislocation of small and large bowel | 2
dislocation of duodenum and pancreas | 2
intra- and extrahepatic cholestases | 2
congestion of the right kidney | 2
ureter descended into the hernia sac | 2
dilated ureter | 2
stabilization | 5
surgery | 5
exploration of the abdominal cavity | 5
signs of peritonitis | 5
purulent liquid in hernia sac | 5
penis identified intra-abdominally | 5
resection of large bowel | 5
resection of distal parts of ileum | 5
resection of hernia sac | 7
inability to close the fascia | 7
inflammatory situation | 7
abdominal cavity reconstructed using absorbable mesh grafts | 7
lesion of the nervus peroneus | 7
polyneuropathia | 7
mobilization | 10
discharged from the hospital | 840
regained ability to walk | 840
regained ability to care for himself | 840
refused further plastic reconstruction | 840