13 years old | 0
female | 0
admitted to the hospital | 0
fever | -120
productive cough | -120
hemoptysis | -120
diarrhea | -120
respiratory distress | 0
tachycardia | 0
chest indrawing | 0
decrease lung sound on the right side | 0
lymphopenia | 0
elevated C-reactive protein | 0
elevated procalcitonin | 0
elevated lactate dehydrogenase | 0
COVID-19 diagnosis | 0
chest computed tomography scan | 0
nasopharyngeal swab sample | 0
reverse transcription polymerase chain reaction test | 0
BiPAP | 0
intensive care unit | 0
Atazanavir | 0
interferon beta-1a | 0
plasmapheresis | 24
fresh-frozen plasma | 24
oxygen therapy | 0
hydroxychloroquine | 0
Lopinavir/ritonavir | 0
Ceftriaxone/cefotaxime | 0
Vancomycin | 0
Ciprofloxacin | 0
arterial oxygen saturation improvement | 48
tachypnea disappearance | 120
tachycardia disappearance | 120
respiratory distress disappearance | 168
oxygen therapy change to nasal cannula | 216
discharged from hospital | 336
good condition | 336
normal oxygen saturation | 336
no fever | 336
follow-up | 336 
plasmapheresis second time | 48
plasmapheresis third time | 72
plasmapheresis fourth time | 96
interferon beta-1a second dose | 144
interferon beta-1a third dose | 216
chest X-ray | 48
chest X-ray improvement | 48
elevated WBC count | 168
leukocytosis | 168
chest CT scan improvement | 168
transferred from ICU to ward | 192 
supplemental oxygen tapering | 240 
room air | 288