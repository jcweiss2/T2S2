53 years old | 0
male | 0
hypertension | 0
hypercholesterolemia | 0
admitted to the hospital | 0
bicuspid aortic valve | 0
aortic valve replacement | -672
bioprosthetic aortic valve replacement | -672
acute abdominal pain | 0
lower extremity pain | 0
lower extremity weakness | 0
right neck pain | -672
low-grade fevers | -224
sweats | -224
malaise | -224
dysphagia | -224
febrile | 0
bilateral cold lower extremities | 0
absent femoral pulses | 0
large ascending aortic pseudoaneurysm | 0
mass effect on the left atrium | 0
mass effect on the superior vena cava | 0
embolic occlusions of the aorta | 0
embolic occlusions of the renal arteries | 0
embolic occlusions of the superior mesenteric artery | 0
embolic occlusions of the hepatic artery | 0
embolic occlusions of the splenic artery | 0
intravenous vancomycin | 0
intravenous cefepime | 0
emergency laparotomy | 24
surgical thrombectomies | 24
bilateral lower limb fasciotomies | 24
mechanical ventilation | 144
vasopressors | 144
renal replacement therapy | 144
magnetic resonance imaging of the brain | 144
multiple supra and infratentorial acute infarcts | 144
intraparenchymal hemorrhages | 144
subarachnoid hemorrhages | 144
histopathology from the thrombus | 144
pigmented septate fungal hyphae | 144
Fontana-Masson stain | 144
melanin in the fungal cell wall | 144
broad-spectrum antifungal therapy | 144
liposomal amphotericin B | 144
intravenous voriconazole | 144
intravenous micafungin | 144
Karius test | 144
metagenomic next-generation sequencing test | 144
fungal culture of the aortic thrombus | 240
black colonies | 240
brown, narrow-angle branching, septate hyphae | 240
sympodial growth | 240
brown multiseptate conidia | 240
Curvularia species | 240
ascending aorta and hemi-arch replacement graft | 504
biological Bentall aortic root and valve replacement | 504
intraoperative transesophageal echocardiography | 504
large mycotic aneurysm | 504
fungal balls | 504
fungal cultures of the intraoperative tissue | 504
Curvularia alcornii | 504
standardized susceptibility tests | 504
amphotericin B | 504
voriconazole | 504
fluconazole | 504
itraconazole | 504
ketoconazole | 504
right neck swelling | 744
increased pulsatility | 744
CT angiogram of the neck | 744
right external carotid artery pseudoaneurysm | 744
open right external carotid artery ligation | 996
histopathology demonstrated septate hyphae | 996
L-AmB | 1008
micafungin | 1008
voriconazole | 1008
posaconazole | 1008
progressive left leg pain | 1224
numbness | 1224
fever | 1224
CT angiography | 1224
bilateral iliac artery pseudoaneurysms | 1224
thrombus | 1224
abscesses | 1224
bilateral iliac artery coil embolization | 1248
L-AmB and micafungin restarted | 1248
voriconazole changed to posaconazole | 1248
further arterial pseudoaneurysms | 1300
emboli | 1300
persistent fever | 1300
transitioned to comfort care | 1300
died | 1300