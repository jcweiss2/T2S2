generalized weakness | -72
fever | -72
cough | -72
12-kg weight loss | -72
HIV-antibody test positive | -72
sputum AFB smear positive | -72
anti-tuberculosis medications started | -40
fluconazole and trimethoprim/sulfamethoxazole started | -40
generalized weakness continued | 0
fever continued | 0
oral thrush | 0
hepatosplenomegaly | 0
ascites | 0
hemoglobin 10.6g/dL | 0
white blood cell 2,700/µL | 0
platelet 58,000/µL | 0
total bilirubin 2.4mg/dL | 0
AST/ALT 131/48IU/L | 0
ALP 114IU/L | 0
GGT 133 IU/L | 0
costophrenic angle blunting | 0
fluid shifting in the right hemithorax | 0
mild pneumonic infiltration in left lung | 0
anti-retroviral agents started | 0
pancytopenia progressed | 1
hemoglobin 7.4g/dL | 1
white blood cell 1,070/µL | 1
platelet 13,000/µL | 1
rifampin discontinued | 1
zidovudine discontinued | 1
trimethoprim/sulfamethoxazole discontinued | 1
new pulmonary infiltrates | 5
septic shock | 5
empirical antibiotic therapy with piperacillin/tazobactam started | 5
mechanical ventilator support started | 6
Gram stain and ordinary culture from sputum and blood revealed no pathologic organisms | 6
bone marrow aspiration and biopsy performed | 9
death | 10
Histoplasma capsulatum identified | 10
disseminated histoplasmosis confirmed | 10