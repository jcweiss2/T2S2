72 years old | 0
female | 0
admitted to the emergency department | 0
asthma | 0
congestive heart failure | 0
dyspnea |%0
abdominal examination normal | 0
no abdominal distension | 0
costophrenic sinuses obscured | 0
no free air under diaphragm | 0
standing direct abdominal X-ray normal | 0
admitted to intensive care unit | 0
respiratory failure | 0
asthma attack | 0
hypoxemia | 4
hypotension | 4
intubation decision | 4
abdominal distension | 4
accidental esophageal intubation | 4
orotracheal intubation | 4
nasogastric tube insertion | 4
peritonitis signs | 4
hemorrhagic fluid from nasogastric tube | 4
general surgery consultation | 4
excessive abdominal distension | 4
peritonitis symptoms | 4
active hemorrhage | 4
abdominal CT massive free air | 4
emergency laparotomy | 4
gastric perforation 2 cm | 4
active arterial bleeding | 4
perforation repair | 4
Roseo-Graham omental patch | 4
bleeding cessation | 4
no mass or ulcer | 4
surgical drain placement | 4
methylene blue test | 72
drain removal | 72
intensive care unit follow-up | 840
discharged | 840
no acute complications | 840
