68 years old | 0
male | 0
vomited after consuming alcohol | -96
epigastralgia | -96
brought to the hospital by ambulance | -96
blood pressure 160/100 mm Hg | 0
pulse rate 105 beats/min | 0
respiratory rate 32 breaths/min | 0
body temperature 38.3°C | 0
SpO2 95% (by mask at 3 l/min) | 0
white blood cell count 5,900/μl | 0
red blood cell count 411 × 104/μl | 0
hemoglobin 12.3 g/dl | 0
neutrophils 81.7% | 0
platelets 9.7 × 104/μl | 0
total protein 6.1 g/dl | 0
albumin 2.4 g/dl | 0
blood urea nitrogen 34 mg/dl | 0
creatinine 1.2 mg/dl |8
creatine phosphokinase 111 IU/l | 0
aspartate aminotransferase 28 IU/l | 0
alanine aminotransferase <10 IU/l | 0
total bilirubin 0.6 mg/dl | 0
Na 142 mEq/l | 0
Cl 108 mEq/l | 0
K 4.2 mEq/l | 0
C-reactive protein 40.2 mg/dl | 0
procalcitonin 12.5 ng/ml | 0
left pleural effusion | 0
cardiomegaly | 0
heart failure suspected | 0
spontaneous esophageal perforation diagnosed | 48
chest tube drainage performed | 48
increasing pleural effusion | 48
general condition deteriorated | 48
sepsis diagnosed | 48
transferred to our hospital | 96
emergent surgery performed | 96
perforated lesion covered with necrotic tissue | 96
large amounts of food residue within left thoracic cavity | 96
5-cm-long perforation at left side of lower esophagus | 96
pyothorax | 96
mediastinitis | 96
left thoracic cavity rinsed with 10 l of saline | 96
thoracic drainage performed | 96
nasoesophageal tube inserted | 96
transcervical mediastinal tube inserted | 96
feeding jejunostomy performed | 96
postoperative enteral nutrition | 96
blood laboratory data improved | 96
contrast medium seen from perforated esophagus as fistula | 480
contrast medium diminished | 1392
lesion of esophageal perforation covered with regenerated epithelium | 1728
peroral intake started | 1824
discharged from hospital | 2064
