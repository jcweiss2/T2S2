38 years old | 0
Afro-Brazilian | 0
female | 0
admitted to the hospital | 0
sickle cell disease | -672
Hb SS | -672
acute painful vaso-occlusive crises | -672
bone infarcts | -672
skin ulcer of the lower limb | -672
acute chest syndrome | -672
autosplenectomy | -672
jaundice | -336
choluria | -336
dyspnea on light exertion | -336
pain in the right upper abdominal quadrant | -336
pain in the lower limbs | -336
blood pressure of 140 × 90 mm Hg | 0
heart rate of 81 beats per minute | 0
respiratory rate of 18 breaths per minute | 0
temperature of 36.7 °C | 0
oxygen saturation of 96% | 0
respiratory sounds were normal | 0
painful enlarged liver | 0
anemia | 0
Hb: 6.7 g/dL | 0
hematocrit: 21% | 0
cholestasis | 0
total bilirubin: 16.01 mg/dL | 0
direct bilirubin: 12.11 mg/dL | 0
aspartate aminotransferase (AST): 138 U/L | 0
alanine aminotransferase (ALT): 46 U/L | 0
alkaline phosphatase (ALP) 445 U/L | 0
gamma-glutamyl transferase (GGT) 437 mg/dL | 0
albumin levels: 3.4 g/dL | 0
international normalized ratio (INR): 1.37 | 0
serology tests for hepatitis B and C: negative | 0
serology tests for HIV: negative | 0
serology tests for autoimmune conditions: negative | 0
positive immunoglobulin (Ig)G antibodies for cytomegalovirus | 0
positive immunoglobulin (Ig)G antibodies for Epstein–Barr virus | 0
alpha-fetoprotein: normal | 0
ceruloplasmin: normal | 0
iron metabolism markers: slightly altered | 0
iron: 174 μg/dL | 0
transferrin saturation: 68% | 0
total iron binding capacity: 256 μg/dL | 0
ferritin: 575 ng/dL | 0
renal function: preserved | 0
creatinine: 0.53 mg/dL | 0
blood cultures: negative | 0
chest X-ray: no change of the pulmonary parenchyma | 0
Hb S fraction: 74% | -744
intravenous fluids | 0
analgesia | 0
folate | 0
supplementary oxygen therapy | 0
packed red blood cells: 900 mL | 0
hematocrit: 25% | 0
exchange blood transfusion (EBT) | 0
Hb S fraction: 14.3–20.4% | 24
resolution of respiratory distress | 24
resolution of lower limb pain | 24
jaundice persisted | 24
choluria persisted | 24
abdominal pain persisted | 24
acute respiratory distress | 312
fever | 312
hypoxemia | 312
diffuse lung opacities | 312
acute chest syndrome | 312
mechanical ventilation | 312
meropenem therapy | 312
mental confusion | 312
seizure | 312
posterior reversible encephalopathy syndrome (PRES) | 312
normal levels of ammonia | 312
hepatic encephalopathy: ruled out | 312
increasing levels of direct bilirubin | 312
elevated INR | 312
renal function deterioration | 624
creatinine: 3.31 mg/dL | 768
refractory shock | 768
death | 768