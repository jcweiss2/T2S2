71 years old | 0
Taiwanese | 0
male | 0
presented with nocturia | -17520
presented with incomplete voiding | -17520
nocturia occurred intermittently for 2 years | -17520
incomplete voiding occurred intermittently for 2 years | -17520
digital rectal examination | 0
enlarged prostate | 0
no hard nodule | 0
urinalysis negative for pyuria | 0
urinalysis negative for haematuria | 0
prostate-specific antigen level 7.845 ng/ml | 0
TRUS-measured prostate volume 64 ml | 0
biopsy performed | -24
5-alpha reductase inhibitor administered | -24
preparation included mandatory cessation of anticoagulants | -24
preparation included cleansing of the rectum | -24
preparation included antibiotic consumption | -24
levofloxacin 750 mg prescribed | -48
TRUS revealed homogenous echogenicity | 0
TRUS revealed no hypoechoic lesions | 0
twelve core prostatic tissue samples collected | 0
gross haematuria observed after biopsy | 0
Foley catheter placed for drainage | 24
observed for 24 hours | 24
no fever evident | 24
Foley catheter removed | 24
normal voided volume of 150 ml | 24
discharged | 24
resumed normal activities | 24
fever of 38.5°C | 24
backache | 24
severe myalgia in the right thigh | 24
temperature 38.5°C | 24
heart rate 103 beats/minute | 24
respiratory rate 18 counts/minute | 24
blood pressure 107/63 mmHg | 24
DRE revealed a tender prostate | 24
leucocytosis not observed | 24
white blood cell count 9550/μl | 24
neutrophil predominance (94%) | 24
elevated C-reactive protein 23.36 mg/dl | 24
elevated procalcitonin 23.3 ng/ml | 24
pyuria (white blood cells: >100/high power field) | 24
prostatitis with sepsis considered | 24
intravenous ceftriaxone 2 g once daily started | 24
backache persisted after 3 days of treatment | 72
condition worsened | 72
developed shortness of breath | 72
transferred to intensive care unit | 72
plain radiography of lumbar spine performed | 72
computed tomography of abdomen performed | 72
radiographic images revealed narrowing of L3–L5 vertebrae | 72
cystic lesion 3.3 cm over right psoas muscle observed on CT | 72
cystic lesion could not be drained percutaneously | 72
continued antibiotic treatment with ceftriaxone for 2 days | 96
scheduled for MRI of lumbar spine | 96
MRI revealed abscesses in L3/4 and L4/5 intervertebral disc spaces | 96
MRI revealed narrow enhancement of L3–L5 vertebral bodies | 96
MRI revealed abnormally enhanced lesions involving both psoas muscles | 96
spiking fever up to 39°C | 96
chills | 96
Escherichia coli identified in blood culture | 96
Escherichia coli showed multiple drug resistance in urine culture | 96
resistant to cefazolin | 96
resistant to ceftriaxone | 96
resistant to ciprofloxacin | 96
resistant to levofloxacin | 96
susceptible to flomoxef | 96
susceptible to piperacillin–tazobactam | 96
susceptible to cefepime | 96
susceptible to doripenem | 96
susceptible to imipenem | 96
ceftriaxone switched to doripenem 0.25 g three times daily | 120
neurosurgeons performed total laminectomies of L4/L5 vertebrae | 168
removal of epidural abscesses | 168
pathology revealed chronic inflammation of spine | 168
pathology revealed chronic inflammation of epidural tissue | 168
discharged on seventh postoperative day | 168
returned to normal activities | 168
