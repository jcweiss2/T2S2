70 years old | 0
female | 0
admitted to the hospital | 0
acute epigastric pain | -1
diabetes mellitus | -672
cholecystectomy | -672
heterozygote alpha-1 antitrypsin deficiency | -672
epigastric tenderness | 0
no fever | 0
pulse rate of 82 beats/min | 0
blood pressure of 128/68 mmHg | 0
normal respiratory rate | 0
normal oxygen saturation | 0
total bilirubin of 0.28 mg/dL | 1
glutamic oxaloacetic transaminase of 45 U/L | 1
glutamic pyruvic transaminase of 30 U/L | 1
γ-glutamyltransferase of 91 U/L | 1
alkaline phosphatase of 99 U/L | 1
lipase of 3518 U/L | 1
severe septic shock | 2
mechanical ventilation | 2
aggressive hemodynamic support | 2
computed tomography scan | 2
air-filled cavity in the right liver lobe | 2
broad-spectrum intravenous antibiotics | 2
percutaneous radiologically guided drainage | 3
endoscopic retrograde cholangiopancreatography | 4
cholangiogram | 4
clear bile | 4
endoscopic sphincterotomy | 4
Escherichia coli | 5
Streptococcus anginosus | 5
Klebsiella oxytoca | 5
weaned from the ventilator | 168
transferred to the ward | 336
discharged | 720
colonoscopy | 720
transthoracic echocardiogram | 720
magnetic resonance imaging | 1008
positron emission tomography | 1134
surgical drainage | 2160
laparoscopic deroofing | 2160
debridement of the hepatic collection | 2160
partial hepatectomy | 2160
no malignancy | 2160
sterile microbiological cultures | 2160
antibiotics discontinued | 2016
coronavirus disease 2019 infection | 2448