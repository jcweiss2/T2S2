17 years old | 0
male | 0
admitted to the hospital | 0
poorly-controlled persistent asthma | 0
obesity | 0
hypertension | 0
type II diabetes | 0
presented to the emergency department | 0
shortness of breath | 0
febrile | 0
temperature 40.6°C | 0
tachycardic | 0
heart rate 140 beats/minute | 0
tachypneic | 0
respiratory rate 28 breaths/minute | 0
slightly elevated blood pressure | 0
127/74 mmHg | 0
oxygen saturation 98% | 0
weight 122 kg | 0
BMI 50.1 kg/m² | 0
skin tenderness | -96
warmth in the gluteal area | -96
2 pack-year history of smoking | 0
non-adherent with metformin | 0
non-adherent with insulin glargine | 0
dry mucous membranes | 0
diminished breath sounds bilaterally | 0
no wheezing | 0
soft abdomen | 0
no guarding | 0
no tenderness | 0
left scrotum erythematous | 0
left scrotum indurated | 0
left perineum erythematous | 0
left perineum indurated | 0
bilateral buttocks erythematous | 0
bilateral buttocks indurated | 0
no drainage | 0
no fluctuance | 0
no crepitus | 0
sodium 131 mEq/L | 0
potassium 3 mEq/L | 0
chloride 92 mEq/L | 0
phosphate 2.3 mg/dL | 0
glucose 320 mg/dL | 0
CRP 28.6 mg/dL | 0
ultrasound consistent with cellulitis | 0
no abscess formation | 0
electrolyte abnormalities | 0
uncontrolled type II diabetes | 0
perineal cellulitis | 0
started on oral clindamycin | 0
IV fluids | 0
insulin for hyperglycemia | 0
remained febrile | 0
remained tachycardic | 0
worsening hypertension | 0
perineal cellulitis progressed to fluid-filled blisters | 24
blisters ruptured | 24
drained purulent fluid | 24
repeat ultrasound | 24
no changes on repeat ultrasound | 24
antibiotic regimen broadened to cefepime | 24
antibiotic regimen broadened to vancomycin | 24
signs of sepsis | 24
white blood cell count 11 K/uL | 24
35% bands | 24
CRP 46.4 mg/dL | 24
contrast CT scan of pelvis | 24
scrotal wall edema | 24
fluid within scrotum | 24
extensive fat stranding | 24
air in subcutaneous tissue | 24
Fournier’s gangrene diagnosis | 24
no fluid collections | 24
no extension into peritoneum | 24
general surgery consulted | 24
urgent debridement | 24
IV clindamycin added | 24
underwent extensive surgical debridement | 24
necrotic soft tissue of left perineum | 24
necrotic tissue extending to left thigh | 24
necrotic tissue extending to inguinal region | 24
necrotic tissue extending posteriorly | 24
560 cm² necrotic tissue debrided | 24
post-operative septic shock | 24
post-operative diabetic ketoacidosis | 24
transfer to PICU | 24
required vasopressors | 24
required insulin infusion | 24
second debridement | 48
no evidence of ongoing necrotizing infection | 48
VAC performed | 48
wound culture grew Actinomyces species | 48
initial fungal culture no growth | 48
initial anaerobic culture no growth | 48
repeat debridement fungal culture positive for Candida albicans | 48
blood cultures negative | 48
antimicrobial regimen narrowed to piperacillin-tazobactam | 48
antimicrobial regimen narrowed to fluconazole | 48
total 6 surgical debridements | 48
wound VAC changes | 48
diverting colostomy | 48
Foley catheter placement | 48
reconstructive surgeries | 48
split-thickness skin grafts | 48
fasciocutaneous flaps | 48
discharged | 1440
surgical wounds healing well | 1440
cleared for colostomy takedown | 1440
colostomy takedown delayed | 1440
barriers to follow-up | 1440
continued smoking | 1440
discharged on amoxicillin | 1440
no recurrences | 1440
type II diabetes |8
presented to the emergency department |0
shortness of breath |0
febrile |0
temperature 40.6°C |0
tachycardic |0
heart rate 140 beats/minute |0
tachypneic |0
respiratory rate 28 breaths/minute |0
slightly elevated blood pressure |0
127/74 mmHg |0
oxygen saturation 98% |0
weight 122 kg |0
BMI 50.1 kg/m² |0
skin tenderness |-96
warmth in the gluteal area |-96
2 pack-year history of smoking |0
non-adherent with metformin |0
non-adherent with insulin glargine |0
dry mucous membranes |0
diminished breath sounds bilaterally |0
no wheezing |0
soft abdomen |0
no guarding |0
no tenderness |0
left scrotum erythematous |0
left scrotum indurated |0
left perineum erythematous |0
left perineum indurated |0
bilateral buttocks erythematous |0
bilateral buttocks indurated |0
no drainage |0
no fluctuance |0
no crepitus |0
sodium 131 mEq/L |0
potassium 3 mEq/L |0
chloride 92 mEq/L |0
phosphate 2.3 mg/dL |0
glucose 320 mg/dL |0
CRP 28.6 mg/dL |0
ultrasound consistent with cellulitis |0
no abscess formation |0
electrolyte abnormalities |0
uncontrolled type II diabetes |0
perineal cellulitis |0
started on oral clindamycin |0
IV fluids |0
insulin for hyperglycemia |0
remained febrile |0
remained tachycardic |0
worsening hypertension |0
perineal cellulitis progressed to fluid-filled blisters |24
blisters ruptured |24
drained purulent fluid |24
repeat ultrasound |24
no changes on repeat ultrasound |24
antibiotic regimen broadened to cefepime |24
antibiotic regimen broadened to vancomycin |24
signs of sepsis |24
white blood cell count 11 K/uL |24
35% bands |24
CRP 46.4 mg/dL |24
contrast CT scan of pelvis |24
scrotal wall edema |24
fluid within scrotum |24
extensive fat stranding |24
air in subcutaneous tissue |24
Fournier’s gangrene diagnosis |24
no fluid collections |24
no extension into peritoneum |24
general surgery consulted |24
urgent debridement |24
IV clindamycin added |24
underwent extensive surgical debridement |24
necrotic soft tissue of left perineum |24
necrotic tissue extending to left thigh |24
necrotic tissue extending to inguinal region |24
necrotic tissue extending posteriorly |24
560 cm² necrotic tissue debrided |24
post-operative septic shock |24
post-operative diabetic ketoacidosis |24
transfer to PICU |24
required vasopressors |24
required insulin infusion |24
second debridement |48
no evidence of ongoing necrotizing infection |48
VAC performed |48
wound culture grew Actinomyces species |48
initial fungal culture no growth |48
initial anaerobic culture no growth |48
repeat debridement fungal culture positive for Candida albicans |48
blood cultures negative |48
antimicrobial regimen narrowed to piperacillin-tazobactam |48
antimicrobial regimen narrowed to fluconazole |48
total 6 surgical debridements |48
wound VAC changes |48
diverting colostomy |48
Foley catheter placement |48
reconstructive surgeries |48
split-thickness skin grafts |48
fasciocutaneous flaps |48
discharged |1440
surgical wounds healing well |1440
cleared for colostomy takedown |1440
colostomy takedown delayed |1440
barriers to follow-up |1440
continued smoking |1440
discharged on amoxicillin |1440
no recurrences |1440
