18 years old| 0
male | 0
admitted to the hospital | 0
fever | -72
rash | -72
acne |  -672
minocycline |  -672
increased WBC count | 0
eosinophilia| 0
systemic involvement| 0
diffuse erythematous or maculopapular eruption| 0
pruritis | 0
DRESS syndrome | 0
fever persisted | 0
rash persisted | 0
discharged | 24
Separate conjunctive phrases into its component events and assign them the same timestamp (for example, the separation of 'fever and rash' into 2 events: 'fever' and 'rash')  If the event has duration, assign the event time as the start of the time interval. Attempt to use the text span without modifications except 'history of' where applicable. Include all patient events, even if they appear in the discussion; do not omit any events; include termination/discontinuation events; include the pertinent negative findings, like 'no shortness of breath' and 'denies chest pain'.  Show the events and timestamps in rows, each row has two columns: one column for the event, the other column for the timestamp.  The time is a numeric value in hour unit. The two columns are separated by a pipe '|' as a bar-separated file. Skip the title of the table. Reply with the table only. Create a table from the following case:
<|eot_id|><|start_header_id|>user<|end_header_id|>
<|eot_id|><|start_header_id|>assistant<|end_header_id|>
19 years old|0
woman|0
admitted to the department of internal medicine|0
pancreatitis| -2880
portal vein thrombosis| -2880
tumor mass at pancreatic head| -2880
explorative laparotomy| -2880
multiple biopsies of tumor mass| -2880
portal venous stent placement| -2880
chronic pancreatitis| -2880
dismissed| -2880
abdominal pain|0
diffuse large tumor mass at pancreatic head|0
intrahepatic cholestasis|0
extrahepatic cholestasis|0
occlusion of portal vein stent|0
portal-systemic collateralization|0
varices|0
dislocation of portal vein stent|0
perforation into stomach|0
CA19.9 elevation|0
admitted to surgical clinic|0
pancreatic tumor compression of duodenum|0
cholestasis|0
portal hypertension|0
duodenal compression|0
interdisciplinary meeting discussion|0
surgical approach decision|0
explorative laparotomy|0
exposure of portal vein|0
exposure of mesenteric root|0
mesenterico-caval shunt|0
release of portal hypertension|0
mobilization of mesenteric root structures|0
dissection of hepatoduodenal ligament|0
identification of portal vein|0
identification of hepatic artery|0
identification of central bile duct|0
removal of dislocated stent|0
ligation of portal vein|0
partial duodenopancreatectomy|0
resection of distal stomach|0
hepatico-jejunostomy|0
gastro-jejunostomy|0
closure of pancreatic stump|0
postoperative monitoring on ICU|0
uneventful clinical course|0
pathological analysis of pancreatitis|0
acinar atrophy|0
ductal ecstasy|0
inflammatory exudate|0
granulocytic epithelial lesions|0
type-2 autoimmune pancreatitis|0
postoperative symptom resolution|0
good quality of life|0
steroid treatment initiation|0
steroid treatment response|0
decreasing cholestasis|0
no evidence of malignancy|0
no conflict of interest|0
no funding|0
informed consent obtained|0
SCARAE criteria compliance|0
