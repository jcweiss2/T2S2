27 years old | 0
female | 0
gravid 2 para 0 | 0
admitted to the hospital | 0
abdominal pain | 0
fever | 0
body temperature 38.9°C | 0
blood pressure 110/70 mmHg | 0
heart rate 115 beats per minute | 0
splenomegaly | 0
cytopenia | 0
hemoglobin 7.9 g/dL | 0
absolute neutrophil count 0.92 × 10^9/L | 0
platelet count 25 × 10^9/L | 0
elevated alanine aminotransferase | 0
elevated aspartate aminotransferase | 0
lactate dehydrogenase elevated | 0
C-reactive protein elevated | 0
hypofibrinogenemia | 0
serum ferritin elevated | 0
prothrombin time prolonged | 0
fibrinogen degradation product elevated | 0
abdominal ultrasound showed splenic swelling | 0
splenic thickness 9.8 cm | 0
viral serology for human immunodeficiency virus negative | 0
viral serology for cytomegalovirus negative | 0
viral serology for hepatitis B and C virus negative | 0
emergency cesarean section | 24
fetal distress | 24
male infant delivered | 24
Apgar scores 5 to 8 points | 24
respiratory distress syndrome | 24
disseminated intravascular coagulation | 48
transfused with packed red blood cells | 48
transfused with fresh frozen plasma | 48
hemoglobin dropped to 5.7 g/dL | 48
abdominal ultrasound showed swollen spleen | 48
splenic thickness 6.3 cm | 48
explorative laparotomy | 72
ruptured spleen found | 72
splenectomy performed | 72
degrading liver function | 96
acute respiratory distress | 96
sustained kidney injury | 96
transferred to intensive care unit | 96
pulse contour cardiac output monitor | 96
continuous renal replacement therapy | 96
ventilator support | 96
multiple blood products transfused | 96
bone marrow biopsy | 120
focal hemophagocytosis | 120
atypical lymphoid cells | 120
flow cytometry failed to detect PNH clones | 120
myeloid flow immune-type showed abnormal NK cells | 120
serologic tests for Epstein-Barr virus positive | 120
titer of EBV DNA >1.0 × 10^7 | 120
splenic pathology supported splenic rupture | 120
diffuse lymphoid cell infiltration | 120
immunohistochemical examination | 120
diagnosed with invasive NK/T-cell lymphoma | 120
diagnosed with HLH | 120
immunosuppressive therapy with dexamethasone | 120
immunosuppressive therapy with etoposide | 120
immunosuppressive therapy with rituximab | 120
patient's condition continued to deteriorate | 168
patient died on the 18th day postoperation | 432
multiorgan failure | -672 
NK/T-cell lymphoma | -672 
HLH | -672 
fever | -672 
abdominal pain | -672 
splenomegaly | -672 
cytopenia | -672 
elevated liver enzymes | -672 
low platelet count | -672 
low hemoglobin | -672 
elevated serum ferritin | -672 
prolonged prothrombin time | -672 
elevated fibrinogen degradation product | -672 
respiratory distress syndrome | 24 
premature birth | 24 
low birth weight | 24 
Apgar scores 5 to 8 points | 24 
respiratory distress | 24 
disseminated intravascular coagulation | 48 
hemorrhage | 48 
transfusion | 48 
splenectomy | 72 
acute respiratory distress | 96 
sustained kidney injury | 96 
multiorgan failure | 168 
death | 432