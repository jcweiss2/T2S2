46 years old | 0
male | 0
Caribbean-Black | 0
presented to the emergency department | 0
fever | -48
cough | -48
shortness of breath | -48
systolic blood pressure 140 mm Hg | 0
heart rate 142 beats per minute | 0
respiratory rate 28 breaths per minute | 0
oxygen saturation 88% on room air | 0
hypertension | 0
tachycardia | 0
tachypnea | 0
normal jugular venous pulse | 0
scattered bilateral crackles | 0
no peripheral edema | 0
12-lead electrocardiogram revealed typical atrial flutter | 0
2 to 1 atrioventricular block | 0
rate-related ST-T segment changes | 0
chest radiograph no acute cardiopulmonary disease | 0
bedside transthoracic echocardiogram preserved left ventricular ejection fraction | 0
no regional wall motion abnormalities | 0
D-dimer 357 ng/dL | 0
pro-brain natriuretic peptide 413 pg/mL | 0
CK-MB 15 U/L | 0
troponin I 0.12 ng/mL | 0
arterial blood gas mild hypoxia | 0
alveolar-arterial gradient 17 mm Hg | 0
hemoglobin 9.4 g/dL | 0
white blood cell count 13.2 × 10^9/L | 0
platelet count 201 × 10^3/µL | 0
serum sodium 134 mmol/L | 0
serum potassium 2.8 mmol/L | 0
serum bicarbonate 22 mmol/L | 0
serum creatinine 0.5 mg/dL | 0
serum osmolality 283 mOsm/kg | 0
blood urea nitrogen 8 mg/dL | 0
fasting blood sugar 116 mg/dL | 0
alanine aminotransferase 26 IU/L | 0
aspartate aminotransferase 68 IU/L | 0
total bilirubin 2.2 mg/dL | 0
alkaline phosphatase 101 IU/L | 0
albumin-corrected calcium 7.3 mg/dL | 0
magnesium 1.6 mg/dL | 0
phosphorous 2.3 mg/dL | 0
serum cortisol level 18.3 µg/dL | 0
thyroid-stimulating hormone 1.44 mU/L | 0
urine osmolality 534 mOsm/kg | 0
urine sodium < 20 mEq/L | 0
erythrocyte sedimentation rate 68 mm/h | 0
high-sensitivity C-reactive protein 83 mg/dL | 0
creatine kinase 873 U/L | 0
lactate dehydrogenase 1717 U/L | 0
blood cultures negative | 0
urine culture negative | 0
initiated on amiodarone and digoxin bolus | 0
moderate-intensity beta-blockade | 0
admitted for hospitalization | 0
unsuccessful cardioversion with 100 J | 0
transitioned to atrial fibrillation with rapid ventricular response | 0
COVID-19 test positive | 0
transferred to quarantine facility with ICU capabilities | 0
continued amiodarone infusion | 24
continued atenolol | 24
symptoms ameliorated | 48
decreasing oxygen requirements | 48
reverted to normal sinus rhythm | 48
anticoagulation deferred | 48
discharged to home quarantine | 120
low-dose amiodarone | 120
follow-up visit | 120
1-week Holter monitor | 120
anemia | 0
mild rhabdomyolysis | 0
hypokalemia | 0
hypomagnesemia | 0
hypophosphatemia | 0
judicious intravenous crystalloid hydration | 0
