53 years old | 0
African American female | 0
body mass index of 27.2 kg/m2 | 0
coronary artery disease | 0
end-stage renal disease | 0
cervical carcinoma | 0
right atrial thrombus | 0
admitted to the emergency department | 0
bleeding from rectum | 0
self-expanding nasal tampons placed in rectum | -1
2 units of PRBCs transfused | -1
MTP started | 0
2 g of intravenous tranexamic acid administered | 0
taken to the operating room | 1
surgical efforts failed to control bleeding | 1
proctoscopy performed | 2
total colectomy | 2
balloon fashioned with Penrose drain and Foley catheter | 2
thromboelastography results | 3
coagulopathy secondary to fibrinogen and platelet deficiency | 3
continued to receive fresh frozen plasma, cryoprecipitate and platelets | 3
consultation with interventional radiology service | 4
brought to the Surgical Intensive Care Unit | 4
two rapid transfuser devices assembled | 5
wide-bore central venous catheter inserted | 5
MT continued | 5
goal mean arterial pressure of 50-60 mmHg | 5
administration of blood products, norepinephrine, and vasopressin infusion | 5
intermittent boluses of epinephrine | 5
resuscitation guided by vital signs, bedside echocardiography, serial TEG and perfusion biomarkers | 5
>14 L blood loss recorded | 5
fistula between right common iliac and rectum identified | 6
10 mm x 40 mm covered self-expanding intravascular stent placed | 6
bleeding stopped | 6
received 60 units PRBC, 23 units FFP, 20 packs of platelets, 6 units cryoprecipitate, 2 g TXA, 30 L of crystalloid, and 2 L of albumin | 7
serial focused cardiac ultrasound guided resuscitation | 7
hypothermia, serum lactate, and base deficit improved | 11
patient able to follow commands | 11
required minimal ventilatory support | 11
abdomen closed | 48
extubated | 48
transferred to the floor | 48