47 years old | 0
male | 0
admitted to the hospital | 0
increasing weight loss | -336
dyspnoea | 0
chest pain | 0
micro haemoptysis | 0
low-grade fever | 0
fatigue | 0
fever | 0
skin paleness | 0
mild tachycardia | 0
laterocervical lymphadenopathy | 0
sinus tachycardia | 0
right bundle branch block | 0
negative T waves in V1-V4, DIII and aVF | 0
pulmonary infarctions | 0
renal infarctions | 0
splenic infarctions | 0
bilateral pulmonary thromboembolism | 0
hypodense lesion in the right parietal lobe | 0
mobile echogenic mass on the mitral valve | 0
no signs of deep vein thrombosis in the lower limbs | 0
bacterial endocarditis suspected | 0
treated with intravenous broad-spectrum antibiotics | 0
treated with low-molecular-weight heparin (LMWH) | 0
right-sided hemiparesis | 192
severe motor aphasia | 192
multiple lesions in hypersignal on T2-weighted images | 192
embolic infarctions in the left frontotemporal and the right parietal lobes | 192
normal carotid Doppler ultrasound | 192
vegetation with an uneven surface on the atrial surface of the mitral valve | 192
no mitral stenosis or regurgitation | 192
hereditary thrombophilia panel normal | 192
autoimmune panel normal | 192
tumour markers taken | 192
alpha-fetoprotein normal | 192
carcinoembryonic antigen normal | 192
prostate-specific antigen normal | 192
Cyfra 21-1 elevated | 192
normochromic, normocytic anaemia | 336
progressive decrease in haemoglobin | 336
haematocrit values decreased | 336
ulcerated tumour at the gastric angle | 336
gastric adenocarcinoma | 336
parenteral anticoagulant, antiplatelet, antibiotic, gastric antisecretory therapy | 336
red blood cell transfusion | 336
neurological status worsened | 336
tetraparesis with left hemiplegia | 336
new infarction in the right sylvian artery | 336
impaired level of consciousness | 504
respiratory failure | 504
transferred to the intensive care unit | 504
supportive care measures | 504
progressive deterioration in consciousness | 504
increased intracranial pressure | 504
transtentorial brain herniation | 504
death | 672