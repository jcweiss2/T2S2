58 years old | 0
female | 0
admitted to the emergency department | -72
dyspnea | -72
bilateral flank pain | -72
pallor | -72
clamminess | -72
blood pressure 170/120 mmHg | -72
heart rate 120 beats/min | -72
body temperature 38.2°C | -72
respiration rate 30 breaths/min | -72
oxygen saturation 89% | -72
body mass index 25.1 kg/m² | -72
taking phendimetrazine tartrate | -43920
crackles in right lung field | -72
soft abdomen without tenderness | -72
elevated CRP 29.5 mg/dL | -72
elevated ESR 120 mm/hr | -72
leukocytosis 14.82×10³/μL | -72
hemoglobin 9.9 g/dL | -72
mean corpuscular volume 90.7 fL | -72
normal platelet count | -72
elevated blood urea nitrogen 25 mg/dL | -72
elevated creatinine 1.66 mg/dL | -72
elevated aspartate aminotransferase 179 IU/L | -72
elevated alanine aminotransferase 106 IU/L | -72
arterial blood gas acidosis | -72
elevated lactate 20 mmol/L | -72
chest radiography bilateral diffuse infiltrations | -72
chest CT round mass 3.8 cm | -72
abdominal CT round mass 3.8 cm | -72
sepsis of unknown origin | 0
acute respiratory distress syndrome | 0
sedated | 0
intubated | 0
admitted to ICU | 0
started broad-spectrum antibiotics | 0
mechanical ventilation | 0
chest radiography resolution of lung infiltrations | 24
persistent high fever | 0
uncontrolled hypertension | 0
elevated troponin-I 0.841 ng/mL | 0
elevated creatine kinase 5.3 ng/mL | 0
elevated NT-proBNP 35,000 pg/mL | 0
echocardiogram hypokinetic segments | 0
reduced LVEF 38% | 0
referred to endocrinologist | 24
elevated urinary metanephrine 2.12 mg/day | 24
elevated plasma norepinephrine 1,588 pg/mL | 24
elevated plasma normetanephrine 2.27 nmol/L | 24
normal plasma epinephrine 18 pg/mL | 24
normal plasma metanephrine 0.04 nmol/L | 24
elevated plasma IL-6 16.5 pg/mL | 24
18F-FDG PET/CT increased uptake | 24
diagnosed functional paraganglioma | 24
SDHB mutation c.541-3C>R | 24
initiated doxazosin | 24
body temperature normalized 36.5°C | 24
blood pressure controlled | 24
excised retroperitoneal mass | 408
tumor size 4.3×3.5×3.7 cm³ | 408
histological cell-nesting pattern | 408
chromogranin A positive | 408
discontinued doxazosin | 408
improved inflammatory biomarkers | 96
improved cardiac biomarkers | 96
improved renal biomarkers | 96
improved hepatic biomarkers | 96
urinary metanephrine 0.25 mg/day | 96
diagnosed diabetes | 96
replaced phendimetrazine with GLP-1 agonist | 96
follow-up CT no recurrence | 10200
asymptomatic follow-up visits | 10200
chronic phendimetrazine intake | -43920
IL-6 overproduction | 24
SIRS | 24
anemia related to chronic inflammation | 24
leukocytosis | 24
no family history | 0
SDHB mutation-associated paraganglioma | 24
no metastases | 24
surgical resection curative | 408
alpha-blockers effective | 24
doxazosin anti-inflammatory | 24
postoperative complications absent | 408
false-positive catecholamine tests possible | 24
normalized IL-6 after surgery | 96
genetic testing recommended | 24
elevated normetanephrine likely true positive | 24
acetaminophen use | 0
stress affecting catecholamines | 0
pseudohypoxia-related gene cluster | 24
SDHB mutation aggressive | 24
nonmetastatic paraganglioma | 24
noradrenergic phenotype | 24
ILB immunohistochemistry not performed | 24
chronic inflammation anemia | 24
IL-6 inducing SIRS | 24
paraganglioma crisis | 24
fever of unknown origin | -72
elevated inflammatory markers | -72
acute kidney injury suspected | -72
liver injury suspected | -72
mixed metabolic-respiratory acidosis | -72
bilateral lung infiltrations | -72
paroxysmal hypertension | -72
palpitations | -72
tachycardia | -72
paraganglioma incidental finding | 24
noradrenergic PPGL | 24
postoperative recovery | 96
diabetes management | 96
no tumor recurrence | 10200
asymptomatic status | 10200
IL-6 evaluation recommended | 24
