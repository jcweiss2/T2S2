21 years old | 0
male | 0
admitted to the emergency department | 0
recurrent generalized skin lesions | -24
recurrent pruritic skin lesions | -24
polymyalgia | -24
polyarthralgia | -24
absence of fever | -24
standard biological analyses | -72
significant inflammatory syndrome (CRP: 100 mg/L) | -72
hyperleukocytosis (WBC: 13800/mm3) | -72
negativity of rheumatoid factor | -72
negative viral serology | -72
clinical examination in emergency department | 0
neurologically conscious | 0
well-oriented | 0
generalized papular cutaneous lesions | 0
erythematous pharynx | 0
absence of fever (36.8°C) | 0
absence of headache | 0
absence of photophobia | 0
absence of neck stiffness | 0
vital signs: cardiac frequency 92/min | 0
vital signs: blood pressure 10.5/80 mm Hg | 0
vital signs: saturation 100% | 0
normal pulmonary examination | 0
normal cardiac examination | 0
soft abdomen | 0
painless abdomen | 0
chest radiography: no systematic focus | 0
chest radiography: no pleural effusion | 0
blood analysis: leukocytosis 18.36 103/mm3 | 0
blood analysis: polyneutrophilia 88% | 0
blood analysis: CRP 243 mg/L | 0
normal renal function | 0
normal hepatic function | 0
normal coagulation | 0
negative serologies | 0
dermatological opinion requested | 0
skin biopsy performed | 0
blood cultures performed without fever | 0
hospitalized in internal medicine department | 0
blood cultures positive for Gram negative diplococci | 24
PCR identification as N. meningitidis | 24
intravenous ceftriaxone initiated | 24
transferred to intensive care unit | 24
lumbar puncture performed | 24
CSF: slightly turbid | 24
CSF: 284 leukocytes/mm3 | 24
CSF: 88% neutrophils | 24
CSF: 8% lymphocytes | 24
CSF: 4% mono-macrophages | 24
CSF: protein 0.56 mg/dL | 24
CSF: glucose 68 mg/dL | 24
CSF Gram staining negative | 24
CSF culture negative after 72h | 96
CSF PCR positive for N. meningitidis B | 96
regression of skin lesions | 48
decreasing leukocytosis | 48
decreasing CRP | 48
transferred to medical unit | 48
transesophageal ultrasound normal | 48
otolaryngology examination normal | 48
histologic examination of skin biopsy | 0
dermal ectatic lymph vessels | 0
capillaries with perivascular lymphocytic infiltration | 0
neutrophil granulocytes | 0
PAS staining performed | 0
Gram staining performed | 0
no mycelial elements | 0
no bacterial elements | 0
PCR on skin biopsy positive for N. meningitidis | 0
chronic meningococcemia diagnosis | 0
normal classical complement pathway | 0
normal alternate complement pathway | 0
normal mannose-binding lectin | 0
normal properdin | 0
total IgG slightly low (6.5 g/L) | 0
normal IgG subclasses | 0
ceftriaxone treatment continued for 7 days | 24
ciprofloxacin relay continued for 7 days | 168
favorable evolution | 168
absence of fever preceding admission | -672
absence of nasopharyngeal carriage | 0
absence of complement deficiency | 0
absence of immunoglobulin deficiency | 0
