28 years old | 0
male | 0
peptic ulcer disease | -72
burning epigastric pain | -72
abdominal distention | -72
nausea | -72
vomiting | -72
bloody diarrhoea | -72
fevers | -72
admitted to the hospital | 0
blood pressure 90/60 | 0
heart rate 111 | 0
respiratory rate 34 | 0
oxygen saturation 91% | 0
pale | 0
diaphoretic | 0
collapsing in triage | 0
weak pulses | 0
undetectable blood pressure | 0
respiratory rate 40 | 0
saturation 90% on ten litres of oxygen | 0
rigid and distended abdomen | 0
absent bowel sounds | 0
decreased level of consciousness | 0
irregularly irregular, wide complex tachycardia | 0
IV fluids | 0
IV dextrose | 0
Haemoglobin 15.8 g/dl | 0
haematocrit 50.1% | 0
white blood cell count 24 × 103/mm3 | 0
segmented neutrophils 52.6 % | 0
lymphocytes 17.4% | 0
platelets 175 × 103/mm3 | 0
point-of-care echocardiogram | 0
large hyperechoic, semisolid, mobile mass within the left ventricle | 0
abdominal ultrasound | 0
dilated and thickened loops of bowel | 0
absence of peristalsis | 0
pneumatosis intestinalis | 0
mesenteric thromboembolism | 0
bowel ischaemia | 0
surgery consulted | 0.5
operating room mobilised | 0.5
exploratory laparotomy | 1
antibiotics | 1
aggressive IV fluid resuscitation | 1
laparotomy | 1
gangrenous necrosis of nearly the entire small bowel | 1
extension to the cecum and ascending colon | 1
viable proximal jejunum | 1
normal pancreas | 1
absent distal superior mesenteric artery pulse | 1
foul-smelling haemorrhagic fluid evacuated | 1
copious lavage with warmed saline | 1
bowel resection deferred | 1
intensive care unit | 2
broad spectrum antibiotics | 2
vasopressors | 2
overwhelming sepsis | 48
multi-organ failure | 48
cardiopulmonary arrest | 48
expired | 48