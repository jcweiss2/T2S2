62 years old | 0
    male | 0
    HIV positive | 0
    bioprosthetic aortic valve replacement | -43800
    admitted to an external hospital | 0
    sepsis | 0
    blood cultures positive for Staphylococcus aureus | 0
    septic shock | 0
    respiratory insufficiency | 0
    renal failure | 0
    initial CT-scan of the chest and abdomen | 0
    transesophageal echocardiography (TEE) | 0
    no endocarditis | 0
    treatment with broad-spectrum antibiotics | 0
    clinical condition improved | 0
    discharged from ICU | 168
    symptoms of a stroke | 168
    CT detected thromboembolism in the posterior cerebral artery | 168
    subsequent TEE | 168
    vegetation on the right coronary cusp of the aortic valve bioprosthesis | 168
    aortic root abscess | 168
    hemodynamically stable | 168
    semi-elective surgical treatment planned | 168
    neurological symptoms declined | 168
    acute deterioration of hemodynamic conditions | 288
    urgent transfer to our hospital | 288
    admission to intensive care unit | 288
    high dose vasopressor therapy | 288
    transthoracic echocardiography (TTE) | 288
    hyperdynamic biventricular function | 288
    shunting from the aortic root to the right atrium | 288
    contrast enhanced computed tomography | 288
    cardiac surgery performed immediately | 288
    removal of the bioprosthesis | 288
    large periannular abscess opening into the right atrium | 288
    pericardial patch plasty performed to exclude the abscess | 288
    another patch to seal the right atrium interiorly | 288
    new bioprosthesis implanted | 288
    postoperative clinical status improved | 288
    left the ICU nineteen days after surgical treatment | 912
    discharged eight weeks after surgery | 2688
    immunodeficiency | 0
    presence of an intracardiac abscess | 168
    transient cerebral ischemia | 168
    staphylococcal sepsis | 0
    no cerebral hemorrhage | 288
    in-hospital transfer minimized | 288
    three-dimensional (3D) TEE not available | 288
    written consent obtained | 0