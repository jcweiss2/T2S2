24 weeks + 3 days gestation | 0
    female | 0
    HIV negative mother | 0
    birth weight 645 grams | 0
    Apgar score 4 at 1 minute | -60
    Apgar score 8 at 5 minutes | -300
    mechanical ventilation | 0
    central umbilical catheters | 0
    total parenteral nutrition | 0
    empiric antibiotics | 0
    skin sensors | 0
    late-onset sepsis | 216
    Escherichia coli bacteremia | 216
    cefepime | 216
    antimicrobial therapy for 10 days | 216
    removal of adhesive patch | 480
    skin abrasion | 480
    erythema | 480
    induration | 480
    plaque with necrotic center | 480
    ulcer with subcutaneous extension | 528
    progression of necrotic area | 528
    healings | 528
    hydrating dermal wound dressings | 528
    hydrocolloids | 528
    thermic instability | 528
    metabolic acidosis | 528
    hyperglycemia | 528
    hypotension | 528
    cutaneous mucormycosis suspected | 528
    skin biopsy | 528
    empiric antifungal treatment | 528
    liposomal amphotericin B | 528
    serum galactomannan not performed | 528
    1,3 beta-D-glucan not performed | 528
    refractory shock | 564
    renal failure | 564
    no surgical debridement | 564
    death | 600
    fungal culture growth Rhizopus spp | 528
    histopathology broad aseptate hyphae | 528
    MALDI-TOF MS Rhizopus arrhizus | 528
    PCR identification Rhizopus arrhizus | 528
    negative fungal blood cultures | 528
    prematurity | 0
    low birth weight | 0
    parenteral nutrition use | 0
    antibiotic use | 0
    orogastric tubes | 0
    skin trauma | 480
    no autopsy performed | 600
    necrotizing cellulitis | 528
    necrotic eschar | 528
    differential diagnosis | 528
    culture confirmation | 528
    histopathology confirmation | 528
    PCR and mass spectrometry confirmation | 528
    no grant funding | 0
    ethics committee approval | 0
    no competing interests | 0
    