39 years old | 0
    female | 0
    scheduled for carinal resection and reconstruction | 0
    adenoid cystic carcinoma in the carina | 0
    mild dyspnea | 0
    chest computed tomography | 0
    bronchoscopy | 0
    left mainstem bronchus obstruction | 0
    extension to carina and right mainstem bronchus | 0
    RMB internal diameter 11 mm | 0
    RMB length 12 mm | 0
    distal LMB length 20 mm | 0
    no underlying diseases | 0
    normal preoperative examinations | 0
    moderate obstructive pattern in pulmonary function test | 0
    forced expiratory volume in one second 1.88 liter | 0
    forced vital capacity 2.81 liter | 0
    ratio 67% | 0
    general anesthesia induced | 0
    propofol 4 µg/ml | 0
    remifentanil 4 ng/ml | 0
    rocuronium 40 mg | 0
    tracheal intubation with 35-Fr double-lumen tube | 0
    moved to right lateral position | 0
    left bronchi and vasculature dissection | 0
    thoracoscopic surgery under right OLV | 0
    PaO2 462 mmHg on FIO2 1.0 | 0
    right-sided double-lumen tube replaced with single-lumen tube | 0
    bronchial blocker placed into RMB | 0
    changed to left lateral position | 0
    right thoracotomy under left OLV | 0
    peak airway pressure 28 cmH2O | 0
    tidal volume 300 ml | 0
    PaO2 110 mmHg after 20 min left OLV | 0
    LMB resection | 0
    reinforced endotracheal tube inserted into LMB | 0
    airway pressure increased to 35 cmH2O | 0
    SpO2 decreased to 70% | 0
    RMB resection | 0
    additional endotracheal tube inserted into right bronchus | 0
    differential bilateral lung ventilation | 0
    SpO2 restored to 100% after 2 min | 0
    carina removal | 0
    lower trachea resection | 0
    RMB anastomosed with trachea | 0
    no air leak at 20 cmH2O | 0
    LMB not implanted | 0
    left lung removal | 0
    left endobronchial tube removed | 0
    non-dependent right OLV | 0
    low tidal volume 200-250 ml | 0
    airway pressure lower than 20 cmH2O | 0
    SpO2 decreased below 80% | 0
    tube reinserted into LMB | 0
    both lungs ventilated | 0
    two-lung ventilation for 5 min | 0
    right OLV reattempted | 0
    SpO2 decreased below 90% after 3 min | 0
    left pulmonary artery clamped | 0
    approach to left pulmonary artery difficult | 0
    surgeon compressed left pulmonary artery | 0
    right OLV confirmed SpO2 100% | 0
    left pulmonary artery ligated | 0
    left endobronchial tube removed | 0
    right thoracotomy closed under right OLV | 0
    PaO2 360 mmHg after 1 hour ligation | 0
    moved to right lateral position | 0
    left thoracotomy performed | 0
    left pulmonary artery and veins resected | 0
    left pneumonectomy completed | 0
    shifted to supine position | 0
    chin sutured to chest | 0
    tracheal extubation | 0
    transferred to ICU | 0
    discharged on postoperative day 13 | 0
    no complications | 0
    