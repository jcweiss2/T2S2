21 years old | 0
pregnant woman | 0
admitted to Shalkar Medical Center | 0
primigravida | 0
severe preeclampsia | 0
intrauterine fetal death | 0
32 weeks’ gestation | 0
abruptio placentae | 0
cesarean section | 0
placenta totally separated | 0
Couvelaire uterus | 0
atonic postpartum hemorrhage | 0
B-Lynch suture | 0
intravenous carbetocin | 0
tranexamic acid | 0
misoprostol | 0
blood loss 2000 ml | 0
received 6 units fresh frozen plasma | 0
received 4 pints packed red blood cells | 0
magnesium sulfate for 24 hours | 0
transferred to WKU maternal ICU | 24
severe preeclampsia complicated by IUFD | 24
renal failure | 24
anuria | 24
monitored with central venous pressure | 24
fluid chart | 24
laboratory investigation | 24
coagulation profile | 24
liver function tests | 24
renal function tests | 24
anemia | 24
hemoglobin 7.8 gm/dl | 24
generalized edema | 24
blood pressure 160/110 mmHg | 24
thrombocytopenia | 24
normal coagulation profile | 24
normal bilirubin | 24
normal liver function tests | 24
HELLP syndrome excluded | 24
hemolysis excluded | 24
normal peripheral blood film | 24
normal reticulocyte count | 24
elevated total leucocyte count 15000/mm3 | 24
normal CRP | 24
normal pro-calcitonin | 24
maternal sepsis excluded | 24
multidisciplinary team management | 24
nephrologist | 24
neurologist | 24
obstetrician | 24
correction of anemia | 24
correction of thrombocytopenia | 24
blood pressure control | 24
labetalol 200 mg/12 hourly | 24
renal dialysis | 24
human albumin | 24
hypoalbuminemia | 24
laboratory investigations every 3 days | 24
two attacks of tonic colonic convulsions | 120
first convulsion lasted 3 minutes | 120
second convulsion lasted 5 minutes | 132
comatose | 132
Glasgow coma scale 11-12 | 132
brain CT showed right partial lobe ICH | 132
ICH volume 1.35 cm3 | 132
carbamazepine 100 mg 12 hourly | 132
thrombocytopenia added to diagnosis | 132
anemia added to diagnosis | 132
ICH added to diagnosis | 132
postpartum eclampsia added to diagnosis | 132
transient renal failure | 132
acute tubular necrosis | 132
five sessions of dialysis | 132
urine output normal | 240
normal renal function tests | 240
ICH size decreased | 384
ICH resolved | 384
discharged from hospital | 480
good general condition | 480
