diagnosed to have tropical chronic pancreatitis | -120
maintained on oral pancreatic enzyme therapy | -120
developed non-insulin-dependent diabetes mellitus | -36
prescribed glucotrol | -36
presented to Saint Peter's University Hospital | 0
complaining of a steady midepigastric pain | 0
CT scan performed | 0
admitted for management of pain secondary to chronic pancreatitis | 0
presented to a medical center in India | -72
CT scan of the abdomen | -72
ERCP performed | -72
medically managed and discharged | -72
developed fever | 48
developed chills and rigors | 48
rapidly progressed to severe sepsis and septic shock | 48
transferred to the medical intensive care unit | 48
intubated for hypoxemic respiratory failure | 48
administration of broad-spectrum antibiotics | 48
vasopressor support | 48
activated recombinant human protein C | 48
ultrasound of the abdomen | 48
bedside emergency ERCP performed | 72
major papilla of Vater visualized spontaneously expelling frank pus | 72
probed with the cannula tip | 72
evacuation of more than 5 ml of yellow pus | 72
cholangiogram obtained | 72
pancreatogram showed marked dilatation of the main pancreatic duct | 72
guide wire introduced into the pancreatic duct | 72
evacuation of approximately 20 ml of pus | 72
5-cm-long 5 F stent placed into the pancreatic duct | 72
reevaluation of the pancreas with a contrast enhanced CT scan | 96
showed inflammatory changes within the fat surrounding the body and tail of the pancreas | 96
dilatation of the pancreatic duct had diminished | 96
calculus showing distal migration towards the sphincter of Oddi | 96
no evidence of pancreatic necrosis or fluid collection | 96
bilateral moderate pleural effusions present | 96
dramatic signs of clinical improvement | 120
stabilization of his hemodynamic parameters | 120
blood cultures grew Klebsiella ornithinolytica | 120
extubated | 120
transferred from the intensive care unit | 120
completed his antibiotic course | 168
discharged home | 168
follow-up examinations at 1 month | 720
follow-up examinations at 3 months | 2160
no further complications | 720
no further complications | 2160