50 years old | 0
female | 0
admitted to the hospital | 0
diagnosed with CML | -252
treatment with imatinib | -252
progressive disease | -168
myeloid blastic transformation | -168
7+3 induction chemotherapy | -168
intubated for severe pneumonia | -168
sepsis | -168
stay in the ICU | -168
bone marrow biopsy | -84
complete remission of the leukaemia | -84
febrile | 0
peripheral and central venous port blood cultures | 0
KP grew | 0
venous port infection | 0
tigecycline treatment | 0
meropenem treatment | 0
treatment discontinued | 14
new onset fever | 19
blood cultures revealed KP | 19
tigecycline and imipenem administered | 19
fever resolved | 24
acute-phase parameters returned to normal | 24
treatment discontinued | 33
fever developed | 35
repeated blood cultures grew pan-resistant KP | 35
rectal swabs collected | 35
rectal swabs were negative | 35
transthoracic echocardiogram performed | 35
enlarged right cardiac chambers | 35
moderate tricuspid valve insufficiency | 35
mass on the tricuspid valve | 35
septic vegetation | 35
diagnosis of tricuspid valve endocarditis | 35
imipenem-cilastatin treatment | 35
gentamicin treatment | 35
sulbactam treatment | 35
tricuspid valve repair | 42
nilotinib treatment | 42
PCR for Bcr/Abl remained positive | 42
unmanipulated peripheral blood allo-SCT | 84
full-matched sibling donor | 84
reduced intensity conditioning regimen | 84
fludarabine treatment | 84
busulfan treatment | 84
cyclosporin A treatment | 84
short-course methotrexate treatment | 84
antithymocyte globulin treatment | 84
neutrophil engraftment | 99
thrombocyte engraftment | 98
complete remission | 168
complete chimerism | 168
no evidence of GVHD | 168
PCR of Bcr/Abl negative | 168
discharged | 168