61 years old | 0
Hispanic | 0
male | 0
admitted to the intensive care unit | 0
syncopal episode | 0
agitation | -840
aggressive behavior | -840
undifferentiated schizophrenia | -840
levothyroxine | -840
hypothyroidism | -840
seizure disorder | -840
divalproex sodium extended release | -840
levetiracetam | -840
glaucoma | -840
dorzolamide/timolol eye drops | -840
clozapine | -840
regular diet | -840
plenty of fluids | -840
fibers | -840
no surgical history | -840
temperature 98°F | 0
blood pressure 86/54 mmHg | 0
pulse 127 beats/min | 0
respiratory rate 16 breaths/min | 0
oxygen saturation 100% | 0
intravenous access | 0
normal saline 500 mL bolus | 0
responsive | 0
confused | 0
agitated | 0
unable to provide any history | 0
abdominal distension | 0
hypoactive bowel sounds | 0
hard impacted stool | 0
stool qualitative guaiac test negative | 0
leukocyte count 17,300/mm3 | 0
neutrophil differential 52% | 0
absolute neutrophil count 9,000/mm3 | 0
band neutrophils 12% | 0
leukocyte count 7,100/mm3 | -168
neutrophil differential 45% | -168
absolute neutrophil count 3,195/mm3 | -168
leukocyte count 6,600/mm3 | -336
neutrophil differential 61% | -336
absolute neutrophil count 4,026/mm3 | -336
leukocyte count 5,400/mm3 | -504
neutrophil differential 65% | -504
absolute neutrophil count 3,510/mm3 | -504
leukocyte count 5,200/mm3 | -672
neutrophil differential 60% | -672
absolute neutrophil count 3,120/mm3 | -672
leukocyte count 6,500/mm3 | -840
neutrophil differential 67% | -840
absolute neutrophil count 4,355/mm3 | -840
hemoglobin 18.6 g/dL | 0
elevated blood urea nitrogen/creatinine | 0
low serum bicarbonate | 0
low serum chloride | 0
elevated anion gap | 0
elevated serum lactic acid | 0
sinus tachycardia | 0
no acute ST-T segment changes | 0
normal serum troponin I | 0
high specific gravity | 0
no bacteria | 0
no elevated nitrate | 0
negative urine toxicology | 0
elevated hemidiaphragm | 0
low lung volumes | 0
clear lung fields | 0
large amount of fecal content | 0
dilated small bowel | 0
bowel obstruction | 0
broad spectrum antibiotics | 0
intravenous fluids | 0
worsening hypotension | 12
cardiac arrest | 12
expired | 12
blood culture revealed Escherichia coli | 24
urine culture revealed no growth | 24
no prior history of constipation | -840
no prior history of fecal impaction | -840
no other risk factors for constipation | -840
minimally communicative | -840
mumbling incoherent words | -840
disorganized | -840
aggressive | -840
denied having any pain | 0
denied having any discomfort | 0
constipation | -840
intestinal obstruction | -840
bowel necrosis | 12
fatal sepsis | 12