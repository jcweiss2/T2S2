46 years old | 0 | 0 
male | 0 | 0 
admitted to the hospital | 0 | 0 
arterial hypertension | -10080 | 0 
obesity | -10080 | 0 
fever | -336 | 0 
hypotension | -336 | 0 
asthenia | -336 | 0 
cardiological examination | -672 | -336 
electrocardiogram (ECG) | -672 | -336 
transthoracic echocardiography (TTE) | -672 | -336 
COVID-19 infection | -336 | -168 
rhinitis | -336 | -168 
mild cough | -336 | -168 
alert | 0 | 0 
oriented | 0 | 0 
cooperative | 0 | 0 
asthenic | 0 | 0 
blood pressure (BP) 85/55 mmHg | 0 | 0 
heart rate (HR) 120 bpm | 0 | 0 
arterial oxygen saturation 85% | 0 | 0 
fever 38.3 C° | 0 | 0 
femoral central venous catheter (CVC) | 0 | 0 
sinus tachycardia | 0 | 0 
diffuse low voltages | 0 | 0 
absence of significant repolarization abnormalities | 0 | 0 
neutrophilic leukocytosis | 0 | 0 
C-reactive protein (CRP) elevation | 0 | 0 
Procalcitonin elevation | 0 | 0 
elevated high sensitivity Troponin (hs-Tn) | 0 | 0 
elevated brain natriuretic peptide (BNP) | 0 | 0 
elevated creatinine | 0 | 0 
transaminases and total bilirubin elevation | 0 | 0 
reverse transcription-polymerase chain reaction (RT-PCR) nasopharyngeal swab for COVID-19 negative | 0 | 0 
COVID-19 IgM antibody test positive | 0 | 0 
normal left ventricular (LV) cavitary dimensions | 0 | 0 
diffuse LV parietal thickening | 0 | 0 
increased myocardial echogenicity | 0 | 0 
severely reduced LV global systolic function | 0 | 0 
low output | 0 | 0 
Grade II LV diastolic dysfunction | 0 | 0 
normal cavitary dimensions | 0 | 0 
reduced global right ventricular (RV) systolic function | 0 | 0 
dilated inferior vena cava (IVC) | 0 | 0 
right ventricular systolic pressure (RVSP) 41 mmHg | 0 | 0 
absence of hemodynamically significant valvulopathy | 0 | 0 
pericardial effusion | 0 | 0 
blood cultures | 0 | 24 
broad-spectrum antibiotic therapy | 0 | 24 
INN-daptomycin | 0 | 24 
piperacillin/tazobactam | 0 | 24 
crystalloid hydration | 0 | 24 
nasal cannula ventilatory therapy | 0 | 24 
norepinephrine | 0 | 12 
poor hemodynamic response | 0 | 12 
levosimendan therapy | 12 | 24 
bolus administration | 12 | 12 
continuous maintenance intravenous infusion | 12 | 24 
BP 100/60 mmHg | 12 | 12 
HR 110 bpm | 12 | 12 
further hemodynamic improvement | 24 | 24 
BP 125/70 mmHg | 24 | 24 
HR 95 bpm | 24 | 24 
diuresis 1800 ml | 12 | 24 
control TTE | 12 | 24 
improvement of systolic performance indices | 12 | 24 
LV EF 66% | 24 | 24 
dP/dT ratio 1275 mmHg/sec | 24 | 24 
TAPSE 23 mm | 24 | 24 
tricuspid S-wave velocity at TDI 11.2 cm/sec | 24 | 24 
SVi 27 ml/m2 | 24 | 24 
CI 2.5 l/min/m2 | 24 | 24 
LV diastolic function improvement | 24 | 24 
IVC diameter 18 mm | 24 | 24 
IVC collapse 100% | 24 | 24 
RVSP 28 mmHg | 24 | 24 
cardiac magnetic resonance imaging (CMR) | 24 | 24 
normal LV and RV volumes | 24 | 24 
normal systolic function | 24 | 24 
mild hypokinesia | 24 | 24 
edema | 24 | 24 
endomyocardial biopsy | 48 | 48 
lymphocytic myocarditis | 48 | 48 
coronary arteriography | 48 | 48 
normal coronary circulation | 48 | 48 
discharged | 504 | 504 
excellent hemodynamic compensation | 504 | 504 
normal laboratory | 504 | 504 
normal electrocardiographic | 504 | 504 
normal echocardiographic findings | 504 | 504 
TTE 1 month after discharge | 744 | 744 
TTE 3 months after discharge | 2232 | 2232 
normal findings | 744 | 2232