26 years old | 0
male | 0
admitted to the emergency room | 0
gastrointestinal obstructive symptoms | -24
aspiration pneumonia | -24
septic shock | -24
chronic pancreatitis | -6720
alcoholism | -6720
Type 1 diabetes mellitus | -6720
schizophrenia | -6720
epilepsy | -6720
severely malnourished | 0
body mass index (BMI) of 15.7 kg/m2 | 0
abdomen was softly distended and tympanic but non-tender | 0
diminished breath sounds at the lower base of the right lung | 0
refractory shock | 0
vasopressors | 0
broad-spectrum antibiotics | 0
nasogastric tube | 0
output of approximately 1.8 L of bilious content | 0
hemodynamic stabilization | 12
computed tomography (CT) scan of the abdomen | 12
distended stomach and first and second portion of duodenum | 12
narrow aortomesenteric angle of 14.3° | 12
extrinsic compression of third portion of the duodenum by the SMA | 12
SMA syndrome | 12
extrinsic compression of the left renal vein | 12
Nutcracker phenomenon | 12
Candida esophagitis | 24
antibiotic treatment | 24
post-obstruction Dobhoff tube | 24
improved | 48
discharged | 168
enteric nutrition | 168
oral antibiotics | 168
denied any history of hematuria | 0
denied decreased urine output | 0
denied flank or low back pain | 0
achieved a BMI of 18 kg/m2 | 1440
resolution of gastrointestinal obstructive symptoms | 1440
no recurrence of abdominal pain | 1440
denied any hematuria | 1440
denied oliguria | 1440
denied flank or low back pain | 1440