27 years old | 0
female | 0
acute myeloblastic leukemia | -1552
myelodysplastic syndrome | -1552
normal karyotype | -1552
WT1+ | -1552
CEBPa mutation | -1552
no NMP1 mutation | -1552
induction chemotherapy | -1552
complete response | -1552
high-dose Ara-C | -1552
pegfilgrastim | -1552
relapse | -728
Ara-C | -728
idarubicine | -728
second complete response | -728
haplo-identical allogeneic HSCT | 0
fludarabine | -14
cyclophosphamide | -14
busulfan | -14
antithymocyte globulin | -14
cyclophosphamide post graft infusion | -14
tacrolimus | -14
mycophenolate mofetil | -14
GvHD prophylaxis | -14
peripheral blood stem cells | -14
CMV+ | -14
HSV+ | -14
HHV6+ | -14
TOXO+ | -14
EBV+ | -14
VZV+ | -14
sinusoidal occlusive syndrome | 0
diuretics | 0
ursodeoxycholic acid | 0
schizocytes | 21
tacrolimus stopped | 21
MMF continued | 21
hematological recuperation | 18
chimerism 100% donor | 18
discharged | 27
EBV PCR | 0
HHV6 PCR | 0
Toxoplasmosis PCR | 0
CMV PCR | 0
ADV PCR | 0
monthly serum immunoglobulin | 0
CMV reactivation | 56
valgancyclovir | 56
valgancyclovir stopped | 112
donor lymphocytes | 134
fever | 157
nausea | 157
vomiting | 157
loss of weight | 157
loss of appetite | 157
severe oral candidiasis | 157
Hg: 9.1 g/dL | 157
WC: 2.7 × 10e3/mm3 | 157
Plat: 56 × 10e3/mm3 | 157
CRP: 86 mg/L | 157
Na: 135 mmol/L | 157
K: 3.0 mmol/L | 157
Protein: 67 g/L | 157
creatinine: 1.06 mg/dL | 157
T Bili: 0.2 mg/dL | 157
D Bili <0.1 mg/dL | 157
AST: 228 U/L | 157
ALT: 136 U/L | 157
ALP: 105 U/L | 157
gamma GT: 75 U/L | 157
posaconazole stopped | 157
ursodeoxycholic acid reintroduced | 157
Ceftazidim | 157
Caspofungin | 157
gastric fibroscopy | 157
biopsies | 157
diarrhea | 159
bacteriological stool analyses | 159
viral stool analyses | 159
fungal stool analyses | 159
Ceftazidim replaced by Tazocillin and Metronidazole | 159
MMF discontinued | 159
steroids started | 159
Foscavir | 159
CMV PCR | 159
GvHD excluded | 159
oral candidiasis confirmed | 159
Chest CT | 159
abdominal CT | 159
pelvic CT | 159
liver biopsy scheduled | 159
sepsis with Staphylococcus hominis | 148
vancomycin | 148
port pulled | 148
diarrhea stopped | 148
steroids decreased | 148
rash | 154
profuse diarrhea | 154
biopsies of gut and skin | 154
steroids increased | 154
hepatomegaly | 157
pain | 157
ascitis | 157
edema | 157
fever | 157
pancytopenia | 158
severe hepatic cytolysis | 158
cholestasis | 158
CMV PCR | 158
EBV PCR | 158
HHV6 PCR | 158
toxoplasmosis PCR | 158
adenovirus PCR | 158
HBV PCR | 158
HCV PCR | 158
BM aspiration | 158
haemophagocytosis excluded | 158
myelotoxicity | 158
liver biopsy | 159
disseminated intravascular coagulation | 159
bleeding in jugular vein | 159
death | 161
hepatic failure | 161
ADV PCR positive | 168
GvHD excluded | 168
viral infection excluded | 168
chimerism 100% donor | 168