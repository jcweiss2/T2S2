6 years old | 0
male | 0
admitted to pediatric emergency department | 0
sudden onset abdominal pain | -1
diffuse abdominal pain | -1
vomited clear fluid | -1
vital sign stable | 0
dehydrated tongue | 0
diffuse abdominal tenderness | 0
elevated white blood cell count | 0
plain abdominal radiograph showed nonspecific small bowel gas | 0
abdominal ultrasound revealed diffuse small bowel wall thickening with ascites | 0
discharged against medical advice | 0
altered mentality | 15
did not respond to painful stimuli | 15
dilated pupils | 15
severe abdominal distension | 15
uncheckable blood pressure | 15
weakly palpable femoral pulse | 15
percutaneous oxygen saturation 77% | 15
blood sugar level 22 mg/dL | 15
pretibial intraosseous cannulation | 15
fluid and medications infused | 15
shock state | 15
arterial blood gas analysis showed pH 7.15 | 15
bicarbonate 7.7 mM | 15
hemoglobin 10.1 g/dL | 15
hematocrit 27.7% | 15
hemoglobin decreased to 4.7 g/dL | 16
hematocrit decreased to 13% | 16
disseminated intravascular coagulopathy | 15
antithrombin III 38.9% | 15
D-dimer 9.18 mg/L | 15
prothrombin time 1.61 international normalized ratio | 15
activated partial thromboplastin time 43.9 seconds | 15
lactic acid 10.9 mmol/L | 15
central venous catheter placed | 15
massive fluid, transfusions, and inotropics delivered | 15
contrast-enhanced abdominal CT scan | 15
large amount of ascites | 15
bowel wall thickening with poor or absent enhancement | 15
serrated beak sign | 15
whirl sign | 15
closed loop obstruction | 15
surgical exploration | 15
congenital transmesenteric hernia | 15
strangulated small bowel | 15
resection of gangrenous small bowel | 15
anastomosis of proximal jejunum and terminal ileum | 15
treatment at pediatric intensive care unit | 15
improved enough to move to general ward | 19
started soft diet | 20
hypertension after renal ischemic injury | 20
short bowel syndrome | 20
cognitive function normal | 20
gradually improving conditions | 20