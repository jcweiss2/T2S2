54 years old | 0
male | 0
admitted to the hospital | 0
acutely discharging sinus | 0
abscess to his right proximal tibia | 0
complex orthopaedic history | 0
infected non-union from an elective right tibial osteotomy | 0
well-controlled asthma | 0
obstructive sleep apnoea | 0
hypertension | 0
deep vein thrombosis | 0
pericarditis | 0
swinging fever | 0
Staphylococcus aureus bacteraemia | 0
flucloxacillin | 0
echocardiogram | 0
non-union of the proximal tibia | 0
sequestrum | 0
CT scan | 0
right tibial exploration and debridement | 0
tissue sampling | 0
CERAMENT G | 0
spanning external fixator | 0
methicillin-sensitive S. aureus | 0
Proteus mirabilis | 0
Enterobacter | 0
oral rifampicin | 0
transthoracic echo | 0
echogenic mobile structure behind the mitral valve leaflet | 0
endocarditis vegetation | 0
flucloxacillin increased | 0
significant pain | 0
acute kidney injury stage III | 0
hypovolaemia | 0
intravenous fluid administration | 0
fever resolved | 0
pregabalin | -120
tapentadol | -120
amitriptyline | -120
sertraline | -120
ketamine | -120
deterioration | 0
hyperthermia | 0
tachycardia | 0
tachypnoea | 0
tremor | 0
hyperreflexia | 0
agitation | 0
bilateral inducible ankle clonus | 0
serotonin syndrome | 0
all serotoninergic medications suspended | 0
critical care involvement | 0
admitted to the critical care unit | 0
blood cultures | 0
P. mirabilis | 0
meropenem | 0
flucloxacillin increased | 0
creatine kinase rose | 24
MRI of the right thigh | 24
myositis ruled out | 24
vital and neurological signs settled | 72
CK dropped | 120
stepped down to the ward | 120
transoesophageal echo | 120
infective endocarditis ruled out | 120
discharged | 336
C-reactive protein | 0
white cell count | 0
neutrophils | 0
lymphocytes | 0
creatinine | 0
alkaline phosphatase | 0
sepsis | 0
infective endocarditis | 0
neuroleptic malignant syndrome | 0
malignant hyperthermia | 0
antibiotics | 336
orthopaedic procedure | 1008
circular fixator | 1008
pin site infections | 1008
pain | 1008
deep vein thrombosis | 1008
walking | 1008
weight bearing | 1008
crutches | 1008
listed for removal of the external fixator | 1008
application of a cast | 1008