66 years old | 0
male | 0
Type II diabetes mellitus | 0
hypertension | 0
hyperlipidemia | 0
acute shortness of breath | -24
cough | -24
fever | -24
recent travel history to Batam, Indonesia | 0
temperature 38.0°C | 0
blood pressure 130/70 mmHg | 0
pulse 140 bpm | 0
respiratory rate 25 per minute | 0
oxygen saturation 92% | 0
placed on 40% Venturi mask | 0
bilateral crepitations | 0
back carbuncle 20 × 20 cm | 0
white blood cell count 31000/µl | 0
hemoglobin level 11.5 g/dl | 0
lactate level 5.92 mmol/L | 0
pro-brain natriuretic peptide level 731 pg/ml | 0
arterial blood gas pH 7.42 | 0
pCO2 35.1 mmHg | 0
pO2 91.9 mmHg | 0
PaO2/FiO2 ratio 230 | 0
chest X-ray bilateral diffuse pulmonary infiltrates | 0
saucerization of the carbuncle | 0
sepsis control | 0
surgery | 0
acute septic | 0
COVID-19 swab test | 0
team huddle | 0
patient transported on plastic-covered trolley | 0
supplemental oxygen via face mask | 0
signage posted | 0
security personnel deployed | 0
plastic cover removed and discarded | 0
airway trolley placed | 0
C-Mac video laryngoscope with disposable blade | 0
drugs and equipment assembled | 0
hand cleansing | 0
glove changing | 0
preoxygenation of 8 vital capacity over 1 minute | 0
FiO2 0.80 | 0
modified rapid sequence induction | 0
propofol 2–3 mg/kg | 0
succinylcholine 1–2 mg/kg | 0
fentanyl 1–2 µg/kg | 0
mask ventilation avoided | 0
muscle paralysis achieved | 0
intubation | 0
desflurane | 0
mechanical ventilation tidal volume 7 ml/kg | 0
normal lung compliance | 0
normal oxygenation | 0
respiratory distress | 0
intubated | 0
tested negative for COVID-19 | 0
patient kept intubated postoperatively | 0
terminal cleaning of OT | 0
OT ventilated for at least one hour | 0
