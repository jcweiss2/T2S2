20 years old | 0
    female | 0
    lactational breast abscess | 0
    pain | -240
    erythema | -240
    edema | -240
    delivered a baby | -792
    pure breastfeeding | -792
    fever | -240
    highest temperature of 38.3 °C | -240
    white blood cell count 14.57 × 109/L | -240
    neutrophil proportion 83.8% | -240
    CRP 13.76 mg/L | -240
    ultrasound showed heterogeneous hypo-echo | -240
    body temperature returned to normal | -240
    antibiotic therapy with Amoxicillin Potassium Clavulanate | -240
    antibiotic therapy with Metronidazole | -240
    symptoms remained poorly controlled | -240
    termination of breastfeeding | 0
    admitted to the hospital | 0
    temperature 36.4 °C | 0
    heart rate 105 beats/min | 0
    respiratory rate 20 breaths/min | 0
    blood pressure 105/69 mmHg | 0
    painful mass 8 cm × 6 cm | 0
    fluctuant skin | 0
    ultrasonography showed anechoic mass with internal heterogeneous hypo-echo | 0
    white blood cell count 15.43 × 109/L | 0
    neutrophil proportion 85.3% | 0
    CRP 11 mg/L | 0
    normal liver function | 0
    normal renal function | 0
    normal coagulation function | 0
    ultrasound-guided needle aspiration failed | 0
    milk agglutination | 0
    necrotic tissue within breast abscess | 0
    milk sent for bacteria test | 0
    pus sent for bacteria test | 0
    Amoxicillin Potassium Clavulanate ineffective | 0
    Metronidazole ineffective | 0
    Cefmetazole administrated | 0
    body temperature rose to 38.6 °C | 0
    surgically removed 150 mL of pus | 0
    surgically removed necrotic tissue | 0
    placed 16G indwelling needle for irrigation | 0
    placed catheter for drainage | 0
    general anesthesia | 0
    body temperature rose to 41.2 °C | 0
    white blood cell count 23 × 109/L | 0
    neutrophil proportion 96.6% | 0
    CRP 138 mg/L | 0
    antibiotic changed to Levofloxacin | 0
    heart rate 150 beats/min | 0
    blood pressure 75/40 mmHg | 0
    septic shock | 0
    norepinephrine initiated at 1 mg/kg/min | 0
    transferred to ICU | 0
    white blood cell count 40.56 × 109/L | 0
    neutrophil proportion 97.4% | 0
    CRP 186 mg/L | 0
    PCT 4.99 | 0
    lactic acid 3.98 mmol/L | 0
    alkaline phosphatase 164.5 U/L | 0
    aspartate aminotransferase 38.7 U/L | 0
    alanine aminotransferase 46.3 U/L | 0
    albumin 23.7 g/L | 0
    total bilirubin 24.1 μmol/L | 0
    activated partial thromboplastin time 55.8 s | 0
    prothrombin time 24.3 s | 0
    INR 2.08 | 0
    cultures of blood negative for microbial agents | 0
    cultures of stool negative for microbial agents | 0
    cultures of urine negative for microbial agents | 0
    chest X-ray negative | 0
    COVID-19 negative | 0
    arterial blood gas pH 7.421 | 0
    lactic acid 3.98 mmol/L | 0
    intensive care | 0
    placement of central venous catheter | 0
    fluid resuscitation | 0
    norepinephrine to maintain blood pressure | 0
    transfusion of plasma | 0
    continuous irrigation of breast abscess | 0
    drainage of breast abscess | 0
    local erythema improved | 24
    edema improved | 24
    culture showed Staphylococcal aureus | 0
    culture showed MRSA | 0
    vancomycin prescribed | 24
    vitals stable | 168
    transferred to department | 168
    erythema disappeared | 168
    edema disappeared | 168
    pain disappeared | 168
    pus disappeared | 168
    drainage extubated | 168
    fluid culture no bacteria | 168
    cured | 240
    discharged | 240
    asymptomatic during follow-up | 240
    asymptomatic at one week follow-up | 336
    asymptomatic at two week follow-up | 480
    asymptomatic at one month follow-up | 672
    <|eot_id|>