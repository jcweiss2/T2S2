35 years old | 0
female | 0
helmeted female bicyclist | 0
no past medical or surgical history | 0
brought in by emergency medical services | 0
level 1 trauma code | 0
struck by a motor vehicle | -1
loss of consciousness | -1
Glasgow Coma Scale (GCS) was 15 | 0
severe respiratory distress | 0
shortness of breath | 0
pulse rate of 125 beats per minute | 0
BP 67/20 | 0
respiratory rate of 45 breaths per minute | 0
ecchymoses around her left eye | 0
facial laceration | 0
decreased breath sounds on her right side | 0
no other obvious external signs of trauma | 0
Focused Assessment with Sonography for trauma (FAST) | 0
negative FAST | 0
isotonic fluid | 0
normalization of her blood pressure | 1
chest X-ray | 1
large right pneumothorax | 1
successful re-expansion of the lung | 1
chest tube | 1
vitals normalized | 2
intubated for agitation | 2
CT head/C-spine | 2
CT Chest/Abdomen/Pelvis with IV contrast | 2
grade 5 liver laceration | 2
grade 5 right kidney laceration | 2
grade 1 splenic laceration | 2
left clavicle fracture | 2
bilateral small pneumothoraces | 2
hypotensive | 3
operating room | 3
large amount of blood | 3
evacuated | 3
four-quadrant packing | 3
right medial visceral rotation | 3
large hematoma in the retroperitoneum | 3
shattered inferior portion of the kidney | 3
superior portion of the kidney was bleeding significantly | 3
renal vessels doubly ligated | 3
nephrectomy | 3
right ureter was unable to be located | 3
hemostasis of the spleen and liver | 3
other abdominal injuries were excluded | 3
repacked | 3
Barker vac | 3
Intensive Care Unit (ICU) | 4
7 units of packed red blood cells | 4
3 units of fresh frozen plasma | 4
4 l of crystalloid | 4
Interventional Radiology | 6
no active extravasation | 6
hepatic or splenic artery | 6
re-exploration | 48
active bleeding over the dome of the liver | 48
repacked | 48
hemostasis | 48
third laparotomy | 120
packs were removed without any bleeding | 120
right ureterectomy | 120
abdomen was closed primarily | 120
ICU | 120
extubated | 168
persistently elevated WBC | 168
CT abdomen/pelvis with IV contrast | 312
right kidney remnant isolated from the collecting system | 312
large, well-defined rim-enhancing collection | 312
urinoma | 312
ultrasound-guided drainage | 384
8 French drainage catheter | 384
cultures sent front the collection were without growth | 384
persistent drainage | 408
IR angioembolization of the remnant right kidney | 408
completion nephrectomy | 408
embolization of the right kidney remnant | 456
traumatic pseudoaneurysms | 456
embolized with 300–500 micron embospheres | 456
lower renal artery was completely occluded | 456
2 × 3 mm tornado microcoil | 456
completion arteriogram | 456
successful occlusion | 456
zero blood flow within the kidney remnant | 456
febrile | 456
severe flank pain | 456
antibiotics | 456
afebrile | 480
resolution of her pain | 480
drain was removed | 600
stable for discharge home | 600
BUN/Cr was 17/1.16 | 600