28 years old | 0
male | 0
insulin-dependent diabetes mellitus | 0
admitted to the ED | 0
urinary incontinence | -8760
dysuria | -8760
shortness of breath | -8760
cachexia | 0
suprapubic tenderness | 0
diffuse lung crackles | 0
decreased breath sounds on the right | 0
blood pressure 150/91 | 0
pulse 84 | 0
temperature 97.5 | 0
respiratory rate 16 | 0
urinalysis revealed white blood cells | 0
leukocyte esterase | 0
blood | 0
10000 mg/dL of glucose | 0
admitted to the Intensive Care Unit | 0
concern over respiratory status | 0
Chest CT scan | 0
multiple bilateral densities and nodules | 0
large consolidated cavitated mass occupying all three lobes of the right lung | 0
Abdominal CT | 0
bilateral hydroureteronephrosis | 0
large fluid collection at the bladder base | 0
suspicious for an abscess causing post-renal obstructive nephropathy | 0
Urology and infectious disease were consulted | 0
bronchoalveolar lavage | 0
urine culture grew Coccidioides immitus | 0
Coccidioidal serology was reactive for both IgG and IgM | 0
complement fixation titer was 1:128 | 0
severe disseminated coccidioidal infection | 0
treated with intravenous amphotericin B | 0
Urology consult recommended CT-guided drainage of the prostatic abscess | 0
drained pus cultured C. immitis | 0
closely monitored in the ICU | 0
follow up CT scan | 336
resolution of the abscess | 336
downtrending serum creatinine values | 336
symptomatic improvement | 336
transferred to the medicine wards | 336
course of amphotericin B was completed | 336
symptoms resolved | 336
discharged | 336