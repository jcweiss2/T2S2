63 years old | 0
male | 0
admitted to the hospital | 0
history of altered sensorium | -72
diabetic | -7200
below-knee amputation | -336
hypoglycemic | 0
pallor | 0
afebrile | 0
febrile | 72
urine sent for routine examination | 72
pus cells in urine | 72
Klebsiella spp. in urine culture | 72
sensitive to colistin | 72
sensitive to meropenem | 72
sensitive to cefoperazone + sulbactam | 72
sensitive to doxycycline | 72
sensitive to tigecycline | 72
resistant to nalidixic acid | 72
resistant to nitrofurantoin | 72
resistant to amikacin | 72
resistant to cefotaxime | 72
resistant to cefepime | 72
resistant to cefoperazone | 72
resistant to piperacillin + tazobactam | 72
ESBL producer | 72
Total leukocyte count 24,100/mm3 | 72
neutrophils 88% | 72
lymphocytes 8% | 72
eosinophils 3% | 72
basophils 1% | 72
hemoglobin 8.4 gm% | 72
platelet count 424,000/mm3 | 72
Serum sodium 137 meq/L | 72
Serum potassium 3.5 meq/L | 72
urea 33 mg/dL | 72
creatinine 0.87 unit/L | 72
blood sugar 119 mg/dL | 72
urinary bladder wall thickening | 72
sludge in urinary bladder | 72
started on intravenous meropenem | 72
afebrile | 120
electrolyte imbalance | 168
Na+ 123 meq/L | 168
K+ 3.9 meq/L | 168
Cl- 8.9 meq/L | 168
fever | 216
pus cells in urine | 216
red blood cells in urine | 216
Stenotrophomonas maltophilia in urine culture | 216
catalase positive | 216
oxidase negative | 216
motile | 216
gram negative rods | 216
reduced nitrates | 216
oxidized glucose | 216
oxidized lactose | 216
oxidized mannitol | 216
oxidized maltose | 216
hydrolyzed gelatin | 216
lysine decarboxylase test positive | 216
arginine hydrolysis negative | 216
susceptible to polymyxin B | 216
susceptible to cefoperazone | 216
susceptible to gatifloxacin | 216
susceptible to piperacillin + tazobactam | 216
susceptible to levofoxacin | 216
susceptible to colistin | 216
resistant to doxycycline | 216
resistant to cotrimoxazole | 216
resistant to meropenem | 216
resistant to amoxicillin + clavulanic acid | 216
resistant to cefotaxime | 216
resistant to ceftazidime | 216
resistant to ticaricillin + clavulanic acid | 216
resistant to nalidixic acid | 216
resistant to amikacin | 216
started on piperacillin + tazobactam | 216
clearance of pyuria | 240
discharged | 288