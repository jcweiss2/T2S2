60 years old | 0
male | 0
admitted to the hospital | 0
fever | -216
cough | -216
chills | -216
fever, cough, and chills did not respond to treatment with clarithromycin | -144
febrile | 0
tachycardic | 0
normotensive | 0
tachypneic | 0
basal rales | 0
perioral grouped blisters | 0
leukocytosis | 0
elevated C-reactive protein | 0
elevated total protein | 0
low albumin | 0
moderate hyponatremia | 0
community-acquired pneumonia | 0
started on empirical antimicrobial therapy with piperacillin/tazobactam plus clarithromycin | 0
blood cultures were positive for S. pneumoniae | 24
sputum cultures were positive for S. pneumoniae | 24
de-escalated to intravenous benzylpenicillin | 24
later to oral amoxicillin | 24
treated for a total duration of 14 days | 168
cutaneous herpes simplex type 1 infection | 0
treated with valaciclovir | 0
positive HSV-1 polymerase chain reaction result | 24
night sweats | -96
weight loss of 4 kg | -96
HIV test was negative | 24
elevated total protein and low albumin levels | 0
pneumococcal bacteremia | 0
suspected MM | 48
serum electrophoresis | 48
immunofixation identified an IgG kappa monoclonal gammopathy | 48
bone marrow biopsy revealed a plasma cell infiltration of >60% | 72
whole-body low-dose computed tomography scan demonstrated 4 lytic lesions in the pelvis and 1 in the cervical spine | 72
diagnosis of MM IgG kappa | 72
standard induction treatment with bortezomib, lenalidomide, and dexamethasone | 168
autologous hematopoietic stem cell transplantation | 168
treatment with intravenous immunoglobulin | 720
13-valent pneumococcal vaccination | 720
discharged | 168