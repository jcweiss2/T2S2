79 years old | 0
male | 0
severe septic shock | 0
urosepsis | 0
multi-organ failure | 0
acute on chronic renal failure | 0
acute respiratory distress syndrome | 0
Arterial hypotension | 0
drowsy mentation | 0
APACHE II score on admission | 0
APACHE II score of 32 | 0
CytoSorb therapy | 0
sustained low effusion dialysis | 0
SLED | 0
citrate | 0
flow rate of 100 ml/min | 0
standard surviving sepsis guidelines treatment | 0
improved hemodynamic parameters | 72
improved ventilator requirements | 72
increasing urine output | 72
APACHE II score of 8 | 72
IL-6 levels | 0
IL-6 level of 1356.3 pg/ml | 0
IL-6 level of 26.12 pg/ml | 72
deteriorated clinically | 120
immunosuppression | 120
removal of helpful anti-inflammatory cytokines | 120
