52 years old | 0
male | 0
colicky upper abdominal pain | -168
nausea | -168
vomiting | -168
pneumonia (2 episodes) | 0
thoracic empyema | 0
chronic pancreatitis | -17520
acute exacerbation of chronic pancreatitis | -17520
hypertension | 0
stage IV chronic renal disease | 0
pneumobilia | 0
tobacco smoker | 0
heavy drinker | 0
denied illicit drugs use | 0
not taking antibiotics | 0
not taking antiemetics | 0
not taking painkillers | 0
critically ill | 0
emaciated (BMI 18) | 0
dehydrated | 0
tachypneic | 0
tachycardic | 0
poor peripheral perfusion | 0
blood pressure 70/50 mmHg | 0
room air oximetry 88% | 0
Glasgow coma scale 15 | 0
cardiac examination unremarkable | 0
pulmonary examination unremarkable | 0
distended abdomen | 0
diffusely painful abdomen | 0
rebound tenderness | 0
normal bowel sounds | 0
mild anemia | 0
leukocytosis with marked left shift | 0
acute renal failure | 0
metabolic acidosis | 0
increased hepatic enzymes | 0
normal amylase | 0
normal lipase | 0
normal bilirubin | 0
normal clotting tests | 0
clinical diagnosis of peritonitis | 0
exploratory laparotomy | 0
free purulent effusion in abdominal cavity | 0
edema of intestinal loops | 0
edema of great omentum | 0
abscess in retro-cavity of epiplon | 0
peritoneal lavage | 0
abscess drainage | 0
closure of abdominal wound with Bogotá bag | 0
referred to intensive care unit | 0
mechanical ventilatory support | 0
vasoactive drugs | 0
hemodynamic instability | 0
death | 24
Escherichia coli culture positive | 0
Group F β-hemolytic Streptococcus culture positive | 0
Raoultella planticola culture positive | 0
median xipho-pubic surgical incision | 0
Bogotá bag closure of abdomen | 0
pleural adhesion in left hemithorax | 0
sero5.hemorrhagic effusion (400 mL) | 0
swollen viscera of peritoneal cavity | 0
fibrinoid material coating peritoneal cavity | 0
pancreas weight 183 g | 0
distorted pancreatic shape | 0
increased pancreatic fat tissue | 0
effaced pancreatic lobulation | 0
mousy pancreatic color | 0
white areas of hardened consistency in pancreas | 0
3 cm pseudocyst | 0
pseudocyst rupture | 0
pancreatic fibrosis | 0
acinar atrophy | 0
intraductal eosinophilic protein plugs | 0
chronic inflammatory infiltration | 0
fibrin coating peripancreatic tissue | 0
peritonitis (histological confirmation) | 0
acute inflammatory infiltration in pseudocyst | 0
venules thrombosis | 0
granulation tissue in pseudocyst | 0
lung atelectasis | 0
respiratory bronchiolitis | 0
tracheal squamous metaplasia | 0
myocardial hypertrophy | 0
bone marrow hypercellularity | 0
myeloid hyperplasia | 0
hepatocyte centrilobular trabeculation loss | 0
hepatocyte vacuolation | 0
acute tubular necrosis | 0
acute splenitis | 0
polymicrobial infection | 0
carbapenem-resistant strain (R. planticola) | 0
malnutrition | 0
immunologic disturbance | 0
pneumobilia as risk factor | 0
fatal outcome | 24
pancreatic pseudocyst co-infection | 0
antimicrobial sensitivity to cephalosporins | 0
antimicrobial sensitivity to fluoroquinolones | 0
antimicrobial sensitivity to carbapenems | 0
