50 years old | 0
male | 0
admitted to the hospital | 0
chest pain | -48
shortness of breath | -48
pulmonary emboli | -48
pulmonary infarction | -48
intubated | 144
severe respiratory distress | 144
progressive necrosis of the RLL infarction | 168
thoracotomy with partial decortication | 168
right thoracoscopy with 3 chest tubes placed | 168
piperacillin-tazobactam | 168
intravenous vancomycin | 168
bronchoalveolar lavage | 216
meropenem-susceptible A. baumannii | 288
antibiotics switched to meropenem | 288
thoracotomy with RLL resection and complete decortication | 288
new large multiloculated pleural effusion | 288
pleural tissue culture demonstrated XDR A. baumannii | 432
intermediate susceptibility to colistin | 432
tigecycline MIC of 2 mg/L | 432
switched from meropenem to tigecycline | 456
vasoactive agents | 624
RLL pyopneumothorax | 624
tigecycline switched to colistin and meropenem | 624
persistent purulent chest tube drainage | 672
bronchoscopy | 672
right bronchopleural fistula | 672
acute tubular necrosis | 672
serum creatinine increasing | 672
infectious diseases service requested eravacycline and cefiderocol susceptibilities | 696
eravacycline and cefiderocol susceptibilities resulted | 696
colistin and meropenem switched to renally adjusted cefiderocol | 696
significant chest tube output continued | 696
bronchial washings collected for culture | 960
XDR A. baumannii | 1080
cefiderocol-resistant | 1080
cefiderocol switched to eravacycline | 1176
eravacycline E-test MIC increased | 1296
eravacycline discontinued | 1296
combination therapy with cefiderocol and tigecycline initiated | 1296
chest tube output remained persistent | 1296
sulbactam–durlobactam susceptibility testing | 1296
SUL-DUR MIC | 1296
meropenem reduced the MIC | 1296
cefiderocol and tigecycline combination therapy discontinued | 1488
sulbactam–durlobactam plus meropenem started | 1488
resolution of chest tube output | 1800
antibiotics discontinued | 1800
discharged | 1872
followed up with ID as an outpatient | 1872
at prehospital baseline | 1872