27 years old | 0
female | 0
decompensated liver cirrhosis | 0
Model for End-Stage Liver Disease score of 30 | 0
primary biliary cholangitis | 0
autoimmune hepatitis overlap | 0
admitted to the intensive care unit | 0
septic shock | 0
acute kidney injury | 0
multidrug-resistant Escherichia coli urinary tract infection | 0
propranolol | -672
primary variceal prophylaxis | -672
chronic normocytic anemia | -672
baseline hemoglobin 8.5 mg/dL | -672
local admission for hematochezia | -144
esophagogastroduodenoscopy (EGD) | -144
nonbleeding grade I esophageal varices | -144
moderate portal hypertensive gastropathy | -144
flexible sigmoidoscopy | -144
mild, nonbleeding, internal hemorrhoids | -144
no rectal varices | -144
negative for spontaneous bacterial peritonitis | 0
hematochezia | 48
worsening anemia | 48
hemoglobin 5.7 mg/dL | 48
EGD | 48
severe portal hypertensive gastropathy | 48
nonbleeding, grade III esophageal varices | 48
esophageal varices banded 4 times | 48
flexible sigmoidoscopy | 48
bleeding rectal varix | 48
placement of 1 band | 48
worsening anemia | 72
hemoglobin 6.7 mg/dL | 72
packed red blood cells | 72
fresh frozen plasma | 72
repeat flexible sigmoidoscopy | 72
large blood clot | 72
ulceration | 72
mild oozing | 72
dislodgement of the band | 72
placement of 2 bands | 72
persistent hematochezia | 120
drop in hemoglobin | 120
hemoglobin 9 mg/dL | 120
hemoglobin 6.7 mg/dL | 120
packed red blood cells | 120
colonoscopy | 120
medium-sized, bleeding rectal varix | 120
stigmata of prior banding | 120
overlying clot | 120
necrotic ulcer base | 120
hot snare with soft coagulation | 120
resection of the protuberant part of the clot | 120
bleeding vessel | 120
over-the-scope clip (OTSC) | 120
placement of OTSC | 120
complete hemostasis | 120
transfer to a transplant center | 144
liver transplant evaluation | 144
death from septic shock | 168