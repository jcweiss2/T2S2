60 years old | 0
male | 0
admitted to the hospital | 0
fever | -48
abdominal pain | -48
edema of the scrotum | -48
edema of the penis | -48
edema of the perineum | -48
edema of the right gluteal region | -48
hypertension | -672
osteoporosis | -672
hemorrhoids | -672
blood pressure 103/62 mmHg | 0
heart rate 135/min | 0
oxygen saturation 88% | 0
white blood cell count 13.11/μL | 0
C-reactive protein level 61.4 mg/dL | 0
serum creatinine 4.3 mg/dL | 0
blood urea 157 mg/dL | 0
blood sugar 142 mg/dL | 0
procalcitonin 8.53 ng/mL | 0
SARS-CoV-2 infection suspected | 0
RT-PCR test for SARS-CoV-2 negative | 0
CT of the abdomen and the pelvis | 0
inflammatory infiltration of the subcutaneous tissues of the hypogastrium and the penis | 0
liquefaction and presence of gas in the subcutaneous tissues of the scrotum | 0
liquefaction and presence of gas in the subcutaneous tissues of the perineum | 0
liquefaction and presence of gas in the subcutaneous tissues of the right gluteal region | 0
Fournier's gangrene | 0
qualified to undergo surgery | 0
antibiotic therapy started | 0
meropenem 1 g thrice daily | 0
metronidazole 500 mg thrice daily | 0
linezolid 600 mg twice daily | 0
resection of the necrotic tissues | 24
bilateral orchiectomy | 24
excision of the penile and scrotal skin | 24
transferred to the intensive care unit | 24
mechanical ventilation | 24
broad-spectrum antibiotics | 24
supportive and nutritional therapies | 24
colostomy | 48
wound debridement | 48
negative pressure wound therapy | 48
sedation discontinued | 72
recovered consciousness | 72
extubated | 72
breathing on his own with oxygen on low flow | 72
hemodynamically stable | 72
diuresis stimulated using furosemide | 72
inflammatory markers decreased | 72
culture of the pus material showed Escherichia coli | 72
culture of the pus material showed Pseudomonas aeruginosa | 72
antibiotic therapy modified | 72
cephazolin 1g twice daily | 72
NPWT discontinued | 72
transferred to the Department of Plastic Surgery | 120
free-skin grafts applied | 168
discharged | 1104
testosterone supplementation 80 mg twice daily | 1104
physiotherapy | 1104
follow-up | 1104