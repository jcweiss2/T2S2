85 years old | 0
    male | 0
    melena | -3624
    weakness | -3624
    dizziness | -3624
    lower abdominal aortic dissecting aneurysm | -2376
    right common iliac arterial pseudoaneurysm | -2376
    lower abdominal aorta–common iliac artery bifurcated stent implantation | -2376
    melena | -2376
    tiredness | -2376
    dizziness | -2376
    hemoglobin decline from 11.5 to 7.0 g/dL | -2376
    superficial gastritis | -2376
    no definite bleeding source | -2376
    gastrointestinal bleeding attributed to aspirin-induced mucosal injury | -2376
    aspirin stopped | -2376
    blood transfusion | -2376
    proton pump inhibitors administered | -2376
    discharged | -2376
    hemoglobin level 7.8 g/dL | -2376
    progressive fatigue | -1464
    loss of appetite | -1464
    weight loss | -1464
    intermittent palpitation | -1464
    intermittent fever | -1464
    leukocytosis | -1464
    anemia | -1464
    diagnosed with pneumonia | -1464
    antibiotics prescribed | -1464
    discharged without significant improvement | -1464
    right back pain | -336
    right knee movement restriction | -336
    right leg swelling | -336
    pale | -336
    skinny | -336
    body temperature 38.2°C | -336
    pulse rate 96/min | -336
    respiratory rate 18/min | -336
    blood pressure 120/96 mm Hg | -336
    soft abdomen | -336
    nontender abdomen | -336
    no palpable masses | -336
    normal bowel sounds | -336
    severe anemia (hemoglobin 5.8 g/dL) | -336
    white blood cell count 8130/mm3 (82.3% granulocytes) | -336
    blood transfusion | -336
    antibiotics administered | -336
    CT showing gas shadow in right external iliac artery | -336
    gas shadow around lower abdominal aorta and common iliac artery | -336
    thrombosis in right common iliac artery | -336
    thrombosis in right external iliac artery | -336
    thrombosis in right common iliac vein | -336
    encapsulated fluid around right psoas | -336
    SAEF diagnosed | -336
    duodenoscopy revealing fistula in third part of duodenum | -336
    open surgery with extraanatomic bypass | 0
    exploratory laparotomy | 0
    aortic stent graft excision | 0
    infrarenal abdominal aortic suture | 0
    left common iliac artery ligation | 0
    extensive surgical debridement | 0
    retroperitoneal abscess resolution | 0
    drainage | 0
    duodenal defect repair | 0
    jejunal feeding tube placement | 0
    operation time 7 hours | 0
    transferred to intensive care unit | 0
    broad-spectrum intravenous antibiotics (imipenem/cilastatin) administered | 0
    multiorgan function monitoring | 0
    Enterococcus faecium in retroperitoneal abscess | 0
    Candida albicans in retroperitoneal abscess | 0
    vancomycin administered | 0
    fluconazole administered | 0
    hospital-acquired pneumonia | 240
    bilateral pleural effusion | 240
    heart failure | 240
    wide-spectrum intravenous antibiotics (imipenem/cilastatin) administered | 240
    cefoperazone/sulbactam administered | 240
    fluconazole continued | 240
    fluid intake restricted | 240
    condition improved | 240
    antibiotic administration terminated | 240
    progressive abdominal distension | 240
    partial small-bowel obstruction | 240
    postoperative intestinal adhesions | 240
    fasting | 240
    parenteral nutrition | 240
    gastrointestinal decompression | 240
    inhibition of gastric acid secretion | 240
    oral paraffin fluid | 240
    enema | 240
    recovered | 240
    no recurrent infection | 240
    no anemia | 240
    well for 15 months | 240