71 years old | 0
female | 0
admitted to the hospital | 0
fever | -3
chills | -3
peak temperature of 39 °C | -3
no cough | -3
no expectoration | -3
no pharyngeal pain | -3
no abdominal pain | -3
no diarrhea | -3
no increased urination frequency | -3
no increased urination urgency | -3
no perianal pain | -3
hypertension | -1092
valsartan | -1092
anemic | 0
wet rales in the right lung | 0
regular heart rhythm | 0
no obvious tenderness or rebound pain in the abdomen | 0
no obvious masses in the abdomen | 0
no edema in the limbs | 0
WBC count 13.2 × 10^9/L | 0
neutrophil percentage 88.5% | 0
hemoglobin 66 g/L | 0
platelet count 11 × 10^9/L | 0
blood glucose 33 mmol/L | 0
inflammation in both lungs | 0
bilateral pleural thickening | 0
thickening of the local intestinal wall in the ascending colon | 0
fever of undetermined origin | 0
pneumonia | 0
hypertension | 0
anti-inflammatory therapy | 0
meropenem | 0
human immunoglobulin | 0
erythrocyte suspension | 0
platelets | 0
insulin micropumps | 0
cold | 24
chills | 24
temperature reached 40 °C | 24
blood pressure dropped to 85/53 mmHg | 24
Escherichia coli in blood culture | 24
Aeromonas hydrophila in blood culture | 24
Aeromonas caviae in blood culture | 24
transferred to the intensive care unit | 24
meropenem micropump | 24
tetracycline | 24
fluid resuscitation | 24
vasoactive drugs | 24
decrease in platelets | 24
decrease in Hb | 24
decrease in WBC count | 24
recombinant human granulocyte colony-stimulating factor | 24
recombinant human PLT growth factor | 24
erythrocyte suspensions | 24
platelets | 24
supportive treatments | 24
infection controlled | 168
blood pressure returned to normal | 168
body temperature returned to normal | 168
blood culture was negative | 168
WBC count returned to normal | 168
Hb levels returned to normal | 168
platelets remained low | 168
bone marrow biopsy | 168
malignant cells in bone marrow smear | 168
cancer metastasis to the bone marrow | 168
18F-FDG PET/CT examination | 168
high metabolic signals in the ascending colon | 168
ascending colon malignant tumor | 168
conservative medical treatment | 168
tumor progressed | 504
patient died | 504
colon adenocarcinoma | 504
autopsy | 504
pathological results | 504