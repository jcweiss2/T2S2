39 years old | 0
female | 0
palpable mass on right breast | -168
Hodgkin lymphoma | -6336
chemotherapy | -6336
mantle field radiation | -6336
inflammatory colitis | -6336
mesalazine | -336
breast cancer | -168
invasive ductal carcinoma | -168
triple-negative phenotype | -168
MIB1 85% | -168
staging CT scan | -168
neoadjuvant chemotherapy | -112
paclitaxel | -112
carboplatin | -112
port-à-cath insertion | -84
subcutaneous cellulitis | -56
colliquative necrosis | -56
fever | -56
elevated white blood cell count | -56
neutrophilia | -56
elevated C-reactive protein | -56
broad-spectrum i.v. antibiotic therapy | -56
piperacillin/tazobactam | -56
daptomycin | -56
PORT rimotion | -56
necrosectomy | -56
defervescence | -48
improvement in subcutaneous cellulitis | -48
improvement in blood works | -48
febrile seizure | -40
WBC rise | -40
worsening of skin lesion | -40
second necrosectomy | -40
peripheral blood cultures | -40
skin plug | -40
i.v. catheter tip | -40
Klebsiella pneumoniae | -40
meropenem | -40
levofloxacin | -40
antibiotic therapy | -40
chest/abdomen CT scan | -40
mediastinitis | -40
bilateral pleural effusion | -40
left pulmonary atelectasis | -40
thoracoscopy | -32
pleural and mediastinal drainage | -32
sepsis | -32
broad-spectrum antibiotic | -32
antifungal therapy | -32
hemodynamic support | -32
non-invasive ventilation | -32
intensive inflammatory infiltrate | -32
neutrophils | -32
PG | -32
systemic methylprednisolone | -32
topical cyclosporine | -32
seriate chest X-ray | -24
progressive resolution of mediastinitis | -24
progressive resolution of pleural effusion | -24
wound improvement | -24
scar | -24
progressive normalization of blood count | -24
progressive normalization of flogosis index | -24
breast ultrasound | -16
no change in the dimension of the lump | -16
multidisciplinary meeting | -16
right mastectomy | -16
axillary dissection | -16
breast surgical wound healing | -16
fibroelastosis | -16
chronic inflammation | -16
isolated neoplastic cells | -16
restaging brain/chest/abdomen CT | -16
no distant metastasis | -16
BRCA | -16
p53 mutation tests | -16
autologous skin graft | 0
no further complications | 0
PICC implant | 0
chemotherapy | 0
carboplatin | 0
paclitaxel | 0
dose reduction | 0
good tolerance | 24
follow-up | 168
TILs | -168
moderate infiltrate | -16