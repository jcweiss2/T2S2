59 years old | 0
male | 0
Asian | 0
migrant worker | 0
admitted to the hospital | 0
diagnosed with COVID-19 | -336
severe COVID-19 | -336
acute disseminated encephalomyelitis (ADEM) | -294
encephalopathy | -294
generalised motor weakness | -294
multifocal magnetic resonance (MR) imaging findings | -294
intravenous immunoglobulin | -294
-67
-241
-190
septic shock | -294
inotropic support | -294
acute kidney injury | -294
haemodialysis | -294
deranged liver function | -294
provoked segmental pulmonary embolism | -294
polyarticular gout flare | -294
history of polyarticular gout | -8760
transferred out of intensive care | -286
minimal neurological recovery | -286
Glasgow Coma Scale (GCS) score of E4VTM1 | -286
no consistent visual pursuit | -286
vocalisations | -286
functional communication | -286
encephalopathy improved | -210
Coma Recovery Scale-Revised (CRS-R) score 9/23 | -210
follow instructions inconsistently | -198
CRS-R score improved to 10/23 | -157
nerve conduction study | -121
axonal sensorimotor polyneuropathy | -121
critical illness polyneuropathy | -121
transferred to inpatient rehabilitation facility | 0
GCS of E4V4M6 | 0
physiatrist-led transdisciplinary rehabilitation programme | 0
three hours per day of rehabilitation therapies | 0
physiotherapy | 0
occupational therapy | 0
speech therapy | 0
psychology reviews | 0
fortnightly dietician reviews | 0
weekly multidisciplinary conferences | 0
functional goal setting | 0
Functional Independence Measure (FIM) | 0
cognitive and behavioural impairments | 0
global and severe cognitive deficits | 0
sustained attention for 10–15 minutes | 0
disoriented | 0
slow information processing speed | 0
follow one-step commands only | 0
immediate information recall impaired | 0
Abbreviated Mental Test (AMT) score 1/10 | 0
participation limited | 0
attentional deficits | 0
slow processing speed | 0
impaired short-term memory | 0
therapy conducted in a quiet environment | 0
coaxing required | 0
cognitive demands reduced | 0
task simplification | 0
increased time for information processing | 0
episodes of irritability and agitation | 0
fatigue | 0
pain | 0
giddiness | 0
time-out-on-the-spot techniques | 0
redirection | 0
unable to use cognitive remediation strategies | 0
errorless learning | 0
repetition | 0
visual memory aids | 0
schedule reminders | 0
daily reality orientation | 0
flexibility of therapy timings | 0
sleep wake regulation | 0
AMT improved to 3/10 | 72
motivation and cooperation improved | 72
supportive counselling | 0
mobile digital media tools | 0
quadriparesis | 0
disproportionate spastic weakness | 0
lower limbs | 0
Medical Research Council (MRC) grade 2/5 | 0
upper limbs | 0
MRC scale 3/5 | 0
periventricular lesions | 0
motor recovery complicated | 0
critical illness polyneuropathy (CIP) | 0
steroid myopathy | 0
dependent in bed mobility | 0
poor sitting balance | 0
maximum assistance for activities of daily living (ADLs) | 0
physical therapy | 0
sitting balance | 0
sitting tolerance | 0
verticalisation via a tilt table | 0
task-specific training for ADLs | 0
mirror visual feedback | 0
grooming tasks | 0
orthostatic hypotension | 0
symptomatic postural hypotension | 0
severe deconditioning | 0
prolonged immobilisation | 0
blood pressure dropped | 0
fluids per day | 0
fluid boluses | 0
bilateral thigh-length elastic compression stockings | 0
abdominal binders | 0
passive increase venous return | 0
tolerated sitting at the edge of the bed | 80
mobilised in a tilt-in-space wheelchair | 80
swallowing and communication | 0
mild oropharyngeal dysphagia | 0
prolonged intubation | 0
tracheostomy | 0
ceased feeding through the nasogastric tube | -244
tolerated a blended diet | -244
video fluoroscopic swallowing study | -147
no aspiration | -147
regular diet consistency | -147
thin fluids | -147
controlled cup drinking | -147
resumed a normal diet | -147
functional communicative ability | 0
expressive speech | 0
receptive speech | 0
nutritional/metabolic parameters | 0
lost 14.4 kg | 216
body mass index (BMI) 21.6 kg/m2 | 216
premorbid weight of 84 kg | -336
BMI 26.5 kg/m2 | -336
nadir albumin level of 24 g/L | -222
improved to 30 g/L | 0
high caloric diet | 0
2,000 Kcal per day | 0
70 g of protein | 0
oral nutritional supplements | 0
nadir anaemia of 6.3 mg/L | -222
improved to 10.2 mg/L | 0
mild immobilisation-related hypercalcemia | -283
normalised during rehabilitation | 0
decubitus ulceration | -147
severe immobility | -147
prolonged recumbency | -147
6-cm × 4-cm Grade 3 sacral ulcer | -147
limited adjunctive mobilisation efforts | -147
electromechanical training | -147
automated body weight-supported treadmills | -147
contraindicated | -147
strict 2–3 hourly bed-turning | -147
pressure relief mattresses | -147
pressure offloading | -147
progressive increases in sitting duration | -147
meticulous skin dressing | -147
wound checks | -147
wound healing | 72
urinary incontinence | 0
indwelling urinary catheter | -147
skin hygiene | -147
regained spontaneous voiding | 72
dependent on diapers | 72
recurrent nosocomial infections | 0
catheter-associated urinary tract infections | 0
Clostridium difficile diarrhoea | 0
responded to appropriate antibiotics | 0
recurrent polyarticular gout flares | 0
left hip | -290
both knees | -290
ankles | -290
first metatarsal phalangeal joints | -290
hindered rehabilitation | 0
right knee aspiration | -290
left hip aspiration | -162
turbid straw-coloured fluid | -290
negatively birefringent crystals | -290
no evidence of septic arthritis | -290
treated with oral prednisolone | -290
uric acid-lowering therapy | -290
febuxostat | -290
renal impairment | -290
serum uric acid levels decreased | 0
acute and chronic lower body pain | 0
intermittent lower limb pain | 0
back pain | 0
impaired sensory discrimination | 0
severe cognitive deficits | 0
multifactorial pain | 0
polyarticular gout flares | 0
decubitus ulcer | 0
joint stiffness | 0
prolonged ICU immobilisation | 0
axonal sensorimotor polyneuropathy | 0
primary neurological insult | 0
central neuropathic pain | 0
spinal-thalamic-cortical pathways | 0
bilateral adductor spasticity | 0
restricted hip abduction | 0
flexion | 0
pain managed | 0
simple analgesia | 0
acetaminophen | 0
NSAIDS | 0
gabapentin | 0
physical modalities | 0
superficial heat | 0
electrical stimulation | 0
contraindicated | 0
insensate skin | 0
cognitive impairment | 0
FIM data | 0
low FIM efficiency | 0
slow progress | 0
high dependency | 0