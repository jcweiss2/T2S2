73 years old | 0
    male | 0
    admitted to the hospital | 0
    lower back pain | 0
    severe fatigue | 0
    20-kg weight loss | 0
    early-stage transitional cell bladder cancer | -105120
    invasion of the submucosa | -105120
    transurethral resection | -105120
    intravesical mitomycin | -105120
    recurrence of disease | -101088
    transurethral resection | -101088
    low-grade non-muscle-invasive tumor | -101088
    adjuvant therapy with intravesical BCG solution | -101080
    once weekly for 6 weeks | -101080
    no adverse events | -101080
    no immunocompromising conditions | -101080
    peripheral edema of the lower extremities | 0
    pain on palpation cranial to the left iliac crest | 0
    no abnormalities on abdomen | 0
    no abnormalities on spine | 0
    occult metastatic disease | 0
    positron emission tomography scan | 0
    pathologic activity of the abdominal aorta | 0
    pathologic activity of the left iliopsoas muscle | 0
    thoracoabdominal computed tomography scan | 0
    pseudoaneurysm of the abdominal aorta | 0
    surrounding infiltration | 0
    mycotic aneurysm | 0
    no septic episodes | 0
    not acutely ill | 0
    mildly elevated infection indicators | 0
    elective open aorta reconstructive surgery | 0
    no preoperative antibiotics | 0
    intravenous perioperative antibiotic prophylaxis | 0
    cephalosporin | 0
    metronidazole | 0
    postoperative antibiotic treatment dependent on culture | 0
    aneurysm began caudal to renal arteries | 0
    neoaortoiliac system bypass considered | 0
    reconstructive repair with bovine tube graft | 0
    infected aneurysmal segment excised | 0
    softened infected mushy tissue on left side | 0
    culture samples taken | 0
    biopsy specimens taken | 0
    excised infected tissue | 0
    resorbable sponge with gentamicin left | 0
    rifampicin applied to cavity | 0
    graft sutured conventionally | 0
    greater omentum wrap plasty | 0
    para-aortic tissue cultured | 0
    M. bovis cultured | 0
    extensive granulomatous inflammation | 0
    necrotizing inflammation | 0
    negative Ziehl-Neelsen staining | 0
    DNA analysis confirmed BCG strain | 0
    source of M. bovis infection | 0
    notified manufacturer | 0
    initial antimicrobial treatment | 0
    rifampicin | 0
    ethambutol | 0
    isoniazid | 0
    pyrazinamide | 0
    pyrazinamide discontinued | 24
    severe inflammatory response syndrome | 24
    admitted to intensive care unit | 24
    acute-on-chronic renal insufficiency | 24
    hemodialysis | 24
    paralytic ileus | 24
    chylous ascites | 24
    paracentesis | 24
    total parenteral nutrition | 24
    octreotide | 24
    condition improved | 72
    hemodialysis stopped | 72
    chylous ascites diminished | 72
    ileus resolved | 72
    transferred to general surgery ward | 72
    condition improved | 72
    transferred to rehabilitation center | 1440
    antimicrobial treatment continued | 1440
    readmitted with fever | 2160
    generalized weakness | 2160
    malaise | 2160
    fever | 2160
    tachycardia | 2160
    elevated C-reactive protein | 2160
    leukocytosis | 2160
    CT scan showed fluid collection | 2160
    CT-guided drainage | 2160
    fluid cultured | 2160
    mycobacterium in aspirated fluid | 2160
    unclear active infection or paradoxical abscess | 2160
    treatment for active infection | 2160
    treatment for paradoxical abscess | 2160
    antibiotic regimen changed | 2160
    rifampicin | 2160
    ethambutol | 2160
    moxifloxacin | 2160
    dexamethasone | 2160
    condition improved | 2160
    follow-up CT scan | 2160
    collection decreased | 2160
    discharged | 2160
    outpatient monitoring | 2160
    