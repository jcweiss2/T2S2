14 years old | 0
    female | 0
    upper left teeth pain | -504
    bulging of the maxillary region | -504
    prescribed cephalexin | -504
    behavioral alterations | -168
    auditory hallucination | -168
    sleep disturbances | -168
    aggression | -168
    frontal headache | -168
    headache (14-day history) | -336
    agitation | 0
    aggressiveness | 0
    somnolence | 0
    mental confusion | 0
    vomiting | 0
    paranasal sinuses CT scan | 0
    brain CT scan | 0
    right maxillary sinuses opacification | 0
    frontal sinuses opacification | 0
    frontal sinus osseous erosion | 0
    subdural empyema | 0
    slight cerebral edema | 0
    inflammatory alterations (lab work-up) | 0
    no acid-base imbalance | 0
    no electrolytes imbalance | 0
    hemoglobin 10.9 | 0
    hematocrit 33.6 | 0
    leukocytes 20,400 | 0
    bands 0 | 0
    segmented 82.8 | 0
    lymphocyte 6.7 | 0
    monocytes 10.5 | 0
    platelets 363,000 | 0
    urea 18 | 0
    creatinin 0.55 | 0
    CRP 174 | 0
    blood culture negative | 0
    referred to pediatric ICU | 0
    empirical antibiotics (ceftriaxone, levofloxacin, vancomycin, acyclovir) | 0
    neurologic deterioration | 0
    sudden cardiopulmonary arrest | 0
    resuscitation maneuvers | 0
    recovered sinus rhythm | 0
    GCS 3 | 0
    new CT scan | 0
    diffuse cerebral edema | 0
    brain herniation | 0
    left internal jugular vein thrombosis | 0
    death | 48
    CSF analysis | 48
    clear CSF appearance | 48
    CSF protein 385.7 | 48
    CSF WBC count 250 | 48
    CSF erythrocytes 50 | 48
    CSF neutrophils 49 | 48
    CSF lymphocytes 30 | 48
    CSF monocytes 21 | 48
    CSF glucose 54 | 48
    CSF lactate 82.7 | 48
    CSF Pandy positive | 48
    CSF culture negative | 48
    negative serology (cytomegalovirus, Epstein Barr virus, HSV-1, HSV-2, varicella-zoster virus, human enteroviruses) | 48
    autopsy performed | 48
    meningeal purulent exudate | 48
    frontal bone erosion | 48
    acute meningitis (neutrophils) | 48
    acute osteomyelitis (frontal, mastoid bones) | 48
    neuronal necrosis | 48
    glial necrosis | 48
    diffuse encephalic ischemia | 48
    left internal jugular vein thrombosis | 48
    thrombophlebitis (superior vena cava, left brachiocephalic vein) | 48
    pneumonia | 48
    alveolar edema | 48
    neutrophilic infiltration (liver, spleen, heart, lymph nodes, bone marrow) | 48
    sepsis | 48
    acute tubular necrosis | 48
