75 years old | 0
male | 0
admitted to the hospital | 0
dyspnoea | -96
chronic heart insufficiency | -0
atrial fibrillation | -0
arterial hypertension | -0
type 2 diabetes mellitus | -0
chronic renal insufficiency | -0
polyneuropathy | -0
dual chamber pacemaker implanted | -1920
started on antibiotics | 0
furosemide | 0
elevated inflammatory markers | 0
C reactive protein | 0
leucocytes | 0
high admission brain natriuretic peptide | 0
transferred to the intensive care department | 0
tachypnoeic | 0
peripheral saturation of 85% | 0
on 10 L/min O2 | 0
via Hudson mask | 0
normotensive | 0
atrial fibrillation | 0
VVI pacing to 70 bpm | 0
cardiac biochemistry negative | 0
troponin I | 0
CK-MB mass | 0
myoglobin | 0
transthoracic echocardiography | 0
congestive heart failure | 0
hypokinetic anteroseptal left ventricular wall | 0
ejection fraction of 38% | 0
moderate mitral regurgitation | 0
dilated left atrium | 0
mild aortic regurgitation | 0
moderately dilated right ventricle | 0
tricuspid annular plane systolic excursion of 23 mm | 0
moderate tricuspid regurgitation | 0
estimated right-sided pleural effusion of 300–400 mL | 0
VVI pacing reset to 90 bpm | 0
limited aeration of the right lower lobe | 36
bronchial breathing | 36
intubated | 36
bronchoscopy | 36
norepinephrine infusion | 36
PSV of 14 cmH2O | 36
PEEP of 8 cmH2O | 36
FiO2 0.50 | 36
tachypnoeic | 36
increasing requirements for oxygen | 36
decreased blood pressure | 36
decreased urine output | 36
elevated left ventricular end-diastolic pressure | 36
moderate-to-severe MR | 36
dilated LA | 36
estimated pulmonary artery systolic pressure of 57 mm Hg | 36
right pleural tap | 36
12F drain | 36
closed collection system | 36
850 mL of transudate evacuated | 36
dobutamine 5.0 µg/kg/min | 36
positive effect on CO | 36
oxygenation | 36
weaned off the mechanical ventilation | 60
extubated | 60
continued on Hudson mask | 60
FiO2 of 0.6 | 60
discharged to a high dependency unit | 168
sufficient expectoration | 168
on antibiotics | 168
NAD 0.08 µg/kg/min | 168
VVI 90 bpm | 168
discharged on day 19 | 456