56 years old | 0
female | 0
cirrhosis | -672
chronic hepatitis C | -672
esophagogastroduodenoscopy | 0
esophageal varices | 0
varix ruptured | 0
TIPS procedure | 0
GORE VIATORR covered stent | 0
transfusion of packed red blood cells | 0
admitted to medical intensive care unit | 0
jaundiced | 72
increased total and direct bilirubin | 72
stable transaminases | 72
stable INR | 72
abdominal ultrasound | 72
patent stent | 72
no biliary obstruction | 72
rising bilirubin | 96
stable alkaline phosphatase | 96
stable transaminases | 96
stable INR | 96
abdominal CT | 120
patent TIPS | 120
no hepatic ischemia | 120
no biliary duct dilatation | 120
ERCP | 360
no biliary-venous fistula | 360
common bile duct stent | 360
sphincterotomy | 360
rising bilirubin | 360
venogram | 360
no biliary-venous fistula | 360
resistant Klebsiella bacteremia | 360
sepsis | 360
renal failure | 360
transferred to intensive care unit | 360
discharged home with hospice care | 720
liver transplantation | 720 
hepatic encephalopathy | -672
hemolytic anemia | -672
hepatic ischemia | -672
stent thrombosis | -672
biliary tree stricture | -672
biliary obstruction | -672
post-TIPS hemolysis | -672
Enterobacteriaceae bacteremia | 360
fat embolism | 360
bile thromboembolism | 360
percutaneous biliary drainage | 720
endoscopic nasobiliary drainage | 720
venous balloon occlusion | 720 
spontaneous closure of biliary-venous fistula | 720