27 years old | 0
female | 0
grade III lesion of pancreas | 0
fell from bicycle | 0
landed on handlebar | 0
pancreatic contusion | 0
trauma CT scan | 0
referred to level 1 trauma center | 0
reassessment of CT scan | 0
complete rupture of pancreatic neck | 0
retroperitoneal hematoma | 0
no other abdominal injuries | 0
MRCP confirmed rupture of main duct | 0
diastasis measuring 2 cm | 0
conservative approach | 0
nasogastric tube | 0
continuous suction | 0
intravenous proton pump inhibitor | 0
pantoprazole 40 mg b.i.d. | 0
subcutaneous octreotide 100 microgram t.i.d. | 0
intravenous cefuroxime 1500 mg t.i.d. | 0
metronidazole 1500 mg q.d. | 0
parenteral nutrition | 0
ERCP | 72
papillotomy of pancreatic duct | 72
no attempt to insert bridge prosthesis | 72
patient's condition deteriorated | 96
increasing abdominal pain | 96
inflammatory parameters | 96
free intraperitoneal fluid | 96
ultrasonography | 96
laparotomy | 96
removal of 2000 ml ascites | 96
no resection of distal part of gland | 96
placement of two external 18 Fr tubes | 96
abdomen closed | 96
general condition improved | 96
no need for pain killers | 96
systemic inflammatory response decreased | 96
started eating regular food | 96
one abdominal tube discontinued | 96
stable fluid level in remaining tube | 96
discharge | 384
follow-up once a week | 384
intermittent retraction of drain | 384
drain removed | 1344
discharge ceased from fistula | 1344
increasing discomfort | 1344
abdominal pain | 1344
CT scan revealed pseudocyst | 1344
MRCP | 1344
MR angiography | 1344
severed pancreatic duct with diameter 6 mm | 1344
both halves of gland with arterial perfusion | 1344
endoscopic ultrasonography | 1344
HOT AXIOSTM stent inserted | 1344
stent deployed | 1344
patient ate normally | 1344
abdominal pain ceased | 1344
discharged | 1368
CT scan revealed collapsed cyst | 1368
stent removed | 2160
CT scan showed no recurrence of cyst | 2160
pancreatic duct still measured 6 mm | 2160
both halves of pancreas had blood supply | 2160
patient doing well | 2160
no signs of malabsorption | 2160
no diabetes | 2160
follow-ups terminated | 2160
open contact to department | 2160
