87 years old | 0
male | 0
atrial fibrillation | 0
CHA2DS2-VASc score of 5 | 0
heart failure with preserved ejection fraction | 0
hypertension | 0
admitted to the hospital | 0
weakness | 0
decreased oral intake | 0
mild cough | 0
dabigatran etexilate 150 mg twice-daily | -3600
thromboembolic prophylaxis of atrial fibrillation | -3600
increased lower extremity edema | -168
atrial fibrillation with a rapid ventricular response averaging 120 beats per minute | -168
serum creatinine 1.20 mg/dL | -168
eGFR 57 mL/min/1.73 m² | -168
verapamil increased from 120 to 240 mg | -168
metoprolol increased from 25 to 100 mg | -168
furosemide increased from 40 to 60 mg | -168
fell while getting out of bed | -48
too weak to stand | 0
vomited three times | 0
last dose of dabigatran taken | -48
axillary temperature 95.7 °F | 0
blood pressure 102/48 mmHg | 0
ventricular rate 36 beats/min | 0
oxygen saturation 96% on 2 L/min supplemental oxygen | 0
jugular venous distension with monophasic waves | 0
hepatojugular reflux | 0
bibasilar crackles | 0
bradycardic irregular rhythm | 0
systolic murmur III/VI | 0
benign abdomen | 0
3+ pitting edema of extremities | 0
normal pulses bilaterally | 0
atrial fibrillation with ventricular response rate ~36 beats/min | 0
right lower lobe infiltrate on chest X-ray | 0
acute renal failure | 0
hepatic dysfunction | 0
septic shock from pneumonia | 0
increased diuretic therapy | 0
bradycardia | 0
electrolyte disturbances | 0
elevated serum lactate | 0
profound coagulopathy | 0
hyperkalemia | 0
received insulin | 0
received dextrose | 0
received calcium gluconate | 0
received sodium bicarbonate | 0
no acute hemorrhage | 0
no fracture | 0
received IV normal saline | 0
received IV glucagon | 0
cultures obtained | 0
treatment with ceftriaxone | 0
treatment with levofloxacin | 0
sodium 137 mmol/L | 0
potassium 6.6 mmol/L | 0
chloride 100 mmol/L | 0
total CO2 10 mmol/L | 0
blood urea nitrogen 45 mg/dL | 0
creatinine 3.05 mg/dL | 0
glucose 102 mg/dL | 0
magnesium 2.6 mg/dL | 0
ALT 546 U/L | 0
AST 422 U/L | 0
alkaline phosphatase 111 U/L | 0
total bilirubin 1.4 mg/dL | 0
direct bilirubin 0.5 mg/dL | 0
CK 170 U/L | 0
CKMB 5.9 ng/mL | 0
troponin T 0.08 ng/mL | 0
NT-proBNP 3,695 pg/mL | 0
white blood cell count 18.52 K/μL | 0
hemoglobin 14.0 g/dL | 0
hematocrit 43.5% | 0
platelet count 214 K/μL | 0
PT 54.4 s | 0
PTT 100.6 s | 0
INR 6.0 | 0
fibrinogen 279 mg/dL | 0
diluted TT 125.0 s | 24
diluted TT 113.1 s | 26
heart rate 48 beats/min | 24
blood pressure 90/50 mmHg | 24
worsening hypoxia | 24
placed on high flow nasal cannula | 24
became acutely unresponsive | 24
loss of palpable pulses | 24
progressive bradycardia <30 beats/min | 24
received chest compressions | 24
return of spontaneous circulation | 24
intubated | 24
mechanical ventilation | 24
no overt signs of active bleeding | 24
hematocrit 33.9% | 24
received FFP | 24
received vitamin K | 24
received PCC | 24
PT and PTT returned to normal | 72
thrombin time >150 s | 24
ALT 4,590 U/L | 24
AST 4,965 U/L | 24
creatinine 3.07 mg/dL | 24
eGFR ≤20 mL/min/1.73 m² | 24
stabilized in ICU | 168
extubated | 120
discharged home | 456
INR 1.8 | 120
PTT 46.9 s | 120
started heparin infusion | 120
started warfarin | 168
creatinine 0.70 mg/dL | 456
PTT 41.3 s | 456
INR 1.8 on warfarin | 456
ALT 271 U/L | 240
AST 32 U/L | 240
