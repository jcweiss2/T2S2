62 years old | 0
male | 0
non-smoker | 0
admitted to the hospital | 0
complaint of worsening pain in the left groin | 0
subjective fevers | 0
second dose of the ChAdOx1 nCoV-19 vaccine | -336
experienced one episode of diarrhoea | -240
total replacement of the left hip | -13140
arthrosis secondary to hip dysplasia | -13140
hypertension | 0
paroxysmal atrial fibrillation | 0
rivaroxaban | 0
admitted to a hospital with diarrhoea, haematochezia, and Bacteroides vulgatus bacteremia | -4380
treated successfully with antibiotics | -4380
no significant gastrointestinal abnormality | -4380
afebrile | 0
mild tachycardia | 0
hypotensive | 0
left hip joint showed irritability to passive movements | 0
elevated levels of inflammatory markers | 0
normal levels of blood metal ion | 0
pelvic x-ray showed no new changes to the prosthesis | 0
aspiration of the hip performed | 0
yielded 20 mL of haemoserous fluid | 0
250,200 white blood cell count (WBC)/µL | 0
gram-negative and positive bacilli detected on microscopy | 0
started on empirical intravenous antibiotic therapy (cefazolin) | 0
transferred to the intensive care unit | 0
light growth of tiny, grey, translucent colonies isolated on an anaerobic agar plate | 48
identified as F. plautii | 96
antibiotic regimen changed to include amoxycillin-clavulanate, gentamicin, metronidazole, and vancomycin | 96
underwent a first-stage revision hip arthroplasty | 168
exploration of the hip performed using the posterior approach | 168
detection of extensive abscess formation and destruction of soft tissue deep to the fascia | 168
debridement of extensive erosion of pericapsular soft tissue performed | 168
pulse lavage and intermittent irrigation with hydrogen peroxide performed | 168
extraction of all hardware followed by implantation of an antibiotic cement articulating spacer | 168
thickened ascending colon observed on a postoperative computed tomography of the abdomen | 168
colonoscopic biopsy showed a single sigmoid tubular polyp and diverticular disease | 168
conservative management administered | 168
received 24-hour intravenous administration of ceftriaxone | 0
received oral amoxicillin/clavulanic acid and metronidazole | 1008
normalisation of the C-reactive protein occurred | 1008
aspiration of the hip performed after completion of oral antibiotics | 1008
yielded 832 WBC/µL, 20% polymorphonuclear cells and negative cultures | 1008
second stage revision arthroplasty performed | 2160
extraction of the antibiotic cement and all spacer implants performed | 2160
no macroscopic evidence of infection or bone necrosis observed | 2160
multiple swabs and tissue cultures sent from both acetabular and femoral sites showed no growth on extended culture | 2160
administration of routine intraoperative surgical antibiotic prophylaxis performed | 2160
preparation of acetabular and femoral sides performed with implantation of uncemented components | 2160
discharged on day 7 | 2160
recovery was uncomplicated | 2160
remains in good health without ongoing infective issues at 12-month follow-up | 8760
remains off antibiotics | 8760
normal, pain free gait with near normal hip range of movement observed by physical examination | 8760