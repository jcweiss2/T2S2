15 years old | 0
male | 0
admitted to the hospital | 0
fever | -24
confusion | -24
eating meat in a fast food restaurant | -24
sweating | -24
vomiting | -24
myalgias | -24
cutaneous rash | -24
mild confusion | 0
body temperature 38.6 °C | 0
blood pressure 60/30 mmHg | 0
heart rate 170 bpm | 0
oxygen saturation 98% | 0
diffuse cutaneous exanthema | 0
chest exanthema | 0
upper limbs exanthema | 0
moderate abdominal tenderness | 0
elevated inflammatory markers | 0
WBC 21000/mm³ | 0
neutrophils 92% | 0
CRP 250 mg/L | 0
coagulopathy | 0
acute renal failure | 0
transferred to Intensive Care Unit | 0
stabilized with intravenous fluids | 0
vasopressors | 0
empirical amoxicillin-clavulanate initiated | 0
blood cultures positive for staphylococci | 24
Staphylococcus aureus identified | 24
PBP2a test negative | 24
multi-sensitive bacterial strain confirmed | 24
follow-up blood cultures negative | 24
stool culture negative | 24
trans-esophageal echocardiography normal | 24
intravenous antibiotics treatment for 7 days | 0
discharged | 168
oral antibiotics for one more week | 168
hand desquamation | 336
feet desquamation | 336
tsst-1 gene presence confirmed | 336
eta toxin absence | 336
etb toxin absence | 336
t2509 Staphylococcus aureus strain | 336
food poisoning suspected | 336
no risk factors for TSS | 336
initial digestive symptoms | 336
- 15 years old | 0
- male | 0
- admitted to the hospital | 0
- fever | -24
- confusion | -24
- eating meat in a fast food restaurant | -48
- sweating | -24
- vomiting | -24
- myalgias | -24
- cutaneous rash | -24
- mild confusion (noted by mother) | 0 (upon admission)
- body temperature 38.6 °C | 0
- blood pressure 60/30 mmHg | 0
- heart rate 170 bpm | 0
- oxygen saturation 98% | 0
- diffuse cutaneous exanthema | 0
- chest exanthema | 0
- upper limbs exanthema | 0
- moderate abdominal tenderness | 0
- mild confusion (on exam) | 0
- elevated inflammatory markers | 0
- WBC 21000/mm³ | 0
- neutrophils 92% | 0
- CRP 250 mg/L | 0
- coagulopathy | 0
- acute renal failure | 0
- transferred to Intensive Care Unit | 0
- stabilized with intravenous fluids | 0
- vasopressors | 0
- empirical amoxicillin-clavulanate initiated | 0
- blood cultures positive for staphylococci | 24
- Staphylococcus aureus identified | 24
- PBP2a test negative | 24
- multi-sensitive bacterial strain confirmed | 24
- follow-up blood cultures negative | 24
- stool culture negative | 24
- trans-esophageal echocardiography normal | 24
- intravenous antibiotics treatment for 7 days | 0 (start time)
- discharged | 168 (after 7 days)
- oral antibiotics for one more week | 168
- hand desquamation | 336 (2 weeks after onset)
- feet desquamation | 336
- tsst-1 gene presence confirmed | 336
- eta toxin absence | 336
- etb toxin absence | 336
- t2509 Staphylococcus aureus strain | 336
- food poisoning suspected | 336 (when PCR results available)
- no risk factors for TSS | 0 (noted during admission)
- initial digestive symptoms | -24 (vomiting, etc.)
+ emesis | -44
+ diarrhea | -44
+ fever | -24
+ confusion | -24
+ sweating | -24
+ vomiting | -24
+ myalgias | -24
+ cutaneous rash | -24
- emesis | -44
# diarrhea | -44
- emesis | -44 (four hours after eating)
- diarrhea | -44
- fever | -24 (one day after eating)
