46 years old | 0
male | 0
benign prostatic hyperplasia | -672
end-stage renal disease requiring hemodialysis | -672
presented to the emergency department with peritonitis and septic shock | -24
computed tomography revealed pneumoperitoneum | -24
taken to the operating room for diagnostic laparoscopy | -24
gross bilious contamination of the entire peritoneal cavity found | -24
perforation of the anterior duodenal bulb identified | -24
modified Graham patch fashioned using a well-vascularized tongue of the greater omentum | -24
endoscopic leak test performed with positive results | -24
procedure converted to an open approach via midline laparotomy | -24
Graham patch reconstructed | -24
repeat endoscopic leak test negative | -24
abdomen irrigated | -24
drains placed by the repair | -24
abdomen closed in standard fashion | -24
intra-abdominal abscess developed | -144
percutaneous drainage on postoperative day 7 | -144
positive test result for Helicobacter pylori | 0
triple therapy (proton pump inhibitor, clarithromycin, and amoxicillin or an imidazole) started | 0
discharged on postoperative day 9 | 216
returned to the emergency room with hematochezia and symptomatic anemia requiring transfusion | 720
computed tomography angiography demonstrated inferior vena cava thrombus with intraluminal air formation concerning for duodenal-caval fistula | 720
upper endoscopy revealed clots and bleeding in the posterior wall of the second portion of the duodenum | 720
diagnosis of duodenal-caval fistula confirmed | 720
taken to the operating room for repair of the duodenal-caval fistula | 720
exploratory laparotomy performed | 720
prior Graham patch assessed and appeared intact | 720
Kocher maneuver performed to mobilize the duodenum | 720
duodenal-caval fistula identified | 720
proximal and distal control obtained of the supra% and infrahepatic IVC, left renal artery and vein | 720
Pringle maneuver performed | 720
right renal artery, vein, and ureter ligated to improve exposure | 720
control distal from the IVC thrombus verified using transesophageal echocardiography and intraoperative ultrasound | 720
duodenum completely dissected off the anterior wall of the IVC | 720
full extent of the fistula revealed with large thrombus identified | 720
clamps placed at the central IVC, renal vein, and peripheral IVC | 720
thrombectomy performed using transesophageal echocardiography to confirm complete evacuation of the thrombus and right ventricular integrity | 720
venorrhaphy performed using running 2-0 Prolene suture | 720
repair of the duodenal perforation using 4-0 Prolene suture | 720
vena cava inflamed but defect small enough for primary repair without narrowing lumen | 720
patch angioplasty avoided to prevent infectious complications | 720
nasogastric tube placed in the stomach for decompression | 720
abdomen temporarily closed using AbThera wound vacuum device | 720
transferred to intensive care unit postoperatively | 720
returned to the operating room for re-exploration on postoperative day 2 | 768
temporary abdominal closure removed | 768
peritoneal cavity inspected | 768
open cholecystectomy performed to prevent future biliary complications | 768
right nephrectomy performed | 768
abdominal cavity closed temporarily with AbThera device | 768
transferred to intensive care unit | 768
returned to the operating room the next day | 792
abdomen opened | 792
inspection of previous duodenal repair showed small opening | 792
small opening closed using 3-0 PDS | 792
omental patch placed on duodenal repair and IVC repair | 792
pyloric exclusion performed via gastrostomy created along the greater curvature of the stomach | 792
pylorus closed with two purse string sutures using 2-0 PDS | 792
enterolysis performed to mobilize enough intestine for gastrojejunostomy | 792
gastrojejunostomy created using 30-cm afferent jejunal limb from the ligament of Treitz | 792
decompressing nasojejunal tube placed in the proximal limb | 792
distal feeding tube placed in the efferent limb | 792
drains placed | 792
abdomen closed in standard fashion | 792
transferred to intensive care unit | 792
hemorrhagic shock on postoperative day 6 | 864
intraluminal bleeding from anomalous duodenal artery originating from the abdominal aorta | 864
emergent angioembolization by interventional radiology | 864
required percutaneous drainage of subhepatic fluid collection on postoperative day 13 | 936
experienced another episode of bleeding from the same anomalous duodenal artery | 1080
underwent repeat angioembolization on postoperative day 23 | 1080
discharged home on postoperative day 40 | 2160
doing well at latest outpatient follow-up | 2160
