53 years old | 0
female | 0
history of multiple cosmetic surgeries | 0
liposculpture surgery | -24
fever | 168
disabling pain at the surgical site | 168
extensive bullae formation | 168
septic shock | 96
vasopressor support | 96
mechanical ventilation | 96
acute renal failure | 96
admitted to the intensive care unit | 96
multiple and extensive lesions | 0
subcutaneous emphysema | 0
leakage of purulent material | 0
erythema | 0
necrosis at the wound edges | 0
CT scan of the abdomen | 0
cutaneous dehiscence | 0
extensive generalized soft tissue emphysema | 0
diagnosis of necrotizing soft tissue infection | 0
surgical wound cleansing | 0
mechanical scrubbing | 0
debridement | 0
prophylactic antibiotics | 0
identification of the pathogen involved | 0
surgical intervention for drainage | 24
debridement of necrotic tissue | 24
placement of a negative pressure therapy system | 24
metabolic acidosis | 0
hyperlactatemia | 0
leukocytosis with a left shift | 0
thrombocytopenia | 0
elevated CRP | 0
elevated ESR | 0
hyperlactatemia | 0
intensive care unit | 0
source of infection controlled | 168
hemodynamic stabilization | 168
hospitalized | 0
15 surgical interventions | 0
multiple wound cleansing | 0
debridement | 0
placement of a negative pressure therapy system | 0
advancement of flaps | 0
lesions reconstruction | 0
procurement and placement of grafts | 0
secretion cultures | 0
E. Coli | 0
Finegoldia magna | 0
Streptococcus mitis | 0
antibiotic management | 0
Vancomycin | 0
Meropenem | 0
Clindamycin | 0
discharged | 1008
intensive rehabilitation program | 1008
no further complications | 1008