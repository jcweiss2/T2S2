57 years old | 0
female | 0
menopausal | 0
admitted to the gynecological emergency unit | 0
left lower quadrant abdominal pain | -1008
pelvic heaviness | -1008
urinary frequency | -1008
past history of 5 miscarriages | -1008
tubal ligation | -1008
active smoker | 0
no medication | 0
large and painful mass | 0
pelvic MRI | 0
mass measuring 18 × 17 × 12 cm | 0
no lymphadenopathy | 0
no ascites | 0
no peritoneal implants | 0
uterus and adnexa were normal | 0
serum tumor markers were negative | 0
surgical pelvic exploration | -672
30-centimeter mass of the left broad ligament | -672
no ascites | -672
no peritoneal carcinomatosis | -672
uterus and right adnexa were normal | -672
total hysterectomy with adnexectomy | -672
removal of the mass | -672
definitive histological diagnosis was leiomyosarcoma | -672
isolated fever | 48
laboratory evaluation | 48
major inflammatory syndrome | 48
leukocytes 15,000/μL | 48
C-reactive protein 317 mg/dL | 48
contrast-enhanced computed tomography scan | 48
bilobed air and fluid collection | 48
abscess | 48
blood pressure dropped | 48
vasopressor therapy | 48
noradrenaline | 48
emergency revision surgery | 48
peritoneal cavity exploration | 72
moderately abundant non-purulent serosanginous peritoneal fluid | 72
adhesions to the Douglas pouch | 72
peritonitis | 72
antibacterial treatment with piperacillin/tazobactam and gentamicin | 72
microbiological samples | 72
extubated | 96
hemodynamic support with noradrenaline | 96
transferred to the intensive care unit | 96
noradrenaline requirement decreased | 120
discontinuation of noradrenaline | 120
decrease in inflammatory markers | 120
microbiological analysis of the peritoneal fluid | 120
Gardnerella vaginalis | 120
gentamicin discontinued | 120
metronidazole added | 120
Atopobium vaginae | 168
antibacterial susceptibility testing | 168
Gardnerella vaginalis resistant to metronidazole | 168
Gardnerella vaginalis susceptible to penicillin G | 168
Gardnerella vaginalis susceptible to amoxicillin/clavulanate | 168
Gardnerella vaginalis susceptible to cefotaxim | 168
Gardnerella vaginalis susceptible to clindamicin | 168
Gardnerella vaginalis susceptible to vancomycin | 168
Atopobium vaginae susceptible to metronidazole | 168
piperacillin/tazobactam active against both bacteria | 168
final diagnosis | 168
early postoperative peritonitis-induced septic shock | 168
caused by Gardnerella vaginalis and Atopobium vaginae | 168
discharged from the intensive care unit | 240
antibacterial therapy stopped | 336