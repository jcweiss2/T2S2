65 years old | 0
male | 0
allergic rhinitis | 0
eczema | 0
dyslipidemia | 0
benign prostatic hyperplasia | 0
blurring of vision | -2628
left visual field quadrantanopia | -2628
no papilloedema | -2628
no other neurological deficit | -2628
pituitary macroadenoma | -2628
low cortisol | -2628
low growth hormone | -2628
low testosterone | -2628
other neuroendocrine hormones normal | -2628
admitted for TSH | 0
TSH | 0
excision of tumor | 0
intraoperatively dura not breached | 0
extubated postoperatively | 0
transferred to ward | 0
polyuria | 24
treated for cranial diabetes insipidus | 24
desmopressin | 24
febrile | 168
tachypneic | 168
tachycardic | 168
minimal cough | 168
no neurological symptoms | 168
no CSF rhinorrhea | 168
air entry equal | 168
no adventitious sound | 168
minimal perihilar haziness | 168
WBC count 9000 cells/cm3 | 168
C-reactive protein 200 mg/L | 168
IV Tazosin | 168
complained of headache | 168
complained of neck pain | 168
Glasgow Coma Scale dropped | 216
pupils reactive | 216
neck stiffness | 216
positive Kernig’s sign | 216
positive Brudzenski sign | 216
blood sepsis parameter increased | 216
WBC count 14000 cells/cm3 | 216
CRP >200 mg/L | 216
blood culture preliminary report | 216
E. meningoseptica | 216
Carbapenam Resistance Enterobacteriaceae | 216
intubated | 216
septic shock | 216
meningitis | 216
transferred to neurocritical care unit | 216
IV Meropenem | 216
IV Ciprofloxacin | 216
lumbar puncture | 216
CSF results | 216
total WBC increased | 216
polymorphs cell | 216
RBC nil | 216
glucose 2.2 mmol/L | 216
protein 0.57 g/L | 216
positive culture E. meningoseptica | 216
CRE | 216
diagnosed with bacteremia | 216
diagnosed with meningitis | 216
did not improve neurologically | 216
contrast-enhanced CT brain | 216
short-segment superior sagittal sinus thrombosis | 216
SC clexane | 216
tracheal aspirate culture | 312
grew Acinetobacter baumannii | 312
XDR | 312
IV Polymyxin B | 312
completed IV Polymyxin | 504
completed IV Meropenem | 504
completed IV Ciprofloxacin | 504
T. Levofloxacin | 504
extubated | 408
repeated CTV Brain | 504
venous sinus thrombosis resolving | 504
septic parameter normalized | 504
WBC 7000 cells/cm3 | 504
CRP negative | 504
discharged | 504
follow-up clinic | 504
full neurological recovery | 504