26 years old | 0
female | 0
sickle cell trait | 0
altered mental status | 0
recovered from viral illness | -336
shortness of breath | -168
diffuse pain | -168
unresponsive | 0
pulseless electrical activity arrest | 0
return of spontaneous circulation | 0
transferred to higher acuity facility | 0
multisystem organ failure | 0
acute respiratory distress syndrome | 0
acute renal failure | 0
bone marrow failure | 0
low hemoglobin | 0
low platelets | 0
high leukocytes | 0
MRI of brain | 24
diffuse scattered areas of restricted diffusion | 24
transcranial Doppler | 168
increased velocity of left middle cerebral artery | 168
increased pulsatility indices | 168
echocardiography | 0
global hypokinesis | 0
low left ventricular ejection fraction | 0
schistocytes on peripheral blood smear | 0
started on broad-spectrum antimicrobials | 0
started on plasma exchange | 0
started on methylprednisolone | 0
hemoglobin electrophoresis | 120
HbSC disease | 120
ADAMSTS activity | 120
peripheral blood smear | 120
schistocytes | 120
neutrophil-containing morulae | 120
bone marrow biopsy | 120
normocellular marrow | 120
trophozoites in RBCs | 120
started on clindamycin | 120
started on atovaquone | 120
started on doxycycline | 120
anaplasmosis-induced sickle cell crisis | 120
Babesia coinfection | 120
PCR for anaplasmosis | 120
PCR for babesiosis | 120
treatment for babesiosis stopped | 120
neurologic examination | 144
decerebrate posturing | 144
not following commands | 144
started on eculizumab | 264
worsening renal function | 264
suspected atypical hemolytic uremic syndrome | 264
transferred out of intensive care | 744
discharged to skilled nursing facility | 1008
tracheostomy | 1008
percutaneous endoscopic gastrostomy | 1008