28 years old | 0 | 0 
female | 0 | 0 
8 weeks pregnant | 0 | 0 
acute severe asthma | -10 | 0 
short non-infective prodrome | -10 | 0 
hypoxic cardiac arrest | -10 | 0 
ventricular fibrillation | -10 | 0 
resuscitation to sinus tachycardia | -10 | -10 
endotracheal intubation | -10 | -10 
therapeutically cooled to 33°C | 0 | 24 
salbutamol | 0 | 48 
ipratropium | 0 | 48 
aminophylline | 0 | 48 
hydrocortisone | 0 | 48 
magnesium | 0 | 48 
ketamine | 0 | 48 
inhalation anesthesia with 1 MAC isoflurane | 0 | 48 
severe hypercapnic acidosis | 0 | 24 
neuromuscular blockade | 0 | 24 
generalised status myoclonus | 48 | 240 
absent motor response to painful stimulus | 96 | 240 
preserved pupillary reflexes | 96 | 240 
preserved corneal reflexes | 96 | 240 
preserved cough reflexes | 96 | 240 
preserved gag reflexes | 96 | 240 
spontaneously breathing | 96 | 240 
severe GSM | 96 | 240 
refractory to three antiepileptic medications | 96 | 240 
generalised periodic discharges | 96 | 240 
no discernable background rhythm | 96 | 240 
reversible causes of coma eliminated | 96 | 240 
plasma neuron-specific enolase | 240 | 240 
somatosensory-evoked potential | 240 | 240 
brain magnetic resonance imaging | 240 | 240 
bilateral basal ganglia and frontoparietal cortex infarction | 240 | 240 
severe hypoxic encephalopathy | 240 | 240 
extubated | 240 | 240 
died | 264 | 264 
comfort measures | 240 | 264