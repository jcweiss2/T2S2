80 years old | 0
female | 0
hypertension | 0
asthma | 0
hypothyroidism | 0
laceration to the right lower extremity | -96
boating on a freshwater river | -96
remained in wet pants for multiple hours | -96
increased edema | -48
erythema | -48
pain to the affected leg | -48
bullae developed | -24
drained the lesions | -24
expression of clear fluid | -24
sloughing of the epidermis | -24
admitted to the hospital | 0
erythematous and edematous right lower extremity | 0
ecchymosis | 0
superficial erosions | 0
clear drainage | 0
WBC count of 7400 cells/mcL | 0
50% band neutrophils | 0
elevated lactate of 3.0 mmol/L | 0
blood cultures obtained | 0
1 g ceftriaxone IVPB given | 0
cellulitis of the right lower extremity | 0
bandemia | 0
lactic acidosis | 0
acute hypoxic respiratory failure | 12
altered mentation | 12
hypotension | 12
transferred to the Intensive Care Unit | 12
severe sepsis | 12
cefepime and metronidazole started | 12
returned to the medical floor | 24
blood cultures grew Plesiomonas shigelloides | 48
antimicrobial susceptibilities displayed | 48
sensitive to ceftriaxone | 48
sensitive to ciprofloxacin | 48
sensitive to ertapenem | 48
sensitive to meropenem | 48
ciprofloxacin added to treatment regimen | 48
changes in stool | 120
ciprofloxacin discontinued | 120
concerns for Clostridium difficile infection | 120
general surgery consulted | 120
wound debridement | 168
condition continued to improve | 168
discharged to inpatient rehab | 336
10-day course of 500 mg metronidazole TID | 336
one month course of 2 g ceftriaxone IVPB | 336
discharged from inpatient rehab | 504
follow up with family doctor | 504