39 years old | 0
female | 0
admitted for elective cardiac surgery | -24
cadaveric renal transplant | -87600
renal transplant failed | -70080
chronic end-stage renal disease | 0
chronic renal dialysis | 0
chronic vesicoureteral reflux | 0
secondary hyperparathyroidism | 0
secondary arterial hypertension | 0
chronic anemia | 0
iron supplements | 0
atorvastatin | 0
aspirin | 0
amlodipine | 0
erythropoietin | 0
vitamin D supplements | 0
worsening dyspnea over 6-12 months | -720
malnourished | 0
cachectic | 0
faint diastolic murmur | 0
bibasal lung crepitations | 0
severe mitral stenosis | 0
severely calcified mitral annulus | 0
sub-valvular apparatus | 0
mean gradient of 10 mmHg | 0
mitral valve area of 0.8 cm2 | 0
severe tricuspid regurgitation | 0
preserved biventricular ejection fraction | 0
no flow-limiting coronary lesions | 0
urea 111 mg/dL | 0
creatinine 4.7 mg/dL | 0
phosphorus 10 mg/dL | 0
calcium 8.6 mg/dL | 0
parathormone hormone (PTH) 725 pg/mL | 0
underwent mitral valve replacement | 0
mechanical prosthesis | 0
tricuspid valve repair | 0
annuloplasty ring | 0
intraoperative severe calcification | 0
extensive tissue debridement | 0
decalcification | 0
transfusion of red blood cells | 0
transfusion of plasma concentrates | 0
transfusion of platelets | 0
transfusion of fibrinogen | 0
significant coagulopathy | 0
bleeding | 0
admitted to intensive care unit | 0
more blood transfusions | 0
continuous renal replacement therapy | 0
metabolic optimization | 0
fluid off-loading | 0
extubated | 48
warfarin started | 72
chest drains removed | 72
transferred to floor | 96
hemodynamically stable | 96
developed skin lesions | 168
multiple ulcerative lesions inner thighs | 168
ulcerative lesions calves | 168
painful ulcers | 168
necrotic base | 168
erythematous borders | 168
ured 10x7 cm lesion | 168
necrotic ulcers fingertips | 168
tissue biopsies | 168
calcium deposition small vessels | 168
necrotic changes | 168
histopathological diagnosis calciphylaxis | 168
conservative wound care | 168
enzymatic debridement | 168
collagenase-based ointment | 168
frequent dressings | 168
empirical prophylactic antibiotics | 168
repeated swab cultures | 168
negative bacterial growth | 168
normal inflammatory markers | 168
warfarin continued | 168
transferred to local hospital | 456
clinical stability | 456
deterioration | 1080
worsening wound infection | 1080
sepsis | 1080
deceased | 1080
