49 years old | 0
    man | 0
    Guangxi, China | 0
    cough | -5040
    fever | -5040
    emaciation | -5040
    mass on the left side of his neck | -5040
    ceftazidime | -5040
    fever resolved | -5040
    mass on the neck had grown | -5040
    no history of previous medical illness | 0
    no history of medication | 0
    body temperature of 38°C | 0
    palpable masses on the left side of his neck | 0
    palpable mass below the right side of his chin | 0
    larger mass was 8 cm in diameter | 0
    masses were inflamed | 0
    masses were sensitive to touch | 0
    moist rales in the upper lobe of the left lung | 0
    white blood cell count of 14,200 cells/µL | 0
    neutrophil count of 12,200 cells/µL | 0
    lymphocyte count of 1.39 cells/µL | 0
    platelet count of 167,000/µL | 0
    hemoglobin of 124 g/L | 0
    C-reactive protein level of 167.04 mg/L | 0
    erythrocyte sedimentation rate of 70 mm/h | 0
    procalcitonin of 0.61 ng/mL | 0
    total CD3+ T-lymphocyte count of 1,137 cells/L | 0
    total CD4+ T-lymphocyte count of 470 cells/L | 0
    total CD8+ T-lymphocyte count of 620 cells/L | 0
    liver function test results normal | 0
    kidney function test results normal | 0
    total immunoglobulin level within normal limit | 0
    galactomannan index of 0.35 | 0
    HIV negative | 0
    computed tomography of the neck | 0
    mixed-density lesions on the left side of the neck | 0
    mixed-density lesions in the right submental area | 0
    started on ceftazidime | 0
    started on levofloxacin | 0
    resection of the neck masses | 0
    pus | 0
    large amount of hemopurulent necrotic material | 0
    pus sample sent for culture | 0
    B. cepacia cultured from the mass on the neck | 168
    B. cepacia cultured from submental pus | 168
    drug sensitivity test results | 168
    sensitive to meropenem | 168
    sensitive to ceftazidime | 168
    sensitive to levofloxacin | 168
    sensitive to cotrimoxazole | 168
    sensitive to minocycline | 168
    continued administration of ceftazidime | 168
    continued administration of levofloxacin | 168
    fever resolved | 168
    masses decreased in size | 168
    productive cough | 336
    CT showed neck masses shrank | 336
    large exudative consolidation shadow in the left upper lobe | 336
    left hilar lymphadenopathy | 336
    bronchofibroscopy | 336
    bronchial nodules in the left upper lobe | 336
    bronchial nodules in the left lower lobe | 336
    obstructing the lumen | 336
    mucosal hyperplasia | 336
    mucosal hypertrophy | 336
    left hilar lymph nodes biopsied | 336
    tracheal nodules biopsied | 336
    samples sent for culture | 336
    TM cultured from bronchial nodule | 336
    TM cultured from left hilar lymph node | 336
    TM cultured from bronchoalveolar lavage fluid | 336
    left hilar lymph node sent for next-generation sequencing | 336
    next-generation sequencing results TM | 336
    diagnosed with disseminated TM infection | 336
    diagnosed with B. cepacia infection | 336
    amphotericin B added as antifungal therapy | 336
    discontinued ceftazidime | 672
    discontinued levofloxacin | 672
    neck mass improved | 672
    cough improved | 672
    febrile again | 1176
    new mass on the right side of the neck | 1176
    chest CT scan | 1176
    significant improvement in the pulmonary lesions | 1176
    CT of the neck | 1176
    abscess in the posterior pharyngeal wall | 1176
    fracture of the 4th cervical vertebra | 1176
    mass on the right side of the neck | 1176
    ceftazidime added as antibacterial treatment | 1176
    levofloxacin added as antibacterial treatment | 1176
    no obvious treatment effect | 1176
    antibiotics switched to meropenem | 1176
    antibiotics switched to cotrimoxazole | 1176
    B. cepacia infection remained uncontrolled | 1176
    acute-onset quadriplegia | 1176
    emergency subtotal resection of the 4th cervical vertebra | 1176
    widening and decompression of the spinal canal | 1176
    transferred to the intensive care unit | 1176
    treated with meropenem | 1176
    treated with tigecycline | 1176
    treated with voriconazole | 1176
    B. cepacia cultured repeatedly from the blood | 1176
    B. cepacia cultured repeatedly from the pus | 1176
    pulmonary lesions improved | 1176
    neck abscess could not be contained | 1176
    abscess disseminated widely to multiple body parts | 1176
    hepatorenal dysfunction | 1848
    cardiac insufficiency | 1848
    hypotension | 1848
    hypoxia | 1848
    repeated immune function test | 1848
    CD3+ T-lymphocyte count of 158 cells/L | 1848
    CD4+ T-lymphocyte count of 48 cells/L | 1848
    CD8+ T-lymphocyte count of 99 cells/L | 1848
    disseminated intravascular coagulation | 2016
    died of B. cepacia sepsis | 2016
    measured the nAIGAs in the peripheral blood | 168
    serum AIGA determined | 168
    high positive titer (11,025 ng/mL) | 168
    antibody titer increased gradually to 50,566 ng/mL | 1344
    positive nAIGA titer | 168
    progressive increase in serum nAIGA titer | 1344
    