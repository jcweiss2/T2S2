66 years old | 0
female | 0
admitted to the hospital | 0
type II diabetes mellitus | 0
chronic obstructive pulmonary disease | 0
severe pulmonary hypertension | 0
schizophrenia | 0
fatigue | 0
shortness of breath | 0
denies fevers | 0
denies rigors | 0
denies changes in quality or color of sputum | 0
denies chest pain | 0
denies palpitations | 0
dizziness | 0
black stool | 0
no history of acute epigastric pain | 0
no lower abdominal pain | 0
no rectal bleeding | 0
no recent bowel habits changes | 0
confused | 0
ill-looking | 0
oxygen saturation 81% on room air | 0
oxygen saturation 95% on 4 L/min oxygen | 0
afebrile | 0
blood pressure 110/60 mm Hg | 0
pulse rate 100 beats/min | 0
reduced breathing sounds over both lung fields | 0
crackles | 0
scattered wheezes | 0
nasopharyngeal swab for SARS-CoV-2 positive | 0
commenced on dexamethasone | 0
commenced on remdesivir | 0
passed a large amount of melena | 24
became hypotensive | 24
responded to 1 L of intravenous fluids bolus | 24
transferred to the intensive care unit | 24
gastroenterology services recommended pantoprazole | 24
gastroenterology services recommended esophagogastroscopy | 24
esophagogastroscopy revealed bleeding duodenal ulcer | 48
controlled by epinephrine injection and bipolar cauterization | 48
surgical consultation recommended an emergent laparotomy | 72
operative intervention performed | 96
perforated sigmoid diverticulitis | 96
Hartmann’s procedure performed | 96
remained on vasopressors support | 96
repeat blood cultures grew C. tertium | 120
switched to intravenous meropenem and metronidazole | 120
histology of the resected colon biopsy confirmed perforated diverticulitis | 120
no evidence of neoplasia | 120
continued on parenteral meropenem and metronidazole | 168
serial blood cultures confirmed clearance of C. tertium bacteremia | 240
challenging postoperative course | 240
difficult weaning from the mechanical ventilator | 240
intensive care unit-acquired weakness | 240
transition into tracheostomy | 240
transferred into a long-term acute care facility | 336
discharged on oral metronidazole and amoxicillin-clavulanate | 336
high-grade fever | 72
hypotensive | 72
tachycardic | 72
requiring vasopressors support | 72
inspiratory crackles over the left lower lung zone | 72
vague generalized abdominal tenderness | 72
blood cultures obtained | 72
C. tertium isolated | 96
commenced on empiric broad-spectrum antibiotics | 96
CT of the abdomen performed | 96
extensive free intraperitoneal gas | 96
thickened distal sigmoid colon wall | 96
adjacent free fluids | 96
concerning for colonic perforation | 96
C. tertium bacteremia | 96
septic shock | 96
COVID-19 | 0
perforated colonic diverticular disease | 96
bacterial translocation | 96
gastrointestinal tract perforation | 96
corticosteroids | 0
poorly controlled diabetes | 0
immunosuppressive status | 0
persistence of Clostridial growth | 168
prolonged course of targeted antibiotics | 168
C. tertium species | 96
aerotolerant | 0
slowly growing | 0
traditional culturing methods | 0
underdiagnoses | 0
inaccurate identification | 0
inappropriate antibiotics selection | 0
modern bacterial identification diagnostics | 96
direct MALDI-TOF mass spectrometry | 96
rapid isolation | 96
accurate isolation | 96
targeted antibiotic therapy | 120
susceptibility results | 120
resistance to antibiotics | 120
third and fourth generation cephalosporins | 0
molecular biology techniques | 0
16S rRNA sequencing | 0
pathogenesis | 0
non-exotoxin-producing | 0
neutropenia | 0
gastrointestinal mucosal injury | 0
bacterial translocation | 0
end-stage liver disease | 0
recent use of broad-spectrum antibiotics | 0
intestinal colonization | 0
chemotherapy | 0
innate immune response | 0
intestinal mucosal injury | 0
translocation | 0
systemic circulation | 0
aggressive treatment | 120
targeted antibiotic therapy | 120
non-highly virulent organism | 0
low direct mortality rate | 0
one-month mortality rate | 0
advanced stage of malignancies | 0
associated medical comorbidities | 0
underlying poor baseline status | 0
limited data | 0
standard duration of directed antibiotic therapy | 0
prolonged course of targeted antibiotics | 168
persistence of Clostridial growth | 168
immunosuppressive status | 168
poorly controlled diabetes | 0
corticosteroids use | 0