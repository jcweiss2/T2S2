24 years old | 0
female | 0
admitted to the hospital | 0
atraumatic right groin pain | -720
nightly pain | -168
sweating | -168
no prior history of hip pathology | 0
otherwise healthy | 0
played contact sports | 0
took no medications | 0
no history of intravenous drug use | 0
no smoking | 0
no immune suppression | 0
afebrile | 0
vital signs stable | 0
antalgic gait | 0
preferred leg in slight flexion and external rotation | 0
internal rotation of hip tender and restricted | 0
normal serum white cell count | 0
elevated C-reactive protein levels | 0
CT scan of right hip suggestive of pyomyositis | 0
no evidence of osseous destruction | 0
MRI of pelvis revealed multiple complex fluid collections | 0
abscess within obturator internus, obturator externus, and pectineus muscles | 0
small right hip joint effusion | 0
synovial enhancement suggestive of intra-articular septic process | 0
antibiotic therapy withheld | 0
intraoperative synovial samples collected for culture | 0
purulence and inflamed synovia identified | 0
synovectomy performed | 0
capsulotomy extended medially to psoas muscle | 0
psoas muscle released | 0
debridement continued medially and posteriorly | 0
obturator membrane encountered | 0
obturator membrane pierced with blunt switching stick | 0
intrapelvic space accessed and debrided | 0
hip joint copiously irrigated | 0
capsulotomy left open | 0
no drains inserted | 0
postoperative weight bearing | 24
abduction brace | 24
afebrile and stable | 24
no need for pressors or ICU stay | 24
CRP level 188 | 24
intraoperative cultures no pathogen | 24
cefazolin IV for 3 weeks | 24
discharged home on postoperative day 4 | 96
residual surgical pain at 3-week follow-up | 504
brace discontinued | 504
referred to physiotherapy | 504
nontender and 4/5 weakness of right hip flexor at 6-week follow-up | 1008
good right hip range of motion | 1008
CRP levels normalized | 1008
completely asymptomatic at 6-month follow-up | 2016
regained 5/5 strength of right hip flexors | 2016
internal rotation improved | 2016
CRP levels remained normal | 2016
scored 88.6/100 on International Hip Outcome Tool questionnaire | 2016
recurrence of abscess at 10 months | 7440
presented to emergency department with atraumatic right buttock pain | 7440
antalgic gait | 7440
limited right hip range of motion | 7440
CRP level 70 | 7440
MRI showed recurrence of intrapelvic abscess | 7440
open irrigation and debridement | 7440