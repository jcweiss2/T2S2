63 years old | 0
female | 0
hypertension | 0
hyperlipidemia | 0
type II diabetes mellitus | 0
HbA1c 6.5% | 0
admitted to the hospital | 0
right neck pain | -168
subjective fevers | -168
rapid strep test | -72
CT head | -72
CT neck | -72
CT temporal bones | -72
amoxicillin-clavulanic acid | -72
recurrent fevers | -24
pulsatile right sided temporal headache | -24
odynophagia | -24
difficulty breathing | 0
stridor | 0
changes in voice | 0
neck stiffness | 0
photophobia | 0
phonophobia | 0
focal neurologic deficits | 0
night sweats | 0
weight loss | 0
catheters | 0
trauma | 0
lesions to the neck | 0
upper respiratory tract infection | 0
dental infection | 0
mouth sores | 0
traveled to the Philippines | -720
sick contacts | 0
animal exposures | 0
outdoor activities | 0
registered nurse | 0
alcohol | 0
cigarette smoking | 0
illicit drug use | 0
febrile | 0
hypotensive | 0
respiratory distress | 0
tenderness | 0
induration | 0
firm nodule | 0
bulging of the right lateral pharyngeal wall | 0
neutrophil-predominant leukocytosis | 0
blood cultures | 0
Gram-negative bacilli | 0
CT neck with and without IV contrast | 0
thrombosis | 0
retromandibular vein | 0
fluid in the retropharyngeal space | 0
inflammatory stranding | 0
suppurative lymphadenopathy | 0
ultrasound of the right neck | 0
complete occlusion of the right internal jugular vein | 0
cystic structures | 0
reactive lymphadenopathy | 0
CT head | 0
intracranial metastases | 0
fluid resuscitation | 0
piperacillin-tazobactam | 0
Fusobacterium species | 0
anaerobic organisms | 0
meropenem | 24
extended-spectrum β-lactamases | 24
rivaroxaban | 48
persistent fevers | 48
increased swelling | 48
increased work of breathing | 48
CT imaging of the neck | 72
septic emboli | 72
ampicillin-sulbactam | 72
discharged | 168
oral amoxicillin-clavulanic acid | 168
rivaroxaban | 168
follow-up | 336
follow-up | 840
Klebsiella pneumoniae | 0
string test | 0
whole genome sequencing | 0
comparative genomic analysis | 0
virulence factors | 0
antimicrobial resistance genes | 0
genomic characterization | 0
phylogenetic relationships | 0
MLSTcheck tool | 0
Sequence Type (ST)-65 | 0
hypervirulent strain | 0
capsular serotype K2 | 0
iron acquisition systems | 0
aerobactin | 0
salmochelin | 0
rmpA | 0
mucoid phenotype | 0
genetic markers | 0
hypervirulence | 0
hyperviscosity | 0
septic metastases | 0
drainable abscesses | 0
antibiotic therapy | 0
prognostic information | 0
Lemierre’s syndrome | 0
Klebsiella-associated Lemierre’s syndrome | 0
diabetics | 0
septic intracranial metastases | 0
biomarkers | 0
clinical decision-making | 0
virulent phenotypes | 0
genotypes | 0