55 years old | 0
female | 0
height 151cm | 0
weight 61kg | 0
return from the Philippines | -168
presentation at regional hospital | 0
fever | -168
cough | -168
lethargy | -168
myalgia | -168
febrile | 0
temperature 42°C | 0
mild asthma | 0
sleep apnoea | 0
Type 2 diabetes mellitus | 0
oral hypoglycaemics prescribed | 0
non-smoker | 0
nasopharyngeal swabs SARS CoV-2 PCR positive | 0
CT chest scan bilateral air-space infiltrates | 0
ground glass density | 0
COVID-19 diagnosis | 0
transfer to quaternary hospital | 0
respiratory deterioration | -96
ICU transfer | -96
semi-elective intubation | -96
lung-protective ventilation initiation | -96
septic shock | -96
multi-organ dysfunction | -96
oxygenation deterioration | -120
metabolic derangements | -120
high PEEP | -120
deep sedation | -120
paralysis with cisatracurium | -120
FiO2 90% | -240
PEEP 20 cmH2O | -240
P/F ratio 62 | -240
echocardiography normal LV function | -240
mild RV dysfunction | -240
mild RV dilatation | -240
mild to moderate tricuspid regurgitation | -240
RESP score 1 | -240
VV ECMO initiation | -240
femoral-femoral cannulation | -240
tidal volume 2ml/kg | -240
PEEP 10 cmH2O | -240
respiratory rate 10 bpm | -240
TOE thrombus in right atrium | -240
haemodynamic improvement | -240
RV function improvement | -240
ECMO dependency | -336
loss of tidal volumes | -336
HRCT minimal recruitable lung | -480
lung consolidation | -480
lung collapse | -480
HRCT bilateral consolidation | -816
ground glass changes | -816
transition to pressure support ventilation | -816
airway bleeding | -336
complete proximal airway occlusion | -336
anticoagulation with heparin | -336
coagulation profile mild heparinization | -336
APTT 1.5x normal | -336
nebulised tranexamic acid | -336
heparin cessation | -336
bronchoscopic thrombus removal | -336
fibrous tissue strands in bronchi | -336
cryotherapy | -336
tranexamic acid injection | -336
epinephrine injection | -336
bronchial cell cytology | -336
ongoing oozing right lower lobe | -336
lung isolation | -336
double-lumen endotracheal tube | -336
reduced bleeding | -408
bronchial mucosa sloughing | -408
argon plasma coagulation | -408
fibrin debris removal | -408
lung recruitment | -408
prone ventilation initiation | -432
CXR improved lung aeration | -432
prone ventilation tolerated | -432
elevated D-dimer | -888
haemolysis evidence | -936
oxygenator change | -936
hypercalcaemia | -768
calcium 3.26 mmol/L | -768
parathyroid hormone normal | -768
serum phosphate normal | -768
1,25-dihydroxy vitamin D normal | -768
thyroid hormone normal | -768
pamidronate disodium | -792
calcitonin | -792
calcium normalization | -1080
ECMO weaning trials | -960
stable gas exchange | -984
ECMO decannulation | -1224
femoral vein repair | -1224
post-ECMO improvement | -1272
surgical tracheostomy | -1320
ventilator weaning | -1344
phonation via tracheostomy | -1344
neurological improvement | -1440
obeying commands | -1440
family interaction | -1440
