75 years old | 0
female | 0
hypertension | -8760
hyperlipidemia | -8760
referred to clinic for evaluation of leukocytosis | -8760
white blood cell count 16.3 × 10^9/L | -8760
weight loss of 6 lbs in 1 year | -8760
fatigue for the past 3 months | -2160
no fever | -2160
no chills | -2160
no night sweats | -2160
WBC count 461 × 10^9/L | 0
hemoglobin 6.9 gm/dL | 0
admitted to the hospital | 0
flow cytometry peripheral blood T-PLL | 0
hyperleukocytosis | 0
bone marrow biopsy | 0
90% atypical T-cells | 0
flow cytometric analysis aspirate T-PLL | 0
cytogenetic analysis inversion chromosome 14 | 0
trisomy 8 | 0
karyotype analysis 47, XX, add(4)(q35), +8, inv(14)(q11.2q32), add(20)(P13) | 0
gross cytomorphologic review marked lymphocytosis | 0
prominent cytologic atypia | 0
T-cell percent 85% | 0
clonal T-cell gamma receptor rearrangement | 0
computed tomography chest, abdomen, pelvis | 0
moderate splenomegaly | 0
no masses | 0
no lymphadenopathy | 0
next-generation sequencing JAK1 p(His374Tyr) | 0
no microsatellite instability | 0
low tumor mutation burden 3.1 mutations/MB | 0
diagnosed T-PLL | 0
treated with alemtuzumab | 0
3 cycles of 3-mg alemtuzumab subcutaneously | 0
WBC persistently elevated | 0
alemtuzumab dose increased to 10 mg | 0
pentostatin added | 0
10 cycles of 10-mg alemtuzumab | 0
2 cycles of pentostatin 4 mg/m² | 0
WBC >500 × 10^9/L | 0
alemtuzumab increased to 30 mg | 0
cycle 13 alemtuzumab | 0
cycle 7 pentostatin | 0
WBC trend down to 300 × 10^9/L | 0
18 cycles alemtuzumab | 0
7 cycles pentostatin | 0
completed chemotherapy | 0
postchemotherapy CBC WBC 2.7 × 10^9/L | 0
Hgb 11 gm/dL | 0
flow cytometry postchemotherapy monoclonal TCR gamma rearrangement | 0
no significant circulating blasts | 0
no abnormal lymphoid population | 0
no abnormal myeloid population | 0
asymptomatic | 0
presented to emergency department with rash | 5040
facial swelling | 5040
sore throat | 5040
dysphagia | 5040
conjunctivitis | 5040
rash entire body | 5040
trunk involvement | 5040
extremities involvement | 5040
face involvement | 5040
edema bilateral lower extremities | 5040
afebrile | 5040
WBC 41 × 10^9/L | 5040
absolute lymphocyte count 28 × 10^9/L | 5040
cytomegalovirus DNA PCR negative | 5040
T-PLL relapse confirmed | 5040
flow cytometry analysis relapse | 5040
peripheral blood smear atypical lymphocytes | 5040
uric acid 13.70 mg/dL | 5040
creatinine 2.52 mg/dL | 5040
tumor lysis syndrome | 5040
rasburicase given | 5040
rash worsened | 5040
anasarca developed | 5040
edema progressed | 5040
dyspnea developed | 5040
partially relieved with steroids | 5040
epinephrine | 5040
antihistamines | 5040
white counts continued to rise | 5040
restarted alemtuzumab | 5040
restarted pentostatin | 5040
CMV prophylaxis valganciclovir | 5040
PCP prophylaxis Bactrim | 5040
peripheral blood smear same morphology | 5040
flow cytometry same CD4/CD3+/CD7+ T-cells | 5040
skin biopsy admission time | 5040
atypical perivascular lymphocytic infiltrate | 5040
CD7+ | 5040
CD2+ | 5040
CD3+ | 5040
CD4+ | 5040
CD5+ | 5040
CD8− | 5040
CD30− | 5040
CD56− | 5040
computed tomography neck lymphadenopathy mediastinal | 5040
cervical chains lymphadenopathy | 5040
white counts began to drop | 5040
respiratory status worsened | 5040
evaluation otolaryngologists airway edema lymphocytic infiltration | 5040
tachypneic | 5040
oxygen saturation 82% | 5040
anasarca worsened | 5040
profound hypotension | 5040
shock | 5040
racemic epinephrine | 5040
Benadryl | 5040
methylprednisolone | 5040
respiratory status did not improve | 5040
emergently intubated | 5040
ventilated | 5040
intravenous pressor support | 5040
white cell counts trended up to 50 × 10^9/L | 5040
lactate increased 12 mmol/L | 5040
creatinine 3.28 mg/dL | 5040
infectious workup sepsis suspected | 5040
transferred to medical ICU | 5040
passed away | 5040
