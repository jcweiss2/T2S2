78 years old | 0
female | 0
abdominal pain | -672
diagnosed with HCC | -672
hypertension | -672
liver cirrhosis | -672
antibodies for hepatitis C virus | -672
advanced HCC | -672
portal invasion | -672
daughter nodules | -672
computed tomography | -672
lenvatinib initiated | 0
lenvatinib 8 mg/day | 0
proteinuria | -128
lenvatinib interrupted | -128
lenvatinib resumed | -128 + 720
lenvatinib 4 mg/day | -128 + 720
unsteady on feet | -168
vomiting after eating | -168
respiratory distress | -168
urge incontinence | -168
night sweats | -168
dehydration | -168
shock | -168
blood pressure not measurable | -168
heart rate 137 beats/min | -168
respiratory rate 33 breaths/min | -168
body temperature 36.4°C | -168
abdomen soft and nontender | -168
no guarding | -168
white blood cells 15,700/μL | -168
hemoglobin 16.0 g/dL | -168
platelets 216,000/μL | -168
creatinine 2.90 mg/dL | -168
C-reactive protein 18.2 mg/L | -168
free air bubbles in abdomen and pelvis | -168
emergency exploratory laparotomy | -168
peritonitis | -168
purulent exudate | -168
focally necrotic perforation | -168
sigmoid colon perforation | -168
Hartmann's procedure | -168
sigmoid resection | -168
end colostomy | -168
transferred to intensive care unit | -168
died 48 h after surgery | 48
sepsis | 48
macroscopic examination | 48
histopathological examination | 48
infiltration of neutrophils | 48
hemorrhage | 48
mitotic arrest | 48
mitotic spindles | 48
lenvatinib-related bowel perforation | 48
apoptosis | 48
crypt hyperplasia | 48