14 years old | 0
male | 0
Joubert syndrome | -2160
chronic renal failure | -2160
peritoneal dialysis | -2160
vomiting | -168
intolerance to food intake | -168
hyponatremia | -168
hypopotassemia | -168
hospitalized | -168
supplementation treatment | -168
blood cultures | -168
urine cultures | -168
peritoneal fluid cultures | -168
IV antibiotherapy with tazobactam-ampicillin | -168
febrile episodes | -168
Candida spp. in peritoneal culture | -144
liposomal amphotericin B | -144
peritoneal dialysis catheter removal | -144
anuric | -144
volume overload | -144
intermittent hemodialysis | -144
abdominal ultrasound | -120
complicated, lobulated, fluid-filled cystic lesions | -120
pseudocyst in the pancreatic loge | -120
multiple cortical cysts in both kidneys | -120
abdominal CT scan | -96
large cystic lesions in the anterior abdominal region | -96
loculated fluid collections in the peripancreatic area | -96
surgery planned | -96
cyst on the anterior abdominal wall | -72
cyst rupture | -72
serohemorrhagic fluid aspirated | -72
cardiac arrest | -72
erythrocyte suspension transfused | -72
fluid support provided | -72
adrenaline and noradrenaline infusions started | -72
transferred to intensive care unit | -72
hypotensive state | -72
bilateral dilated pupils | -72
absent light reflex | -72
capillary refill time 6-7 seconds | -72
arterial blood gas pH 7.15 | -72
PaCO2 41.8 mmHg | -72
PaO2 82.8 mmHg | -72
base excess -13.2 mmol/L | -72
HCO3 14 mmol/L | -72
lactate 16 mmol/L | -72
BUN 87 mg/dL | -72
creatinine 2.7 mg/dL | -72
mechanical ventilation | -72
saline solution given | -72
dopamine, dobutamine, adrenaline, and noradrenaline infusions started | -72
erythrocyte suspension infused | -72
thrombocyte suspension transfused | -72
prothrombin time 24 seconds | -72
international normalized ratio 2.16 | -72
IV fresh frozen plasma administered | -72
combined antibiotherapy with meropenem, vancomycin, and amikacin | -72
metronidazole added | -72
single dose of IV steroid administered | -72
3-F catheter inserted into the femoral vein | -72
cardiac output monitored using PiCCO pulse contour monitor | -72
cardiac index 6.5 L/minute | -72
systemic vascular resistance index 338 dynes/second/cm5/m2 | -72
global end-diastolic index 780 mL/m2 | -72
extravascular lung water index 15 mL/kg | -72
systolic blood pressure 67 mmHg | -72
diastolic blood pressure 32 mmHg | -72
mean arterial blood pressure 46 mmHg | -72
pulse rate 106/minute | -72
TP administered as an IV bolus dose | 0
increase in blood pressure | 0.17
SBP 94 mmHg | 0.17
DBP 45 mmHg | 0.17
MAP 60 mmHg | 0.17
TP treatment changed to infusion | 0.17
noradrenaline dose reduced | 0.17
decrease in cardiac index and heart rate | 0.17
increase in SVRI, GEDI, and EVLWI | 0.17
continuous venovenous hemodiafiltration initiated | 1
ultrafiltrate aspirated | 12
control BUN and creatinine values | 12
decrease in GEDI and ELWI values | 12
ischemic manifestations on the right big toe | 9
TP infusion discontinued | 9
SBP 69 mmHg | 10
DBP 46 mmHg | 10
MAP 54 mmHg | 10
cardiac arrest | 12
cardiopulmonary resuscitation applied | 12
patient lost | 12