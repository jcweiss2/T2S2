60 years old | 0
female | 0
admitted to the hospital | 0
diabetes mellitus | -8760
chronic renal failure | -8760
severe pain in upper lip | -96
bullous lesion in upper lip | -96
cellulitis in upper lip | -96
no trauma history | -96
zoster infection suspected | 0
antiviral treatment initiated | 0
non-adherence to diabetes medication | -96
serum glucose level of 346 mg/dL | 0
hemoglobin A1c of 7.8% | 0
white blood cell count of 12,000/μL | 0
C-reactive protein level of 93.7 mg/L | 0
chest pain | 12
electrocardiography | 12
cardiac enzyme measurements | 12
NSTEMI diagnosed | 12
transferred to intensive care unit | 12
transferred to department of internal medicine | 12
high fever | 12
hypotension | 12
mental status deteriorated to stupor | 12
general condition worsened | 12
swelling and inflammation of upper lip increased | 12
ulcerative lesion on oral mucosa of upper lip | 12
foul odor with purulent discharge | 12
white blood cell count of 23,000/μL | 12
C-reactive protein level of 385.8 mg/L | 12
septic shock | 12
coronary angiography | 24
3-vessel disease | 24
severe stenosis | 24
intravenous broad-spectrum antibiotics initiated | 24
boosters and adjunctive treatment measures commenced | 24
upper lip gangrene and necrosis progressed | 48
contrast-enhanced facial computed tomography | 48
diffuse gaseous necrosis and cutaneous fistula | 48
chest CT | 48
abscess-like lung nodule in right upper lobe | 48
Laboratory Risk Indicator for Necrotizing Fasciitis score of 10 | 48
septic shock due to upper lip NF | 48
surgical intervention planned | 48
debridement under general anesthesia | 48
full-layer necrosis of upper lip | 48
K. pneumoniae confirmed in blood and pus cultures | 120
antibiotic regimen consisting of ceftriaxone and metronidazole | 120
serial debridement | 120
follow-up pus culture confirmed K. pneumoniae and MRSA | 312
full-layer skin and soft tissue defect with scar contracture | 312
discharged | 1200
scar release and Abbe flap coverage | 2160
Abbe flap surgery | 2160
flap detachment | 2208
flap division | 2376
follow-up revealed favorable correction of upper lip drooling | 2376