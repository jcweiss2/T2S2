42 years old | 0
male | 0
referred to emergency department | 0
testicular pain | -192
testicular pain migrated into abdomen | -192
testicular pain migrated into back | -192
testicular pain migrated into chest | -192
fever | -48
denied respiratory symptoms | 0
diffuse abdominal tenderness | 0
CT abdomen captured lung bases | 0
pulmonary ground-glass opacification | 0
consolidation consistent with pneumonia | 0
possible colitis | 0
notified COVID-19-positive status | 48
attended biotechnology conference | -336
COVID-19-impacted area | -336
healthcare workers accidental exposure to SARS-CoV-2 | 0
