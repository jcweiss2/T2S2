29 years old | 0
woman | 0
presented for inpatient continuous epidural infusion | 0
worsening CRPS of the left upper extremity | 0
sports-related injury to left shoulder | -2160
over a dozen surgical revisions | -2160
recurrent shoulder infections | -2160
prolonged shoulder infections | -2160
isolated microorganisms | -2160
Pseudomonas aeruginosa | -2160
Sphingomonas paucimobilis | -2160
Candida colliculosa | -2160
Staphylococcus aureus | -2160
left shoulder tendon release | -720
revision performed | -720
development of CRPS | -720
severe pain | 0
allodynia | 0
edema | 0
muscle spasms | 0
temperature changes of LUE | 0
EMG evaluation | 0
brachial plexus injury | 0
past medical history of asthma | -1752
selective IgG3 deficiency diagnosed | -1752
recurrent joint infections | -1752
CRPS symptoms refractory to oral medical management | 0
opioids | 0
antidepressants | 0
antispasmodics | 0
significant symptom relief with left stellate ganglion blockade | 0
favorable response to sympathectomy | 0
2 prior admissions for continuous cervical epidural infusions | 0
decreased pain | 0
improved participation with physical therapy | 0
reduction in oral opioid requirements | 0
placement of left C6–C7 interlaminar epidural catheter | 0
fluoroscopic guidance | 0
transferred to PACU | 0
preprocedure labs normal | 0
complete blood count | 0
complete metabolic panel | 0
creatinine phosphokinase | 0
history of selective IgG subclass deficiency | 0
atypical infections in the past | 0
received antibiotic prophylaxis | 0
intravenous vancomycin | -1
ruled out for intrathecal placement | 0
ruled out for intravascular placement | 0
epidural infusion started | 0
0.25% bupivacaine | 0
hydromorphone 10 mcg per mL | 0
clonidine 1 mcg per mL | 0
continuous rate of 4 mL per hour | 0
oral home medications continued | 0
methadone 10 mg twice a day | 0
hydromorphone 4 to 8 mg as needed | 0
diazepam 10 mg 4 times a day | 0
baclofen 20 mg 4 times a day | 0
amitriptyline 100 mg once a day | 0
tolerated therapy well | 0
decrease in pain from 9/10 to 7/10 on VAS | 0
less muscle spasms | 0
continuous infusion increased to 6 mL per hour | 24
demand dose of 2 mL every 15 minutes started | 24
improved sleep | 24
further decrease in LUE spasms | 24
further decrease in edema | 24
VAS of 5/10 | 24
prophylactic vancomycin continued | 24
dosed according to trough levels | 24
febrile to 38.1°C | 120
decision to wean infusion rapidly | 120
decision to remove epidural catheter | 120
epidural catheter removed | 126
developed progressive headache | 126
developed neck pain | 126
further increase in temperature to 40.0°C | 126
neurological examination unchanged | 126
epidural site nontender to palpation | 126
no signs of active infection | 126
blood cultures sent | 126
urine cultures sent | 126
chest x-ray negative | 126
increase in white count to 9.7×103/μL | 126
addition of cefepime to vancomycin | 126
abatement of fever | 126
decrease in white count to 5.9×103/μL | 126
underwent MRI of cervical spine | 126
epidural collection from C3 to T1 | 126
compression of left C5 and C6 nerve roots | 126
effacement of thecal sac | 126
no cord deformity | 126
interstitial edema in left paraspinal muscles | 126
transfer to NSICU | 126
suspected epidural abscess | 126
hourly neurological examination | 126
intractable nausea and vomiting | 150
left arm weakness | 150
taken to operating room for decompression | 150
evacuation via C3 to C7 cervical laminectomies | 150
C4–C5 and C5–C6 left foraminotomies | 150
epidural space filled with inflammatory mass | 150
pockets of purulent material | 150
intraoperative cultures positive for P aeruginosa | 150
urine cultures negative | 126
blood cultures negative | 126
vancomycin stopped | 150
cefepime continued | 150
resolution of arm weakness | 150
uneventful postoperative course | 150
discharged home | 174
continued intravenous cefepime | 174
total of 6 weeks | 174
