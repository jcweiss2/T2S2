13 years old | 0
male | 0
admitted to the hospital | 0
uncontrolled bleeding at the operation site | 0
swelling of the right thenar muscle | -168
fall | -168
no improvement for over 5 months | -672
excision of the lesion | -24
marginal excision | -24
no history of bleeding tendency | -24
normal coagulation screening tests | -24
two additional operations | -48
bleeding at the operation site continued | -48
pathologic finding of the mass suggested a diagnosis of malignancy | -24
transferred to our hospital | 0
poor general state | 0
pallor | 0
weakness | 0
bruising at the intravenous site | 0
purpura on the operation site | 0
continuous bleeding | 0
2×2 cm-sized lymph node in the right axillary area | 0
1 cm-sized hepatosplenomegaly | 0
laboratory tests revealed markedly decreased platelet and hemoglobin levels | 0
features suggestive of DIC | 0
white blood cell, 9,900 /µL | 0
hemoglobin, 4.8 g/dL | 0
platelets, 28,000 /µL | 0
prothrombin time, 1.47 international normalized ratio | 0
activated partial thromboplastin time, 45.4 sec | 0
fibrinogen, 87 mg/dL | 0
fibrin/fibrinogen degeneration product, 656.4 µg/mL | 0
D-dimer, 16.17 mg/L | 0
coagulation factors II, VII, IX, fibrinogen, and von willebrand factor were all normal | 0
factors V and VIII were 30% and 40% | 0
18-Fluoro-2-deoxy-D-glucose positron emission tomography scan | 0
hypermetabolic lesions | 0
post-operative inflammation in the right thenar muscle | 0
metastatic lymphadenopathy in the right axillary space | 0
massive bleeding from the operation site and the intravenous access site worsened | 72
gross hematuria developed | 72
pathologic findings of the mass were reported as alveolar rhabdomyosarcoma | 96
immunohistochemical stains of myognesin, desmin, and MyoD | 96
negative resection margin | 96
transferred to the intensive care unit | 96
chemotherapy consisting of vincristine, doxorubicin, and cyclophosphamide | 96
repeated transfusions | 96
synthetic protease inhibitor | 96
substitution of antithrombin-III | 96
massive epistaxis | 240
hematemesis of approximately 1.5 L of blood | 240
transfusions of 4 units of red blood cells | 240
9 units of platelet concentrates | 240
1 unit of fresh frozen plasma | 240
8 units of cryoprecipitate | 240
two times of cauterization | 240
laboratory findings of DIC showed improvement | 336
BM section biopsy | 336
axillary LN biopsy | 336
histologic finding of BM | 336
involvement of rhabdomyosarcoma | 336
total blood transfusions of 311 units | 672
discharged | 672
combination chemotherapy consisting of VAC every 3 weeks | 672
size of right axillary LN decreased | 6048
BM showed disappearance of rhabodyosarcoma | 15120
negative immunostaining for desmin or myogenin | 15120
two rounds of APBSC collections | 15120
nodule in the right forearm | 18972
biopsy revealed it as an alveolar rhabdomyosarcoma | 18972
salvage chemotherapy | 18972
ifosfamide, carboplatin, etoposide | 18972
palliative radiation therapy | 18972
died 5 months later | 21600
disease progression to the liver and the brain | 21600