87 years old | 0
male | 0
admitted to the hospital | 0
fever | 0
general fatigue | 0
denies a history of trauma | 0
denies a history of falls | 0
endoscopic sphincterotomy | -720
choledocholithiasis | -720
percutaneous coronary intervention | -6720
ischemic heart disease | -6720
warfarin potassium | 0
aspirin | 0
antidiabetic | 0
diuretics | 0
heart rate of 115 per minute | 0
blood pressure of 92/61 mmHg | 0
respiratory rate of 13 per minute | 0
body temperature of 36.2°C | 0
Glasgow coma scale was E4, V4, and M4 | 0
height was 164 cm | 0
body weight was 70 kg | 0
body mass index was 26.0 kg/m2 | 0
moderate abdominal pain | 0
tenderness in the epigastrium | 0
hemoglobin of 9.6 g/dL | 0
white blood cell count of 23170/µL | 0
platelet count of 13.6 × 104/µL | 0
total bilirubin of 1.0 mg/dL | 0
alanine transaminase of 843 IU/L | 0
aspartate aminotransferase level of 339 IU/L | 0
lactate dehydrogenase of 1278 U/L | 0
alkaline phosphatase of 947U/L | 0
blood urea nitrogen of 40.5 mg/dL | 0
creatinine of 3.06 mg/dL | 0
prothrombin time of 18.3 seconds | 0
prothrombin time % of 44% | 0
international normalized ratio of 1.6 | 0
activated partial thromboplastin time of 38.4 seconds | 0
procalcitonin of 251 ng/mL | 0
C-reactive protein of 17.4 mg/dL | 0
lactate of 33 mg/dL | 0
brain natriuretic peptide of 1206 ng/mL | 0
α-Fetoprotein of 0.7 ng/mL | 0
sepsis | 0
anemia | 0
liver dysfunction | 0
renal dysfunction | 0
heart failure | 0
coagulopathy | 0
plain abdominal CT | 0
swelling and wall thickening of the gallbladder were not detected | 0
subcapsular high density area of the liver | 0
free fluid around the spleen | 0
initial diagnosis of sepsis due to cholangitis or liver damage | 0
intravenous antibiotics | 0
meropenem hydrate | 0
endoscopic retrograde cholangiography | 24
no stone in the bile duct | 24
endoscopic nasobiliary drainage | 24
noradrenaline | 24
dobutamine hydrochloride | 24
shock | 24
blood culture positive for klebsiella oxytoca | 24
sensitive to meropenem hydrate | 24
meropenem hydrate administered for 6 days | 24
anemia progressed | 72
required 2 units of blood transfusion | 72
renal damage slightly improved | 72
infection could not be controlled | 72
inflammatory markers remained high | 72
contrast-enhanced abdominal CT | 72
intrahepatic and subcapsular low density areas | 72
wall defect seen in coronal and sagittal - sections | 72
free fluid around the liver and spleen | 72
fluids obtained through paracentesis were hemorrhagic | 72
transhepatic perforation of acute cholecystitis suspected | 72
emergency interventional radiology | 72
percutaneous transhepatic gallbladder drainage attempted | 96
abdominal ultrasonography before PTGBD | 96
high echogenic debris in the gallbladder | 96
no gallbladder swelling, wall thickening and defect | 96
7 Fr. drainage tube inserted into the gallbladder | 96
90 mL of bad smelling red-yellow pus aspirated | 96
cholangiography revealed an orifice of fistula | 96
fistula drained into the intrahepatic secondary abscess | 96
fistula drained into the intraperitoneal cavity | 96
percutaneous abscess drainage attempted | 96
150 mL of hemorrhagic fluid aspirated | 96
abdominal angiography attempted | 96
no evidence of extravasation, hepatic artery aneurysm or cystic artery aneurysm | 96
diagnosis of transhepatic gallbladder perforation confirmed | 96
general condition dramatically improved | 120
emergency laparotomy avoided | 120
culture of red-yellow pus positive for enterococcus avium, enterococcus gallinarum, and klebsiella oxytoca | 120
culture of intrahepatic abscess positive for enterococcus gallinarum | 120
repeat blood culture negative | 120
antibiotics changed to sulbactam sodium/ampicillin sodium | 120
administered for 7 days | 120
contrast-enhanced CT showed reduction in size and localization of intrahepatic abscess and subcapsular hematoma | 408
cholangiography via PTGBD tube revealed recanalization of cystic duct | 408
orifice of fistula not detected | 408
stone in the gallbladder and bile duct not detected | 408
discharged | 792