36 years old | 0
female | 0
admitted to the hospital | 0
loss of consciousness | -2
head trauma | -2
fall from own height | -2
loss of strength in lower extremities | -2
impaired ambulation | -2
holocranial headache | -336
aggressive behavior | -336
vertigo | -336
somatoform disorder | -432
depressive episode | -432
major depression | -1296
suicide attempts | -1296
Glasgow coma score of 11 | 0
mutism | 0
horizontal nystagmus | 0
oculogyric crises | 0
stereotyped movements in all four extremities | 0
normal plantar and other deep tendon reflexes | 0
mass in the right axillar line | 0
blood pressure of 94/60 mm Hg | 0
heart rate of 77 bpm | 0
respiratory rate of 20 rpm | 0
temperature of 36.5°C | 0
body-weight of 60 kg | 0
height of 158 cm | 0
BMI of 24.0 | 0
olanzapine | 0
sertraline | 0
alprazolam | 0
magnesium valproate | 0
urinary tract infection | 0
intravenous ceftriaxone | 0
Acinetobacter baumannii | 72
invasive artificial airway with an endotracheal tube | 72
admittance to the Intensive Care Unit | 72
purulent bronchial secretions | 72
body temperature of 39°C | 72
increase in leucocyte count | 72
intravenous colistimethate and meropenem | 72
extreme bradycardia | 312
asystole | 312
advanced life support protocol | 312
cardiac arrest | 312
necropsy examination | 312
hemorrhagic lesions at the corpus callosum level | 312
multiple paratracheal and perihilar lymph nodes | 312
poorly differentiated malignant neoplastic lesion | 312
melanoma metastasis from an occult primary cancer | 312
axillary ganglion biopsy | 24
high-grade and poorly differentiated malignancy | 24
immunohistochemical staining | 24
HMB-45 staining positive | 24
melan-A staining positive | 24
vimentin staining positive | 24
S-100 staining positive | 24
magnetic resonance imaging | 24
computed tomography | 24
tumor markers screening | 24
electroencephalogram | 24
autoimmune etiology screening | 24
cytoplasmic antineutrophil cytoplasmatic antibodies | 24
perinuclear antineutrophil cytoplasmatic antibodies | 24
anti-double-stranded deoxyribonucleic acid | 24
anti-cardiolipin IgG | 24
anti-cardiolipin IgM antibody | 24
anti-N-methyl-D-aspartate receptor | 24
procalcitonin serum levels | 24
urinalysis | 24
antibodies for hepatitis B virus | 24
antibodies for hepatitis C virus | 24
antibodies for HIV | 24
urinalysis for benzodiazepines | 24
urinalysis for barbiturates | 24
urinalysis for cannabis | 24
urinalysis for cocaine | 24
urinalysis for methamphetamines | 24
urinalysis for opiates | 24
type one respiratory insufficiency | 72
discharged | - 
Note: The event "discharged" is not applicable in this case as the patient passed away.