75 years old | 0
male | 0
admitted to the hospital | 0
painful right scrotal swelling | 0
scrotal swelling increased | -48
scrotal pain increased | -48
fever | -48
rigor | -48
history of diabetes mellitus | -6720
diabetes mellitus controlled with medications | -6720
diabetes mellitus controlled with dietary modifications | -6720
pulse rate 110 beats/minute | 0
blood pressure 100/60 mmHg | 0
temperature 39 Celsius | 0
central abdominal tenderness | 0
suprapubic tenderness | 0
scrotal redness | 0
scrotal tenderness | 0
increased scrotal temperature | 0
elevated white blood cells count | 0
neutrophils | 0
parenteral antibiotics | 0
little improvement | 48
anorexia | 72
nausea | 72
severe abdominal pain | 72
backache | 72
fever | 72
rigor | 72
tenderness all over the abdomen | 72
guarding all over the abdomen | 72
mild bilateral pleural effusions | 72
dilated loops of the small bowel | 72
collection of fluid at the pelvic cavity | 72
normal serum amylase | 72
normal serum lipase | 72
large amount of air collection in the retroperitoneal space | 72
air collection displacing the right kidney toward the midline | 72
air collection extending to the right scrotum | 72
tracking of the contrast media to the retroperitoneum | 72
tracking of the contrast media to the right scrotum | 72
laparotomy | 96
large amount of thin pus in the peritoneal cavity | 96
air and fluid collection in the retroperitoneal space | 96
perforation in the posterior wall of the duodenum | 96
suturing with slowly absorbable suture material | 96
peritoneal cavity washed with warm normal saline | 96
2 drains left in the abdomen | 96
admitted to the intensive care unit | 96
clinical condition improved | 120
drains removed | 120
complete abdominal dehiscence | 192
right scrotal abscess | 192
anther surgery | 192
abdomen closed with tension sutures | 192
drainage of the scrotal abscess | 192
general clinical situation improved | 240
discharged | 240
tension sutures removed | 504
improvement of both the clinical and the imaging studies | 504