57 years old | 0
female | 0
menopausal | 0
admitted to the gynecological emergency unit | 0
left lower quadrant abdominal pain | -336
pelvic heaviness | -336
urinary frequency | -336
miscarriages | -10080
tubal ligation | -10080
active smoker | 0
no medication | 0
large and painful mass | 0
pelvic MRI | 0
mass | 0
no lymphadenopathy | 0
no ascites | 0
no peritoneal implants | 0
uterus and adnexa were normal | 0
serum tumor markers were negative | 0
surgical pelvic exploration | 672
mass of the left broad ligament | 672
no ascites | 672
no peritoneal carcinomatosis | 672
uterus and right adnexa were normal | 672
total hysterectomy with adnexectomy and removal of the mass | 672
leiomyosarcoma | 672
fever | 48
major inflammatory syndrome | 48
leukocytes 15,000/μL | 48
C-reactive protein 317 mg/dL | 48
contrast-enhanced computed tomography scan | 48
abscess | 48
blood pressure dropped | 48
vasopressor therapy | 48
noradrenaline | 48
emergency revision surgery | 72
peritoneal cavity exploration | 72
non-purulent serosanginous peritoneal fluid | 72
adhesions to the Douglas pouch | 72
peritonitis | 72
antibacterial treatment | 72
piperacillin/tazobactam | 72
gentamicin | 72
microbiological samples | 72
extubated | 72
hemodynamic support | 72
noradrenaline | 72
transferred to the intensive care unit | 72
clinically improved | 96
noradrenaline requirement decreased | 96
discontinuation of noradrenaline | 96
decrease in inflammatory markers | 96
microbiological analysis of the peritoneal fluid | 96
Gardnerella vaginalis | 96
gentamicin discontinued | 96
metronidazole | 96
Atopobium vaginae | 120
antibacterial susceptibility testing | 120
Gardnerella vaginalis resistant to metronidazole | 120
Gardnerella vaginalis resistant to ciprofloxacin | 120
Gardnerella vaginalis susceptible to penicillin G | 120
Gardnerella vaginalis susceptible to amoxicillin/clavulanate | 120
Gardnerella vaginalis susceptible to cefotaxim | 120
Gardnerella vaginalis susceptible to clindamicin | 120
Gardnerella vaginalis susceptible to vancomycin | 120
Atopobium vaginae susceptible to metronidazole | 120
piperacillin/tazobactam active against both bacteria | 120
discharged from the intensive care unit | 168
antibacterial therapy stopped | 168