29 years old | 0
primigravida | 0
32-week gestation | 0
presented to the emergency department | 0
acute history of sore throat | -240
high-grade fever | -240
abdominal pain | -240
cough | -240
progressive shortness of breath | -240
poor urine output | -48
decreased fetal movements | -48
uneventful pregnancy | -168
ultrasonography at 30 weeks | -672
single live fetus | -672
normal biometry parameters | -672
symptoms suspicious for COVID-19 | 0
tested by RT-PCR assay | -240
worsening clinical condition | 0
referred to our hospital | 0
strong suspect for COVID-19 | 0
residence in containment zone | 0
investigated for COVID-19 with RT-PCR assay | 0
COVID-19 RT-PCR test negative | 0
previous COVID-19 RT-PCR test negative | 0
chest X-ray | 0
minimal bilateral basal haziness | 0
prominent interstitial markings | 0
acute hypoxemic respiratory failure | 0
hypotension | 0
admitted to the respiratory intensive care unit | 0
community-acquired pneumonia | 0
septic shock | 0
inhaled oxygen supplementation | 0
intravenous fluids | 0
vasopressors | 0
broad-spectrum antibiotics | 0
fundal height corresponding to gestational age | 0
fetal movements not perceived | 0
fetal heart rate not perceived | 0
anemia | 0
leucocytosis | 0
elevated CRP levels | 0
elevated serum procalcitonin levels | 0
acute kidney injury | 0
deranged liver function tests | 0
USG showed intrauterine fetus | 0
no cardiac activity | 0
informed intrauterine death | 0
high-risk consent obtained | 0
induction of labor | 0
stillborn male fetus | 0
no intrapartum adverse events | 0
no postpartum adverse events | 0
Haemoglobin 11.2 gm/dl | 0
total leucocyte counts 20,300/mm3 | 0
platelet counts 2.15 lac/mm3 | 0
serum bilirubin 2.0 mg/dl | 0
SGOT 93 U/L | 0
SGPT 70 U/L | 0
serum creatinine 2.5 mg/dl | 0
CRP 9.8 mg/L | 0
serum sodium 132 mmol/l | 0
serum potassium 4.3 mmol/l | 0
prothrombin time 12.5 s | 0
INR 1.01 | 0
d-dimers 235 ng/ml |.0
blood culture sterile | 0
urine culture sterile | 0
high vaginal swab culture sterile | 0
work-up for Malaria negative | 0
work-up for Dengue negative | 0
work-up for Typhoid negative | 0
work-up for Leptospira negative | 0
work-up for H1N1 Influenza negative | 0
general condition stabilized | 24
reduction in vasopressor requirements | 24
reduction in oxygen requirements | 24
continued febrile | 48
work-up for tropical fevers | 48
peripheral smear for malaria negative | 48
antigen-based assays for malaria negative | 48
serology for dengue negative | 48
serology for leptospira negative | 48
serum Widal tests negative | 48
Scrub typhus IgM-ELISA positive | 48
eschar on right thigh | 48
doxycycline therapy started | 48
clinical response seen | 168
clinical parameters improved | 168
radiological parameters improved | 168
leukocyte counts normalized | 168
serum creatinine normalized | 168
maintaining vitals without oxygen | 168
discharged | 168
