9 months old | 0
male | 0
born by normal vaginal delivery | -26160
healthy parents | 0
presented to Paediatric Emergency Department | 0
four-week history of intermittent pyrexia | -672
irritability | -672
coryzal symptoms | -672
upper respiratory tract infection | -672
urticarial rash | -336
food allergy | -336
vomiting | -336
pallor | -336
loss in weight | -336
received a seven-day course of oral Augmentin | -336
admitted to the hospital | 0
febrile | 0
oxygen saturation 95% in air | 0
pulse rate 152 beats per minute | 0
grade 2/6 ejection systolic murmur | 0
tachypnoeic | 0
respiratory rate 65 breaths per minute | 0
bilateral subcostal recessions | 0
4cm tender hepatomegaly | 0
full sepsis screen | 0
commenced on intravenous ceftriaxone | 0
normocytic normochromic anaemia | 0
haemoglobin level 7.6g/dl | 0
leucocytosis 21.8×10^9/l | 0
lymphocytosis 12×10^9 | 0
normal platelet count | 0
cerebrospinal fluid sterile | 0
mild pleocytosis | 0
normal protein concentration | 0
blood and urine cultures sterile | 0
raised C-Reactive Protein 144 | 0
Erythrocyte Sedimentation Rate 115mm/hr | 0
marked inflammatory response | 0
liver and renal function tests normal | 0
no evidence of disseminated intravascular coagulation | 0
abdominal ultrasound showed homogenous hepatomegaly | 0
no other focal abnormalities | 0
Chest X-ray showed small right pleural effusion | 0
no cardiomegaly | 0
trans-thoracic echocardiogram | 0
giant aneurysm of the left anterior descending artery | 0
thrombus formation in-situ | 0
left main coronary dilated | 0
left circumflex artery dilated | 0
right coronary artery dilated | 0
started on 2g/kg of intravenous immunoglobulin | 0
high dose aspirin therapy | 0
supporting transfusion of crossmatched packed red cells | 0
worsening anaemia | 0
transferred to Neonatal Intensive Care Unit | 0
stringent monitoring | 0
remained febrile | 0
treated with IVIG | 0
responded to methylprednisolone | 0
magnetic resonance angiographic study | 0
excluded concomitant aneurysms | 0
started on regular diuretics | 0
aspirin | 0
heparinisation | 0
weaned onto warfarin | 0
clinical condition resolving steadily | 0
discharged home | 432
treatment regimen consisted of Prednisolone 12mg daily | 432
Aspirin 80mg every 6 hours | 432
Furosemide 8mg twice a day | 432
Spironolactone 8mg twice a day | 432
Warfarin 1mg daily | 432
monitored clinically | 432
repeated trans-thoracic echocardiography | 432
normal development | 8760
developmental milestones satisfactory | 8760
weight 12.0 kg | 8760
serial echocardiograms | 8760
increase in size of aneurysm | 8760
left main and left anterior descending coronary arteries dilated | 8760
Montreal Z-Score 28.1 | 8760
left main coronary artery dilated | 8760
Z-Score 5.6 | 8760
right main coronary artery dilated | 8760
Z-score 2.1 | 8760
proximal aneurysm | 8760
Z-score 13.6mm | 8760
good systolic function | 8760
decent pulsatility of abdominal aorta | 8760
no diastolic tail or reverse flow | 8760
interventricular septum intact | 8760
coronary dilatation confirmed on high resolution CT scan | 8760