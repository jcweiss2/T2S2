36 years old | 0
    female | 0
    admitted to the hospital | 0
    abdominal pain | 0
    constipation | 0
    jaundice | 0
    hypertension | 0
    pre-eclamptic toxaemia | -48
    emergency lower segment caesarean section (LSCS) | -48
    triplet delivery | -48
    elevated alanine amino transferase (ALT) 228.1 IU/L | -24
    elevated aspartate amino transferase (AST) 604.2 IU/L | -24
    hyperbilirubinaemia (356.7 umol/L) | -24
    tachycardia (140/minute) | 0
    blood pressure 176/100 mmHg | 0
    peripheral oxygen saturation 92% (4 L/minute oxygen) | 0
    conscious | 0
    alert | 0
    no neurological deficits | 0
    tachypnoea | 0
    decreased air entry in bilateral lower lung fields | 0
    tender abdomen | 0
    distended abdomen | 0
    tense abdomen | 0
    oliguria | 0
    right-sided consolidation (chest X-ray) | 0
    pleural effusion (ultrasound confirmed) | 0
    massive intraperitoneal collection (CT abdomen) | 0
    thickened bowel loops (CT abdomen) | 0
    severe thrombocytopenia (platelets 20 × 10^9/L) | 0
    haemoglobin 10.2 g% | 0
    white blood cells 11.2 × 10^9/L | 0
    normal coagulation profile | 0
    diagnostic ascites tapping (480/mm3 white blood cells) | 0
    transudative ascites | 0
    bowel injury suspected | 0
    exploratory laparotomy | 24
    ascitic fluid drained (5.7 L) | 24
    haemorrhagic liver parenchyma | 24
    no bowel injury | 24
    no uterus injury | 24
    no abdominal organ injury | 24
    platelet transfusion (12 units) | 24
    intubation | 24
    admission to ICU | 24
    metabolic acidosis (pH 7.17, pCO2 5.1, pO2 8.4, HCO3– 13.9, BE −13.8) | 24
    urine culture negative | 24
    sputum culture negative | 24
    blood culture negative | 24
    negative septic screening | 24
    negative hepatitis viral markers | 24
    negative HIV | 24
    fragmented red cells (peripheral smear) | 24
    anaemia (dimorphic cells) | 24
    polychromatic cells | 24
    burr cells | 24
    thrombocytopenia (peripheral smear) | 24
    leucocytosis (absolute neutrophilia) | 24
    hyperbilirubinaemia (postoperative) | 24
    elevated liver enzymes (postoperative) | 24
    hypoalbuminaemia (postoperative) | 24
    thrombocytopenia (postoperative) | 24
    negative ANA | 24
    negative ANCA | 24
    plasmapheresis initiated | 30
    plasmapheresis (8 times) | 30
    haemodialysis (4 times) | 30
    packed red cells transfusion (5 units) | 48
    packed red cells transfusion (1 unit) | 144
    thrombocytopenia improvement | 240
    liver function improvement | 240
    renal function improvement | 240
    lung condition improvement | 240
    right-side pneumonia | 264
    synpneumonic effusion | 264
    successful extubation | 264
    urine output increased (2.5 L/day) | 312
    shifted to ward | 360
    discharged home | 600