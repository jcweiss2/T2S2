69 years old | 0
man | 0
gastroesophageal reflux | -120
aspiration | -120
dysphagia | -120
intractable esophageal dysmotility | -120
distorted gastroesophageal anatomy | -120
distended intrathoracic post-Collis gastroplasty gastric segment | -120
failed fundoplication | -120
endoscopic esophageal dilations | -120
underwent Ivor Lewis esophagectomy | 0
upper midline abdominal incision | 0
right posterolateral thoracotomy | 0
sixth intercostal space | 0
postoperative anastomotic leak | 48
mediastinitis | 48
sepsis | 48
required return to operating theatre | 48
40 days in intensive care unit | 48
10 days on surgical ward | 48
discharged from hospital | 2160
represented with swelling | 4464
erythema | 4464
pain over right costal margin | 4464
below and medial to end of right thoracotomy wound | 4464
costal osteomyelitis suspected | 4464
noncontrast CT ordered | 4464
osteomyelitis and/or osteochondritis suspected | 4464
bacterial cause assumed | 4464
clindamycin 300 mg 3 times a day prescribed | 4464
surgical options initially declined | 4464
no change in symptoms after 2 months antibiotics | 7296
medical and surgical options discussed again | 7296
elected surgical intervention after 2 weeks | 8736
preoperative MRI demonstrated enhancing collection over sixth rib | 8736
phlegmonous changes involving anterior and lateral right chest wall | 8736
oblique sinus tract extending from collection to seventh costal cartilage | 8736
associated rib fracture | 8736
elective surgical debridement and washout of right costal cartilage | 8736
inflamed soft tissue debridement | 8736
tissue samples showed growth of C. albicans | 8736
C. albicans initially thought to be contaminant | 8736
discharged with oral clindamycin for 6 weeks | 8736
surgical wound remained tender | 11256
swelling | 11256
warmth | 11256
microbiology results re-evaluated | 11256
oral fluconazole 400 mg commenced | 11256
marginally improved after 1 week | 12096
readmitted for intravenous fluconazole and clindamycin | 12096
developed skin breakdown | 12096
cellulitis over affected area | 12096
taken back to theatre for further debridement | 12096
washout | 12096
resection of right anterior fifth and sixth ribs | 12096
tissue samples again showed C. albicans | 12096
made good recovery | 12096
6-month course of oral 400 mg fluconazole | 12096
69 years old|0
man|0
gastroesophageal reflux|-120
aspiration|-120
dysphagia|-120
intractable esophageal dysmotility|-120
distorted gastroesophageal anatomy|-120
distended intrathoracic post-Collis gastroplasty gastric segment|-120
failed fundoplication|-120
endoscopic esophageal dilations|-120
underwent Ivor Lewis esophagectomy|0
upper midline abdominal incision|0
right posterolateral thoracotomy|0
sixth intercostal space|0
postoperative anastomotic leak|48
mediastinitis|48
sepsis|48
required return to operating theatre|48
40 days in intensive care unit|48
10 days on surgical ward|48
discharged from hospital|2160
represented with swelling|4464
erythema|4464
pain over right costal margin|4464
below and medial to end of right thoracotomy wound|4464
costal osteomyelitis suspected|4464
noncontrast CT ordered|4464
osteomyelitis and/or osteochondritis suspected|4464
bacterial cause assumed|4464
clindamycin 300 mg 3 times a day prescribed|4464
surgical options initially declined|4464
no change in symptoms after 2 months antibiotics|7296
medical and surgical options discussed again|7296
elected surgical intervention after 2 weeks|8736
preoperative MRI demonstrated enhancing collection over sixth rib|8736
phlegmonous changes involving anterior and lateral right chest wall|8736
oblique sinus tract extending from collection to seventh costal cartilage|8736
associated rib fracture|8736
elective surgical debridement and washout of right costal cartilage|8736
inflamed soft tissue debridement|8736
tissue samples showed growth of C. albicans|8736
C. albicans initially thought to be contaminant|8736
discharged with oral clindamycin for 6 weeks|8736
surgical wound remained tender|11256
swelling|11256
warmth|11256
microbiology results re-evaluated|11256
oral fluconazole 400 mg commenced|11256
marginally improved after 1 week|12096
readmitted for intravenous fluconazole and clindamycin|12096
developed skin breakdown|12096
cellulitis over affected area|12096
taken back to theatre for further debridement|12096
washout|12096
resection of right anterior fifth and sixth ribs|12096
tissue samples again showed C. albicans|12096
made good recovery|12096
6-month course of oral 400 mg fluconazole|12096
