25 years old | 0
male | 0
congenital macrocephaly with hydrocephalus | -8760
behavioral changes | -2
insomnia | -2
language impairment | -2
admitted to the hospital | 0
abundant stereotypies | 0
tics | 0
discharged | 4
prescription of benzodiazepine | 4
prescription of antipsychotic drug | 4
returned to the hospital | 4
worsening of symptoms | 4
decreased level of consciousness | 4
high fever | 4
non-collaborative | 4
eyes closed | 4
miotic pupils | 4
no conjugated eye deviation | 4
dysarthria | 4
low production of speech | 4
auricular temperature of 39.9 ºC | 4
blood pressure of 103/54 mmHg | 4
HR of 127 bpm | 4
blood gas analysis | 4
blood workup | 4
mild leukocytosis with neutrophilia | 4
slight lymphopenia | 4
normal C-reactive protein | 4
normal procalcitonin | 4
lumbar puncture (LP) | 4
ceftriaxone | 4
ampicillin | 4
acyclovir | 4
CSF showed a slight increase in total proteins | 4
CSF showed 38 cells/mm3 | 4
presumed episodes of focal onset impaired awareness seizures | 24
levetiracetam | 24
sodium valproate | 48
repeated LP for antibody testing | 120
acyclovir stopped | 120
methylprednisolone | 120
EEG showed marked bi-hemispherical cerebral activity disorganization | 120
brain contrasted MRI showed no remarkable signal changes | 120
presence of Anti-NMDAR antibodies in both CSF and serum | 168
admitted to the ICU | 168
respiratory distress | 168
decreased level of consciousness | 168
fluctuating heart rate | 168
low arterial blood pressure profile | 168
vasopressors | 168
severe bradycardia | 168
pauses of up to 5 seconds | 168
severe dystonia | 168
dyskinesia | 168
sialorrhea | 168
IVIg | 240
rituximab | 240
recovery hindered by several infectious complications | 720
discharged from hospital to a rehabilitation facility | 720
decreased level of consciousness | 720
no verbal response | 720
no collaboration on physical exam | 720
bilateral stereotypical movements of the upper limbs | 720
discrete oro-mandibular dyskinesia | 720
recovered well in the next 6 months | 2160
capable of executing everyday activities | 2160
memory lapses of the time he was admitted to the hospital | 2160