66 years old | 0
male | 0
DM | 0
benign prostatic hyperplasia | 0
fatigue | -1008
suprapubic tenderness | -72
urinalysis | 0
protein 1+ | 0
glucose 3+ | 0
blood 3+ | 0
no nitrites | 0
no leukocyte esterase | 0
ultrasound | 0
moderate hydronephrosis of the right kidney | 0
urinary retention | 0
Foley catheter | 0
improved symptoms | 0
returned one week later | 168
lethargy | 168
hyperglycemia | 168
blood glucose 840 mg/dL | 168
continued dysuria | 168
urine culture positive for multidrug-resistant E. coli | 168
blood culture positive for multidrug-resistant E. coli | 168
hemoglobin A1c 13.6% | 168
CT | 168
extensive gas within the bilateral renal parenchyma | 168
gas within the left renal sinus | 168
perinephric fat stranding | 168
thickening of Gerota's fascia | 168
septic shock | 168
bilateral radical nephrectomy | 168
post-operative dialysis-dependent | 168
readmitted for recurrent MDR E. coli pyocystitis | 168
anemia | 168
persistent urinary retention | 168
required intravenous antibiotics | 168
required red blood cell transfusions | 168
required iron supplementation | 168
suprapubic catheter placement | 168
drainage of defunctionalized bladder | 168
EPN diagnosis | 168
bilateral perinephric fat stranding | 168
gas within left renal sinus | 168
mild perivesical fat stranding | 168
mural thickening not visualized | 168
hemorrhage | 168
necrosis | 168
air spaces in subcapsular and perinephric spaces | 168
acute pyelonephritis with abscesses | 168
foci of infarction | 168
abscesses filled with neutrophils | 168
necrotic tissue | 168
bacterial colonies | 168
gas-filled cysts | 168
vasculitis | 168
diabetic nephropathy | 168
RPS class IIB | 168
diffuse thickening of glomerular and tubular basement membranes | 168
severe mesangial expansion | 168
diffuse acute tubular injury/necrosis | 168
loss of proximal tubule brush border | 168
simplified tubular epithelium | 168
sloughed epithelial cells in tubular lumen | 168
mild to moderate intimal fibrosis | 168
thickening of arteriolar walls | 168
dialysis-dependent | 168
recurrent MDR E. coli pyocystitis | 168
readmitted on several occasions | 168
complications requiring antibiotics and transfusions | 168
Foley catheter in bladder | 168
perivesical fat stranding | 168
lack of distention | 168
absence of intravenous contrast | 168
gas in periphery of renal parenchyma | 168
gas in left renal pelvis | 168
bilateral nephrectomy | 168
post-operative complications | 168
readmitted for recurrent infections | 168
suprapubic catheter | 168
defunctionalized bladder drainage | 168
EPN | 168
emphysematous pyelonephritis | 168
gas-forming microorganisms | 168
urinary tract obstruction | 168
septic complications | 168
bilateral EPN | 168
thrombocytopenia | 168
acute renal impairment | 168
altered consciousness | 168
shock | 168
mortality risk factors | 168
lifesaving intervention | 168
infection source control failure | 168
post-operative MDR E. coli pyocystitis | 168
urinary retention | 168
dialysis dependence | 168
readmissions | 168
