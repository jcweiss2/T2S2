73 years old | 0
male | 0
admitted to the hospital | 0
acute on chronic COPD exacerbation | 0
Type 2 respiratory failure | 0
noninvasive ventilation | 0
noradrenaline infusion | 0
continuous veno-venous hemodiafiltration | 0
hemodynamic monitoring | 0
pH 7.057 | 0
base excess -7.5 | 0
PCO2 11.23 kPa | 0
PaO2 13.7 kPa | 0
FiO2 50% | 0
P: F ratio 200 | 0
total leukocyte count 26 × 10^9/L | 0
procalcitonin 11.2 mcg/L | 0
C-reactive protein 104 mg/L | 0
oliguric | 0
acidotic | 0
raised PaCO2 10.86 kPa | 12
failure to remove CO2 | 12
vasopressors requirements increased | 12
Extracorporeal carbon dioxide removal | 12
pump flow 0.56 L/min | 12
sweep flow 10 L/min | 12
sweep FiO2 1.0 | 12
CO2 removal 6-10 L | 12
activated partial thromboplastin time ratio 1.2-1.6 | 12
platelets monitored | 12
fibrinogen monitored | 12
Hb monitored | 12
sweep flows adjusted | 12
heparin infusions avoided | 12
pH improved to 7.30 | 12
PaCO2 normalized to 6.5 kPa | 12
non-invasive ventilation continued | 12
bi-level positive airway pressure MODE | 12
Sats >90% | 12
pH >7.3 | 12
R/R <30 | 12
inflammatory markers improved | 12
TLC 16 × 10^9/L | 12
CRP 46 mg/L | 12
procalcitonin 0.9 mcg/L | 12
enteral nutrition continued | 12
sepsis relapse | 24
acidotic | 24
work of breathing worsened | 24
sweep flows adjusted | 24
Extracorporeal carbon dioxide removal continued | 24
continuous veno-venous hemodiafiltration turned off | 48
renal function recovered | 48
Extracorporeal carbon dioxide removal turned off | 480
sweep flows gradually taken down | 480
critical illness related weakness | 480
prolonged weaning | 480
rehabilitation | 480
physiotherapy | 480
decannulated | 480
discharged from the intensive care unit | 480