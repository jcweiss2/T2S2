27 years old | 0
male | 0
admitted to the hospital | 0
car crash | -1
severe respiratory distress | 0
cyanosis | 0
hemodynamic instability | 0
right pneumothorax | 0
thoracic drainage | 0
bilateral pneumothorax | 0
rib fractures | 0
multiple pulmonary contusions | 0
sacral wing fractures | 0
right tibial plateau fractures | 0
no traumatic brain injury | 0
intubation | 0
mechanical ventilation | 0
left chest drainage | 0
conscious sedation | 0
dexmetomidine | 0
Remifentanil | 0
RASS-2 | 0
pulmonary contusions | 0
bronchial toilet | 0
systemic antimicrobial treatment | 0
amikacin | 0
cefazolin | 0
plate osteosynthesis | 24
septic episode | 96
no shock | 96
microbiological sampling | 96
blood cultures | 96
bilateral broncoalveolar lavage | 96
empiric antimicrobials | 96
piperacillin-tazobactam | 96
linezolid | 96
Pseudomonas spp | 96
Staphylococcus spp | 96
XDR Pseudomonas aeruginosa | 120
high-dose meropenem | 120
colistin | 120
nebulized colistin | 120
intense headache | 144
neck rigidity | 144
lumbar puncture | 144
cerebrospinal fluid cloudy | 144
neutrophils >500/microL | 144
glucose 19 mg/dL | 144
protein 279 mg/dL | 144
Gram-negative bacteria | 150
Pseudomonas spp | 150
high-dose Ceftolozane-tazobactam | 150
high-dose Fosfomycin | 150
Rifampicin | 150
Dexamethasone | 150
right middle-ear suppurative infection | 150
mastoid suppurative infection | 150
meningeal syndrome resolved | 192
right mastoidectomy | 192
tympanoplasty | 192
extubated | 192
transferred to Infectious Diseases Unit | 192
sterile CSF | 216
normalized parameters | 216
fosfomycin discontinued | 216
ceftolozane-tazobactam discontinued | 288
control head bone CT-scans | 288
complete resolution of otomastoiditis | 288
discharged | 288
no clinically relevant neurological sequelae | 288
chronic otitis media | -1000
recurring otitis | -1000
quinolones | -1000
cephalosporins | -1000
XDR-PA selection | -1000
skull fractures | 0
CNS complication | 144
bloodstream infections | 96
pulmonary infections | 96
meningitis | 144
CNS isolates | 150
MICs for colistin | 150
CNS breakthrough infection | 150
insufficient colistin penetration | 150
blood brain barrier | 150
inefficient CNS meropenem concentrations | 150
XDR-PA CNS infections | 150
off-label prescription | 150
Ethics Committee | 150
urgent procedure | 150
pharmacy department | 150
off-label use of C-T | 150
Professor P. Viale | 150
Dr. C. Tascini | 150
urgent discussion | 150
therapeutic option | 150
meningitis | 150