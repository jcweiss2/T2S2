56 years old | 0
    woman | 0
    admitted to the urology department | 0
    undergone ureteroscopy for left ureter | 0
    laparoscopy for lysis of adhesion around left ureter | 0
    abdominal discomfort | 48
    abdominal distension | 48
    oliguria | 48
    irritable | 48
    body temperature of 39.4°C | 48
    pulse rate at 114 beats per minute | 48
    blood pressure declined to 86/59 mm Hg | 48
    respiratory rate at 28 breaths per minute | 48
    oxygen saturation of 89% | 48
    white blood cell count of 15.4 ×10^9/L | 48
    neutrophils 95% | 48
    lymphocytes 5% | 48
    platelet count of 33 ×10^9/L | 48
    blood lactate level of 3.6 mmol/L | 48
    base excess of −11.4 | 48
    serum creatinine increased to 365.7 μmol/L | 48
    ALT of 224U/L | 48
    AST of 858U/L | 48
    prothrombin time extended to 24.2 second | 48
    C-reactive protein of 180.3 mg/L | 48
    procalcitonin of 49.17 ng/mL | 48
    qSOFA score of 3 | 48
    transferred to the ICU | 48
    APACHE II score of 32 | 48
    SOFA score of 17 | 48
    sepsis | 48
    septic shock | 48
    Primaxin (imipenem/cilastatin) | 48
    norepinephrine | 48
    hydrocortisone | 48
    supplemental fluids | 48
    continuous renal replacement therapy | 48
    acute kidney injury (stage 3) | 48
    respiratory distress | 72
    oxygenation index of 184 mm Hg | 72
    endotracheal intubation | 72
    mechanical ventilation | 72
    white blood cell count peaked at 45.3 ×10^9/L | 120
    neutrophils 91.5% | 120
    lymphocytes 1.8% | 120
    blood culture negative | 120
    urine culture negative | 120
    abdominal drainage fluid culture negative | 120
    TB of 245.5 μmol/L | 168
    DB of 196.6 μmol/L | 168
    liver failure | 168
    abdominal ultrasound examination | 168
    gallbladder wall edema | 168
    plasma exchange | 168
    TB dropped | 216
    mechanical ventilation stopped | 216
    endotracheal tube withdrawn | 216
    hemodialysis continued | 216
    transferred back to the urology department | 288
    ALT of 23 U/L | 288
    AST of 39 U/L | 288
    TB of 99.4 μmol/L | 288
    DB of 69.8 μmol/L | 288
    liver function returned to normal | 360
    