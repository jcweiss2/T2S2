45 years old | 0
male | 0
admitted to the hospital | 0
hepatic echinococcosis | -2880
pulmonary echinococcosis | -1800
surgery | -2160
right abdominal distension pain | -2880
pulmonary hypertension | 0
enoxaparin | 0
torsemide | 0
spironolactone | 0
albendazole | 48
praziquantel | 144
diarrhea | 240
stomachache | 240
increased bilirubin | 168
febrile | 240
hair loss | 240
severe myelosuppression | 240
WBC 1.35 × 10^9/L | 240
NEUT 0.73 × 10^9/L | 240
Hgb 97 g/L | 240
WBC 0.46 × 10^9/L | 264
NEUT 0.13 × 10^9/L | 264
Hgb 88 g/L | 264
parenteral nutrition | 264
omeprazole | 264
glutathione | 264
meropenem | 264
granulocyte colony-stimulating factor | 264
gastrointestinal tract reaction recovered | 312
WBC 0.86 × 10^9/L | 312
NEUT 0.25 × 10^9/L | 312
PLT 78 × 10^9/L | 312
Hgb 92 g/L | 312
blood cells began to return to normal levels | 432
discharged | 720