60 years old | 0
male | 0
presented to the emergency department | 0
bilateral wrist pain | 0
left ankle swelling | 0
left ankle pain | 0
pain | 0
pain increased with movement | 0
pain not relieved by ibuprofen | 0
history of gout attack | -72
denied intravenous drug abuse | 0
denied fever | 0
denied recent illness | 0
HIV status | 0
CD4 count 604 | -720
HIV RNA PCR quantity 120000 | -720
low grade fever 37.5°C | 0
tachycardia 120 bpm | 0
non-toxic appearance | 0
no rash | 0
limitation of active movement bilateral wrists | 0
limitation of active movement left ankle | 0
warmth | 0
tenderness to palpation | 0
trace edema left ankle | 0
treated with colchicine 1.2 mg | 0
treated with colchicine 0.6 mg (4 doses) | 0
treated with ibuprofen 800 mg | 0
treated with hydrocodone/acetaminophen 5/325 mg | 0
discharged | 0
prescription for ibuprofen | 0
prescription for hydrocodone/acetaminophen | 0
diagnosed with HIV | 0
diagnosed with acute gout attack | 0
returned 3 days after discharge | 72
worsening pain left ankle | 72
erythema left ankle | 72
swelling left ankle | 72
new right ankle pain | 72
new right ankle erythema | 72
new right ankle edema | 72
new left knee pain | 72
new left knee erythema | 72
new left knee edema | 72
normal vitals | 72
tachycardia 122 bpm | 72
labs obtained | 72
arthrocentesis left knee | 72
treated with ketorolac | 72
peripheral WBC 9.4 | 72
uric acid 6.9 mg/dL | 72
joint aspirate WBC 8.7×10³ cells/μL | 72
no crystals in joint aspirate | 72
discharged | 72
nonsteroidal anti-inflammatory drugs | 72
rheumatology follow up | 72
diagnosed with inflammatory arthritis | 72
found 2 days after second discharge | 168
unresponsive | 168
entire left lower extremity edema | 168
purpura left leg | 168
purpura right ankle | 168
CT left leg edema only | 168
head CT negative | 168
acute renal failure Cr 2.2 | 168
peripheral WBC 6.6 | 168
17% bands | 168
knee cultures growing gram negative coccobacilli | 168
taken to OR for washout | 168
admitted to ICU | 168
intubated for airway protection | 168
blood cultures grew N. meningitides | 168
cerebral spinal fluid cultures grew N. meningitides | 168
required xigris | 168
required levophed | 168
prolonged hospital course | 168
multiple surgical procedures for debridement/washouts | 168
I&Ds bilateral lower extremities | 168
infected wounds from purpura fulminans | 168
wound vac management | 168
skin grafts left lower extremity | 168
acute renal failure due to urinary retention | 168
hydronephrosis | 168
urology consult | 168
taught in-and-out catheterizations | 168
diagnosed with mild SIADH | 168
fluid restriction | 168
left-sided hearing loss due to meningitis | 168
deep vein thrombosis right upper extremity | 168
bridged from enoxaparin to warfarin | 168
treated for hospital-acquired UTI | 168
required multiple blood transfusions | 168
nutritional supplementation for malnourishment | 168
neurology consult | 168
negative brain MRI | 168
negative EEG | 168
infectious disease consult | 168
treated with ceftriaxone 14 days | 168
treated with vancomycin | 168
treated with meropenem | 168
discharged after 62 days | 1488
