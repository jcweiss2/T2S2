75 years old | 0
female | 0
left THA | -4320
osteoarthritis | -4320
complication free for 2 years postoperatively | -4320
three dislocations | -17520
most recent dislocation 3 years prior | -25920
left hip pain | 0
inability to ambulate | 0
posterosuperior prosthetic hip dislocation | 0
left leg internally rotated | 0
left leg shortened | 0
detailed neurovascular examination | 0
closed reduction attempted under general anesthesia | 0
paralytic agent used | 0
reduction techniques: axial traction with 90 degrees flexion | 0
internal rotation |0
adduction | 0
flexion | 0
axial traction with alternating external rotation | 0
internal rotation | 0
radiographs showing posterior-superior dislocation | 0
anterior-inferior-medial dislocation | 0
anterior-lateral dislocation | 0
failed closed reduction | 0
decision to transfer to tertiary referral center | 0
dense sciatic nerve motor injury | 0
no motor function below knee | 0
decreased sensation | 0
paresthesia | 0
florid acute pulmonary edema | 0
Takotsubo cardiomyopathy | 0
intensive care unit admission | 0
transfer delayed for 3 days | 72
successful closed reduction with specialized traction table | 72
bone fragment from ischium | 72
nerve exploration considered | 72
patient's medical condition prevented nerve exploration | 72
sciatic nerve no recovery | 72
discharged home with ankle foot orthosis | 72
recurrent dislocation 3 weeks later | 600
revision indicated | 600
sciatic nerve exploration | 600
laceration of 60% of sciatic nerve | 600
neurolysis performed | 600
revision to dual-mobility liner | 600
retention of primary cup | 600
added 7 mm head length | 600
implanted device: 22 + 7-mm inner-diameter ball | 600
41-mm polyethylene sphere | 600
decision against intraoperative nerve repair consult | 600
peripheral nerve consult obtained postoperatively | 600
decision to forgo nerve repair | 600
diminished sensation | 600
abnormal sensation | 600
0/5 motor function in sciatic nerve distribution | 600
dislocation event 2 weeks post revision | 600
spinopelvic immobility | 600
stable for 6 months postoperatively | 4320
ambulating with walker | 4320
slap foot/steppage gait | 4320
no pain | 4320
0/5 motor function | 4320
diminished sensation | 4320
discontinued ankle foot orthosis | 4320
heel ulcer | 4320
