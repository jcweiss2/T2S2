50 year old | 0
    female | 0
    visited the emergency department | 0
    epigastric pain | -360
    fever | -360
    chill | -360
    nausea | -360
    abdominal surgery for multiple biliary stones | -175200
    acute continuous dull-like pain | 0
    epigastrium pain without radiation | 0
    abdomen soft | 0
    tender on right upper quadrant | 0
    no rebound tenderness | 0
    white blood cell count 14760/mm3 | 0
    hemoglobin level 10.0 g/dL | 0
    erythrocyte sedimentation ratio 140 mm/hr | 0
    c-reactive protein level 23.89 mg/dL | 0
    aspartate aminotransferase level 101 IU/L | 0
    alanine aminotransferase level 114 IU/L | 0
    total bilirubin 4.6 mg/dL | 0
    amylase level 48 U/L | 0
    abdominal computed tomographic scan | 0
    multiple stones in common bile duct | 0
    multiple stones in intra-hepatic duct | 0
    biliary obstruction | 0
    multifocal liver abscesses | 0
    air-biliarygram | 0
    emergency ERCP performed | 0
    opening of choledochoduodenostomy observed | 0
    cholangiogram confirmed multiple filling defects in CBD | 0
    wide ostomy orifice | 0
    marked dilatation of CBD | 0
    extraction of brown-pigmented mud stones | 0
    suddenly became hypoxic | 0
    suddenly became bradycardic | 0
    comatose | 0
    cardiac arrest developed | 0
    procedure terminated | 0
    cardio-pulmonary resuscitation commenced | 0
    prompt intubation | 0
    transferred to intensive care unit | 0
    resuscitation continued | 0
    died without restoration | 0
    chest X-ray suggested massive systemic air embolism | 0
    death caused by massive cardiac and pulmonary air embolism | 0
    multiple liver abscesses | 0
    history of choledochoduodenostomy | -175200
    sphincterotomy during ERCP | 0
    ERCP following liver biopsy | 0
    ERCP following PTBD | 0
    high intraluminal air pressure | 0
    biliary-hepatic venous fistulas | 0
    insufflated air | 0
    pathological state of hepatobiliary tissues | 0
    deteriorated vital signs | 0
    deteriorated neurologic signs | 0
    <|eot_id|>
    