21 years old | 0
male | 0
admitted to the hospital | 0
febrile urinary tract infection | 0
no significant medical history | 0
physical examination was normal | 0
mild thrombocytopenia | 0
elevated liver enzymes | 0
primary EBV infection | 0
MRI of the kidneys revealed no abnormalities | 0
splenomegaly | 0
multiple hepatic lesions | 0
antibiotic therapy was stopped | 0
paracetamol was replaced by metamizole | 0
no microbiological urine culture | 0
no blood culture | 0
liver function had decreased dramatically | 96
acute liver failure | 96
acute renal failure | 96
leucopenia | 96
thrombopenia | 96
elevated ferritin level | 96
severe immune dysregulation | 96
transferred to the University Hospital Vienna | 96
genital lesions suggestive of HSV infection | 96
intravenous acyclovir was started | 96
patient's condition rapidly deteriorated | 100
multiorgan failure | 100
died | 144
EBV DNA was detected by PCR | 120
primary EBV infection was confirmed by serology | 120
HSV1 PCR was highly positive | 120
HSV IgG antibody seroconversion | 120
postmortem analysis of liver, spleen, kidney and gallbladder | 144
HSV1 and EBV DNA in all samples | 144
histopathology of liver samples | 144
necrosis pattern of HSV hepatitis | 144
mixed reactive inflammatory infiltrate | 144
immunoperoxidase staining confirmed HSV1 hepatitis | 144
characteristic features of EBV-hepatitis | 144
EBV LMP1 detected by alkaline phosphatase staining | 144
EBV by PCR after extraction of EBV DNA | 144
haemophagocytosis in liver tissue | 144
SHLH was suspected | 96
SHLH was diagnosed | 144
soluble CD25 was elevated | 144
fulminant hepatitis | 0
severe disease in immunocompetent persons | 0
secondary haemophagocytic lymphohistiocytosis | 0 
fever | 0
splenomegaly | 0
cytopenia in two blood cell lines | 96
elevated ferritin | 96
elevated sCD25 | 144 
virological diagnosis | 120
antiviral therapy | 96
immunosuppressive treatment | 96 
supportive intensive care | 96