32 years old | 0
female | 0
Hispanic | 0
admitted to the hospital | 0
fever | -72
chills | -72
generalized weakness | -72
malaise | -72
body aches | -72
tachycardia | -72
heart rate of 120 beats per minute | -72
blood pressure of 128/82 mmHg | -72
respiratory rate of 18 breaths per minute | -72
oxygen saturation of 99% | -72
denies chest pain | -72
denies cough | -72
denies shortness of breath | -72
denies abdominal pain | -72
resided in a rural community in coastal South Texas | 0
had dogs and cats at home | 0
no recent exposure to communicable diseases | 0
no recent travel outside of the country | 0
no tobacco use | 0
no alcohol use | 0
no illicit drug use | 0
white blood cells 4300 cells/mm3 | -72
neutrophils 85% | -72
lymphocytes 11.4% | -72
monocytes 3% | -72
hemoglobin 12.4 g/dL | -72
hematocrit 37.2% | -72
platelets 230,000 per cubic mm | -72
aspartate aminotransferase 38 U/L | -72
alanine aminotransferase 28 U/L | -72
alkaline phosphatase 62 U/L | -72
rapid influenza A and B test normal | -72
urinalysis normal | -72
lactic acid normal | -72
thyroid-stimulating hormone normal | -72
chest radiograph indicated mild peribronchial cuffing | -72
received one liter of 0.9% normal saline intravenously | -72
received one oral dose of ibuprofen 800 mg | -72
diagnosed with viral bronchitis | -72
discharged home | -72
returned to the Emergency Department | 96
temperature of 101.2 °F | 96
tachycardia with a heart rate of 125 beats per minute | 96
respiratory rate of 17 breaths per minute | 96
blood pressure of 118/56 mmHg | 96
oxygen saturation of 99% | 96
diminished breath sounds to bilateral lung fields | 96
dry mucous membranes | 96
decreased skin turgor | 96
white blood cells 3600 cell/mm3 | 96
neutrophils 82.8% | 96
lymphocytes 11% | 96
monocytes 5% | 96
hemoglobin 11.6 g/dL | 96
hematocrit 33.2% | 96
platelets 64,000 per cubic mm | 96
aspartate aminotransferase 226 U/L | 96
alanine aminotransferase 138 U/L | 96
alkaline phosphatase 182 U/L | 96
D-dimer >5000 ng/mL | 96
lactic acid 2.4 mmol/L | 96
fibrinogen normal | 96
chest radiograph identified bilateral alveolar infiltrates | 96
computed tomographic angiogram of the chest negative for pulmonary embolism | 96
bilateral lower lobe consolidation | 96
admitted to the medical-surgical floor | 96
diagnosis of sepsis secondary to community-acquired pneumonia | 96
sepsis protocol initiated with meropenem and voriconazole | 96
resuscitation with 3 liters of intravenous 0.9% normal saline fluid | 96
became hypotensive | 102
blood pressure of 87/53 mmHg | 102
heart rate of 137 beats per minute | 102
respiratory rate of 36 breaths per minute | 102
transferred to the Intensive Care Unit | 102
received two more liters of intravenous fluid of 0.9% normal saline | 102
developed a dry cough | 108
acute hypoxemic respiratory failure | 108
heart rate of 144 beats per minute | 108
respiratory rate of 33 breaths per minute | 108
oxygen saturation of 82% | 108
echocardiogram revealed mild right heart chamber dilatation | 108
normal left ventricular systolic function | 108
ejection fraction of 65% | 108
arterial blood gases showed PaO2/FiO2 of 102 | 108
managed with non-invasive positive pressure ventilation | 108
voriconazole discontinued | 108
meropenem and doxycycline continued | 108
nontender pink maculopapular rash to the bilateral lower extremities | 144
without associated lymphadenopathy | 144
zoonoses serology panel confirmed acute infection of murine typhus | 168
Typhus Fever group IgM titer of 1:128 | 168
murine typhus IgG titer of 1:258 | 168
meropenem discontinued | 168
antimicrobials deescalated to doxycycline monotherapy | 168
weaning process from non-invasive positive pressure ventilation | 168
high flow oxygen nasal cannula | 168
low flow oxygen nasal cannula at 2 liters per minute | 168
discharged home without oxygen supplementation | 192
treatment completed with minocycline for 11 additional days | 192
generalized weakness at the moment of discharge | 192
no other complaints | 192