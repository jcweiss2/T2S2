57 years old | 0
male | 0
heavy consumption of alcohol | 0
lumbar spinal epidural abscess | 0
dental infection | -240
lumbar torsion | -240
low back pain | -240
loss of balance | -240
rough ground | -240
lumbar pain | -240
fever | -240
systemic inflammatory syndrome | 0
erythrocyte sedimentation rate of 60 mm/hour | 0
C-reactive protein of 111 mg/L | 0
white cell count of 23 G/L | 0
segmented neutrophils 91% | 0
blood cultures collected | 0
lumbar radiographs showing degenerative signs | 0
lumbar MRI showing epidural abscess | 0
L3-L4 epidural abscess | 0
L4-L5 epidural abscess |$0$
L5-S1 epidural abscess | 0
L5-S1 discopathy | 0
psoas abscess | 0
emergency surgery | 0
decompressive laminectomy | 0
posterior approach | 0
L3 to S1 decompression | 0
collections visualized | 0
microbiological studies | 0
intravenous amoxicillin-clavulanic acid | 0
abscess cultures positive for Streptococcus mitis/oralis | 0
blood cultures positive for Streptococcus mitis/oralis | 0
fragment of ligamentum flavum analyzed | 0
transoral echocardiography performed | 0
BARD 5f picc-line placed | 0
penicillin-G treatment | 0
lumbar pain decreased | 0
no fever during hospital stay | 0
CRP decreased | 0
WCC normalized | 0
discharged | 264
surgical wound healing well | 264
antibiotic treatment changed to ceftriaxone | 264
infected teeth treated | 264
asymptomatic at 6-week follow-up | 1008
CRP of 6 mg/L at 6-week follow-up | 1008
lumbar MRI showing resolved infection | 1008
L5-S1 collapse | 1008
asymptomatic at 1-year follow-up | 8760
no persistent infection | 8760
no recurrent infection | 8760
L5-S1 collapse stable | 8760
surgical wound appearance postoperatively | 0
local peripheral redness | 0
wound swelling | 0
wound resolved | 240
spondylodiscitis diagnosis confirmed | 0
no neurological deficit | 0
reflexes normal | 0
reflexes symmetrical | 0
Lasègue manoeuvre negative | 0
Bragard manoeuvre negative | 0
no endocarditis | 0
no chest pain | 0
no shortness of breath | 0
denies chest pain | 0
no vertebral erosion | 0
no evidence of spondylolisthesis | 8760
peripheral inflammatory pannus resolved | 8760
