67 years old | 0
    male | 0
    referred to hepatobiliary surgical team | 0
    obstructive jaundice | -720
    anorexia | -720
    weight loss (10 kg over several months) | -720
    raised serum bilirubin (93 μmol/l) | 0
    elevated serum AST (50 IU/l) | 0
    elevated serum ALP (454 IU/l) | 0
    ultrasound confirmed biliary obstruction | 0
    CT scan showing intraluminal filling defect in mid common bile duct | 0
    endoscopic retrograde cholangiopancreatography | 0
    biliary stenting | 0
    high-grade dysplastic cells | 0
    no invasive malignancy | 0
    provisional diagnosis of cholangiocarcinoma | 0
    pylorus-preserving pancreatoduodenectomy | 24
    Roux-en-Y reconstruction | 24
    pancreatojejunostomy | 24
    hepaticojejunostomy | 24
    gastrojejunostomy | 24
    two foci of high-grade biliary dysplasia in cystic duct | 24
    high-grade biliary dysplasia in intrapancreatic segment of common bile duct | 24
    low-volume pancreatic leak | 168
    sepsis | 168
    Hb level 8.5 g/dl | 168
    white cell count 21.3 × 10^9/l | 168
    neutrophil count 18.1 × 10^9/l | 168
    platelet count 293 × 10^9/l | 168
    bilirubin 31 μmol/l | 168
    AST 45 IU/l | 168
    ALP 63 IU/l | 168
    CRP 73 mg/l | 168
    pleural drain placement | 168
    peritoneal drain placement | 168
    nasojejunal tube for feeding | 168
    in-patient stay of nearly 3 weeks | 504
    discharged | 504
    haematemesis | 576
    collapse | 576
    hemodynamic instability | 576
    Hb level 5 g/dl | 576
    platelets 113 × 10^9/l | 576
    transfusion with packed red blood cells | 576
    platelet transfusion | 576
    coagulation products administered | 576
    intensive care unit admission | 576
    angiogram revealing gastro-duodenal artery stump hemorrhage | 576
    covered stent placement over gastro-duodenal artery origin | 576
    bile leak from old drain site | 672
    retrievable covered stent across hepaticojejunostomy | 672
    percutaneous transhepatic cholangiography | 672
    CT-guided drainage of collection | 672
    broad-spectrum antibiotics | 672
    Enterococcus faecalis infection | 672
    appropriate antibiotics for Enterococcus faecalis | 672
    discharge after 4 weeks | 1344
    jaundice | 10368
    biliary sepsis | 10368
    bilirubin 54 μmol/l | 10368
    AST 52 IU/l | 10368
    ALP 320 IU/l | 10368
    CRP 91 mg/l | 10368
    CT scan showing 9 cm central liver mass | 10368
    multiple smaller liver lesions | 10368
    no evidence of malignancy on liver biopsy | 10368
    antibiotics treatment | 10368
    percutaneous transhepatic cholangiogram | 10368
    biliary drains | 10368
    repeat CT showing no change in liver lesions | 1344
    repeat cholangiography | 1344
    repeat biliary stenting | 1344
    repeat liver biopsy | 1344
    moderately differentiated adenocarcinoma | 1344
    metastatic cholangiocarcinoma | 1344
    deterioration of liver function tests | 1440
    bilirubin 234 μmol/l | 1440
    alanine aminotransferase 80 IU/l | 1440
    AST 200 IU/l | 1440
    ALP 364 IU/l | 1440
    gamma-glutamyl transferase 563 IU/l | 1440
    palliative care referral | 1440
    death due to biliary sepsis | 1440
    