18 years old | 0
male | 0
Asian-Indian | 0
tropical chronic pancreatitis | -720
oral pancreatic enzyme therapy | -720
non-insulin-dependent diabetes | -720
glucotrol | -720
midepigastric pain | -6
dull pain | -6
radiating pain | -6
exacerbated by food intake | -6
recurrent pain | -720
pain control with narcotics | -720
epigastric pain | -48
increased intensity | -48
nausea | -48
vomiting | -48
no fever | -48
CT scan | -48
fatty atrophy of pancreatic head and uncinate process | -48
pancreatic duct filled with large calcifications | -48
obstruction at the level of the neck | -48
upstream ductal dilatation | -48
1.5 cm | -48
hospitalized for pain control | -48
similar pain and fever | -144
CT scan of the abdomen | -144
chronic atrophic calcific pancreatitis | -144
dilated pancreatic duct | -144
intraductal calculi | -144
ERCP | -144
pancreatography | -144
medically managed | -144
discharged | -144
removal of ductal stones | -144
fever | -48
chills | -48
rigors | -48
severe sepsis | -48
septic shock | -48
intubated for hypoxemic respiratory failure | -48
acute respiratory distress syndrome | -48
multiorgan failure | -48
broad-spectrum antibiotics | -48
vasopressor support | -48
activated recombinant human protein C | -48
ultrasound of the abdomen | -48
markedly dilated pancreatic duct | -48
8.7 × 7.6 mm calculus | -48
diffusely echogenic pancreas | -48
prominent common bile duct | -48
bedside emergency ERCP | -48
Olympus TJF-160 side viewing video duodenoscope | -48
major papilla of Vater | -48
frank pus | -48
no papillitis | -48
no tumor | -48
no previous sphincterotomy | -48
cannula tip | -48
evacuation of pus | -48
yellow pus | -48
viscous fluid | -48
cholangiogram | -48
normal biliary tree | -48
no stones | -48
pancreatogram | -48
marked dilatation of the main pancreatic duct | -48
single distal calculus | -48
guide wire | -48
pancreatic duct | -48
total of approximately 20 ml of pus | -48
duct manipulation | -48
5-cm-long 5 F stent | -48
failed to show any more pus draining | -48
pulled out | -48
contrast enhanced CT scan | -48
inflammatory changes within the fat surrounding the body and tail of the pancreas | -48
edema | -48
diminished dilatation of the pancreatic duct | -48
calculus showing distal migration towards the sphincter of Oddi | -48
no evidence of pancreatic necrosis or fluid collection | -48
bilateral moderate pleural effusions | -48
24 hours after the endoscopic intervention | -24
dramatic signs of clinical improvement | -24
stabilization of hemodynamic parameters | -24
blood cultures | -24
Klebsiella ornithinolytica | -24
sensitive to the antibiotics given | -24
extubated | -24
transferred from the intensive care unit | -24
completed his antibiotic course | -24
discharged home | -24
11 days after admission | -24
follow-up examinations | -24
no further complications | -24