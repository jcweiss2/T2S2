66 years old | 0
female | 0
endometrial cancer | -192
chemotherapy | -192
doxorubicin | -192
cisplatin | -192
neutropenic fever | 0
pancytopenia | 0
admitted to the hospital | 0
broad-spectrum antibiotics | 0
hypoxic respiratory failure | 72
intubation | 72
endotracheal tube diameter 8.0 mm | 72
acute pulmonary edema | 72
septic shock | 72
minute ventilation suddenly dropped | 84
suctioning endotracheal tube | 84
mildly blood-tinged material | 84
chest radiography no change | 84
chest radiography completely opacified left hemithorax | 96
no breath sounds over left chest | 96
platelets 38,000/µL | 96
flexible bronchoscopy | 96
large blood clot obstructing left main bronchus | 96
bronchoscopic lavage | 96
forceps extraction | 96
unsuccessful removal attempts | 96
cryoprobe application | 96
frozen for 10 seconds | 96
blood clot attached to probe | 96
successful removal in four pieces | 96
follow-up chest X-ray significant improvement | 96
fifteen minutes required for removal | 96
no further obstructive events | 96
repeat bronchoscopic evaluation | 528
no evidence of clot | 528
airways patent | 528
recovered from septic shock | 528
discharged from hospital | 576
