60 years old | 0
male | 0
ischemic cardiomyopathy | 0
admitted for VT storm | 0
anteroseptal myocardial infarction | -10800
treated with thrombolytic medication | -10800
primary-prevention subcutaneous implantable cardioverter-defibrillator | -3600
VT episodes | -3600
medication adjustments | -3600
S-ICD explant | -240
cardiac resynchronization therapy | -240
cardiac magnetic resonance imaging | -240
LV thrombus | -240
treatment via vitamin K antagonist | -240
VT storm | -240
transferred to academic hospital | -240
hypotensive | -240
external electrical cardioversions | -240
high-dose antiarrhythmic drugs | -240
amiodarone | -240
beta-blockers | -240
mexiletine | -240
quinidine | -240
septic | -240
antibiotic therapy | -240
Staphylococcus aureus bacteremia | -240
antibiotics adjusted | -240
physical examination | -240
echocardiography | -240
positron emission tomography | -240
endocarditis protocol | -240
no signs of endocarditis | -240
antibiotics continued | -240
catheter ablation considered | -240
apical thrombus | -240
unsuitable for catheter ablation | -240
sedation | -240
intubation | -240
adjustment of antiarrhythmic medication | -240
VTs recurred | -240
percutaneous left stellate ganglion blockade | -240
cardiac radioablation considered | -240
therapeutic options discussed | -240
patient opted for cardiac radioablation | -240
written informed consent | -240
cardiac radioablation | 0
targeting guided by American Heart Association Segmented Model | 0
electro-anatomic alterations | 0
VT exit sites | 0
delayed enhancement on cardiac MRI | 0
wall-thinning on cardiac CT | 0
semiautomatically segmented treatment-planning 4D-CT-scan | 0
myocardial scar | 0
echocardiographic deformation imaging | 0
abnormal strain percentages | 0
basal inferior segment | 0
normal shortening | 0
VT morphologies | 0
inferred exit sites | 0
basal anterior | 0
inferolateral apex | 0
clinical target volume | 0
internal target volume | 0
planning target volume | 0
dose of 25 Gy | 0
volumetric-modulated arc therapy plan | 0
patient treated on Agility | 0
77 sustained VT-episodes | -888
mean of 2.1 VT-episodes/day | -888
25 VT episodes required termination by electrical cardioversion | -888
VT recurred 4 hours after cardiac radioablation | 4
no further VTs occurred | 4
patient transferred back to secondary hospital | 312
patient discharged home | 672
no further episodes of VT | 1008
COVID-19 infection | 1008
no VT episodes | 1008
cardiac rehabilitation therapy | 1008
antiarrhythmic drugs tapered off | 1008
no signs of myocardial injury | 0
hs-Troponin-T levels unchanged | 0
echocardiographic ejection fraction unchanged | 0
electrocardiogram unchanged | 0
NT-ProBNP reduced by 77% | 24
no pericardial effusion | 24
nausea and vomiting | 48
antiemetic medication | 48
no adverse events or complications | 0
whole body [18F]FDG-PET/CT-scan | 720
no signs of endocarditis | 720
increased metabolic activity | 720
left ventricle showed extensive 18F-FDG uptake | 720
actual treatment target not metabolically active | 720
LV thrombus evaluated with follow-up CT-scans | 720