75 years old | 0
male | 0
admitted to the hospital | 0
fever | -168
chills | -168
dizziness | -168
remission after fever | -168
no headache | -168
no abdominal pain | -168
no diarrhea | -168
no sputum | -168
no nasal congestion | -168
no runny nose | -168
hypertension | -672
highest body temperature 39.0 °C | -168
body temperature 39 °C | 0
heart rate 98 bpm | 0
respiratory rate 20 breaths per minute | 0
blood pressure 139/75 mmHg | 0
oxygen saturation 98% | 0
clear breath sounds | 0
uniform heart rhythm | 0
negative neurological tests | 0
white blood cell count 7.1 × 10^9/L | 0
neutrophils 58.6% | 0
monocytes 24.4% | 0
hemoglobin 83 g/L | 0
C-reactive protein 111.20 mg/L | 0
interleukin-6 279.22 pg/mL | 0
interleukin-10 3653.30 pg/mL | 0
procalcitonin 0.19 ng/mL | 0
blood amyloid A 509.5 mg/L | 0
erythrocyte sedimentation rate 71 mm/L | 0
lactate dehydrogenase 694 U/L | 0
creatine kinase 19 U/L | 0
albumin 27 g/L | 0
K+ 2.99 mmol/L | 0
Na+ 135.1 mmol/L | 0
Cl- 98.5 mmol/L | 0
calcium 1.87 mmol/L | 0
phosphorus 0.65 mmol/L | 0
normal creatinine level | 0
anti-nuclear antibody titer 1:100 | 0
anti-SSA- | 0
anti-SCL70 positive | 0
normal TORCH test | 0
normal Plasmodium test | 0
normal fungal D-glucan test | 0
normal coronavirus disease 2019 | 0
normal hemorrhagic fever IgM antibody | 0
normal Widder test | 0
normal Weil Felix reaction | 0
bilateral blood culture test positive for L. monocytogenes | 0
cerebrospinal fluid nucleated cell count 420 × 10^6/L | 0
cerebrospinal fluid lymphocyte 75% | 0
cerebrospinal fluid lactate dehydrogenase 472 U/L | 0
cerebrospinal fluid total protein 261.3 mg/dL | 0
cerebrospinal fluid glucose 1.51 mmol/L | 0
cerebrospinal fluid chloride content 111.0 mmol/L | 0
cerebrospinal fluid adenosine deaminase 16 U/L | 0
cerebrospinal fluid cryptococcal smear negative | 0
cerebrospinal fluid cryptococcal capsular antigen test negative | 0
cerebrospinal fluid culture negative | 0
cerebrospinal fluid metagenomic test positive for L. monocytogenes | 0
pleural effusion | 0
nodules in pleura and under pleura | 0
sepsis | 0
lung infection | 0
respiratory failure | 0
electrolyte imbalance | 0
hyponatremia | 0
hypokalemia | 0
autoimmune disease | 0
Listeria monocytic meningoencephalitis | 0
levofloxacin 0.5 g qd | 0
body temperature above 39.0 °C | 72
Staphylococcus capital subspecies | 72
Vancomycin injection 500000 U q6h | 72
body temperature normal | 120
discharged | 168
high fever | 168
chills | 168
cough | 168
sputum | 168
thick sputum | 168
no chest pain | 168
no limb twitching | 168
sluggish pupils | 168
confusion | 168
mental softness | 168
diarrhea | 168
hospitalized in ICU | 168
high-frequency oxygen inhalation | 168
piperacillin and tazobactam 4.5 g q8h | 168
methylprednisolone 40 mg | 168
repeated fever | 192
body temperature above 38.3 °C | 192
levofloxacin 0.5 g qd | 192
body temperature normal | 216
CRP 76.4 mmol/L | 216
transferred to general ward | 216
atrial fibrillation | 216
unresponsiveness | 216
slurred speech | 216
shortness of breath | 216
slow light reflexes | 216
stiff neck | 216
increased muscle tone | 216
wet rales | 216
septic shock | 216
norepinephrine micropump | 216
vancomycin injection 1 million units q12h | 216
meropenem injection 1.0 g q8h | 216
methylprednisolone reduced to 20 mg | 216
methylprednisolone stopped | 216
unconsciousness | 240
base of tongue fell back | 240
shortness of breath | 240
stiff neck | 240
tremor of limbs | 240
heart rate 40 beats per minute | 240
tracheal intubation | 240
ventilator-assisted ventilation | 240
deteriorating condition | 240
multiple organ failure | 240
discontinuation of treatment | 240