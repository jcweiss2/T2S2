64 years old | 0
white | 0
male | 0
presented to the hospital | 0
ground-level fall | 0
episode of dizziness | 0
episode of lightheadedness | 0
hypoglycemia | 0
hemodynamically stable | 0
alert | 0
oriented | 0
bilateral lower extremity pitting edema | 0
small superficial forehead abrasion | 0
stage 2 sacral decubitus ulcer | 0
ruptured skin blister on the left medial calcaneus | 0
leukocytosis | 0
white blood cell count of 14.7 × 103 cells/μl | 0
neutrophil count of 12.2 × 103 cells/μl | 0
serum creatinine concentration of 1.33 mg/dl | 0
optimal medical therapy | 0
signs and symptoms of evolving sepsis | 0
septic shock | 24
exacerbation of congestive heart failure | 24
admission to the intensive care unit | 24
bacteremia | 24
methicillin-sensitive Staphylococcus aureus infection | 24
acute tubular necrosis | 264
dialysis | 264
persistently positive blood cultures | 264
evaluated for infective endocarditis | 264
heart failure with preserved ejection fraction | -1464
symptomatic bradycardia | -1464
status-post pacemaker placement | -1464
hypertension | -1464
hyperlipidemia | -1464
controlled type 2 diabetes mellitus | -1464
dental procedure | -1344
computed tomography of the chest | 0
large bilateral pleural effusions | 0
pulmonary vascular congestion | 0
blood cultures obtained on admission | 0
MSSA bacteremia | 0
repeated blood cultures | 24
multiple thoracentesis | 24
transudative effusions | 24
no evidence of bacteria | 24
cultures of urine | 24
cultures of sputum | 24
cultures of bronchial washings | 24
no bacterial growth | 24
transthoracic echocardiogram | 24
moderate pulmonic valve regurgitation | 24
no vegetation visualized on the valves | 24
transesophageal echocardiogram | 264
mobile 7- × 8-mm mass on the ventricular surface of the pulmonic valve | 264
moderate regurgitation | 264
differential diagnoses for the mass | 264
papillary fibroelastoma | 264
bacterial vegetation | 264
severe illness | 264
deemed not a surgical candidate | 264
AngioVac mass debulking | 384
ultrasonography-guided approach | 384
accessed right common femoral vein | 384
accessed left common femoral vein | 384
therapeutic anticoagulation with heparin | 384
serial dilation | 384
18-F cannula inserted | 384
attached to the return of the cardiopulmonary bypass | 384
26-F sheath advanced to the inferior vena cava | 384
pigtail catheter advanced to the pulmonary artery | 384
Amplatz Super Stiff guidewire advanced through the pigtail | 384
fluoroscopic guidance | 384
TEE guidance | 384
AngioVac cannula advanced to the right ventricular outflow tract | 384
steered into the side of the mass | 384
right heart bypass initiated by the AngioVac system | 384
flow up to 3 l/min | 384
successful extraction of the mass | 384
repeat TEE imaging indicated complete removal of the mass | 384
no damage to the valve | 384
no worsening of moderate regurgitation | 384
tolerated the procedure well | 384
no complications | 384
mass confirmed to be cardiac papillary fibroelastoma | 384
MSSA bacteremia | 384
culture of the PFE revealed Streptococcus salivarius | 384
culture of the PFE revealed Rothia spp | 384
source of MSSA infection suggested to be the skin | 384
treated with linezolid | 384
treated with meropenem | 384
follow-up blood cultures resulted in no bacterial growth | 384
opted to pursue comfort care | 480
elected to continue care under hospice services | 480
overall functional decline from multisystem organ failure | 480
discharged to hospice | 480
no relationships relevant to the contents of this paper to disclose | 480
