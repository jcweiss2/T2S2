44 years old | 0
male | 0
alcoholic liver cirrhosis | -672
decompensated liver cirrhosis | -672
chronic left leg wound | -672
chronic thrombocytopenia | -672
anemia of chronic disease | -672
portal hypertensive gastropathy | -672
esophageal varices grade 1 | -672
recurrent ascites | -672
low total protein ascites | -672
admitted to the hospital | 0
worsening jaundice | 0
diffuse abdominal pain | 0
subjective fevers | 0
progressive erythema in left leg | 0
dull right shoulder pain | 0
denies recent trauma | 0
denies prolonged immobilization | 0
regular bowel movements | 0
denies insomnia | 0
denies confusion | 0
resided in Wisconsin | 0
lived with one dog | 0
lived with three cats | 0
no animal bites | 0
no animal scratches | 0
temperature 38.4 | 0
blood pressure 160/65 | 0
heart rate 114 | 0
respiratory rate 22 | 0
oxygen saturation normal | 0
alert | 0
pale | 0
icteric | 0
distressed due to abdominal pain | 0
mucous membranes dry | 0
neck supple | 0
no neck rigidity | 0
heart exam normal | 0
lung exam normal | 0
abdomen distended | 0
positive ascitic wave | 0
diffuse tenderness to palpation | 0
no guarding | 0
no rebound | 0
bilateral pitting edema | 0
open wound with yellowish secretion | 0
surrounding erythema | 0
distal pulses palpable | 0
right shoulder non-tender | 0
no limitation for flexion and extension | 0
hemoglobin 9.3 | 0
platelet count 86 | 0
leukocytosis 17.0 | 0
neutrophilia | 0
lactic acid 6.5 | 0
ammonia 43 | 0
INR 2.2 | 0
C-reactive protein 45.5 | 0
magnesium 2.2 | 0
potassium 5.2 | 0
sodium 136 | 0
bicarbonate 14 | 0
anion gap 20 | 0
creatinine 1.19 | 0
glucose 93 | 0
AST 66 | 0
ALT 26 | 0
alkaline phosphatase 48 | 0
total serum protein 6.5 | 0
serum albumin 3.0 | 0
LDH 273 | 0
total bilirubin 5.1 | 0
lipase 18 | 0
SARS-Coronavirus-2 PCR negative | 0
urinalysis negative for infection | 0
ascitic fluid yellow cloudy | 0
total nucleated cells 20,375 | 0
neutrophils 86% | 0
lymphocytes 14% | 0
LDH 86 | 0
total protein 1.0 | 0
albumin 0.5 | 0
glucose 61 | 0
amylase 20 | 0
Gram stain no organisms | 0
CT abdomen and pelvis negative | 0
chest x-ray no infiltrates | 0
x-ray left tibia and fibula soft tissue edema | 0
ultrasound left lower extremity no deep venous thrombosis | 0
treated with IV fluids | 0
treated with Ceftriaxone | 0
treated with Vancomycin | 0
admitted to ICU | 0
diagnosis of sepsis | 0
received IV albumin | 24
blood cultures grew Pasteurella multocida | 24
ascitic fluid culture grew Pasteurella multocida | 24
abdominal pain improved | 48
afebrile | 48
right shoulder pain | 72
limitation for flexion and extension | 72
MRI right shoulder osteolytic change | 72
edema at AC joint | 72
septic arthritis | 72
debridement and irrigation of right shoulder | 96
acute osteomyelitis | 96
purulence and necrotic tissue | 96
abdominal pain improved | 120
right shoulder pain improved | 120
discharged to rehabilitation facility | 336
antibiotic therapy | 336
SBP prophylaxis | 336