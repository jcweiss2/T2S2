21 months old | 0
female | 0
admitted to secondary care hospital | -744
isolated fever | -744
treated as bacterial pulmonary infection | -744
discharged | -720
put on long-term course of oral antibiotics | -720
presented to health facility with worsening abdominal pain | -672
fever | -672
abdominal ultrasound | -672
angio-computed tomography (CT) | -672
abdominal aortic aneurysm (AAA) measuring 40 mm in diameter | -672
referred to hospital for surgical management | -672
admitted to hospital | 0
hemodynamic shock | 0
pale | 0
tachycardiac | 0
hypotensive | 0
admitted to intensive care unit | 0
emergency CT scan | 0
ruptured infrarenal aortic aneurysm | 0
giant retroperitoneal hematoma | 0
underwent urgent surgery | 0
surgical exploration | 0
giant AAA compressing on approximate organs | 0
signs of inflammation and rupture | 0
aorta ligated below the origin of the renal arteries | 0
aorta ligated above the iliac bifurcation | 0
collateral circulation verified on angio-CT | 0
aortic aneurysm sac resected | 0
abdominal cavity rinsed and closed | 0
put on intravenous (IV) antibiotics | 0
amoxicillin | 0
clavulanic acid | 0
gentamicin | 0
anemia | 0
hemoglobin at 10.5 mg/dL | 0
white blood cell count at 30,000 cells/µL | 0
erythrocyte sedimentation rate at 52 mm/hh | 0
C-reactive protein at 142.78 mg/L | 0
electrocardiography (EKG) normal | 0
echocardiography showed no signs of endocarditis | 0
postoperative angio-CT | 24
persistent retroperitoneal hematoma | 24
no signs of lower limb ischemia | 24
hypertension | 24
treated with beta-blockers | 24
treated with angiotensin-converting enzyme (ACE) inhibitors | 24
treated with calcium channel blockers (CCBs) | 24
discharged home | 432
put on pain medication | 432
put on beta-blockers for 3 months | 432
pathologic examination of aortic tissue | 432
inflammatory signs with suppuration | 432
mycotic aneurysm | 432
microbiological cultures of aortic tissue sterile | 432
blood cultures sterile | 432