70 years old | 0
female | 0
gastric malignancy | 0
oxaliplatin | -84
tiggio | -84
sintilimab | -240
erythematous maculopapular rash | -240
methylprednisolone | -228
rash deterioration | -225
new rashes | -225
blistering | -225
skin denudation | -225
outpatient clinic visit | -225
systemic widespread rashes | -225
epidermolysis | -225
Nikolsky’s sign | -225
epidermal detachment | -225
palpation tenderness | -225
TEN diagnosis | -225
refused treatment | -225
refused hospitalization | -225
intravenous immunoglobulin | -222
no improvement | -219
adalimumab | -216
rash resolution | -192
no new epidermal detachment | -192
no new bullae | -168
negative Nikolsky’s sign | -168
body temperature 37°C | -168
bullae scabbed | -120
skin lesions subsided | -120
desquamation | -120
adalimumab again | -120
follow-up visit | 45
no rash recurrence | 45
discharged | 0