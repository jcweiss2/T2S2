84 years old | 0
male | 0
admitted to the hospital | 0
chronic constipation | -8760
referred to gastroenterologist | -8760
scheduled for diagnostic barium enema | -24
barium enema | 0
lower abdominal discomfort | 0
pain during barium enema | 0
vague pain in lower abdomen | 0
increased pain during procedure | 0
history of chronic heart failure | 0
history of atrial fibrillation | 0
stable and normal vital signs | 0
generalized abdominal tenderness | 0
rebound tenderness in hypogastric region | 0
loose, bloody stool | 0
digital rectal exam | 0
emergent supine plain abdominal x-ray | 0
contrast extravasation | 0
rectal perforation | 0
barium extravasation | 0
adequate fluid replacement | 0
resuscitation | 0
prophylactic antibiotics | 0
emergent exploratory laparotomy | 2
midline incision | 2
no visible perforation in distal colon | 2
no visible perforation in sigmoid and upper rectum | 2
barium on posterior wall of peritoneum | 2
barium around sigmoid mesocolon and mesoileum | 2
barium penetration into intraperitoneal cavity | 2
barium extraction | 2
massive irrigation and lavage | 2
diverting ileostomy | 2
tissue sample from mesenteric tissue | 2
fat necrosis | 2
foreign-body reaction | 2
broad-spectrum intravenous antibiotics | 2
intensive care unit | 2
signs and symptoms of sepsis | 48
rigid proctoscopy | 48
massive inflammation and blood clots on posterior wall of rectum | 48
open, corrugated, presacral drain | 48
general condition improved | 120
sepsis resolved | 120
generalized abdominal pain | 336
high fever | 336
abdominopelvic computed tomography scan | 336
extensive hyperdense area within retroperitoneal space | 336
second laparotomy | 336
massive dissemination of barium | 336
barium up to inferior pole of both kidneys | 336
barium in mesentery of colon and small intestine | 336
retroperitoneal tissues fragile and inflamed | 336
proper irrigation | 336
massive debridement of necrotic tissues | 336
two open, corrugated drains | 336
stable vital signs | 432
fever disappeared | 432
regained appetite | 432
presacral and abdominal drains removed | 432
oral diet | 432
discharged | 480
referred to stoma care center | 480
biweekly visits | 480
diversion ileostomy closed | 1344
monthly visits | 1344
bimonthly visits | 1344
normal life | 1344
x-rays show residual barium | 1752
good general and health condition | 1752