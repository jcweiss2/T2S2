5 years old | 0
male | 0
weight 20 kg | 0
admitted to the hospital | 0
scheduled for emergency craniotomy | 0
decompression of right parieto-occipital glioma | 0
Glasgow coma scale (GCS) of E2 V2 M3 | 0
bilateral crackles | 0
sensorium worsening | -72
weakness of the left side of the body | -72
operated 3 months earlier | -2160
lost to follow-up | -2160
presented to the neurosurgery outpatient department | -72
blood grouping and cross matching performed | 0
blood products arranged | 0
sedative premedication not given | 0
fentanyl 40 mcg intravenously | 0
injection thiopental 100 mg intravenously | 0
loss of eye lash reflex | 0
bag-mask ventilation confirmed | 0
vecuronium 2 mg intravenously | 0
trachea intubated | 0
arterial line placed in the left radial artery | 0
central line deferred | 0
venous access attained through two peripheral veins | 0
Foley's catheter inserted | 0
anesthesia maintained with oxygen and air mixture | 0
isoflurane and vecuronium | 0
propofol infusion started | 0
noncontrast computed tomography showed significant midline shift and edema | 0
baseline arterial blood gas done | 0
Mannitol 100 ml given | 0
furosemide 10 mg intravenously | 0
phenytoin given | 0
dexamethasone given | 0
antibiotics given | 0
surgery lasted 3 h | 180
total blood loss 400 ml | 180
crystalloids replaced | 180
200 ml of packed red blood cells transfused | 180
central venous access attempted | 180
subclavian approach attempted | 180
guidewire not inserted into the subclavian vein | 180
internal jugular vein (IJV) approach attempted | 180
guidewire inserted | 180
no ECG changes | 180
free flow of blood from two ports | 180
line secured with sutures | 180
patient shifted to ICU | 180
chest X-ray advised | 180
central venous line totally out of place | 180
no evidence of pneumothorax | 180
line removed | 180
Triple lumen B Braun Central Line inserted through the left IJV | 24
postoperative course marked by cardiovascular instability | 24
sepsis | 24
patient recovered well | 240
removed from ventilatory support | 240
shifted to the surgical ward | 336