76 years old | 0
female | 0
admitted to the hospital | 0
dyspnea | 0
cerebrovascular disease | -8760
inability to ambulate | -8760
hypertension | -6480
type 2 diabetes mellitus | -6480
subarachnoid hemorrhage | -6120
endobronchial tuberculosis | -5040
intracerebral hemorrhage | -1440
pneumonia | -1440
recovered from pneumonia | -1440
blood pressure 140/54 mmHg | 0
pulse rate 90 beats/min | 0
body temperature 36.1°C | 0
respiratory rate 14 breaths/min | 0
crackle breathing sounds | 0
indwelling urinary catheter | 0
white blood cell count 361,000/µL | 0
hemoglobin level 7.2 g/dL | 0
platelet count 76×103/µL | 0
C-reactive protein level 41.7 mg/L | 0
blood urea nitrogen 61 mg/dL | 0
creatinine 0.8 mg/dL | 0
Na 130 mEq/L | 0
total protein 3.4 g/dL | 0
albumin 2.2 g/dL | 0
pro B-natriuretic peptide 3,669 pg/mL | 0
arterial blood gas analysis | 0
pH level 7.3999 | 0
arterial carbon dioxide partial pressure 53.1 mmHg | 0
arterial oxygen partial pressure 61.9 mmHg | 0
peripheral oxygen saturation 99% | 0
fractional inspired oxygen 60% | 0
Candida tropicalis in blood culture | 0
Candida tropicalis in urine culture | 0
Klebsiella pneumoniae in sputum culture | 0
pneumonia | 0
acute respiratory failure | 0
candidemia | 0
meropenem treatment | 0
colistimethate sodium treatment | 0
fluconazole treatment | 0
high-flow nasal cannula oxygen therapy | 0
flexible bronchoscopy | 24
narrowing of the right main bronchus | 24
anthracotic pigmentation | 24
bronchial washing | 24
acid-fast bacilli staining | 24
Mycobacterium tuberculosis PCR | 24
cytology | 24
worsening hypoxia | 33
dyspnea | 33
endotracheal intubation | 33
mechanical ventilation | 33
urinalysis | 72
microscopic hematuria | 72
urine cytology test | 72
HSV serology | 72
IgM negative | 72
IgG positive | 72
HSV type 1-positive cells | 168
intranuclear inclusions | 168
multinucleation | 168
acyclovir treatment | 168
repeat bronchoscopy | 168
percutaneous dilatational tracheostomy | 168
HSV type 1-infected cells in urine cytology | 168
absence of HSV infection in urine cytology | 336
stable vital signs | 336
no fever | 336
white blood cell count 4,400/µL | 336
hemoglobin level 8.6 g/dL | 336
platelet count 65×103/µL | 336
C-reactive protein level 78.1 mg/L | 336
stable right upper lobe atelectasis | 336
vancomycin-resistant Enterococci in urine culture | 480
vancomycin-resistant Enterococci in stool culture | 480
sepsis | 480
linezolid treatment | 480
decreased urine output | 480
acute renal failure | 480
refused hemodialysis | 480
refused cardiopulmonary resuscitation | 480
death | 672