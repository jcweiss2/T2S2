26 years old | 0
male | 0
admitted to the hospital | 0
height: 180 cm | 0
weight: 74 kg | 0
kidney transplant | -5916
end-stage kidney disease | -8784
immunosuppression | 0
mycofenolate sodium | 0
methylprednisolone | 0
estimated glomerular filtration rate (eGFR) 35.9 mL/min/1.73 m2 | 0
proteinuria 117 mg/d | 0
chronic kidney transplant disease stage 3bA1 | 0
status post vascular rejection | -5916
chronic calcineurin-inhibitor toxicity | -5916
new-onset headache | 0
blurred vision | 0
cranial CT- and MRI scans | 0
several contrast-enhancing intracerebral lesions | 0
perifocal edema | 0
methylprednisolone therapy stopped | 0
dexamethasone administered | 0
brain edema | 0
transmitted to the university department of Nephrology | 24
transmitted to the department of Neurosurgery | 48
brain biopsy | 72
diagnosis of cerebral PTLD | 72
diffuse large B-cell lymphoma | 72
positive for Ebstein-Barr virus | 72
initial chemotherapy regime | 120
high-dose cytarabin | 120
Rituximab | 120
MRI scan confirmed complete remission of PTLD | 240
impairment of the transplant function aggravated | 240
eGFR 25.4 mL/min/1.73 m2 | 240
cytomegalovirus (CMV) reactivated | 672
pneumocystis jirovecii pneumonia | 672
chemotherapy changed to Rituximab | 672
antiviral and antibiotic therapy | 672
dose of mycofenolate sodium tapered | 672
generalized seizure | 960
cerebral MRI scan demonstrated the recurrence of PTLD | 960
HDMTX administered | 960
Leukovorine administered | 960
Rituximab administered | 960
vigorous hydration | 960
alkalinization of the urine | 960
HFHD started | 984
dialysis procedures | 984
MTX-level measurements | 984
nadir of leucocytes | 1008
severe CMV- and E.coli pneumonia | 1056
sepsis | 1056
acute kidney transplant failure | 1056
transmission to an intensive care unit | 1056
invasive ventilation | 1056
sepsis managed | 1080
follow-up cerebral MRI scan | 1104
small regredience of PTLD | 1104
cerebral radiation | 1104
no relevant response of the disease | 1128
dialysis sessions | 984
Gambro machine AK 200 | 984
high-flux dialyser | 984
dialysate SelectBag One AX 450 G | 984
unfractionated heparin | 984
MTX-level measurements | 984
fluorescence polarization immunoassay | 984
TDx analyser | 984
HFHD for MTX elimination | 984
successful elimination of MTX | 1104
no significant rebound of MTX level | 1104
no changes in the estimated glomerular filtration rate | 1104
hematological toxicities limited | 1104
leucocytes dropped to 1.1/nL | 1008
no granulocyte colony-stimulating factor required | 1008
preexisting anemia did not impair significantly | 1008
no changes in the number of thrombocytes | 1008
infection developed | 1056
leucopenia | 1008
CMV-colonization | -5916
frequent relapses of CMV-activation | -5916
high risk of a new CMV reactivation | 0
posttransplant immunosuppressive therapy | 0
impaired kidney function | 0
rituximab | 0
contribution to the development of the infection | 1056
unique case | 0
HDMTX in a patient with a preliminary significantly impaired kidney function | 0
feasibility of administering HDMTX | 0
add-on HFHD for MTX clearance | 984
no major hematological toxicity | 1104
no onset of an acute on chronic kidney failure | 1104
limited evidence of a successful elimination of MTX with HFHD | 1104
administration of HDMTX did not achieve a remission of PTLD | 1128
ultima ratio | 960
last chemotherapy option | 960
recurrent PTLD | 960
administration of HDMTX possible in a transplant kidney with already preliminary impaired function | 960
comorbidities limit tolerance of an aggressive therapy | 0
question about the right time to start the dialysis after HDMTX administration | 0
question about the appropriate duration of dialysis sessions | 0
requires further research | 0