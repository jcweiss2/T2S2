76 years old | 0
female | 0
admitted to the hospital | 0
sore throat | -288
dry cough | -288
fever | -288
diabetes mellitus | 0
hypertension | 0
glaucoma | 0
smoker | 0
visited Japan | -672
arrived at Yokohama Harbor | -672
aboard the Diamond Princess cruise ship | -672
COVID-19 outbreak | -672
quarantine inspection | -672
RT-PCR test | -288
positive result for SARS-CoV-2 | -288
lopinavir-ritonavir | -24
moxifloxacin | -24
transferred to hospital | 0
body temperature 38.3 °C | 0
oxygen saturation 93% | 0
coarse crackles in the upper chest | 0
peripheral blood lymphopenia | 0
elevated BUN | 0
elevated creatinine | 0
elevated CRP | 0
elevated LDH | 0
chest CT scan | -216
ground-glass opacities | -216
consolidation | -216
piperacillin-tazobactam | 0
peramivir | 0
endotracheal intubation | 24
endotracheal aspirate positive for SARS-CoV-2 | 24
intravenous immune globulin | 72
low gamma-globulin level | 72
respiratory failure | 168
dyspnea | 168
fever alleviation | 168
venous-venous extracorporeal membrane oxygenation | 168
compression ultrasound | 168
deep vein thrombosis | 168
ventilator settings | 168
PaO2/FiO2 | 168
vancomycin | 240
viral testing negative | 240
tracheotomy | 264
ECMO discontinued | 288
intravenous meropenem | 288
ventilator-associated pneumonia prophylaxis | 288
chest CT scan | 312
organizing pneumonia | 312
methylprednisolone | 360
improvement of organizing pneumonia | 360
taken off respirator | 480
condition stable | 480