71 years old | 0
male | 0
Taiwanese | 0
admitted to the hospital | 0
nocturia | -1728
incomplete voiding | -1728
digital rectal examination | 0
enlarged prostate | 0
no hard nodule | 0
urinalysis | 0
negative for pyuria | 0
negative for haematuria | 0
prostate-specific antigen level | 0
7.845 ng/ml | 0
TRUS-measured prostate volume | 0
64 ml | 0
biopsy | 0
5-alpha reductase inhibitor | -24
mandatory cessation of anticoagulants | -24
cleansing of the rectum | -24
antibiotic consumption | -24
Levofloxacin | -24
750 mg | -24
TRUS | 0
homogenous echogenicity | 0
no hypoechoic lesions | 0
twelve core prostatic tissue samples | 0
gross haematuria | 0
Foley catheter | 0
fever | 24
backache | 24
severe myalgia | 24
right thigh | 24
temperature | 24
38.5°C | 24
heart rate | 24
103 beats/minute | 24
respiratory rate | 24
18 counts/minute | 24
blood pressure | 24
107/63 mmHg | 24
tender prostate | 24
leucocytosis | 24
white blood cell count | 24
9550/μl | 24
neutrophil predominance | 24
neutrophil | 24
94% | 24
elevated C-reactive protein | 24
23.36 mg/dl | 24
elevated procalcitonin | 24
23.3 ng/ml | 24
pyuria | 24
white blood cells | 24
>100/high power field | 24
prostatitis | 24
sepsis | 24
ceftriaxone | 24
2 g | 24
once-daily intravenous | 24
shortness of breath | 72
intensive care unit | 72
plain radiography | 72
lumbar spine | 72
computed tomography | 72
abdomen | 72
narrowing of the L3–L5 vertebrae | 72
cystic lesion | 72
3.3 cm | 72
right psoas muscle | 72
percutaneous approach | 72
magnetic resonance imaging | 120
lumbar spine | 120
abscesses | 120
L3/4 intervertebral disc spaces | 120
L4/5 intervertebral disc spaces | 120
narrow enhancement | 120
L3–L5 vertebral bodies | 120
abnormally enhanced lesions | 120
psoas muscles | 120
spiking fever | 120
39°C | 120
chills | 120
Escherichia coli | 120
blood culture | 120
multiple drug resistance | 120
urine culture | 120
resistant | 120
cefazolin | 120
ciprofloxacin | 120
levofloxacin | 120
susceptible | 120
flomoxef | 120
piperacillin–tazobactam | 120
cefepime | 120
doripenem | 120
imipenem | 120
doripenem | 144
0.25 g | 144
intravenous | 144
three times daily | 144
total laminectomies | 168
L4/L5 vertebrae | 168
removal of the epidural abscesses | 168
pathology | 168
chronic inflammation | 168
spine | 168
epidural tissue | 168
discharged | 168
seventh postoperative day | 168
normal activities | 168