65 years old | 0
male | 0
hypertension | -86400
persistent atrial fibrillation | -86400
antiarrhythmic drug therapy | -86400
catheter-based radiofrequency pulmonary vein isolation procedure | 0
irritative cough | 336
cough attributed to respiratory origin | 336
severe headache | 504
persistent cough | 504
fever | 504
awake | 504
unremarkable vital signs except fever | 504
incessant cough | 504
cough exacerbating when speaking | 504
leukocytosis (21,000 cells/mL) | 504
subarachnoid hemorrhage | 504
excessive coughing on anticoagulant therapy | 504
admitted to intensive care unit | 504
warfarin withheld | 504
broad-spectrum antibiotics | 504
shortness of breath | 504
transthoracic echocardiography ordered | 504
bubbles in left ventricle | 504
bubbles in left atrium | 504
air within heart | 504
communication with esophagus or bronchial tree | 504
decline in consciousness level | 504
cerebral air emboli | 504
mechanical ventilation | 504
endotracheal tube placed in right main bronchus | 504
upper endoscopy | 504
large clot on distal esophageal wall | 504
atrioesophageal fistula | 504
covered stent placed | 504
condition worsening | 504
cardiac arrest | 504
coronary artery air embolization | 504
resuscitation attempts | 504
pronounced dead | 504
autopsy confirming 3mm fistula | 504
