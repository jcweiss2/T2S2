70 years old | 0
male | 0
admitted to the hospital | 0
sudden and severe loss of vision | -96
eye pain | -96
conjunctival injection | -96
swelling | -96
consumed oral diclofenac | -144
viral prodrome | -144
rashes all over the body | -120
oral mucosal ulcerations | -120
macular rash over upper torso | 0
ulcerating lesions over buccal and perioral tissue | 0
diagnosis of toxic epidermal necrolysis (TEN) | 0
supportive treatment initiated | 0
extreme conjunctival congestion | 0
corneal sloughing | 0
corneal thinning | 0
severe anterior chamber reaction | 0
hypopyon | 0
amniotic membrane transplant planned | 0
topical moxifloxacin started | 0
lubricants started | 0
corneal perforation | 2
uveal prolapse | 2
mild proptosis | 2
lid edema | 2
restricted extraocular muscles | 2
systemic steroids started | 2
electrolytes started | 2
antibiotics started | 2
evisceration in both eyes | 24
patient died | 72
multi-organ failure | 72
eviscerated material sent for microbiological examination | 24
blood culture sent for microbiological examination | 24
no bacterial growth | 72