26 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
otherwise healthy | 0 | 0 | Factual
referred to the department | -72 | -72 | Factual
rising levels of human chorionic gonadotropin | -72 | -72 | Factual
intermittent vaginal bleeding | -72 | -72 | Factual
vaginal ultrasound scan | -72 | -72 | Factual
intrauterine pregnancy | -504 | -504 | Factual
legal medical abortion | -504 | -504 | Factual
placental remnants in the uterus | -72 | -72 | Factual
surgical evacuation of the uterus | 0 | 0 | Factual
discharged | 12 | 12 | Factual
readmitted | 24 | 24 | Factual
temperature of 39.5°C | 24 | 24 | Factual
abdominal pain | 24 | 24 | Factual
severe endometritis | 24 | 24 | Possible
metronidazole | 24 | 48 | Factual
benzylpenicillin | 24 | 48 | Factual
gentamicin | 24 | 48 | Factual
deteriorated | 48 | 48 | Factual
saturation fell to 90% | 48 | 48 | Factual
respiratory rate rose to around 40 breaths per minute | 48 | 48 | Factual
oxygen given by mask | 48 | 48 | Factual
temperature peaked at 40.7°C | 48 | 48 | Factual
C-reactive protein rose to around 300 mg/L | 48 | 48 | Factual
leukocytes to around 15 × 10^9/L | 48 | 48 | Factual
moved to the intensive care unit | 48 | 48 | Factual
intubated | 48 | 48 | Factual
CT scan | 72 | 72 | Factual
thrombophlebitis of the internal jugular vein | 72 | 72 | Factual
hepatomegaly | 72 | 72 | Factual
diagnosed with Lemierre's syndrome | 72 | 72 | Factual
benzylpenicillin and gentamicin discontinued | 72 | 72 | Factual
tazocin and clindamycin administered | 72 | 336 | Factual
metronidazole administered | 72 | 336 | Factual
heparin injections | 72 | 336 | Factual
recovered | 336 | 336 | Factual
discharged | 504 | 504 | Factual
infection with F. necrophorum | -72 | 504 | Factual
blood cultures showed infection with F. necrophorum | 72 | 72 | Factual
F. necrophorum cultivated from the patient's cervix | 72 | 72 | Factual
infection originated from the cervix | 72 | 72 | Factual
no symptoms from the oropharyngeal tract | 0 | 504 | Factual