13 years old | 0
male | 0
admitted to the hospital | 0
near-drowning event | -1800
cardiac arrest | -1800
severe aspiration pneumonia | -1800
acute respiratory failure | -1800
acute renal failure | -1800
ventilator support | -1800
extracorporeal membrane oxygenation | -1800
continuous renal replacement therapy | -1800
Acinetobacter baumannii | -1800
Elizabethkingia meningoseptica | -1800
methicillin-resistant Staphylococcus aureus | -1800
antibiotics | -1800
weaned from ventilator | -720
improvement of pneumonia | -720
transferred to general ward | -720
poor oral intake | -720
nausea | -720
general weakness | -720
mental confusion | -480
disorientation | -480
magnetic resonance imaging (MRI) scan | -480
brain MRI scan | -480
contrast-enhancing lesion | -480
cerebrospinal fluid (CSF) examination | -480
red blood cell (RBC) | -480
white blood cell (WBC) | -480
protein | -480
glucose | -480
CSF culture | -480
brain abscess | -480
ventriculitis | -480
antibiotics | -480
vancomycin | -480
cefotaxime | -480
metronidazole | -480
Cotrim | -480
amphotericin B | -480
mental confusion improved | -336
intravenous antibiotics | -336
follow-up MRI | -336
surrounding edema | -336
enhancement of left lateral ventricle | -336
ventriculitis | -336
antibiotic regimen changed | -336
voriconazole | -336
meropenem | -336
Cotrim | -336
CSF culture | -336
stereotactic biopsy | 0
greenish-yellow pus | 0
hyphae | 0
S. apiospermum | 0
intravenous antibiotics | 0
voriconazole | 0
isoconazole | 0
amphotericin B | 0
follow-up MRI | 168
diffuse contrast enhancement | 168
dilation of left lateral ventricle | 168
aggravation of edema | 168
extraventricular drainage | 168
CSF drainage | 168
voriconazole injection | 336
intraventricular injection | 336
drowsy | 360
emergent MRI | 360
acute hydrocephalus | 360
septations | 360
mannitol treatment | 360
alert | 360
minimal headache | 360
repeated EVD | 384
endoscopic septostomy | 384
occipital burr-hole trephination | 384
alert | 384
stable vital signs | 384
sudden hypotension | 408
respiratory distress | 408
acute septic shock | 408
transferred to ICU | 408
expired | 420