13 years old | 0
    female | 0
    admitted to the hospital | 0
    difficult-to-control seizures | 0
    worsening of handwriting | -72
    involuntary, repetitive pill"rolling hand movements | -72
    focal seizures | -72
    generalized tonic-clonic seizures | -72
    facio-brachial dystonic seizures | -72
    periods of agitation | -72
    unresponsiveness | -72
    mutism | -72
    lucid between episodes | -72
    attempting to form words | -72
    no speech production | -72
    bruxism | -72
    dystonic posturing | -72
    full body rigidity | -72
    opisthotonic posturing | -72
    insomnia | -72
    appeared afraid | -72
    agitation | -72
    cried abnormally | -72
    cried spontaneously | -72
    brisk reflexes | -72
    unsustained clonus bilaterally | -72
    waxy catatonia | -72
    opsoclonus | -72
    high-grade fever | 240
    deteriorated sensorium | 240
    orofacial dyskinesia | 240
    autonomic instability | 240
    irregular respiration | 240
    sepsis | 240
    urinary tract infection | 240
    colitis | 240
    modified Rankin Scale score 5 | 240
    normal hemogram | 240
    normal liver function tests | 240
    normal renal function tests | 240
    normal serum electrolytes | 240
    normal thyroid function | 240
    normal viral markers | 240
    normal initial MRI Brain | 240
    normal repeat MRI Brain | 240
    electroencephalogram delta slowing in left hemispheric regions | 240
    normal cerebrospinal fluid cell count | 240
    normal cerebrospinal fluid sugar | 240
    normal cerebrospinal fluid protein | 240
    negative Herpes Simplex virus in CSF | 240
    negative Japanese Encephalitis virus in CSF | 240
    negative serum antinuclear antibody | 240
    no evidence of malignancy on Chest X-ray | 240
    no evidence of malignancy on CECT abdomen | 240
    no evidence of malignancy on ultrasound pelvis | 240
    no evidence of malignancy on skeletal survey X-rays | 240
    tumor markers not done | 240
    empirical Acyclovir started | 240
    multiple antiepileptic drugs | 240
    anti-NMDAR antibody detected | 240
    intravenous methylprednisolone started | 240
    intravenous immunoglobulins started | 240
    oral prednisolone started | 240
    symptoms improvement | 672
    modified Rankin Scale score 4 | 672
    continued improvement on oral prednisolone | 672
    antiepileptic drugs tapered | 672
    modified Rankin Scale score 1 | 2880
    amnesia | 2880
    mild language disintegration | 2880
    occasional agitation | 2880
    advised regular follow-up | 2880
    advised repeat ultrasound/MRI abdomen and pelvis | 2880
    advised screening by tumor markers | 2880
    subacute onset AED resistant seizures at 5 years old | -70080
    abnormal behavior at 5 years old | -70080
    abnormal body movements at 5 years old | -70080
    normal routine investigations at 5 years old | -70080
    unremarkable CSF analysis at 5 years old | -70080
    normal MRI Brain at 5 years old | -70080
    remission of seizures after 3 months | -70080
    remission of abnormal movements after 3 months | -70080
    gradual recovery | -70080
    no immunotherapy recorded | -70080
    fully functional before second attack | -70080
    second attack eight years later | 0
    