79 years old | 0
female | 0
medial femoral neck fracture | -144
low energy trauma | -144
emergency department presentation | 0
right hip pain | 0
arterial hypertension | 0
hypothyreosis | 0
cataract |,0
macular degeneration | 0
hypacusis | 0
multiple eye and hand operations | 0
soft abdomen | 0
no abdominal tenderness | 0
regular peristaltic sounds | 0
dual head prosthesis implantation | 24
postoperative regular course | 24
hemodynamic instability | 144
decreasing hemoglobin levels | 144
serum lactate levels progression | 144
vasopressor dependency | 144
intubation | 144
blood transfusion | 144
free intraabdominal fluid | 144
large intraperitoneal hematoma | 144
suprasplenic coagulum | 144
pleural effusion | 144
pericardial effusion | 144
emergency splenectomy | 144
respiratory failure | 168
pneumonia | 168
septic shock | 168
multiple organ failure | 168
death | 648
