73 years old | 0
male | 0
admitted to the hospital | 0
diabetes mellitus | -8760
Parkinsonism | -8760
trans-urethral resection of the prostate | -8760
laparoscopic cholecystectomy | -105120
dysphagia for solid food | -720
type II achalasia | -720
manometry | -720
water-soluble studies | -720
endoscopic pneumatic dilatation | -120
symptoms worsened | -24
endoscopic pneumatic dilatation | 0
general anesthesia | 0
endotracheal intubation | 0
left lateral position | 0
Rigiflex dilator | 0
gastroesophageal junction dilated | 0
desaturation | 0
esophageal perforations | 0
plain chest radiography | 0
left-sided pneumothorax | 0
pneumomediastinum | 0
chest tube inserted | 0
oxygen saturation improved | 0
thoracic and upper gastrointestinal surgical teams involved | 0
diagnostic laparoscopy | 0
primary esophageal repair attempted | 0
esophageal mucosa dissected | 0
mucosa showed multiple linear tears | 0
unhealthy edges | 0
double-tract reconstruction decided | 0
distal esophagus transected | 0
esophagostomy created | 0
proximal gastrectomy | 0
jejunal loop measured | 0
end-to-side jejuno-jejunostomy | 0
mesenteric defect closed | 0
size 25 circular stapler introduced | 0
anvil and stapler aligned | 0
circular stapler fired | 0
gastrostomy and jejunostomy created | 0
side-to-side gastro-jejunostomy | 0
Blake drain inserted | 0
patient transferred to ICU | 0
extubated | 24
shifted to regular ward | 24
intravenous fluids | 24
nil per os | 24
broad-spectrum antibiotics | 24
antifungal drugs | 24
clear liquid diet | 120
water-soluble study | 120
GI tract continuity confirmed | 120
anastomotic leakage excluded | 120
discharged | 192
follow-up | 4320