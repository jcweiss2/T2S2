54 years old | 0
male | 0
admitted to University of Texas Medical Branch | 0
work up of newly diagnosed acute myeloid leukemia | 0
prostate cancer | -672
hepatitis C virus | -672
non-insulin dependent diabetes mellitus | -672
hypertension | -672
initiation of chemotherapy | 24
neutropenic fevers | 48
pneumonia | 72
respiratory distress requiring intubation | 72
septic shock | 72
blood cultures revealed Serratia marcescens | 72
treated with vancomycin | 72
treated with pipercillin-tazobactam | 72
prophylactic acyclovir | 72
prophylactic fluconazole | 72
condom catheter placed | 72
extubated | 168
condom catheter removed | 168
penile pain | 168
lesion seen | 168
Urology consulted | 528
genitourinary exam | 528
blackened scrotum | 528
penile shaft with crepitus and eschars | 528
Fournier's gangrene | 528
genitourinary debridement | 528
left orchiectomy | 528
left hemiscrotectomy | 528
post-operative stable and afebrile | 552
altered mental status | 552
episodes of confusion | 552
quantitative analysis returned positive for zygomycetes | 592
started on systemic liposomal Amphotericin B | 592
wound mottled with paucity of granulation tissue | 592
second debridement | 592
right orchiectomy | 592
suprapubic tube placement | 592
penectomy | 592
groin debridement | 592
Burn team consulted | 592
amphotericin soaked dressing changes | 592
amphotericin bladder irrigation | 592
third debridement | 624
hypotensive | 784
tachycardic | 784
febrile | 784
green growth on groin | 784
further debridement scheduled | 784
patient's condition worsened | 816
patient's demise | 816