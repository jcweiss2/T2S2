22 years old | 0
    Afghan migrant worker | 0
    male | 0
    admitted to emergency room | 0
    dysphagia | -168
    chest pain | -168
    fever | -168
    chills | -168
    low BMI (16) | 0
    symptoms started 7 days prior to presentation | -168
    worsening symptoms | -168
    prolonged fever | -4320
    weight loss | -4320
    dealing with suspected TB patient | -4320
    febrile | 0
    tachycardic (130/min) | 0
    tachypneic (28/min) | 0
    oxygen saturation 89% | 0
    chest X-ray showing left pleural effusion | 0
    CT scan showing left pleural effusion | 0
    pneumothorax | 0
    pneumomediastinum | 0
    extraluminal contrast in mediastinum | 0
    distal esophageal perforation | 0
    chest tube insertion | 0
    purulent fluid (700 cc) | 0
    aggressive resuscitation | 0
    emergent thoracotomy | 0
    large perforation in distal esophagus | 0
    esophagectomy | 0
    cervical esophagostomy | 0
    gastrostomy | 0
    transfer to surgical ICU | 0
    persistent septic shock | 0
    multi-organ failure | 0
    death | 96
    PCR detection of mycobacterial DNA in pleural fluid | 0
    histopathologic confirmation of TB in esophagus | 0
    esophageal TB diagnosis | 0
    perforation | 0
    septic shock | 0
    no recent upper endoscopy | 0
    no underlying mucosal damage | 0
    no response to conventional antibiotics | 0
    surgical intervention | 0
    no delay in diagnosis beyond 24 hours | 0
    TB coverage antibiotics initiated | 0
    informed consent obtained | 0
    <|eot_id|>
    
  - fever |-168
  - chills |-168
  - chest pain |-168
  - dysphagia |-168
  - weight loss |-4320
  - prolonged fever |-4320
  - dealing with suspected TB patient |-4320
  - symptoms started 7 days prior to presentation |-168
  - low BMI (16) |0
  - admitted to emergency room |0
  - febrile |0
  - tachycardic (130/min) |0
  - tachypneic (28/min) |0
  - oxygen saturation 89% |0
  - chest X-ray showing left pleural effusion |0
  - CT scan showing left pleural effusion |0
  - pneumothorax |0
  - pneumomediastinum |0
  - extraluminal contrast in mediastinum |0
  - distal esophageal perforation |0
  - chest tube insertion |0
  - purulent fluid (700 cc) |0
  - aggressive resuscitation |0
  - emergent thoracotomy |0
  - large perforation in distal esophagus |0
  - esophagectomy |0
  - cervical esophagostomy |0
  - gastrostomy |0
  - transfer to surgical ICU |0
  - persistent septic shock |0
  - multi-organ failure |0
  - death |96
  - PCR detection of mycobacterial DNA in pleural fluid |0
  - histopathologic confirmation of TB in esophagus |0
  - esophageal TB diagnosis |0
  - perforation |0
  - septic shock |0
  - no recent upper endoscopy |0
  - no underlying mucosal damage |0
  - no response to conventional antibiotics |0
  - surgical intervention |0
  - no delay in diagnosis beyond 24 hours |0
  - TB coverage antibiotics initiated |0
  - informed consent obtained |0
  