56 years old | 0
    morbidly obese | 0
    no history of cardiac disease | 0
    feeling poorly | -72
    cough | -72
    fatigue | -72
    found nonresponsive | 0
    no palpable pulse | 0
    chest compressions initiated | 0
    automated external defibrillator used | 0
    automated rhythm analysis | 0
    shock advised | 0
    shock delivered | 0
    awakened the patient | 0
    admitted to medical intensive care unit | 0
    diagnosed with Klebsiella pneumonia | 0
    successfully treated | 336
    echocardiogram demonstrated normal heart | 336
    no arrhythmias during hospital course | 336
    consulted cardiac electrophysiologist | 336
    implantation of implantable cardioverter-defibrillator considered | 336
    rhythm strip not available initially | 336
    rhythm strip obtained after several days | 432
    incorrect interpretation of sinus tachycardia as ventricular arrhythmia | 432
    shock advised and delivered | 432
    shock awakened the patient | 432
    sinus tachycardia | 432
    continued sinus tachycardia postshock | 432