17 years old | 0
male | 0
Caucasian | 0
admitted to the hospital | 0
throat pain | -168
odynophagia | -168
blood tests | 0
Hemoglobin: 7.0 g/dL | 0
Hematocrit: 21% | 0
WBC: 33 x 10^9 cells/L | 0
platelets: 38 x 10^9 cells/L | 0
Acute promyelocytic leukemia (M3) | 0
daunorubicin | 0
vesanoid | 0
necrotic lesion in the M. palatoglossus | 0
necrotic lesion in the soft palate | 0
necrotic lesion in the uvula | 0
necrotic lesion in the right tonsil | 0
unpleasant odor | 0
biopsy | 0
culture | 0
nonspecific chronic diffuse inflammation | 0
necrotic areas | 0
numerous bacteria | 0
Enterococcus spp | 0
Staphylococcus aureus | 0
Candida SP | 0
noma-like lesion | 0
antibiotic therapy | 0
ceftazidime | 0
amicacin | 0
vancomycin | 0
fluconazole | 0
penicillin G | 0
pneumonia | 24
sepsis | 24
treatment in the intensive care unit | 24
total recovery | 1080
extensive loss of soft palate tissue | 1080