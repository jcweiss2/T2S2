60 years old | 0
    female | 0
    presented to the emergency department | 0
    left flank pain | -48
    pain radiating to the groin | -48
    vomiting | -48
    dizziness | -48
    lightheadedness | -48
    coronary artery disease | N/A
    prior angioplasty | N/A
    difficult-to-control type 2 diabetes mellitus | N/A
    insulin glargine 30 units twice a day | N/A
    insulin lispro 30 units thrice a day | N/A
    dulaglutide 1.5 mg weekly injection | N/A
    empagliflozin 25 mg once daily | -2928
    hypertension | N/A
    losartan 50 mg daily | N/A
    hypertriglyceridemia | N/A
    icosapent ethyl 2 g twice a day | N/A
    former smoker | N/A
    quit smoking 7 years ago | N/A
    family history for heart disease | N/A
    family history for hypertension | N/A
    family history for diabetes | N/A
    family history for dyslipidemia | N/A
    body mass index 26 kg/m2 | 0
    costovertebral tenderness | 0
    tachycardia | 0
    hypotension | 0
    did not respond to crystalloids | 0
    required vasopressors | 0
    lactic acidosis 8.4 mmol/L | 0
    leukocytosis 10900 | 0
    left shift (segments 77%, bands 9%) | 0
    platelet count 76000 | 0
    glycosylated hemoglobin A1C 14% | 0
    creatinine 3.5 | 0
    blood urea nitrogen 57 mg/dL | 0
    shock | 0
    severe sepsis | 0
    hypovolemia | 0
    aspartate aminotransaminase 81 U/L | 0
    alanine transaminase 79 U/L | 0
    alkaline phosphatase 160 | 0
    total bilirubin 1.6 | 0
    serum glucose >500 mg/dL | 0
    urine analysis large amount of glucose | 0
    urine analysis rare bacteria | 0
    urine analysis white blood cells <1/HPC | 0
    imaging abdomen showed severe emphysematous pyelonephritis left kidney | 0
    imaging abdomen showed radiological signs of ischemic colitis | 0
    portal venous gas | 0
    air within branches of superior mesenteric vein | 0
    initial antibiotic treatment with cefepime | 0
    initial antibiotic treatment with vancomycin | 0
    initial antibiotic treatment with metronidazole | 0
    emergent nephrectomy | 0
    bowel found viable | 0
    postoperative management in ICU | 0
    successful recovery | 0
    pan-susceptible Escherichia coli isolated | 0
    antibiotics de-escalated | 0
    discharged home | 24
    instructed to take cefpodoxime 200 mg twice daily for 7 days | 24
    empagliflozin discontinued | 24
    admitted to the hospital after near-syncope episode | 1488
    abdominal pain | 1488
    small bowel obstruction | 1488
    decompensated quickly | 1488
    cardiopulmonary arrest | 1488
    massive emesis | 1488
    aspiration of gastric contents | 1488
    full resuscitation | 1488
    ICU stay | 1488
    did not recover | 1488
    anoxic brain injury | 1488
    critical condition following cardiopulmonary collapse | 1488
    surgery never performed | 1488
    family decided to withdraw life support | 1488
    patient died | 1488
    