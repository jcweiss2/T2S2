55 years old | 0  
    Chinese woman | 0  
    referred to the Second Affiliated Hospital | -8760  
    gastric adenocarcinoma | -8760  
    physical examination unremarkable | -8760  
    no abdominal mass | -8760  
    no superficial lymph node | -8760  
    chest CT scan | -8760  
    abdominal CT scan | -8760  
    surgery | -8784  
    white nodules in abdominal cavity | -8784  
    poorly differentiated adenocarcinoma | -8784  
    extensive abdominal metastases | -8784  
    signet-ring cell carcinoma | -8784  
    immunohistochemistry CerbB-2 2+ | -8784  
    Ki67+ | -8784  
    Syn− | -8784  
    CgA− | -8784  
    FISH negative CerbB-2 gene amplification | -8784  
    first-line palliative chemotherapy | -8784  
    oxaliplatin | -8784  
    S-1 | -8784  
    imaging examination | -8784  
    stable disease | -8784  
    maintenance treatment with S-1 | -8784  
    cardiac obstruction | -4320  
    ENFTP | -4320  
    second-line chemotherapy | -4320  
    albumin-bounded paclitaxel | -4320  
    oxaliplatin | -4320  
    obstructive symptoms relieved | -4320  
    feeding tube removed | -4320  
    grade 4 neutropenia | -4320  
    rh-GCSF treatment | -4320  
    disease progression | -1440  
    incomplete gastrointestinal obstruction | -1440  
    apatinib prescribed | 0  
    apatinib administration | 0  
    obstruction symptoms | 0  
    nausea | 0  
    vomiting | 0  
    abdominal pain | 0  
    blood pressure rise | 0  
    spit blood streak | 456  
    clot | 456  
    fecal occult blood positive | 456  
    hematemesis | 456  
    fasting | 456  
    parenteral nutrition | 456  
    PPI prescription | 456  
    apatinib stopped | 456  
    sudden severe abdominal pain | 456  
    emergency erect abdominal plain radiograph | 456  
    gastrointestinal obstruction | 456  
    no subphrenic free air | 456  
    analgesic therapy | 456  
    spasmolytic therapy | 456  
    unstable hemodynamics | 456  
    antishock treatment | 456  
    enhanced abdominal CT scan | 456  
    large amount of ascites | 456  
    gastric mass | 456  
    peritoneal metastatic lesions | 456  
    acute surgical consultation | 456  
    gastrointestinal perforation | 456  
    acute diffuse peritonitis | 456  
    septic shock | 456  
    emergency operation | 456  
    purulent ascites | 456  
    perforated ulcer | 456  
    miliary nodules in abdominal cavity | 456  
    ileal tumor | 456  
    metastatic signet-ring cell carcinoma | 456  
    enterolysis | 456  
    perforated gastric wall repair | 456  
    ileal tumor resection | 456  
    transferred to ICU | 456  
    septic shock continued | 456  
    MODS | 456  
    death | 1176  
