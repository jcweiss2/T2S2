61 years old|0
female|0
type 2 diabetes mellitus|-672
poor glycaemic control|-672
fever|0
headache|0
severe anorexia|0
lethargy|0
apathy|0
dehydration|0
ill appearance|0
erythematous patch over right maxillary bone|0
tenderness over right maxillary bone|0
high neutrophil leukocytosis|0
CRP >200 mg/l|0
opacity in right maxillary sinus on OM view|0
bacterial sinusitis suspected|0
IV ceftriaxone initiated|0
blood culture obtained|0
insulin infusion started|0
basal bolus insulin regime|0
blood sugar 140-180 mg/dl|0
urinary ketones negative|0
referred to ENT for antral washout|0
antral wash samples sent for culture|0
no necrotic material in right maxillary sinus|0
clinical deterioration|0
hypotension|0
admitted to ICU|0
managed as septic shock|0
IV fluids administered|0
noradrenaline administered|0
E. coli in blood culture|0
E. coli in sinus washout culture|0
IV meropenem initiated|0
Rhizopus in sinus washout culture|96
broad folded ribbon-like non-septate hyphae|96
necrotic skin over right maxillary bone|96
IV liposomal amphotericin B started|96
USS abdomen arranged|168
chest x-ray arranged|168
left-sided psoas abscess detected|168
CECT abdomen confirmed abscess|168
asymptomatic psoas abscess|168
abscess aspirated under USS guidance|168
samples sent for culture and AFB|168
recollection of abscess|192
repeat USS psoas abscess|192
repeat aspiration under USS guidance|192
repeat flexible rhinoscopy|192
necrotic debris removed|192
maxillary bone erosion including orbital cavity|336
amphotericin B dose increased to 5 mg/kg/day|336
surgical drainage of psoas abscess|336
clinical improvement|336
biochemical improvement|336
hematological improvement|336
sudden deterioration of consciousness|672
normal metabolic screening|672
NCCT brain showing pneumocephalus|672
high-flow oxygen initiated|672
conscious level improved|672
repeat NCCT brain after 6 days|672
pneumocephalus improved by >50%|672
oxygen continued for another week|672
amphotericin B continued to cumulative 5g|0
meropenem continued for 6 weeks|0
complete clinical recovery|0
complete biochemical recovery|0
complete hematological recovery|0
final flexible rhinoscopy|0
no necrotic material|0
referred for facial reconstruction|0
