26 years old | 0
woman | 0
Vietnamese descent | 0
presented to the emergency department | 0
widespread symmetric erythematous and pustular eruption | 0
outbreak initially affected waistline | -96
outbreak initially affected axillary folds | -96
outbreak initially affected inguinal folds | -96
outbreak initially affected inframammary folds | -96
eruption spread to neck | -72
eruption spread to wrists | -72
eruption spread to areolae | -72
eruption spread to antecubital fossae | -72
eruption spread to popliteal fossae | -72
superficial flaccid nonfollicular pustules | -72
pustules evolved to confluent purulent lakes | -72
sparing of lower aspect of legs | 0
sparing of palms | 0
sparing of soles | 0
sparing of upper aspect of back | 0
Nikolsky sign absent | 0
mucous membrane involvement absent | 0
no target lesions | 0
no blisters | 0
diffuse burning sensation | -72
facial swelling | -72
subjective fevers | -72
malaise | -72
consumed 10 mg mifepristone | -96
emergency contraception | -96
not taken other medications | -96
not previously ill | -96
mifepristone purchased without prescription | -96
pharmacy in Vietnam | -96
used medication once prior | -96
tachycardic | 0
heart rate 150 beats/min | 0
elevated temperature 37.7°C | 0
total lymphocyte count 18,000/mm3 | 0
absolute neutrophils 17,800/mm3 | 0
albumin 2.3 g/dL | 0
calcium 6.5 mg/dL | 0
alkaline phosphatase 31 U/L | 0
sodium 131 mmol/L | 0
potassium 3.2 mmol/L | 0
bicarbonate 19 mmol/L | 0
phosphorus 1.8 mg/dL | 0
glucose 179 mg/dL | 0
renal function tests unremarkable | 0
liver function tests unremarkable | 0
skin swab cultures negative | 0
blood cultures negative | 0
skin swab PCR for varicella zoster virus negative | 0
skin swab PCR for herpes simplex virus negative | 0
quantitative hCG 1982.0 mIU/mL | 0
last menstrual period approximately 5 weeks prior | -840
unaware of pregnancy | 0
treated with 125 mg methylprednisolone | 0
treated with 1 g ceftriaxone | 0
admitted to hospital | 0
received second 125 mg methylprednisolone | 24
received four 600 mg clindamycin | 24
punch biopsy specimen | 24
extensive subcorneal pustules | 24
neutrophil spongiosis | 24
prominent papillary dermal edema | 24
hemorrhage | 24
brisk perivascular mixed inflammatory infiltrate | 24
many neutrophils | 24
eosinophils | 24
focal small-vessel vasculitis | 24
diagnosis of AGEP | 24
treatment with oral diphenhydramine | 24
triamcinolone 0.1% cream | 24
admitted to critical care service | 48
hypotension | 48
tachycardia not responsive to 5 L IV normal saline | 48
central line placed | 48
arterial line placed | 48
fluid resuscitation continued | 48
blood pressure recovered | 72
tachycardia resolved | 72
lines removed | 72
transferred to family medicine | 72
discharged | 72
complete recovery | 72
no sequela | 72
pregnancy electively terminated | 72
