75 years old | 0
female | 0
recurrent urinary tract infections | -672
hypothyroidism | -672
chronic pain | -672
depression | -672
opioid dependence | -672
altered mental status | 0
Temperature 100°F | 0
Heart rate 130 bpm | 0
Blood Pressure 114/60 mmHg | 0
Pulse Oximetry 86% on room air | 0
using accessory muscles | 0
diminished air entry | 0
scattered rhonchi and wheezes bilaterally | 0
bilateral lower extremity edema | 0
alert and awake | 0
oriented only to self | 0
White Blood Cell (WBC) Count of 19,000 | 0
neutrophilic predominance | 0
BUN 43 mg/dl | 0
Creatinine of 2.1 mg/dl | 0
albumin of 3 g/dl | 0
Lactic acid of 2.2 mg/dL | 0
acute hypoxic respiratory failure | 0
bilateral infiltrates on chest X-ray | 0
Bilevel Positive Airway Pressure (BiPAP) ventilation | 0
improvement within 24-48 hours | 24
worsening respiratory status | 72
inability to maintain oxygen saturation | 72
sinus tachycardia | 72
new onset paroxysmal atrial fibrillation | 72
S1QIIITIII pattern on EKG | 72
ceftriaxone and azithromycin | 0
prophylactic low molecular weight heparin | 0
saddle PE on Chest Computed Tomography Angiography (CTA) | 72
lethargic | 72
intubated for respiratory support | 72
Mycoplasma titers positive | 72
IgM greater than 950 U/mL | 72
IgG greater than 320 U/mL | 72
WBC count improved | 120
lactic acid normalized | 120
negative cultures | 120
hypercoagulable workup | 120
decreased protein C activity | 120
increased cold agglutinin titers | 120
catheter directed thrombolysis with tissue plasminogen activator (tPA) | 120
heparin drip | 120
intubated for about three days | 120
weaned off mechanical ventilation | 168
taken off antibiotics | 168
maintaining oxygen saturation | 168
severely hypoxic | 216
reintubated | 216
possible intraalveolar haemorrhage | 216
bedside bronchoscopy | 216
serosanguinous secretions | 216
full dose anticoagulation | 216
cefepime, vancomycin and fluconazole | 216
negative cultures from bronchoalveolar lavage | 216
extubated again | 240
downgraded from ICU to medical telemetry floor | 264
discharged to a rehabilitation facility | 336