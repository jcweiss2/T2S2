61 years old | 0
female | 0
admitted to the hospital | 0
breathing difficulties | -48
vomiting | -48
diarrhea | -48
right hemithoracic pain | -48
arterial hypertension | 0
hypercholesterolemia | 0
arthritis | 0
type 2 diabetes | 0
allergy to molds | 0
metformin | 0
co-lisinopril | 0
tramadol | 0
atorvastatin | 0
allopurinol | 0
ranitidine | 0
quinine sulfate | 0
naproxen | -240
arthritis (current) | 0
chest pain | 0
restless | 0
pale | 0
hypotensive | 0
sinus tachycardia | 0
pH 7.27 | 0
pCO2 23 mm Hg | 0
paO2 154 mm Hg | 0
base excess -17.5 | 0
serum bicarbonate 11 mEq/L | 0
potassium 3.14 mEq/L | 0
lactate 55 mg/dL | 0
marbled legs and thorax | 0
thirst | 0
admitted to ICU | 0
fluid resuscitation | 0
central venous pressure 14 mm Hg | 0
ScVO2 52% | 0
low urine output | 0
bradycardic | +few
cardiac arrest | +few
multiple organ failure | +few
respiratory failure | +few
renal failure | +few
liver failure | +few
coagulopathy | +few
inotropes | +few
amoxicillin-clavulanic acid | +few
amikacin | +few
meropenem | +few
vancomycin | +few
fluconazole | +few
SOFA score 21 | +few
APACHE II score 38 | +few
marbled skin pattern on thorax | 0
petechial lesions | +6
confluent petechial lesions | +24
erythematous eruptions | +24
bullous eruptions | +24
Nikolsky sign positive | +24
body surface involvement 80% | +24
epidermal necrosis | +24
muscle necrosis | +24
chest x-ray | 0
electrocardiogram | 0
lumbar puncture | 0
urine culture | 0
blood culture | 0
thoracoabdominal CT scan | 0
skin swab | 0
LTT positive for naproxen | +24
LTT negative for co-lisinopril | +24
LTT negative for allopurinol | +24
LTT negative for quinine | +24
LTT negative for amikacin | +24
LTT negative for metronidazole | +24
LTT negative for meropenem | +24
LTT negative for amoxicillin-clavulanic acid | +24
LTT negative for fluconazole | +24
anti-skin antibodies absent | +24
anti-skeletal muscle antibodies absent | +24
antineutrophil cytoplasmic antibody absent | +24
anti-glomerular basement membrane antibody absent | +24
anti-Jo1 antibody absent | +24
anti-scl70 antibody absent | +24
Mycoplasma pneumoniae serology negative | +24
Chlamydia pneumoniae serology negative | +24
hepatitis A virus serology negative | +24
hepatitis B virus serology negative | +24
hepatitis C virus serology negative | +24
naproxen discontinued | +24
methylprednisolone 1200 mg | +24
death | +48
So, rhabdomyolysis | 0, AKI |0.
AKI | 0
Rhabdomyolysis | 0
TEN | 0
naproxen 500 mg TID | -240
naproxen 1.5 g | 0
naproxen (500 mg TID) | -240
naproxen (1.5 g) | 0
bradycardic | +6
cardiac arrest | +6
multiple organ failure | +6
respiratory failure | +6
renal failure | +6
liver failure | +6
coagulopathy | +6
inotropes | +6
amoxicillin-clavulanic acid | +6
amikacin | +6
meropenem | +6
vancomycin | +6
fluconazole | +6
SOFA score 21 | +6
APACHE II score 38 | +6
