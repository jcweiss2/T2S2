11 years old | 0
male | 0
admitted to the hospital | 0
construction iron bar entered body | -1
iron bar entered from the right site of the anus | -1
iron bar exited from the loin | -1
waited for the fire department | -1
fire department arrived | -1
fire department cut the iron bar | -1
cut into a 140 cm piece | -1
taken to the nearest state hospital | -1
transferred to the emergency service | 0
slightly hypothermic | 0
intermediate overall condition | 0
no active hemorrhaging | 0
normal abdomen | 0
difficulty in breathing | 0
chest and abdominal x-ray examinations | 0
Pediatric Surgery, Orthopedics, Brain Surgery, Anesthesiology, and Radiology departments | 0
pain increased | 1
breathing difficulty increased | 1
intubated | 1
computed tomography (CT) | 1
no abdominal or chest injury detected | 1
possibility of rectosigmoid/retroperitoneal injury | 1
laparotomy | 2
tetanus vaccination | 2
antibiotic treatment started | 2
ampicillin/sulbactam, amikacin, ornidazole | 2
abdominal region opened | 2
hematoma at the sigmoid colon mesentery | 2
abdominal skin closed | 2
placed in the face-down position | 2
fire department called to cut the iron bar | 2
scissor-type cutter not suitable | 2
spiral cutter not suitable | 2
spiral-type cutter used | 2
cold water poured to prevent burning | 2
iron bar shortened and removed | 3
oxygen and nitrous oxide container tubes removed | 3
light exudate containing bone pieces | 3
wound washed and cleaned | 3
lumbar exit hole closed with a suture | 3
long Penrose drain placed | 3
abdominal cavity examined and closed | 3
intensive care unit | 4
discharged on the 11th day | 240
control lumbar spinal magnetic resonance image | 240
subcutaneous degenerative changes at L4-L5 levels | 240
degenerative changes in the nerve roots at S2–S5 levels | 240
electromyography findings normal | 240
no problems while walking, defecating, and urinating | 240
follow-up continued | 336
no problems after the 14th postoperative month | 672