25 years old | 0
woman | 0
obesity | 0
body mass index 40.1 kg/m² | 0
polycystic ovary syndrome | 0
iodine allergy | 0
gastritis | 0
admitted to receive LAGB procedure | 0
band placed laparoscopically via pars flaccida technique | 0
discharged on third day | 72
weight dropped to 95 kg | 168
occasional malaise | 168
feverishness | 168
recurrent upper respiratory tract infections | 168
readmitted to surgery department | -2160
fever | -2160
signs of port site infection | -2160
port removed | -2160
discharged after a day | -2160
occasional malaise | -2160
feverishness | -2160
gastroscopy | -2088
no signs of functioning band | -2088
no band erosion | -2088
readmitted to another surgical department | -2112
suspicion of band infection | -2112
laparoscopy | -2112
conversion to laparotomy | -2112
band removed | -2112
bacterial culture revealed E. coli infection | -2112
targeted antibiotics administered | -2112
minimal surgical wound infection | -2112
discharged on 8th day | -2112
returned after 2 weeks | -2112
hectic fever | -2112
elevated WBC | -2112
elevated CRP | -2112
abdominal CT scan | -2112
peritoneal adhesions | -2112
abdominal lymphadenopathy | -2112
mediastinal lymphadenopathy | -2112
left pleural effusion | -2112
broad-spectrum antibiotics administered | -2112
cilastatin | -2112
linezolid | -2112
no improvement | -2112
chest CT scan | -2112
increased parenchymal density | -2112
referred to pulmonology department | -2112
elevated Ca-125 | -2112
elevated GGTP | -2112
elevated D-dimer | -2112
elevated procalcitonin | -2112
hypoalbuminemia | -2112
IgA deficiency | -2112
bone marrow biopsy | -2112
reactive changes due to infection | -2112
no parasite infection confirmed | -2112
broad-spectrum antibiotics continued | -2112
antifungal agents continued | -2112
immunoglobulin therapy | -2112
prepared for surgery | -2112
sudden abdominal pain | -2112
signs of septic shock | -2112
urgent laparotomy | -2112
massive peritoneal adhesions | -2112
moderate ascites | -2112
swabbed for culture | -2112
parietal peritoneum covered in small nodules | -2112
visceral peritoneum covered in small nodules | -2112
greater omentum covered in small nodules | -2112
liver biopsy | -2112
omental biopsy | -2112
peritoneal biopsy | -2112
histopathological examination ruled out cancer | -2112
ruled out lymphoma | -2112
chronic granulomatous inflammation | -2112
Ziehl-Neelsen stain negative | -2112
transferred to intensive care unit | -2112
bronchial lavage tested for M. tuberculosis DNA | -2112
peritoneal effusion tested for M. tuberculosis DNA | -2112
test negative | -2112
suspecting atypical mycobacteriosis | -2112
ethambutol introduced | -2112
clarithromycin introduced | -2112
amikacin introduced | -2112
posaconazole introduced | -2112
antiparasitic agents introduced | -2112
total parenteral nutrition introduced | -2112
status stabilized | -2112
CRP levels normalized | -2112
WBC levels normalized | -2112
persisting fever | -2112
corticosteroids administered | -2112
fever lowered | -2112
enteral nutrition introduced | -2112
discharged | -2112
postoperative specimen tested genetically | -2112
revealed M. tuberculosis DNA | -2112
corticosteroids discontinued | -2112
isoniazid administered | -2112
rifampicin administered | -2112
pyrazinamide administered | -2112
streptomycin administered | -2112
therapy completed | -2112
abdominal CT scan no pathological findings | -2112
fever withdrew | -2112
malaise withdrew | -2112
no symptoms | -2112
