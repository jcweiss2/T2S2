62 years old | 0
female | 0
Caucasian | 0
weight 84 kg | 0
BMI 34 | 0
admitted to the hospital | 0
reno-vascular hypertension | -8760
type 2 diabetes | -8760
dyslipidemia | -8760
non-STEMI | -8760
end stage renal disease | -8760
kidney transplant | -8760
immunosuppressive regimen | -8760
mycophenolate | -8760
tacrolimus | -8760
prednisolone | -8760
acute pancreatitis | 0
pseudocyst formation | 0
tigecycline | -24
urinary tract infection | -24
carbapenem-resistant KP | -24
fosfomycin | -24
fever | 144
leukocytosis | 144
urine culture positive for KP | 144
meropenem | 144
fosfomycin | 144
abdominal pain | 288
hemorrhagic pancreatic pseudocyst | 288
ERCP | 432
EUS | 432
FNA | 432
presumed sepsis | 432
vancomycin | 432
ciprofloxacin | 432
amikacin | 432
caspofungin | 432
tacrolimus halted | 432
mycophenolate halted | 432
coagulase-negative Staphylococci | 432
ciprofloxacin replaced by meropenem | 504
amikacin discontinued | 504
CRE KP | 504
gastrointestinal bleeding | 1008
hypoxia | 1064
lung consolidation | 1064
BAL | 1104
KP resistant to antibiotics | 1104
ceftazidime/avibactam | 1104
blood cultures grew KP | 1152
Enterococcus faecium | 1152
vancomycin added | 1152
abdominal CT scan | 1152
pancreatic-pseudocyst-related soft tissue inflammatory changes | 1152
necrotic abscess | 1152
cardiac arrest | 1408
ertapenem and meropenem | 1408
cyst drainage | 1608
KP with same resistance profile | 1608
necrosectomy | 1764
Candida parapsilosis fungemia | 1764
fluconazole | 1764
abdominal fluid cultures grew KP | 1764
combination therapy continued | 1764
fever | 2112
resistant KP from urine | 2112
combination ertapenem and meropenem | 2112
discharged | 2520
rectal swab showed KP producing carbapenemases | 2520
NDM and OXA | 2520
Second admission | 4560
dysuria | 4560
left costovertebral angle tenderness | 4560
urine culture grew KP | 4560
ertapenem and meropenem | 4560
repeat urine culture negative | 4656
completed treatment course | 4710
Third admission | 5040
fever | 5040
chills | 5040
abscess on the right buttock | 5040
drained | 5040
Streptococcus sp | 5040
E. Coli | 5040
susceptible K. oxytoca | 5040
blood cultures grew KP | 5040
double carbapenem regimen | 5040
discharged | 5184
Fourth admission | 5616
fever | 5616
respiratory symptoms | 5616
Chest X-ray | 5616
computed tomography scan | 5616
necrotizing pneumonia | 5616
ertapenem and meropenem | 5616
sputum culture grew MSSA | 5616
KP of the same phenotype | 5616
carbapenem combination continued | 5616
discharged | 6048
Fifth admission | 6624
fever | 6624
thigh abscess | 6624
urinary symptoms | 6624
abscess drained | 6624
fluid and urine culture grew KP | 6624
combination therapy with ertapenem and meropenem | 6624
discharged | 6832
recent urine culture negative | 7256