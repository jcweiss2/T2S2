history of stage IIIA lung cancer | -648
history of smoking | -648
history of hypertension | -648
history of hypothyroidism | -648
history of dyslipidemia | -648
abdominal pain | 0
pancreatic head lesion | 0
spiculated suprahilar 4.5 × 2.6 cm right upper lobe (RUL) nodule | -648
multiple sub-centimeter left lung nodules | -648
augmented activity in the RUL mass | -648
NSCLC | -648
adenocarcinoma | -648
lymph node sampling was negative for nodal involvement | -648
stage IIIA lung adenocarcinoma (T4N0M0) | -648
program death ligand-1 expression was 15% | -648
surgical resection of the mass was planned | -648
surgical resection of the mass was aborted | -648
carboplatin and paclitaxel | -648
radiation therapy | -648
decrease in the RUL mass | -120
adjuvant immunotherapy with durvalumab | -90
pneumonitis | -60
steroid taper | -60
increase in the RUL mass | -30
stable lung nodules | 0
stable post-radiation changes | 0
epigastric pain | 0
constipation | 0
loss of appetite | 0
weight loss | 0
mass in the head of the pancreas | 0
pancreatic ductal dilatation | 0
endoscopic ultra-sound-guided biopsy of the pancreatic head mass | 0
tumor cells with nuclear pleomorphism | 0
tumor cells with prominent nucleoli | 0
tumor cells with irregular nuclear contours | 0
tumor cells with coarse chromatin | 0
CK7 positivity | 0
TTF-1 positivity | 0
Napsin-A positivity | 0
CDX-2 negativity | 0
KOC negativity | 0
synaptophysin negativity | 0
Smad-4 mixed staining pattern | 0
lung adenocarcinoma metastasized to the pancreas | 0
normal liver enzymes | 0
normal total bilirubin | 0
normal direct bilirubin | 0
CA 19.9 | 0
PET/CT scan | 30
fluorodeoxyglucose-avid mass in the pancreatic head | 30
increased uptake in the porta hepatis | 30
brain MRI scan | 30
no intracranial metastasis | 30
palliative radiation therapy to the pancreatic mass | 90
combination chemotherapy with carboplatin and pemetrexed | 90
generalized weakness | 120
dyspnea at rest | 120
electrolyte derangements | 120
acute anemia | 120
hemoglobin nadir of 6.9 g/dL | 120
transfusion | 120
new 9 mm left lower lobe nodule | 120
staging PET/CT scan | 180
decreased metabolic activity in the pancreatic mass | 180
metabolic activity in the new left lower lobe nodule | 180
fatigue | 180
no further treatments | 180
increased dyspnea | 210
cough | 210
generalized weakness | 210
right lung consolidation | 210
loculated pleural effusion | 210
broad-spectrum antibiotics | 210
oxygen supplementation | 210
bilevel-positive airway pressure | 210
altered mentation | 216
worsening hypoxemia | 216
vasopressor support | 216
palliative medicine team | 216
inpatient hospice care | 216
death | 216