5 years old | 0
male | 0
admitted to the hospital | 0
fever | -144
night sweats | -144
weight loss | -144
cough | -144
bilateral anterior cervical lymph nodes enlargement | 0
peripheral cyanosis in digits | 0
hemoglobin concentration: 128 g/L | 0
white blood cell count: 9.12×10^9/L | 0
neutrophils: 30.1% | 0
lymphocytes: 57.3% | 0
eosinophils: 6.61% | 0
monocytes: 4.54% | 0
basophils: 1.45% | 0
platelet count: 329×10^9/L | 0
liver enzymes normal | 0
serum bilirubin normal | 0
creatinine normal | 0
blood urea nitrogen normal | 0
blood culture showed no bacterial growth | 0
bilateral airway narrowing | 0
multiple bilateral anterior cervical as well as supraclavicular and infraclavicular lymphadenopathy | 0
cystic degeneration suggestive of central necrosis | 0
heterogenous density of thyroid gland | 0
bilateral nodular and micronodular lung densities | 0
hilar lymphadenopathy | 0
mild hepatomegaly | 0
paraaortic lymph node enlargement | 0
excisional biopsy of a single cervical lymph node | 24
bone marrow trephine biopsy | 24
histopathological examination of the lymph node showed proliferation of malignant thyroid glands | 48
diagnosis of metastatic papillary thyroid carcinoma | 48
bone marrow biopsy was negative for metastasis | 48
total thyroidectomy and cervical lymph nodes excision | 168
radioactive iodine therapy | 168
respiratory symptoms | 2160
CT scan revealed multiple bilateral pulmonary nodules consistent with metastasis | 2160
unstable vital signs | 2232
admitted to intensive care unit | 2232
septicemia by methicillin-resistant Staphylococcus aureus | 2280
death | 2280