26 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
height 180 cm | 0 | 0 | Factual
weight 74 kg | 0 | 0 | Factual
kidney transplant | -18960 | -18960 | Factual
end-stage kidney disease | -29040 | -18960 | Factual
immunosuppression | 0 | 0 | Factual
mycofenolate sodium | 0 | 0 | Factual
methylprednisolone | 0 | 0 | Factual
headache | -24 | 0 | Factual
blurred vision | -24 | 0 | Factual
estimated glomerular filtration rate 35.9 mL/min/1.73 m2 | 0 | 0 | Factual
proteinuria 117 mg/d | 0 | 0 | Factual
chronic kidney transplant disease stage 3bA1 | 0 | 0 | Factual
chronic transplant nephropathy | 0 | 0 | Factual
status post vascular rejection | -18960 | -18960 | Factual
chronic calcineurin-inhibitor toxicity | -18960 | -18960 | Factual
cranial CT scan | 0 | 0 | Factual
cranial MRI scan | 0 | 0 | Factual
contrast-enhancing intracerebral lesions | 0 | 0 | Factual
perifocal edema | 0 | 0 | Factual
methylprednisolone therapy stopped | 0 | 0 | Factual
dexamethasone administered | 0 | 24 | Factual
brain edema | 0 | 24 | Factual
transmitted to university department of Nephrology | 24 | 24 | Factual
transmitted to department of Neurosurgery | 24 | 24 | Factual
brain biopsy | 48 | 48 | Factual
cerebral PTLD diagnosed | 48 | 48 | Factual
diffuse large B-cell lymphoma | 48 | 48 | Factual
Epstein-Barr virus positive | 48 | 48 | Factual
CT scan of thorax | 48 | 48 | Factual
abdomen sonography | 48 | 48 | Factual
bone marrow biopsy | 48 | 48 | Factual
chemotherapy regime | 72 | 168 | Factual
high-dose cytarabin | 72 | 168 | Factual
Rituximab | 72 | 168 | Factual
MRI scan confirmed complete remission | 168 | 168 | Factual
impairment of transplant function aggravated | 168 | 168 | Factual
eGFR 25.4 mL/min/1.73 m2 | 168 | 168 | Factual
cytomegalovirus reactivated | 504 | 504 | Factual
pneumocystis jirovecii pneumonia | 504 | 504 | Factual
chemotherapy changed | 504 | 504 | Factual
Rituximab dose increased | 504 | 504 | Factual
antiviral therapy | 504 | 504 | Factual
antibiotic therapy | 504 | 504 | Factual
mycofenolate sodium dose tapered | 504 | 504 | Factual
leukopenia | 504 | 504 | Factual
infections | 504 | 504 | Factual
generalized seizure | 1008 | 1008 | Factual
cerebral MRI scan demonstrated recurrence of PTLD | 1008 | 1008 | Factual
HDMTX administered | 1032 | 1032 | Factual
leukovorine administered | 1032 | 1032 | Factual
Rituximab administered | 1032 | 1032 | Factual
vigorous hydration | 1032 | 1032 | Factual
alkalinization of urine | 1032 | 1032 | Factual
high-flux hemodialysis | 1056 | 1104 | Factual
MTX-level measurements | 1056 | 1104 | Factual
dialysis parameters | 1056 | 1104 | Factual
nadir of leucocytes | 1140 | 1140 | Factual
CMV- and E.coli pneumonia | 1188 | 1188 | Factual
sepsis | 1188 | 1188 | Factual
acute kidney transplant failure | 1188 | 1188 | Factual
transmission to intensive care unit | 1188 | 1188 | Factual
invasive ventilation | 1188 | 1188 | Factual
sepsis managed | 1200 | 1200 | Factual
mycofenolate sodium discontinued | 1200 | 1200 | Factual
antiviral therapy | 1200 | 1200 | Factual
antibiotic therapy | 1200 | 1200 | Factual
follow-up cerebral MRI scan | 1296 | 1296 | Factual
small regredience of PTLD | 1296 | 1296 | Factual
cerebral radiation | 1296 | 1296 | Factual
no relevant response to radiotherapy | 1296 | 1296 | Factual