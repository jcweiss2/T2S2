10 years old | 0
male | 0
admitted to the hospital | 0
fever | -168
impetigo | -144
diarrhea | -120
medical history unremarkable | 0
family history unremarkable | 0
acutely ill | 0
uncomfortable | 0
irritable | 0
unable to stand | 0
unable to converse normally | 0
heart rate 147 beats/min | 0
blood pressure 101/61 mmHg | 0
temperature 40.5˚C | 0
respiratory rate 42 breaths/min | 0
oxygen saturation 100% | 0
no nuchal rigidity | 0
lung fields clear | 0
cheek erythema | 0
pharyngeal erythema | 0
impetigo on forehead and jaw | 0
abdominal tenderness | 0
swelling left elbow | 0
redness left elbow | 0
tenderness left elbow | 0
swelling left ankle | 0
redness left ankle | 0
tenderness left ankle | 0
rapid antigen detection test positive | 0
blood culture positive for Streptococcus pyogenes | 0
throat culture positive for Streptococcus pyogenes | 0
impetigo pus culture positive for Streptococcus pyogenes | 0
ampicillin/sulbactam administered | 0
clindamycin administered | 0
intravenous immunoglobulins administered | 0
blood cultures negative | 72
fever persisted | 0
rhTM administered | 0
antithrombin-III administered | 0
danaparoid administered | 48
DIC score increased | 48
general condition poor | 48
fever persisted | 48
DIC score decreased | 72
swelling left lower leg worsened | 120
redness left lower leg worsened | 120
pain left lower leg worsened | 120
contrast-enhanced CT scan performed | 168
inflammation left popliteal vein | 168
coagulopathy left popliteal vein | 168
LRINEC score 8 | 168
skin biopsy performed | 168
spongiotic dermatitis diagnosed | 168
suppurative panniculitis diagnosed | 168
magnetic resonance imaging performed | 216
inflammatory findings left soleus | 216
inflammatory findings left gastrocnemius | 216
no arthritis | 216
no osteomyelitis | 216
condition improved | 240
discharged | 480
no sequelae | 480
no medication-related adverse events | 480