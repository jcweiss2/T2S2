86 years old | 0
male | 0
dementia | 0
hypertension | 0
cough | -168
shortness of breath | -168
no chest pain | -168
acute hypoxic respiratory failure | -24
mechanical ventilation | -24
anteroseptal ST-segment elevation | -24
blood pressure 85/57 mmHg | 0
sedated and intubated | 0
no abnormalities on cardiopulmonary exam | 0
elevated troponin | 0
elevated creatinine | 0
elevated lactate dehydrogenase | 0
elevated C-reactive protein | 0
bilateral infiltrates on chest radiography | 0
ST-segment elevations in leads V2 and V3 | 0
ejection fraction 50-55% | 0
no significant regional wall motion abnormalities | 0
no signs of cardiac tamponade | 0
admitted to intensive care unit | 0
requiring mechanical ventilation | 0
requiring vasopressor support | 0
troponin increased to 7.84 ng/mL | 24
COVID-19 test positive | 72
respiratory status worsened | 120
required increased oxygen | 120
required positive end-expiratory pressure | 120
renal function worsened | 120
lymphopenia | 120
inflammatory biomarker abnormalities | 120
required higher amounts of oxygenation | 168
loss of R waves on electrocardiogram | 168
transient T wave inversions on electrocardiogram | 168
deepened Q waves on electrocardiogram | 168
worsening kidney injury | 192
rise in D-dimer level | 192
pursue comfort care measures | 192
died | 192