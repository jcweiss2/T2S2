54 years old | 0
female | 0
admitted to the hospital | 0
altered mental status | -672
weakness | -672
elevated blood pressure | 0
moon facies | 0
weakness in bilateral lower extremities | 0
reduced strength in bilateral hip flexors | 0
inability to ambulate independently | 0
diabetes mellitus | -672
hypertension | -672
breast cancer | -10080
bilateral total mastectomy | -10080
adjuvant hormonal therapy | -10080
profund hypokalemia | 0
alkalemia | 0
elevated serum cortisol | 0
elevated serum ACTH | 0
abnormal dexamethasone suppression testing | 0
elevated serum chromogranin | 0
bilateral pulmonary lesions | 0
intraabdominal lymphadenopathy | 0
bilateral diffuse adrenal gland thickening | 0
multiple hepatic metastases | 0
2.5 cm lesion at the pancreatic tail | 0
severe proximal myopathy | 0
severe generalized myofiber atrophy | 0
metastatic NET | 0
NET, G1 | 0
Ki-67 proliferative index <3% | 0
mitotic rate not reported | 0
neoplastic cells positive for synaptophysin | 0
neoplastic cells positive for chromogranin | 0
neoplastic cells positive for caudal-type homeobox 2 (CDX2) | 0
neoplastic cells negative for calretinin | 0
neoplastic cells negative for inhibin | 0
neoplastic cells negative for S100 | 0
neoplastic cells negative for cytokeratin-7 (CK7) | 0
neoplastic cells negative for GATA binding protein 3 (GATA-3) | 0
neoplastic cells negative for thyroid transcription factor-1 (TTF-1) | 0
started on octreotide acetate | 24
started on ketoconazole | 48
received a total of 38 days of oral ketoconazole | 120
started on abiraterone acetate (AA) | 120
effects of serum cortisol reduction were immediate | 120
serum cortisol levels completely normalized | 130
underwent bilateral adrenal artery embolization | 130
AA was stopped | 134
discharged to a rehabilitation facility | 144
admitted to the medical intensive care unit | 168
septic shock secondary to pneumonia | 168
succumbed | 168