77 years old | 0
male | 0
benign prostatic hyperplasia | 0
nocturia | 0
increased frequency | 0
hypertension | 0
fatty liver | 0
hemiparesis due to acute infarction of the basal ganglia | 0
cilostazol discontinued | -336 (2 weeks before surgery)
holmium laser enucleation of the prostate | 0
prostate biopsy | 0
general anesthesia induced with propofol and rocuronium | 0
remifentanil infusion | 0
laryngeal mask airway insertion | 0
sevoflurane maintenance | 0
mechanical ventilation | 0
anesthesia time 85 minutes | 85
arrival in recovery room | 85
shivering | 85 + 10 minutes = 95 minutes (timestamp: 95)
severe anxiety | 95
pethidine injection | 95
fentanyl injection | 95
mental status deterioration to stupor | 95
masseter muscle rigidity | 95
arm rigidity | 95
sudden hyperventilation | 95
oxygen mask applied | 95
blood pressure 220/168 mmHg | 95
heart rate 134 beats/minute | 95
respiratory rate 30 breaths/minute | 95
body temperature 38.1°C | 95
oxygen saturation 98% | 95
body temperature increased to 39.8°C | 95 + 10 minutes = 105 (timestamp: 105)
worsened masseter muscle rigidity | 105
MH clinical classification score 53 | 105
dantrolene sodium administration | 105
aggressive cooling | 105
esmolol administration | 105
arterial blood gas analysis | 105
compensated metabolic acidosis | 105
creatine phosphokinase increased | 105
lactate dehydrogenase increased | 105
myoglobin increased | 105
body temperature decreased to 36.8°C | 105 + 10 minutes = 115 (timestamp: 115)
systemic muscle rigidity resolved | 115
ICU admission | 115
consciousness restored | 115
general weakness | 115
stable respiratory pattern | 115
body temperature between 36.7°C and 37.5°C | 115
urinalysis | 115
sanguineous urine | 115
postoperative day 1 mild fever (37.2°C to 38.2°C) | 24
chest radiograph mild pulmonary edema | 24
white blood cell count 28,700/µL | 24
hemoglobin 10.3 g/dL | 24
hematocrit 31% | 24
platelet count 74,000/µL | 24
C-reactive protein 10.51 mg/dL | 24
arterial blood gas analysis pH 7.48 | 24
PaCO2 28 mmHg | 24
PaO2 66 mmHg | 24
bicarbonate 20.9 mmol/L | 24
oxygen saturation 94% | 24
antibiotics started | 24
postoperative day 2 body temperature 37.7°C to 38.6°C | 48
blood urea nitrogen 19.3 mg/dL | 48
creatinine 1.15 mg/dL | 48
sanguineous urine | 48
postoperative day 4 oral diet started | 96
Klebsiella pneumoniae identified in blood | 96
transferred to general ward | 144
discharged | 288
MH recurrence warning | 288
dantrolene sodium rapid reversal of symptoms | 115
MH almost certain diagnosis | 105
no residual sevoflurane exposure | 95
delayed-onset MH | 95
clinical grading scale MH | 105
no cola-colored urine | 115
ruled out sepsis and other differentials | 24
MH resolved | 115
muscle weakness after dantrolene | 115
confirmation test not performed | 288
dantrolene administration once | 105
morbidity due to MH | 288
continuous education importance | 288
prompt diagnosis importance | 288
