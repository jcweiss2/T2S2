69 years old | 0
male | 0
hypertension | 0
coronary artery disease | 0
stage 4 chronic kidney disease | 0
diarrheal illness | -1440
fever | -1440 (absence noted in the history of diarrheal illness)
nausea | -1440 (absence noted in the history of diarrheal illness)
abdominal pain | -1440 (absence noted in the history of diarrheal illness)
jaundice | -1440 (absence noted in the history of diarrheal illness)
admitted to the hospital | 0
septic shock | 12
transferred to Medical Intensive Care Unit | 12
intravenous ceftriaxone | 12
escalated to meropenem | 24 (after blood cultures returned positive)
blood cultures positive for P. aeruginosa | 24
sharply defined erythematous plaques on left anterior leg | 24 (second day of admission)
spread to right anterior leg | 24 (second day of admission)
involvement of lateral aspects of both thighs | 24 (second day of admission)
patchy involvement over posterior aspects of both legs | 24 (second day of admission)
tense bullae formation | 24 (subsequent hours after plaques developed)
serous fluid in bullae | 24
clinical differential diagnoses | 24
bullous drug reaction | 24
bullous erysipelas | 24
septic vasculitis | 24
biopsy taken from right thigh | 24
histological examination | 24 (after biopsy)
partial necrosis of the epidermis | 24
sub-epidermal blistering | 24
microthrombi in dermal blood vessels | 24
deeper vessels showing neutrophilic infiltrate | 24
nuclear dust | 24
Gram-negative bacilli extruding from vessel wall | 24
fluid culture from bulla aspirate grew P. aeruginosa | 24
aggressive fluid resuscitation | 24 (ongoing after septic shock)
high vasopressor support | 24 (ongoing after septic shock)
appropriate antibiotic therapy | 24 (ongoing after septic shock)
severe sepsis | 24 (ongoing)
evolving ST elevation myocardial infarction | 24 (during ICU stay)
severe disseminated intravascular coagulopathy | 24 (during ICU stay)
intracranial bleeding | 24 (during ICU stay)
passed away | 24 (eventually after complications)
