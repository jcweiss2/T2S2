23 years old | 0
male | 0
retrosternal pleuritic chest pain | -72
low-grade fever | -72
apyretic | 0
normotensive | 0
pericardial rub | 0
sinus tachycardia | 0
widespread ST elevation | 0
PR segment depression | 0
mild pericardial effusion | 0
normal high sensitivity troponin I | 0
mild leukocytosis | 0
very elevated C-reactive protein | 0
cardiac tamponade | 24
pericardiocentesis | 24
profund shock | 24
high noradrenaline doses | 24
methylprednisolone | 24
excellent clinical response | 48
weaning of noradrenaline | 48
resolution of the effusion | 48
childhood asthma | -100000
nonallergic rhinitis | -100000
idiopathic episcleritis | -100000
topical corticosteroids | -100000
septic shock | -720
tonsillitis | -720
Streptococcus mitis | 24
ceftriaxone | 24
constrictive-effusive physiology | 24
autoimmunity workup | 24
colchicine | 168
ibuprofen | 168
prednisolone | 168
idiopathic acute pericarditis | 168
incessant pericarditis | 672
cardiac tamponade | 672
pericardiocentesis | 672
pleuro-pericardial window | 672
pericardial biopsy | 672
diastolic paradoxical septal movement | 672
diffuse pericardial late gadolinium enhancement | 672
hyperkalemia | 1344
hyponatremia | 1344
adrenal insufficiency | 1344
adrenocorticotropin | 1344
cortisol | 1344
Addison's disease | 1344
hormonal replacement therapy | 1344
fludrocortisone | 1344
prednisolone | 1344
autoimmune polyglandular syndrome type 2 | 1344
anti-intrinsic factor autoantibodies | 1344
primary hypogonadism | 1344
free T4/TSH | 168
γ Interferon | 168
Human immunodeficiency virus serology | 168
Cytomegalovirus | 168
Epstein Barr virus | 168
Parvovirus | 168
Herpes virus 1 | 168
Herpes virus 2 | 168
Coxiella burnetti | 168
Borrelia burgdoferi | 168
Rickettsia conori | 168
Treponema pallidum | 168
Antinuclear antibodies | 168
Anti-dsDNA antibodies | 168
Anti-pANCA/c ANCA | 168
Anti-SSA60, Sm, RNP, Scl70, JO | 168
Rheumatoid factor | 168
discharged | 1344
readmitted | 1344
recurrence | 2016
prednisolone tapering | 2016
new recurrence | 3024