history of primary refractory acute myeloblastic leukemia | -8760
allogeneic bone marrow transplant from cord blood | -648
vancomycin-resistant Enterococcus, Streptococcus viridans and Streptococcus mitis bacteremia | -648
treated with tedizolid, cefepime, Flagyl and daptomycin | -648
on filgrastim | 0
on prophylaxis with acyclovir, Bactrim, and caspofungin | 0
on antibiotics for bacteremia | 0
acute abdominal pain | 0
fever to 38.2°C | 0
tachycardia to 155 | 0
hypotension to 99/81 | 0
tachypnea to 36 | 0
ill appearing with a distended abdomen and localized peritonitis | 0
white cell count was 0.2 x 10^9 /L | 0
absolute neutrophil count (ANC) of zero | 0
anemic with a hemoglobin of 7 g/L | 0
thrombocytopenic with a platelet count of 10 x 10^9 /L | 0
lactic acid of 3.1 mmol/L | 0
CT scan revealed segmental ischemia of the small bowel | 0
exploratory laparotomy | 2
15 cm ischemic bowel segment was identified without perforation | 2
approximately 50 cm of small bowel was resected | 2
primary anastomosis was performed with a stapler device | 2
required norepinephrine and vasopressin for blood pressure support | 2
transesophageal echo was unremarkable | 2
admitted to the intensive care unit | 2
pressors were weaned | 24
extubated | 24
transferred to the floor | 72
diet was advanced | 72
passed flatus | 72
new fevers | 96
increased abdominal pain | 96
lactic acidosis | 96
respiratory decompensation | 96
continued to be neutropenic with white cell count of 0.1x 10^9 /L | 96
ANC 0 | 96
lactic acid at that time was 3.7 mmol/L | 96
amphotericin B (AmBisome) was started | 96
repeat CT scan showed an area of necrotic small bowel | 96
expedited pathology report of the resected small bowel revealed invasive fungal forms | 96
invasive fungal forms in both the omental and small intestinal resection specimens | 96
amphotericin B was added to his antimicrobials | 96
decision was made to proceed to comfort measures | 120
died | 120