59 years old | 0
male | 0
heavy smoker | 0
painless gross hematuria | 0
lower urinary tract symptoms | -1096
α1 blocker medication | -1096
mild pale patient | 0
Blood pressure 120/60 mm/Hg | 0
Pulse = 70 | 0
mild tenderness in the lower abdominal region | 0
hemoglobin of 9 g/dl | 0
white blood cell count of 13 × 10^9/l | 0
platelet count of 390 × 10^9/l | 0
creatinine normal | 0
urea normal | 0
electrolytes normal | 0
excess RBC/HPF | 0
30-50 WBC/HPF | 0
4-5 epithelial cells/HPF | 0
grade 3 right renal hydronephrosis | 0
simple cyst | 0
bladder diverticulum in the right bladder wall | 0
mass with blood supply | 0
CT confirmed diagnosis of right bladder diverticulum with 21.3 × 51.9 mm mass intradiverticulum | 0
cystoscopy | 24
enlarged prostate | 24
severe bladder trabeculation | 24
transurethral resection of the prostate (TUR-P) | 24
partial cystectomy | 48
para-aortic lymph node dissection | 48
papillary transitional cell carcinoma (high grade) PT3 grade | 48
lymph nodes not free | 48
cardiac arrhythmia | 168
right pleural effusion | 168
sepsis | 168
death | 168