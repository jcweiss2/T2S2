60 years old | 0
male | 0
admitted to the hospital | 0
fever | -48
abdominal pain | -48
edema of the scrotum | -48
edema of the penis | -48
edema of the perineum | -48
edema of the right gluteal region | -48
hypertension | 0
osteoporosis | 0
hemorrhoids | 0
blood pressure 103/62 mmHg | 0
heart rate 135/min | 0
oxygen saturation 88% | 0
high white blood cell count | 0
elevated C-reactive protein | 0
serum creatinine 4.3 mg/dL | 0
blood urea 157 mg/dL | 0
blood sugar 142 mg/dL | 0
procalcitonin 8.53 ng/mL | 0
RT-PCR test for SARS-CoV-2 negative | 0
CT abdomen and pelvis findings | 0
Fournier's gangrene diagnosis | 0
meropenem therapy | 0
metronidazole therapy | 0
linezolid therapy | 0
resection of necrotic tissues | 0
bilateral orchiectomy | 0
excision of penile skin | 0
excision of scrotal skin | 0
transferred to ICU | 0
mechanical ventilation | 0
broad-spectrum antibiotics | 0
supportive therapy | 0
nutritional therapy | 0
colostomy | 0
wound debridement | 0
negative pressure wound therapy | 0
condition improvement | 0
sedation discontinued | 0
recovered consciousness | 0
extubated | 0
self-breathing with oxygen | 0
hemodynamically stable | 0
furosemide use | 0
inflammatory markers decreased | 0
pus culture showing Escherichia coli | 0
pus culture showing Pseudomonas aeruginosa | 0
antibiotic therapy modification | 0
cephazolin therapy | 0
NPWT discontinued | 0
transferred to Plastic Surgery | 0
free-skin grafts applied | 0
discharged | 1104
nursing home care | 1104
free-skin graft care | 1104
regular dressing changes | 1104
physiotherapy | 1104
testosterone supplementation | 1104
colostomy reversal planned | 1104
