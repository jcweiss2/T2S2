59 years old | 0
    male | 0
    prostatic cancer | 0
    computed tomography guided percutaneous transhepatic core needle liver mass biopsy | -9
    angio-embolization of hepatic mass | -9
    presented in recovery room | 0
    blood pressure 84/55 | 0
    heart rate 77 | 0
    respiratory rate 26 | 0
    acidotic with pH 7.31 | 0
    base deficit of 6.5 | 0
    INR of 1.6 | 0
    PT 17.8 | 0
    bladder pressure 25 mmHg | 0
    repeat CT of abdomen and pelvis | 0
    increasing bladder pressure | 0
    persistent hypotension | 0
    expansion of perihepatic hematoma | 0
    no evidence of blush | 0
    admission to surgical ICU | 0
    coagulopathy correction | 0
    coagulopathy not corrected despite transfusions | 0
    developed severe intra-abdominal hypertension | 0
    compartment syndrome with bladder pressure 40 mmHg | 0
    taken to operating room | 0
    bleeding liver mass located in segments 7 and 8 | 0
    falciform ligament taken down | 0
    right upper quadrant packed | 0
    stabilized | 0
    packs dry at end of case | 0
    resumed bleeding within 24 hours | 24
    angiography of right hepatic artery | 24
    no blush | 24
    bleeding thought to be venous in origin | 24
    fed by superior right hepatic artery branch | 24
    selective right hepatic artery embolization performed | 24
    returned to OR for continued hemorrhage | 24
    hepatic artery branch ligated | 24
    laparotomy packing performed in right upper quadrant | 24
    stabilized | 24
    post-operative day 2 | 48
    returned for re-exploration | 48
    liver packs removed | 48
    parenchymal bleeding resumed | 48
    Surgicel used | 48
    Argon beam coagulation | 48
    fibrin sealant | 48
    more packing | 48
    insufficient hemostasis | 48
    initiated BOLSA | 48
    intraoperative improvements after BOLSA placement | 48
    BP at surgery start 80/45 | 48
    BP as low as 75/45 | 48
    BP at end 90/50 | 48
    case lasted 19 minutes | 48
    massive transfusion protocol ongoing | 48
    transfusions: 3 units PRBC, 3 units FFP | 48
    EBL 2 liters | 48
    case 2 lasted 32 minutes | 24
    initial BP 100/49 | 24
    BP low 80/40 | 24
    BP at end 125/55 | 24
    case 3 (BOLSA placement) | 120
    BP low 90/45 | 120
    BP at end 110/50 | 120
    vasopressors used | 120
    case lasted 2 hours | 120
    BOLSA creation 10 minutes | 120
    BOLSA placement 10 minutes | 120
    transfusions: 4 PRBC, 3 FFP, 1 10-pack platelets | 120
    case 4 (POD 4) | 168
    cholecystectomy performed | 168
    Wittmann patch placement | 168
    case lasted 2 hours 2 minutes | 168
    BP start 100/60 | 168
    BP end 120/60 | 168
    transfusions: 2 PRBC, 2 FFP, 1 10-pack platelets | 168
    final case (POD 7) | 168
    abdominal closure | 168
    no transfusions | 168
    pathology report returned as hemangioma | 168
    POD 9 | 216
    BOLSA removed | 216
    abdomen closed primarily | 216
    resumed activities of daily living | 216
    discharged home | 216
    ischemic cholecystitis secondary to embolization | 168
    Wittmann patch serial tightening | 168
    mesh sheets sutured | 48
    purse-string sutures created | 48
    right coronary and triangular ligaments taken down | 48
    pro-coagulant material placed | 48
    BOLSA placed around right liver lobe | 48
    gallbladder accommodated without strangulation | 48
    no sutures to ligaments | 48
    cholecystectomy for ischemic cholecystitis | 168
    Wittmann patch due to visceral edema | 168
    liver biopsy pathology hemangioma | 168
    BOLSA removal without bleeding | 216
    abdominal closure | 216
    discharge home | 216
    