59 years old | 0
male | 0
underwent radical cystoprostatectomy | -105984
ileal neobladder (Studer Pouch) reconstruction | -105984
bladder cancer (G2pT2) | -105984
isolated 60 cm distal ileal segment | -105984
left 10 cm proximal ileum intact | -105984
sutured neobladder creation | -105984
standard ureteroileal anastomosis | -105984
post-operative urinary incontinence | -105984
urodynamics at 9 months | -105984
small capacity neobladder | -105984
high pressures (35 cm H2O) | -105984
neobladder augmentation cystoplasty | -7224
increased pouch capacity (550 ml) | -7224
presented to emergency department | 0
dyspnea at rest | 0
right loin pain | 0
polycystic kidney disease | 0
urinary tract infection | 0
oral antibiotics | 0
cachectic | 0
dry mucous membranes | 0
tachypnea (26 breaths/min) | 0
tachycardia (108 beats/min) | 0
hypotension (92/64 mmHg) | 0
well-healed laparotomy incision | 0
leucocytosis (14.1 × 10³/μl) | 0
raised C-Reactive Protein (23.3 mg/dl) | 0
hypokalaemia (3.3 mmol/L) | 0
elevated creatinine (304 μmol/L) | 0
elevated urea (33.1 mmol/L) | 0
normal anion gap (12.1 mEq/l) | 0
microscopic haematuria | 0
sterile pyuria | 0
sinus tachycardia (ECG) | 0
normal chest X-ray | 0
initial diagnosis of severe urosepsis | 0
acute kidney injury | 0
admitted to general medical ward | 0
broad-spectrum antibiotics | 0
urinary catheterization | 0
crystalloid fluid resuscitation | 0
confusion | 48
lethargy | 48
increasing respiratory distress | 48
worsening hyperchloremic metabolic acidosis | 48
deteriorating vital signs | 48
unresponsive (GCS 8/15) | 48
consultation with original surgical team | 48
hyperchloremic metabolic acidosis diagnosis | 48
transfer to intensive care unit | 48
sodium bicarbonate 8.4% infusion | 48
regained consciousness | 52
improving metabolic acidosis | 52
remained in ICU for 3 days | 52
sodium bicarbonate 1.26% infusions | 52
discharged with oral sodium bicarbonate | 168
recuperation period | 168
neobladder excision | 168
ileal conduit formation | 168
no further metabolic acidosis episodes | 672
completed 4 years follow-up | 35040
hyperchloremic metabolic acidosis complication | 0
delayed diagnosis | 0
early referral to surgical team | 0
oral alkalizing agents (sodium bicarbonate) | 0
ileal conduit as alternative diversion | 0
