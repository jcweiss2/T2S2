36 years old | 0
    male | 0
    hospitalized | 0
    low back pain | -96
    bruised hips | -96
    macroscopic hematuria | -96
    gingival bleeding | -96
    conscious | 0
    oriented | 0
    pale | 0
    tachycardic (108 beats per minute) | 0
    blood pressure 120/90 mmHg | 0
    mild edema | 0
    varicose veins of the lower limbs | 0
    chronic malleolar ulcers | 0
    bleeding in pelvic region | 0
    bruising in pelvic region | 0
    denied personal history of bleeding diathesis | 0
    denied family history of bleeding diathesis | 0
    ruled out renal diseases | 0
    ruled out urological diseases | 0
    hemoglobin level 4.8 g/dL | 0
    platelet count 270 × 10^9/L | 0
    incoagulable blood (PT) | 0
    incoagulable blood (APTT) | 0
    transfusion of red blood cells | 0
    transfusion of cryoprecipitate | 0
    transfusion of fresh frozen plasma | 0
    transferred to intensive care unit | 0
    hematuria | 48
    ecchymosis | 48
    incoagulable blood (PT) | 48
    patient-to-control APTT ratio 1.79 | 48
    continued transfusion support | 48
    positive lupus anticoagulant antibodies | 48
    negative anticardiolipin IgM antibodies | 48
    negative anticardiolipin IgG antibodies | 48
    negative anticardiolipin IgA antibodies | 48
    negative antinuclear factors | 48
    negative rheumatoid factors | 48
    factor VII activity 3% | 48
    factor II activity 130% | 48
    factor V activity 150% | 48
    factor VIII activity >200% | 48
    factor IX activity 47% | 48
    factor X activity 75.8% | 48
    started intravenous pulse therapy with methylprednisolone | 48
    administered prothrombin complex concentrate | 48
    recovered well | 408
    no bleeding | 408
    maintained oral prednisone 1 mg/kg/day | 408
    discharged | 408
    referred to outpatient clinic | 408
    reduced corticoid dose | 408
    consecutive PT tests progressive toward normality | 408
    condition stabilized | 408
    no new hemorrhagic episodes | 408
    suspended corticoid treatment | 2160
    PT 83.2% | 2400
    patient-to-control APTT ratio 1.05 | 2400
    fibrinogen level 248.7 mg/dL | 2400
    FVII activity 60.6% | 2400
    <|eot_id|>