57 years old | 0
male | 0
admitted to the hospital | 0
generalized weakness | -336
fatigue | -336
confusion | -336
dizziness | -336
mild jaundice | -336
hypertension | 0
diabetes mellitus | 0
hyperlipidemia | 0
hypothyroidism | 0
former smoker | 0
consumed alcohol occasionally | 0
anemia | 0
thrombocytopenia | 0
acute liver injury | 0
acute renal failure | 0
intermittent hemodialysis | 0
lactic acidosis | 0
sepsis | 0
worsening hepatic encephalopathy | 0
febrile | 0
hemoglobin 7.5 g/dL | 0
platelets 26,000/mm3 | 0
creatinine 4.34 mg/dL | 0
total bilirubin 19 mg/dL | 0
alanine aminotransferase 395 U/L | 0
aspartate aminotransferase 261 U/L | 0
serum lactate 10 mmol/L | 0
serum ferritin >40,000 ng/mL | 0
serum triglycerides 556 mg/dL | 0
coagulopathic | 0
international normalized ratio 4.2 | 0
fibrinogen <70 mg/dL | 0
MELD score >40 | 0
emergent liver transplant evaluation | 0
hepatic steatosis | 0
splenomegaly | 0
multiple splenic infarcts | 0
right axillary and retropectal lymphadenopathy | 0
mechanical ventilation | 24
circulatory shock | 24
vasopressor support | 24
worsening renal failure | 24
continuous renal replacement therapy | 24
bone marrow biopsy | 24
no evidence of leukemia | 24
no evidence of lymphoma | 24
no evidence of HLH | 24
transjugular liver biopsy | 48
diffuse large B-cell lymphoma | 48
fever | 48
bicytopenia | 48
splenomegaly | 48
ferritin level | 48
hypertriglyceridemia | 48
chemotherapy | 72
dexamethasone | 72
ifosfamide | 72
carboplatin | 72
etoposide | 72
worsening metabolic acidosis | 96
hypoglycemia | 96
shock | 96
subdural hemorrhages | 96
generalized tonic-clonic seizures | 96
comfort care measures | 120
death | 120