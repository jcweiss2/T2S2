47 years old | 0
male | 0
alcohol-induced dilated cardiomyopathy | -10000
chronic atrial fibrillation | -10000
excess alcohol consumption | -17520
hospitalized for heart failure | -1000
admitted to the hospital | 0
New York Heart Association class IV dyspnea | 0
dyspnea | 0
azotemia | 0
dobutamine infusion | 0
milrinone infusion | 0
continuous renal replacement therapy | 0
cardiac arrest | 792
ventricular fibrillation | 792
cardiopulmonary resuscitation | 792
transthoracic echocardiography | 0
decreased left ventricular systolic function | 0
decreased right ventricular systolic function | 0
severe mitral regurgitation | 0
severe tricuspid regurgitation | 0
dilated inferior vena cava | 0
pericardial effusion | 0
severe cardiomegaly | 0
elevated serum creatinine | 0
elevated total bilirubin | 0
psychiatric evaluation | 0
psychosocial support | 0
left ventricular assist device insertion | 1176
tricuspid annuloplasty | 1176
surgery | 1176
median sternotomy | 1176
cardiopulmonary bypass | 1176
beating heart tricuspid annuloplasty | 1176
LVAD inflow cannula | 1176
LVAD outflow cannula | 1176
inotropic support | 1176
stable vital signs | 1176
transfer to cardiovascular ICU | 1176
hypotension | 1176
tachycardia | 1176
inotrope infusion | 1176
nitric oxide inhalation | 1176
unstable | 1176
emergent RVAD insertion | 1176
veno-pulmonary artery extracorporeal life support | 1176
percutaneous femoral venous cannulation | 1176
pulmonary artery cannulation | 1176
left anterior mini-thoracotomy | 1176
RVAD initiation | 1176
stable hemodynamics | 1180
inhaled nitric oxide tapered | 1180
RVAD rpm and flow rates decreased | 1180
spontaneous recovery of right ventricular systolic function | 1180
RVAD removal | 1200
thoracotomy closure | 1200
transfer to general ward | 1272
resolution of lower leg pitting edema | 1296
rehabilitation therapy | 1296
discharged | 1296
readmitted for recurrent alcohol abuse | 22752
right ventricular failure | 22752
LVAD turned off | 22752
septic encephalopathy | 22752
coma | 22752