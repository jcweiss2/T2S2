77 years old | 0
male | 0
admitted to the hospital | 0
progressive lethargy | -72
shortness of breath | -72
septic shock | 0
hypotension | 0
hypoxia | 0
ventilatory support | 0
vasopressor support | 0
tube thoracostomy | 0
large left pleural effusion | 0
purulent fluid | 0
splenectomy | -8760
chemotherapy | -8760
non-Hodgkin's B-cell lymphoma | -8760
tumor recurrence | -5040
radiation therapy | -5040
progressive dysphagia | -1008
home TPN | -1008
EGD | -336
bleeding gastric ulcer | -336
cauterization | -336
chest CT | 24
abdominal CT | 24
oral contrast in chest tube | 24
upper gastrointestinal series | 48
gastropleural fistula | 48
diagnostic laparoscopy | 72
bulky tumor | 72
laparoscopic GPF takedown | 72
partial sleeve gastrectomy | 72
intraoperative EGD | 72
fistulous tract patched | 72
bovine pericardium mesh | 72
closed suction drain | 72
feeding jejunostomy tube | 72
malignant B-cell lymphoma | 72
quick initial recovery | 96
early extubation | 96
transfer out of ICU | 96
persistent anorexia | 120
pulmonary complications | 120
left thoracotomy | 240
pulmonary decortication | 240
debridement of empyema | 240
discharged home | 2160
died | 2208