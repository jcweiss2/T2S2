68 years old | 0
male | 0
presented to the emergency room (ER) | 0
progressive bullous and erosive skin lesions involving the whole body | 0
painful oral ulcer | -336
bilateral enlarged supraclavicular lymph nodes | -336
metastatic squamous cell carcinoma | -336
diagnosed with diabetes | -175200
treated with diabetic nephropathy | -70080
blood pressure 93/64 mmHg | 0
heart rate 91/min | 0
respiration rate 20/min | 0
flaccid blisters | 0
exfoliated skin | 0
crusted erosions involving eyelids | 0
buccal mucosa lesions | 0
tongue lesions | 0
trunk lesions | 0
back lesions | 0
extremities lesions | 0
anemia | 0
thrombocytopenia | 0
white blood count 5,170/mm3 | 0
hemoglobin 7.7 mg/dL | 0
platelets 426,000/mm3 | 0
azotemia | 0
blood urea nitrogen 52.3 mg/dL | 0
creatinine 2.98 mg/dL | 0
diabetic nephropathy | 0
multiple cervical lymph node enlargement | 0
mediastinal lymph node enlargement | 0
increased fluorodeoxyglucose uptake | 0
deep ulcerative mass on mid to distal esophagus | 0
moderately differentiated squamous cell carcinoma | 0
suprabasal acantholysis | 0
bullous cleft formation | 0
C3 deposits in the basal layer of mucosa | 0
esophageal cancer stage IVB | 0
rapid aggravation of skin lesion | 0
rapid aggravation of general condition | 0
admitted to the intensive care unit | 0
palliative combination chemotherapy with fluorouracil and carboplatin | 0
intravenous methylprednisolone 40 mg/day | 0
skin lesion worsened | 96
extensive skin defects | 96
progressive exfoliation | 96
increased discharge | 96
neutropenic fever | 144
broad spectrum antibiotics | 144
expired due to overwhelming sepsis | 216
