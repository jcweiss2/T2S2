36 years old| 0
    female | 0
    pregnant | 0
    uterine fibroid | -624
    hypercalcemic crisis | -72
    recurrent vomiting | -72
    epigastric pain | -72
    weight loss (10 kg) | -624
    no change in bowel habits | -72
    no hematemesis | -72
    no rectal bleeding | -72
    no history of hematuria | -72
    no passing stones | -72
    using iron tablets | 0
    ill appearance | 0
    marked dehydration | 0
    drowsiness | 0
    blood pressure 126/76 mmHg | 0
    pulse rate 94 min–1 | 0
    respiratory rate 30 min–1 | 0
    temperature 36.6°C | 0
    no lymphadenopathy | 0
    no thyromegaly | 0
    no edema | 0
    uterus size of 40 weeks | 0
    tender epigastric area | 0
    hypotonia | 0
    brisk deep tendon reflexes | 0
    no focal neurological signs | 0
    down-going plantar reflexes | 0
    chest unremarkable | 0
    cardiovascular system unremarkable | 0
    hemoglobin 8.7 g/dl | 0
    WBCs 7000 μl–1 | 0
    platelets 445000 μl–1 | 0
    ESR 109 mm/h | 0
    toxic granulation of WBCs | 0
    BUN 4.4 mmol/l | 0
    creatinine 59 μmol/l | 0
    HCO3 22 mmol/l | 0
    Na 138 mmol/l | 0
    Ca 4.8 mmol/l | 0
    uric acid 508 μmol/l | 0
    lactic acid 1.2 mmol/l | 0
    phosphorous 0.8 mmol/l | 0
    HIV negative | 0
    calcium at 14 weeks’ gestation 2.43 mmol/l | -1680
    ALT 4 u/l | 0
    AST 11 u/l | 0
    ALP 150 u/l | 0
    total protein 72 g/l | 0
    albumin 30 g/l | 0
    cholesterol 4.05 mmol/l | 0
    triglyceride 3.59 mmol/l | 0
    PTH 3 pg/ml | 0
    TSH 0.68 mIU/l | 0
    free thyroxin 16.6 pmol/l | 0
    cortisol 1849 nmol/l | 0
    vitamin D 15 ng/ml | 0
    normal serum protein electrophoresis | 0
    normal angiotensin-converting enzyme level | 0
    normal saline infusion | 0
    intramuscular calcitonin | 0
    transferred to medical ICU | 0
    diagnosis of humoral hypercalcemia of benignancy (uterine fibroid) | 0
    rupture membrane | 24
    urgent cesarean section | 24
    hypercalcemia | 0
    reduced urine output | 24
    rise in serum creatinine | 24
    hemodialysis | 24
    surgery complicated by bleeding | 24
    hypotension | 24
    blood transfusion | 24
    delivery of baby girl (2.9 kg) | 24
    removal of uterine masses (30 × 25 × 15 cm) | 24
    histopathology consistent with leiomyoma with calcifications | 24
    no evidence of malignancy | 24
    postoperative serum calcium 2.34 mmol/l | 24
    phosphorus 1.1 mmol/l | 24
    BUN 6.2 mmol/l | 24
    Cr 75 mmol/l | 24
    Na 143 mmol/l | 24
    K 4.2 mmol/l | 24
    HCO3 16 mEq/l | 24
    chloride 113 mEq/l | 24
    albumin 21 g/l | 24
    serum lactate 5.19 | 24
    serum PTH 155 pg/ml | 24
    serum amylase 88 u/l | 24
    serum lipase 73 u/l | 24
    Hb 5.8 g/dl | 24
    platelets 125000 μl–1 | 24
    CT scan chest and pelvis (no mass lesion or organomegaly) | 24
    MRI brain (infarcts right cerebellum, lentiform nucleus, frontal, parietal, occipital lobes) | 24
    MRA (vasospasm internal carotid, middle and anterior carotid arteries) | 24
    diffuse ischemic changes secondary to hypoxic insult | 24
    condition improvement | 48
    neurological status requiring physiotherapy | 48
    generalized muscle weakness | 48
    stiffness | 48
    discharged home | 96
    final diagnosis of humoral hypercalcemia associated with uterine fibroid | 96
    serum calcium remained normal over 6 months | 4320
    <|eot_id|>
    