72 years old | 0
woman | 0
admitted to the hospital | 0
general weakness | 0
poor oral intake | 0
bilateral knee joint pain | -2928
symptoms exacerbated | -2928
osteoarthritis | -1344
intra-articular steroid injections | -1344
triamcinolone acetonide (Kenalog-40) | -1344
glucose monitoring not performed | -1344
knee joint pain reduced | -1344
cholecystectomy | -175200
random glucose level normal | -175200
weight gain | -1344
mild systemic edema | -1344
cushing's syndrome | -1344
blood pressure 120/80 mm Hg | 0
pulse 98 beats per minute | 0
respiratory rate 20 breaths per minute | 0
body temperature 37.9℃ | 0
acute ill appearance | 0
constantly sleepy | 0
multiple ulcers | 0
whitish patches in oral mucosa | 0
mild crackle sound in entire lung field | 0
hemoglobin 15.3 g/dL | 0
white blood cell count 13×103/mL | 0
neutrophil 96.3% | 0
lymphocyte 3.1% | 0
monocyte 0.6% | 0
platelet count 349×103/µL | 0
random blood glucose 174 mg/dL | 0
Hb A1C 7.7% | 0
fasting plasma C-peptide 6.1 ng/mL | 0
serum albumin 2.4 g/dL | 0
C-reactive protein 13.37 mg/dL | 0
human immunodeficiency virus test negative | 0
T3 10 ng/dL | 0
free T4 1.2 ng/dL | 0
thyroid stimulating hormone 30 mIU/mL | 0
sick euthyroid state | 0
rapid adrenocorticotropic hormone stimulation test | 0
basal cortisol 0.55 µg/dL | 0
30 minute cortisol 6.3 µg/dL | 0
90 minute cortisol 5.5 µg/dL | 0
adrenal insufficiency | 0
chest X-ray multiple cavitary nodules | 0
chest computed tomography mass and cavitary nodules | 0
percutaneous needle biopsy | 72
fungal hypae with acute angle branching | 72
rare fruit body | 72
invasive aspergillosis involving lungs | 72
diabetes caused by intraarticular corticosteroid injection | 72
amphotericin B intravenous | 120
unconscious | 144
brain MRI | 144
cerebrospinal fluid tapping | 144
MRI numerous thin peripheral enhancing cystic nodules | 144
CSF non-specific findings | 144
invasive aspergillosis involving brain | 144
amphotericin B continued | 144
condition deteriorated | 144
transferred to intensive care unit | 168
ventilator care | 168
voriconazole | 168
condition deteriorated daily | 168
died | 336
respiratory failure | 336
septic shock | 336
