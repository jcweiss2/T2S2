hospitalized for cardiogenic shock | 0
diagnosed with biventricular failure | 0
ejection fraction 5–10% | 0
imaging concerning for myopericarditis and constrictive physiology | 0
PICC line placed | 0
discharged on milrinone | 0
presented to Emergency Department with septic shock | -48
PICC line removed | -48
started on IV vancomycin and piperacillin/tazobactam | -48
transferred to intensive care unit for vasopressor support | -48
Chryseobacterium indologenes grew from his admission PICC line and peripheral blood cultures | -24
antibiotics were changed to ciprofloxacin and piperacillin/tazobactam | -24
weaned off vasopressor support | -24
underwent pericardiectomy | 8
completed 14 days of antibiotics | 14
discharged from the hospital off inotropes with stable vital signs and labs | 21
seen in outpatient cardiology clinic, remains in good health with no evidence of recurrent infection | 365
fevers/chills | -48
tachycardia | -48
blood pressure of 96/57 mmHg | -48
heart that was tachycardic, but normal rhythm without any murmurs, rubs, or gallops | -48
no signs of elevated jugular venous pressure | -48
no lower extremity oedema | -48
bilateral radial and dorsalis pedis pulses were equal and 2+ bilaterally | -48
lungs were clear to auscultation bilaterally | -48
no redness or drainage around the PICC line | -48
chest X-ray showed no abnormalities | -48
electrocardiogram was significant for sinus tachycardia | -48
became febrile to 39.5°C | -48
developed severe rigours | -48
hypotension with blood pressure in 70 s/40s mmHg | -48
elevated lactate level of 5.5 mmol/L | -48
blood cultures were drawn | -48
started on empiric vancomycin and piperacillin/tazobactam | -48
transferred to the cardiac intensive care unit | -48
preliminary report of his blood cultures revealed Gram-negative rods | -24
cultures drawn from the PICC line became positive for growth | -24
infectious disease team was consulted | -24
started on ciprofloxacin | -24
susceptibility testing on the isolated C. indologenes demonstrated sensitivity to ciprofloxacin | -24
improved clinically on treatment with antibiotics | -10
remained afebrile | -10
weaned off vasopressor support | -10
follow-up blood cultures remained negative | -10
interval echocardiogram showed a dilated and hypertrophied left ventricle | -10
diastolic septal bounce consistent with constrictive pericarditis | -10
EF of 30–35% | -10
right ventricle was dilated with reduced systolic function | -10
no evidence of valvular stenosis, regurgitation, or vegetations | -10
simultaneous right and left heart catheterization demonstrated discordance of the right and left ventricular pressures | -10
diastolic equalization of pressures supporting the diagnosis of constrictive pericarditis | -10
pericardiectomy | 8
completed 14 days of antibiotics | 14
discharged from the hospital off inotropes | 21
inotrope independent | 21
guideline-directed medical therapy for heart failure with reduced EF | 21
furosemide 40 mg once daily | 21
metoprolol succinate 12.5 mg once daily | 21
sacubitril-valsartan 24–26 mg every 12 h | 21
follow-up transthoracic echocardiogram performed 5 days after the pericardiectomy | 13
left ventricular EF had increased to 50–55% | 13
right ventricular systolic dysfunction had improved | 13
no evidence of recurrent infection | 365
reported great improvement in his functional status | 365
denied any symptoms of heart failure | 365
classified as NYHA Class I | 365