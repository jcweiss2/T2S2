23 years old | 0
G2P1L1 | 0
28 weeks gestation | 0
previous normal vaginal delivery | -672
admitted to emergency labor room | 0
state of shock | 0
unconscious | 0
unrecordable blood pressure | 0
unrecordable pulse | 0
unrecordable fetal heart sound | 0
history of amenorrhea | -1968
bleeding per vaginam | -24
no history of drug abuse | 0
no history of alcohol intake | 0
large bore intravenous cannula secured | 0
i.v fluids started | 0
Foley's catheter put | 0
urine output measured | 0
urine sent for albumin | 0
albumin test negative | 0
electrolytes within normal limits | 0
blood sugar level 84 mg% | 0
emergency ultrasound | 0
absent fetal heart | 0
shifted to Intensive Care Unit | 0
cardiac arrest | 0
wedge kept under right hip | 0
chest compressions started | 0
intubated with endotracheal tube | 0
rescue breaths given | 0
injection adrenaline given | 0
inotropes started | 0
dopamine started | 0
noradrenaline started | 0
shifted to ICU | 0
put on ventilator | 0
SIMV-VC mode | 0
FiO2 100% | 0
tidal volume 500 ml | 0
PEEP Off | 0
PSV 15 | 0
BP 92/60 mmHg | 0
pulse rate 120 bpm | 0
SPO2 95% | 0
managed with whole blood | 0
vasopressors continued | 0
second bout of bleeding per vaginam | 1
P/A examination done | 1
uterus measured at 28 weeks | 1
oblique lie | 1
ultrasound scan showed Grade 4 placenta previa | 1
shifted to operation theater | 2
emergency lower segment cesarean section | 2
i.v ketamine given | 2
vecuronium given | 2
isoflurane given | 2
dead baby extracted | 2
placenta removed | 2
uterus closed in layers | 2
whole blood transfusions | 2
Ringer lactate transfused | 2
fresh frozen plasma transfused | 2
blood samples taken | 2
shifted back to ICU | 4
put on ventilator | 4
SIMV-VC mode | 4
FiO2 50% | 4
tidal volume 500 ml | 4
PEEP 3 | 4
PSV 15 | 4
stable with vitals | 4
BP 120/72 mm Hg | 4
pulse rate 115 bpm | 4
SpO2 95% | 4
inotropes tapered off | 96
regained consciousness | 168
responded to verbal commands | 168
weaned off from ventilator | 168
shifted to ward | 216
discharged | 216
intact neurological functions | 216