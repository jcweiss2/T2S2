19 years old | 0
nulliparous | 0
mammary ptosis | 0
mammary asymmetry | 0
history of surgery for appendicitis | - (approximated to a prior event but no specific time given; as appendicitis surgery is unrelated to current admission, timestamp remains 0 unless specified)
5 tattoos without complications | 0
mastopexy with placement of 240-mL silicone implants | 0
discharged from hospital | 0
returned to clinic with ulceration and necrosis at incision | 96 (4 days after discharge, discharge time is 0)
no secretions | 96
no fever | 96
tachycardic | 96
arterial hypotension | 96
hemoglobin 7.5 g/dL | 96
hematocrit 23% | 96
leukocytes 64,500/mm³ | 96
C-reactive protein >270 mg/L | 96
low levels of total proteins and fractions (4.10 g/dL) | 96
serum albumin 2.0 g/dL | 96
globulins 2.1 g/dL | 96
transferred to intensive care unit | 96
suspected infection of the surgical site | 96
sepsis | 96
received systemic vancomycin | 96
received meronem for 20 days | 96
received daptomycin (Cubicin) | 96
local wound care with saline solution | 96
local wound care with chlorhexidine antiseptic | 96
alternated between rifampicin and silver sulfadiazine | 96
surgical removal of silicone implants | 216 (9 days after initial surgery; initial surgery was at 0)
rinsed with 2 L saline | 216
garamycin 80 mg | 216
kefazol 1 g | 216
breasts reconstructed using mononylon sutures | 216
samples taken and cultured | 216
no bacterial growth in samples from breast region | 216
no bacterial growth in other areas of the body | 216
no bacterial growth in blood culture | 216
no bacterial growth in surgical instruments, autoclave, etc. | 216
biopsies of edges of surgical wound sent to 2 different labs | 216
dermatitis | 216
diffuse neutrophilic panniculitis | 216
necrosis | 216
new dehiscence of entire surgical wound | 264 (3 days after second surgery; second surgery was at 216)
large area of necrosis | 264
no secretion | 264
rapid and progressive aggravation of lesion | 264
worsening of general clinical condition | 264
dressings changed under analgesia | 264
delimitation of necrotic area achieved | 264
each wound reaching 20×25 cm | 264
wound care using negative pressure VAC | 264
hydrophobic polyurethane foam sponges with silver introduced | 264
4 VAC changes at 2- to 4-day intervals | 264
purplish secretion aspirated by VAC machine | 264
worsening of patient’s clinical condition | 264
anasarca | 264
introduced prednisone 40 mg/d | 312 (6 days after second surgery; second surgery at 216)
prednisone increased up to 125 mg/d | 312
patient’s general condition improved | 312
granulation tissue observed | 312
contraction of wound edges | 312
adherence between pectoralis major muscle and glandular tissue | 312
used hydrophobic polyvinyl alcohol (white) foam | 312
3 VAC foam changes | 312
deep mononylon sutures placed | 312
surgical remodeling of breast cone | 696 (29 days after initial surgery; 29 days *24 = 696)
improved appearance of wound after 4 foam changes | 696
creating symmetry in nipple–areola complex | 744 (31 days *24 = 744)
seventh VAC change | 960 (40 days *24 = 960)
surgical wound improved after 27 days of VAC therapy | (27 days after VAC started at 264; 27*24=648; 264+648=912)
discharged 42 days after original surgery | 1008 (42 days *24 = 1008)
prednisone 60 mg/d at discharge | 1008
outpatient wound care | 1008
progressive improvement in wound’s appearance | 1008
corticosteroids gradually reduced | (over time after discharge, but discharge is timestamp 1008)
corticosteroids suspended after 4 months | (4 months after discharge; 4*30*24=2880; 1008+2880=3888)
initial sensitivity in areola and nipple | 1824 (7 months after procedure; 7*30*24=5040, but procedure was at 0, so 7*30=210 days *24=5040; but in the case, "Seven months after the procedure" would be 7*30*24=5040)
history of surgery for appendicitis | - (prior event but no specific time given, so timestamp remains 0)
returned to clinic with ulceration and necrosis at incision | 96
surgical removal of silicone implants | 216
new dehiscence of entire surgical wound | 264
introduced prednisone 40 mg/d | 312
surgical remodeling of breast cone | 696
creating symmetry in nipple–areola complex | 744
seventh VAC change | 960
surgical wound improved after 27 days of VAC therapy | 912
discharged 42 days after original surgery | 1008
corticosteroids gradually reduced | 1008
corticosteroids suspended after 4 months | 3888
initial sensitivity in areola and nipple | 5040
