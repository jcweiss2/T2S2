43 years old|0
man|0
presented to emergency room|0
history of consuming 12 g aluminum phosphide|-24
history of consuming four tablets aluminum phosphide|-24
aluminum phosphide poisoning|0
abdominal pain|0
bowel incontinence|0
breathlessness|0
heart rate 113/min|0
blood pressure 60 systolic|0
respiratory rate 48/min|0
saturation not recordable|0
profound shock|0
resuscitated with fluid bolus 30 ml/kg|0
initiated on dual inotropes|0
refractory shock|0
point-of-care echocardiogram|0
severe left ventricular dysfunction|0
ejection fraction 15%|0
severe hemodynamic compromise|0
rapid sequence intubation|0
ketamine|0
rocuronium|0
preintubation arterial blood gas|0
severe metabolic acidosis|0
pH 6.98|0
bicarbonate 8|0
lactate levels 146|0
intravenous sodium bicarbonate 100 milli equivalence|0
sodium bicarbonate 50 milliequivalents repeated every 15 min|0
intravenous magnesium sulfate 3 g|0
magnesium sulfate 6 g per 24-h infusion|0
heart rate dropped to 35/min|0
intravenous atropine every 4 min|0
maximum 3 doses atropine|0
transient variable heart blocks|0
planned to proceed with ECMO|0
venoarterial ECMO performed|0
19 French right femoral artery cannula|0
29 French right femoral venous cannula|0
8 French distal perfusion cannula|0
post-ECMO vitals stabilized|24
shifted to intensive care unit|24
decannulated on 3rd day|72
bilateral cerebral infarcts|72
acute kidney injury|72
renal replacement therapy initiated|72
coagulopathy|72
multiple blood transfusions|72
lower respiratory tract infection|72
Elizabethkingia meningoseptica infection|72
minocycline started|72
reactive pleural effusion|72
intercostal drainage placed|72
intercostal drainage removed|72
admitted to hospital for 41 days|0
managed by multidisciplinary team|0
discharged home|984
no neurological deficits|984
improving kidney function|984
