32 years old | 0
female | 0
history of intravenous drug use | -672
attention deficit/hyperactivity disorder | -672
fever | -168
chills | -168
generalized weakness | -168
shortness of breath | -72
non-smoker | 0
no alcohol consumption | 0
abusing fentanyl intravenously | -672
dextroamphetamine/amphetamine | -672
Temperature 102.7 °Fahrenheit | 0
blood pressure 102/56 mmHg | 0
pulse 136 beats per minute | 0
respiratory rate 38 breaths per minute | 0
oxygen saturation 94% on room air | 0
moderate respiratory distress | 0
bilateral rhonchi | 0
tachycardia | 0
no murmur, rub or gallop | 0
WBC 12,200/mm3 | 0
hemoglobin 10.9 g/dL | 0
platelet count 85,000/mm3 | 0
ESR 60 mm/hr | 0
hyponatremia | 0
sodium 124 mmol/L | 0
creatinine level 2.8 mg/dL | 0
BUN 98 mg/dL | 0
NT-proBNP 1028 pg/mL | 0
sinus tachycardia | 0
bilateral lower lobe infiltrates | 0
small pleural effusions | 0
IV fluids | 0
levofloxacin | 0
septic shock | 24
acute respiratory failure | 24
pressors | 24
mechanical ventilation | 24
gram-positive cocci | 24
vancomycin | 24
vegetation at the tip of anterior leaflet of tricuspid valve | 24
moderate-to-severe tricuspid regurgitation | 24
patent foramen ovale | 24
shunt | 24
septic emboli | 24
non-oliguric AKI | 24
renal replacement therapy | 24
acute tubular necrosis | 24
MSSA | 72
oxacillin | 72
improved on supportive and antimicrobial therapy | 168
weaned off pressors | 168
extubated | 168
renal function started to recover | 168
bilateral nontender purpuric papules | 216
bullous lesions | 240
no mucosal or palmar involvement | 216
no abdominal pain | 216
no arthralgias | 216
no paresthesia | 216
no fever | 216
no chills | 216
HIV antibody negative | 216
hepatitis B serology negative | 216
p-ANCA negative | 216
c-ANCA negative | 216
cryoglobulin negative | 216
rheumatoid factor negative | 216
ANA weakly positive | 216
anti-ds DNA antibody negative | 216
Complement C3 low | 216
Complement C4 normal | 216
anti-HCV antibody positive | 216
HCV viral load 4.16 × 105 IU/mL | 216
no significant changes in red blood count | 216
no significant changes in leukocyte count | 216
no significant changes in kidney function | 216
eosinophil count normal | 216
no bacteria in aspirated fluid | 216
no organisms on gram staining | 216
perivascular neutrophil infiltration | 216
fibrinoid necrosis of small vessels | 216
leukocytoclastic vasculitis | 216
vancomycin | 216
resolution of skin lesions | 264
tricuspid valve replacement surgery | 720
no perioperative complications | 720
no recurrence of skin lesions | 744