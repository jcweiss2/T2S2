36 years old | 0
male | 0
admitted to the hospital | 0
IgA nephropathy | 0
hemodialysis | 0
left forearm arteriovenous fistula (AVF) | 0
hepatitis B | 0
hypertension | 0
Charcot-Marie-Tooth disease | 0
sudden onset of left flank pain | 0
constant pain | 0
non-radiating pain | 0
pain aggravated with deep breaths | 0
denied fever | 0
denied chest pain | 0
denied shortness of breath | 0
denied cough | 0
denied vomiting | 0
denied diarrhea | 0
denied dysuria | 0
denied prior problems with the AVF | 0
temperature 98.5°F (36.9°C) | 0
temperature 102.3°F (39.0°C) | 24
pulse 108 beats per minute | 0
respiratory rate 17 cycles per minute | 0
blood pressure 106/64 mmHg | 0
oxygen saturation 99% | 0
mild distress due to pain | 0
soft abdomen | 0
non-tender abdomen | 0
no costovertebral angle tenderness | 0
AVF site not tender | 0
normal sinus rhythm on ECG | 0
white blood cell (WBC) 10.2 k/ul | 0
WBC peak 41.9 k/ul | 192
WBC peak 36.5 k/ul | 192
WBC 10.2 k/ul on day 19 | 456
hemoglobin 10.9 g/dl | 0
platelets 197 k/ul | 0
erythrocyte sedimentation rate 48 | 0
procalcitonin >200 ng/dl | 0
C-reactive protein 4.81 mg/dl | 0
sodium 134 mmol/l | 0
potassium 4.2 mmol/l | 0
chloride 91 mmol/l | 0
bicarbonate 27 mmol/l | 0
blood urea nitrogen 66 mg/dl | 0
creatinine 12.4 mg/dl | 0
urinalysis WBC 1/HPF | 0
absence of bacteria in urinalysis | 0
absence of leukocyte esterase in urinalysis | 0
absence of nitrate in urinalysis | 0
chest x-ray (CXR) clear lungs | 0
CT abdomen and pelvis no acute appendicitis | 0
CT abdomen and pelvis no diverticulitis | 0
CT abdomen and pelvis no mechanical bowel obstruction | 0
CT abdomen and pelvis no ascites | 0
CT abdomen and pelvis no portal hypertension | 0
atrophic kidneys | 0
open wound at AVF noticed | 24
AVF wound swabbed and cultured | 24
AVF wound dressed regularly | 24
AVF wound culture grew Streptococcus group A (GAS) | 24
WBC increased to 12.5 k/ul | 24
hypotension | 24
blood cultures drawn | 24
vancomycin initiated | 24
meropenem initiated | 24
right internal jugular (IJ) hemodialysis catheter inserted | 24
transferred to Medical Intensive Care Unit | 24
blood pressure improved with IV fluids | 24
CXR moderate left pleural effusion | 24
chest CT very large left pleural effusion | 48
chest CT near-complete atelectasis left upper lobe | 48
chest CT complete atelectasis left lower lobe | 48
CXR near-complete opacification left lung | 48
CXR mediastinal shift to the right | 48
pigtail chest tube inserted | 48
CXR resolved large left pleural effusion | 48
1.3 L pleural fluid removed | 48
pleural fluid cloudy | 48
pleural fluid WBC 15,762/cumm | 48
pleural fluid RBC 3,556/cumm | 48
pleural fluid polynuclear white blood cells 84% | 48
pleural fluid glucose 2 mg/dL | 48
pleural fluid total protein 4.2 | 48
pleural fluid LDH 9208 u/L | 48
serum protein 5.1 g/dl | 48
serum LDH 150 u/l | 48
exudative pleural fluid (Light’s criteria) | 48
clindamycin added | 48
CXR small residual left effusion | 168
chest tube removed | 168
pain at chest tube insertion site | 168
CXR re-accumulation of pleural fluid | 192
VATS performed | 192
pleural drainage and decortication | 192
3 chest tubes inserted (anterior, lateral, posterior) | 192
chest CT improved left hemithorax | 240
chest CT loculated pleural effusion/emphysema | 240
chest CT small residual area 1.5 cm | 240
chest CT right-sided pleural effusion | 240
left anterior chest tube removed | 288
left lateral chest tube removed | 288
left posterior chest tube removed | 360
sepsis | 24
intermittent fever spikes | 24
tachycardia | 24
tachypnea | 24
hypotension requiring IV fluids | 24
vital signs improved | 72
negative blood cultures | 0
negative pleural fluid cultures | 48
transthoracic echocardiogram no valvular vegetations | 0
regular dialysis via temporary jugular catheter | 24
discharged with right tunneled permanent catheter | 648
AVF revised and repaired | 192
meropenem discontinued after 12 days | 288
clindamycin discontinued after 11 days | 264
switched to ceftriaxone | 288
ceftriaxone for 14 days | 288
vancomycin continued for 6 weeks | 648
gradual recovery | 648
discharged after 27 days | 648
explosive pleuritis | 48
AVF infection source | 24
no respiratory tract infection | 0
no pneumonia | 0
no endocarditis | 0
negative microbiological evidence of bacteremia | 0
pyrexia | 24
leukocytosis | 24
elevated inflammatory markers | 24
oozing from AVF | 24
GAS identified in AVF culture | 24
explosive pleuritis within 48 hours | 48
fluid reaccumulation | 192
VATS decortication | 192
temporary hemodialysis catheter | 24
permanent tunneled catheter at discharge | 648
antibiotics duration adjusted | 648
rare phenomenon | 0
no identifiable risk factors | 0
no apparent sources of infection | 0
