32 years old | 0
female | 0
admitted to the hospital | 0
JAK2 mutation-negative essential thrombocythemia | -6912
treated by pipobroman | -6912
treated by hydroxyurea | -576
treated by anagrelide | -432
asthenia | -120
gradual decrease in hemoglobin level | -120
anagrelide stopped | -120
bone marrow biopsy | -120
grade 2 myelofibrosis | -120
blastic cells in peripheral blood | -84
acute myeloid leukemia | -84
allogeneic bone marrow hematopoietic stem-cell transplantation | 0
admitted to intensive care unit | 0
acute respiratory distress syndrome | 0
Staphylococcus aureus | 0
Escherichia coli | 0
broad-spectrum antibiotherapy | 0
furosemide | 0
oral fluconazole prophylaxis | 0
readmitted to ICU | 12
septic shock | 12
empirical antibiotherapy | 12
afebrile | 12
Graft-versus-Host Disease | 37
corticosteroids | 37
inolimomab | 37
sirolimus | 37
basiliximab | 37
digestive disorders | 37
hemorrhagic manifestations | 37
new antibiotic regimen | 63
intravenous caspofungin | 63
Candida albicans | 63
Candida kefyr | 63
caspofungin stopped | 192
oral fluconazole | 192
unexplained fever | 216
thoracic computed tomography | 216
pulmonary nodules | 216
pulmonary aspergillosis | 216
voriconazole | 216
serum galactomannan assay | 216
bronchoalveolar lavage | 216
(1→3)-β-d-glucan antigenemia | 234
deep candidiasis | 234
caspofungin | 234
acute renal failure | 240
multiple organ failure | 240
death | 240