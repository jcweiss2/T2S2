43 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
difficult-to-manage bronchial asthma | 0 | 0 | Factual
hospitalized in the last 8 months on 10 occasions | -672 | 0 | Factual
acute exacerbations | -672 | 0 | Factual
asthmatic crisis | -672 | 0 | Factual
24-hour history of dry cough | -24 | 0 | Factual
progressive dyspnea | -24 | 0 | Factual
psychomotor agitation | -24 | 0 | Factual
audible wheezing | -24 | 0 | Factual
salbutamol | -24 | 0 | Factual
ipratropium bromide | -24 | 0 | Factual
critical condition | 0 | 0 | Factual
diaphoretic | 0 | 0 | Factual
tachycardic | 0 | 0 | Factual
dyspneic | 0 | 0 | Factual
supraclavicular retractions | 0 | 0 | Factual
respiratory rate of 30 breaths/minute | 0 | 0 | Factual
ambient oxygen saturation 87% | 0 | 0 | Factual
auscultation with abolished vesicular murmur | 0 | 0 | Factual
Glasgow coma scale 12/15 | 0 | 0 | Factual
arterial blood gases analysis | 0 | 0 | Factual
respiratory acidosis | 0 | 0 | Factual
hypoxemia | 0 | 0 | Factual
invasive ventilatory support | 0 | 0 | Factual
midazolam | 0 | 48 | Factual
propofol | 0 | 48 | Factual
hydrocortisone | 0 | 192 | Factual
magnesium sulfate | 0 | 192 | Factual
antibiotics | 0 | 192 | Factual
piperacillin tazobactam | 0 | 192 | Factual
clarithromycin | 0 | 192 | Factual
neuromuscular blocking agents | 48 | 96 | Factual
cisatracurium | 48 | 96 | Factual
ventilatory weaning | 96 | 96 | Factual
dual sedation | 0 | 96 | Factual
NMB | 48 | 96 | Factual
dexmedetomidine | 96 | 720 | Factual
GCS 15/15 | 144 | 144 | Factual
weakness of the neck flexor muscles | 144 | 144 | Factual
facial paresis | 144 | 144 | Factual
muscular strength 1/5 in lower limbs | 144 | 144 | Factual
muscular strength 2/5 in upper limbs | 144 | 144 | Factual
flaccid hyporeflexia | 144 | 144 | Factual
preserved sensitivity | 144 | 144 | Factual
brain MRI | 144 | 144 | Factual
cervical MRI | 144 | 144 | Factual
cerebrospinal fluid study | 144 | 144 | Factual
MRC score 37 points | 144 | 144 | Factual
electromyography | 144 | 144 | Factual
denervation | 144 | 144 | Factual
irritability | 144 | 144 | Factual
myopathic pattern | 144 | 144 | Factual
polyneuropathic compromise | 144 | 144 | Factual
axonal pattern | 144 | 144 | Factual
ICUAW diagnosis | 144 | 144 | Factual
physiotherapy | 144 | 720 | Factual
comprehensive rehabilitation | 144 | 720 | Factual
ventilator withdrawal | 240 | 240 | Factual
MRC score 55 points | 720 | 720 | Factual
normal ABG control | 720 | 720 | Factual
symptomatic resolution | 720 | 720 | Factual
hospital discharge | 720 | 720 | Factual