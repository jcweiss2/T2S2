74 years old | 0
male | 0
admitted to the hospital | 0
diarrhoea | -72
vomiting | -72
agitated | 0
Glasgow Coma Scale score of 12/15 | 0
pansystolic murmur | 0
evidence of impaired oral hygiene | 0
inflammatory markers elevated | 0
peripheral blood cultures taken | 0
intravenous ceftriaxone started | 0
blood culture grew Staphylococcus aureus | 24
SARS-CoV-2 nasopharyngeal swab negative | 0
transthoracic echocardiogram showed severe mitral regurgitation | 0
vegetations on both mitral and aortic valves | 0
definite IE confirmed | 0
Osler nodes | 0
Janeway lesion | 0
renal failure | 120
anuric | 192
haemodialysis | 192
transferred to a tertiary hospital | 240
admitted to the intensive care unit | 240
continuous venovenous haemofiltration | 240
SARS-CoV-2 nasopharyngeal swab positive | 264
nausea | 576
vomiting | 576
CT imaging of chest showed peripheral ground glass change with bilateral pleural effusions | 576
started on supplementary oxygen | 576
oral dexamethasone | 576
intravenous remdesivir | 576
died from acute respiratory distress syndrome | 744
COVID-19 pneumonia | 744