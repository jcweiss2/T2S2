47 years old | 0
male | 0
visited emergency room | 0
decreased mentality | 0
diabetes mellitus | 0
blood pressure 60/30 mm Hg | 0
body temperature 38.5℃ | 0
white blood cell 13.150×10^9/L | 0
neutrophils 90.7% | 0
lymphocytes 8.5% | 0
hemoglobin 14.3 g/dL | 0
platelet count 507×10^9/L | 0
glucose 443 mg/dL | 0
blood urea nitrogen 52.5 mg/dL | 0
serum creatinine 1.9 mg/dL | 0
aspartate aminotransferase 69 IU/L | 0
alanine transaminase 38 IU/L | 0
sodium 125.7 mmol/L |%0
potassium 5.4 mmol/L | 0
C-reactive protein 19.42 mg/dL | 0
ketone bodies in blood 3 positive | 0
HbA1c 18.20% | 0
arterial blood gas pH 7.032 | 0
pCO2 21.8 mm Hg | 0
pO2 83.3 mm Hg | 0
HCO3 5.8 mmol/L | 0
chest X-ray multiple consolidation | 0
chest CT ground glass opacities | 0
diagnosed diabetic ketoacidosis | 0
severe pneumonia | 0
immediate hydration | 0
insulin therapy | 0
piperacillin and tazobactam sodium | 0
admitted to ICU | 0
mechanical ventilator therapy | 0
ketoacidosis improved | 24
diuretic-resistant pulmonary edema | 48
continuous renal replacement therapy | 48
Klebsiella pneumonia identified | 48
lung lesions regressed | 192
moved to general ward | 192
vague abdominal pain | 240
pain aggravated | 240
severe tenderness | 240
erect abdominal X-ray gaseous distention | 240
stepladder sign | 240
abdominal CT multiple perforation | 240
panperitonitis | 240
emergency laparotomy | 240
necrotic intestines observed | 240
resected specimen septated fungal hyphae | 240
acute angle branching | 240
diagnosed colonic IA | 240
intravenous liposomal amphotericin-B | 240
discharged | 720
oral voriconazole | 720
remaining abdominal discomfort | 720
mildly elevated CRP | 720
voriconazole discontinued | 2400
abdominal discomfort relieved | 2400
CRP normalized | 2400
