34 years old|0
    Chinese man|0
    admitted to the hospital|0
    recurrent fever|-36240
    rigors|-36240
    high fever|0
    chills|0
    right leg pain|0
    lung infection|0
    soft tissue infection|0
    antibiotics given|0
    dyspnea|24
    cough|24
    chest pain|24
    transferred to a hospital in Xi'an City|24
    elevated white blood cell count|0
    high neutrophil percentage|0
    increased procalcitonin level|0
    chest CT showing lung infection with encapsulated effusion|0
    abscess in right lower leg|0
    incision and drainage of abscess|0
    ceftazidime therapy|0
    Proteus vulgaris growth from drainage culture|120
    imipenem infusion|120
    sulbactam/cefoperazone infusion|120
    temperature normalized|120
    respiratory symptoms improved|120
    leg wound coalesced|120
    discontinuation of antibiotics|120
    recurrent fever|168
    cough|168
    chills|168
    hospital stay for 2 weeks|168
    blood culture revealing Morganella morganii|336
    resistant to imipenem|336
    sensitive to cefoperazone/sulbactam|336
    sulperazone infusion|336
    discharged from hospital|336
    discontinuation of antibiotic infusion|336
    fever with chills|336
    cough recurred|336
    antibiotic therapy for 3 months|336
    recurrent high fever|336
    chills|336
    pneumonia persisted|336
    transferred to our hospital|0
    higher fever|0
    chills|0
    chest pain|0
    cough|0
    fatigue|0
    no history of cardiac disease|0
    no invasive procedures|0
    not an intravenous drug abuser|0
    never drank alcohol excessively|0
    HIV negative|0
    no central venous catheterization|0
    tachycardia (110 beats/min)|0
    blood pressure 108/70 mmHg|0
    temperature 40.2°C|0
    respiratory rate 24 breaths/min|0
    oxygen saturation 96%|0
    grade II systolic murmur|0
    no subcutaneous hemorrhagic spot|0
    no undernail linear hemorrhage|0
    no Roth spots|0
    normal leukocyte count|0
    elevated neutrophil percentage|0
    elevated CRP|0
    elevated ESR|0
    normal kidney function|0
    normal liver function|0
    normal procalcitonin level|0
    normal electrolytes|0
    normal NT-proBNP|0
    HIV negative|0
    autoantibodies negative|0
    normal B lymphocyte count|0
    normal immunoglobulin levels|0
    normal lymphocyte subpopulations|0
    CT scan showing bilateral pulmonary inflammatory shadows|0
    ECG showing sinus tachycardia|0
    blood culture revealing Morganella morganii|120
    resistant to piperacillin|120
    resistant to tazobactam|120
    resistant to imipenem|120
    sensitive to cefoperazone/sulbactam|120
    next generation sequencing confirming M. morganii DNA|120
    TTE showing tricuspid vegetation|0
    tricuspid regurgitation|0
    diagnosis of infective endocarditis|0
    cefoperazone/sulbactam therapy|0
    amikacin therapy|0
    episodes of fever with chills during treatment|168
    surgical indications|168
    open-heart surgery performed|504
    vegetation curetted|504
    tricuspid valvuloplasty|504
    bacterial culture of vegetation confirming M. morganii|504
    recovered quickly post-operation|504
    pneumonia resolved|504
    fever resolved|504
    TTE follow-up showing normal heart function|672
    tricuspid valve closure and opening normally|672
    small regurgitation|672
    thoracic CT scan showing cured pulmonary infections|480
    no relapse of infections|480

