63 years old | 0
    female | 0
    hypertension | -1752
    hyperlipidemia | -1752
    type II diabetes mellitus | -1752
    HbA1c 6.5% | -1752
    presented with right neck pain | -168
    presented with subjective fevers | -168
    emergency department presentation | -168
    rapid strep test | -168
    CT head | -168
    CT neck | -168
    CT temporal bones | -168
    discharged with amoxicillin-clavulanic acid | -168
    recurrent fevers | -168
    Tmax 101 °F | -168
    pulsatile right sided temporal headache | -168
    new onset odynophagia | -168
    denied difficulty breathing | -168
    denied stridor | -168
    denied changes in her voice | -168
    denied neck stiffness | -168
    denied photophobia | -168
    denied phonophobia | -168
    denied focal neurologic deficits | -168
    denied night sweats | -168
    denied weight loss | -168
    no preceding catheters | -168
    no trauma | -168
    no lesions to the neck | -168
    no previous upper respiratory tract infection | -168
    no recent dental infection | -168
    no dental procedure | -168
    no mouth sores | -168
    traveled to the Philippines | -1344
    denied sick contacts | -1344
    denied animal exposures | -1344
    denied outdoor activities | -1344
    worked as a registered nurse | -1344
    denied alcohol use | -1344
    denied cigarette smoking | -1344
    denied illicit drug use | -1344
    febrile to 39 °C | 0
    hypotensive | 0
    no signs of respiratory distress | 0
    tenderness of the right sternocleidomastoid border | 0
    induration of the right sternocleidomastoid border | 0
    firm nodule anterior to the right sternocleidomastoid | 0
    bulging of the right lateral pharyngeal wall | 0
    neutrophil-predominant leukocytosis 14.1 × 103/μL | 0
    blood cultures grew Gram-negative bacilli | 0
    CT neck with IV contrast | 0
    CT neck without IV contrast | 0
    occluded right internal jugular vein | 0
    thrombus extended into retromandibular vein | 0
    extensive fluid in the retropharyngeal space | 0
    inflammatory stranding | 0
    suppurative lymphadenopathy | 0
    ultrasound of the right neck | 0
    no color Doppler flow in right internal jugular vein | 0
    cystic structures | 0
    decision not to decompress | 0
    CT head negative for intracranial metastases | 0
    initial hypotension | 0
    fluid resuscitation | 0
    diagnosed with Lemierre’s syndrome | 0
    treatment with piperacillin-tazobactam | 0
    Gram-negative bacillus identified as Klebsiella pneumoniae | 24
    changed to meropenem | 24
    treated with rivaroxaban | 0
    persistent fevers | 24
    increased swelling to the midline | 24
    increased work of breathing | 24
    repeat CT neck | 24
    CT chest revealed subpleural nodules | 24
    improved clinically | 72
    transitioned to ampicillin-sulbactam | 72
    discharged | 168
    completed 6-week amoxicillin-clavulanic acid | 168
    completed 3-month rivaroxaban | 168
    returned to productive life | 240
    no sequelae | 240
    positive string test | 168
    whole genome sequencing | 168
    comparative genomic analysis | 168
    virulence factors identified | 168
    antimicrobial resistance genes identified | 168
    DNA extraction | 168
    PacBio sequencing | 168
    phylogenetic analysis | 168
    species verification analysis | 168
    MLST analysis | 168
    virulence factors iroB and iucA | 168
    antibiotic resistance genes | 168
<|eot_id|>
