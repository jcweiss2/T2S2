40 years old | 0
female | 0
extraction of upper right back tooth | -264
swelling on right side of face | 0
pain | 0
unhealed socket in right maxillary posterior region | -264
decreased mouth opening | 0
referred to medical school | -264
toxic general condition | 0
GCS score 11 | 0
temperature 40℃ | 0
tender swelling | 0
fluctuant swelling | 0
swelling extended from temporal region to inferior border of mandible | 0
swelling extended from angle of mouth to angle of mandible | 0
necrosis over right infraorbital region | 0
diplopia | 0
dilated pupil | 0
proptosis | 0
periorbital ecchymosis | 0
loss of vision | 0
abducens nerve palsy | 0
chemosis of right eye | 0
fractured maxillary tuberosity | 0
necrosis of palatal mucosa | 0
necrosis of upper right vestibule | 0
random blood sugar 311 mg/dL | 0
total leucocyte count 18,200 cubic millimeter | 0
polymorph value 92% | 0
CT scan mucosal thickening bilateral maxillary sinuses | 0
CT scan mucosal thickening right ethmoidal sinuses | 0
CT scan venous dilatation right superior ophthalmic vein | 0
CT scan suggestive of thrombosis | 0
CT scan abscess right buccal space | 0
CT scan abscess right temporal space | 0
intravenous imipenem | 0
intravenous clindamycin | 0
intravenous ceftriaxone | 0
intravenous chloramphenicol | 0
intravenous metronidazole | 0
intravenous furosemide | 0
intravenous mannitol | 0
intravenous dexamethasone | 0
nonsteroidal anti-inflammatory drugs | 0
paracetamol | 0
subcutaneous insulin | 0
subcutaneous low molecular weight heparin | 0
diagnosis of cavernous sinus thrombosis | 0
incision and drainage of right buccal and temporal spaces | 48
admission to intensive care unit | 48
chemosis in left eye | 72
paralysis of contralateral side of body | 72
GCS score 7 | 72
ventilator | 72
meningitis | 96
septic emboli | 96
blindness | 96
cranial nerve palsies | 96
sepsis | 96
shock | 96
death | 96
