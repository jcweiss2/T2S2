toothache | -96
dyspnea | -96
chest pain | -96
sweating | -96
tachyarrhythmia | -96
sore throat | -96
fever | -96
gross swelling of the lower right cheek | -96
gross swelling of the submandibular and mental regions | -96
erythematous and warm on palpation | -96
difficulties in opening the jaw | -96
inflammatory changes of the mucous membrane of the oral cavity | -96
treated with ceftriaxone-steroids-based 3 g once daily | -96
ineffective treatment | -48
worsening of the condition | -48
dyspnea | -48
chest pain | -48
admission to the Emergency Service | 0
increase in the amount of white blood cells | 0
increase in the amount of neutrophils | 0
increase in the level of C-reactive protein | 0
orotracheal intubation | 0
left pleural effusion | 0
mediastinitis | 0
right parapharyngeal abscess | 0
drainage of the right neck | 0
left chest drain | 0
intravenous antibiotic therapy with piperacillin sodium plus tazobactam sodium | 0
worsening of the clinical condition | 48
transfer to an Intensive Care Unit | 48
air collection in the right submandibular | 48
air collection in the left carotid | 48
air collection in the retroesophageal and pretracheal spaces | 48
collections characterized by air and fluids in the upper, anterior, and posterior mediastinum | 48
bilateral pleural effusions | 48
additive pleural drain on the right side | 72
abscesses in the cervical spaces | 72
extensive mediastinal empyema | 72
left pleural effusion | 72
right hydropneumothorax | 72
aggressive mediastinal debridement | 72
VATS | 72
incision and drainage of the neck abscesses | 72
oral tooth extraction | 72
purulent fluid in the cavity below was drained and packed | 72
growth of Streptococcus anginosus | 72
growth of Gemella morbillorum | 72
growth of Staphylococcus lugdunensis | 72
antibiotic therapy with amoxicillin | 72
antibiotic therapy with metronidazole | 72
dismissed in better health conditions | 168