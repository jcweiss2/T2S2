14 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
near-drowning incident | -1 | -1 | Factual
cardiopulmonary resuscitation (CPR) | -1 | -1 | Factual
abdominal pain | 0 | 0 | Factual
diffuse abrasions on torso | 0 | 0 | Factual
pneumoperitoneum | 0 | 0 | Factual
pneumomediastinum | 0 | 0 | Factual
intraabdominal free fluid | 0 | 0 | Factual
hollow viscus perforation | 0 | 0 | Possible
laparotomy | 0 | 0 | Factual
gastroesophageal junction (GEJ) disruption | 0 | 0 | Factual
damage control procedure | 0 | 0 | Factual
distal esophagus stapled closed | 0 | 0 | Factual
proximal stomach stapled closed | 0 | 0 | Factual
mediastinal drain placed | 0 | 0 | Factual
gastrostomy (G) tube placed | 0 | 0 | Factual
nasogastric (NG) tube placed | 0 | 0 | Factual
septic shock | 0 | 24 | Factual
respiratory failure | 0 | 24 | Factual
prolonged intubation | 0 | 432 | Factual
deep venous thrombosis | 0 | 24 | Factual
pulmonary embolism | 0 | 24 | Factual
bilateral pleural effusions | 0 | 24 | Factual
general deconditioning | 0 | 1200 | Factual
parenteral nutrition started | 0 | 0 | Factual
extubated | 432 | 432 | Factual
leak in esophagus | 432 | 432 | Factual
enteral nutrition initiated via G tube | 432 | 432 | Factual
discharged | 1200 | 1200 | Factual
Ivor-Lewis distal esophagectomy | 2160 | 2160 | Factual
gastric pull-up for esophagogastric anastomosis | 2160 | 2160 | Factual
jejunostomy tube placed | 2160 | 2160 | Factual
extubated | 2163 | 2163 | Factual
esophagram showed no leak | 2167 | 2167 | Factual
initiated on liquid diet | 2167 | 2167 | Factual
discharged | 2170 | 2170 | Factual
tolerate regular diet | 2600 | 2600 | Factual
gaining weight and recovering well | 2600 | 2600 | Factual