73 years old | 0
male | 0
presented to the hospital | 0
meteorism | -120
diarrhea | -120
vomiting | -120
fever (T=38.3°C) | -120
low blood pressure (BP=90/50 mm Hg) | -120
ischemic stroke | 0
untreated type II diabetes | 0
enlarged abdomen | 0
slightly painful with palpation in the right iliac fossa | 0
paraumbilical hydroaerial levels | 0
white blood cell count (WBC)=13.1×10^9/L | 0
hemoglobin=116 g/L | 0
glucose=10 mmol/L | 0
creatinine=0.37 mmol/L | 0
urea=28.3 mmol/L | 0
creatine phosphokinase=269 U/L | 0
potassium=5.3 mmol/L | 0
sodium=150 mmol/L | 0
chloride=114.7 mmol/L | 0
bicarbonate=10 mmol/L | 0
procalcitonin (PCT) value >32 µg/L | 0
CRP value=1228.5 nmol/L | 0
septic shock of intra-abdominal origin | 0
empirical intravenous antibiotic therapy with third-generation cephalosporins | 0
emergency surgery | 0
general anesthesia with orotracheal intubation | 0
exploratory laparotomy | 0
agglutinated intestinal loops in the right iliac fossa | 0
false membranes | 0
purulent-appearing fluid | 0
acute gangrenous appendicitis with perforation | 0
suppurative omentitis | 0
overdistended jejunum and ileum with occlusive appearance | 0
appendectomy | 0
segmental omentectomy | 0
lavage and drainage of the peritoneal cavity | 0
neglected peritonitis in the occlusive phase | 0
acute fibrinopurulent peritonitis | 0
acute granulocytic inflammatory infiltrate in the greater omentum | 0
bacterial culture and sensitivity of the peritoneal fluid | 0
Escherichia coli | 0
hospitalized in the intensive care unit | 0
acute pancreatitis | 0
paroxysmal atrial fibrillation (heart rate: 168–190 bpm) | 0
low blood pressure (80/40 mm Hg) | 0
complex drug treatment | 0
antibiotics | 0
anticoagulants | 0
analgesics | 0
corticosteroids | 0
vasopressors | 0
fluid volume replacement | 0
electrolyte and acid-base rebalancing | 0
discharged | 456
good general health at 3-month check-up | 0
resumption of activities of daily living | 0
