recurrent fever | -720
nausea | -168
vomiting | -168
admitted to hospital | 0
neutrophil count 6.96×10^9/L ↑ | 0
monocyte count 0.86×10^9/L ↑ | 0
lymphocyte percentage 14.9% ↓ | 0
red blood cell count 3.17×10^12/L ↓ | 0
hemoglobin content 87 g/L ↓ | 0
hematocrit 0.28 L/L ↓ | 0
average red blood cell hemoglobin concentration 312 g/L ↓ | 0
platelet count 363×10^9/L ↑ | 0
platelet distribution width 8.3 fl ↓ | 0
C-reactive protein (CRP) 52.01 mg/L ↑ | 0
diagnosed with secondary infectious thrombocytopenia | 0
diagnosed with gram-negative bacilli septicemia (Klebsiella pneumoniae) | 0
diagnosed with liver abscess | 0
diagnosed with bilateral lung inflammation | 0
diagnosed with type 2 diabetes | 0
diagnosed with hypertension grade 3 | 0
given vancomycin | 0
given caspofungin | 0
given dexamethasone | 0
given posaconazole oral suspension | 0
liver abscess puncture and drainage treatment | 24
inflammatory indexes decreased | 48
light perception disappeared in the left eye | 72
eyelid redness and pain | 72
purulent secretion | 72
repeated fever | 72
left-sided headache | 72
diagnosed with endogenous endophthalmitis (left) | 72
diagnosed with orbital cellulitis (left) | 72
diagnosed with rubeosis iridis (left) | 72
diagnosed with exudative retinal detachment (left) | 72
diagnosed with diabetic retinopathy (right) | 72
intravitreal injection with vancomycin and ceftazidime | 96
symptoms relieved | 120
left eyeball enucleation | 168
fever again after the operation | 168
given moxifloxacin | 168
given sulperazon | 168
temperature elevated again | 192
CT examination | 192
inflammation of both lungs | 192
pericardial effusion | 192
bilateral pleural thickening and effusion | 192
atelectasis in right inferior lobe | 192
liver cyst | 192
liver abscess | 192
right renal cyst | 192
myoma of the uterus | 192
history of hypertension | -8760
convulsion with unconsciousness | 240
transferred to the respiratory intensive care unit | 240
emergency CT examination | 240
lacunar infarction | 240
encephalomalacia | 240
bilateral pleural effusion | 240
lower lobe of the right lung insufficiently inflated | 240
in a coma | 240
unresponsive | 240
slight neck resistance | 240
weak light response of the eye | 240
uncooperative physical examination of limb muscle strength | 240
low muscle tension | 240
suspicious left Babinski sign (+) | 240
right Babinski sign (−) | 240
impression of intracranial infection | 240
lumbar puncture | 240
cerebrospinal fluid (CSF) sent for biochemistry analysis and microbial metagenomic next-generation sequencing (mNGS) | 240
biochemistry analysis | 246
glucose <1.1 mmol/L ↓ | 246
chlorine 108 mmol/L ↓ | 246
CSF protein >3,000 mg/L ↑ | 246
microbial mNGS results | 246
high sequence of Klebsiella pneumoniae with drug-resistant gene SHV-type beta-lactamases (blaSHV) | 246
administered 2 g meropenem every 8 hours (q8h) prolonged for 3 h | 246
body temperature improved | 264
blood routine improved | 264
CRP improved | 264
CT examination | 408
pulmonary edema and pleural effusion gradually dissipated and absorbed | 408
CSF analyses | 432
chlorine 119 mmol/L ↓ | 432
micro amount of proteins 1,107 mg/L ↑ | 432
microalbumin 816.3 mg/L ↑ | 432
immunoglobulin G 308.5 mg/L ↑ | 432
α2-macroglobulin 18.5 mg/L ↑ | 432
β2-microglobulin 2.67 mg/L ↑ | 432
discharged from the hospital | 504