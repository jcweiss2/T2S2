11 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
fever | -72 | 0 | Factual
vomiting | -72 | 0 | Factual
generalized abdominal pain | -72 | 0 | Factual
no unusual history of drug allergies | 0 | 0 | Factual
no medical history | 0 | 0 | Factual
no surgical procedures | 0 | 0 | Factual
family lives in Rahovec | 0 | 0 | Factual
grandfather diagnosed with COVID-19 | -720 | -720 | Factual
rash on palms and trunk | 0 | 0 | Factual
no conjunctivitis | 0 | 0 | Negated
no lymphadenopathy | 0 | 0 | Negated
severe drowsiness | 0 | 0 | Factual
meningeal signs negative | 0 | 0 | Negated
respiratory rate 25/min | 0 | 0 | Factual
oxygen saturation 93% | 0 | 0 | Factual
harsh breathing with crackles | 0 | 0 | Factual
tachycardic | 0 | 0 | Factual
hypotension | 0 | 0 | Factual
abdomen tender to palpation | 0 | 0 | Factual
white blood cell count 13.5 × 10^3/μL | 0 | 0 | Factual
red blood cell count 3.5–5.8 × 10^6/mm^3 | 0 | 0 | Factual
erythrocyte sedimentation rate increased | 0 | 0 | Factual
C-reactive protein increased | 0 | 0 | Factual
procalcitonin increased | 0 | 0 | Factual
SARS-CoV-2 test negative | 0 | 0 | Factual
abdominal ultrasound showed enlarged appendix | 0 | 0 | Factual
emergency laparotomy appendectomy | 0 | 24 | Factual
postoperative course toxic | 24 | 48 | Factual
tachycardia | 24 | 48 | Factual
hypotension | 24 | 48 | Factual
fractional shortening | 24 | 48 | Factual
oxygen therapy | 24 | 48 | Factual
bronchopneumonia | 24 | 48 | Factual
treatment with ceftriaxone and amikacin | 24 | 48 | Factual
switched to imipenem | 48 | 72 | Factual
positive history of contact with COVID-19 | 0 | 0 | Factual
serologic test positive for SARS-CoV-2 | 48 | 48 | Factual
ferritin elevated | 48 | 48 | Factual
IL6 elevated | 48 | 48 | Factual
high-sensitivity troponin elevated | 48 | 48 | Factual
D-dimer elevated | 48 | 48 | Factual
enoxaparin initiated | 48 | 72 | Factual
IV immunoglobulin administered | 48 | 72 | Factual
aspirin administered | 48 | 120 | Factual
general condition worsened | 72 | 72 | Factual
febrile | 72 | 96 | Factual
anemic | 72 | 96 | Factual
toxic | 72 | 96 | Factual
red blood cell transfusion | 72 | 72 | Factual
pulse dosage of systemic corticosteroids | 96 | 96 | Factual
re-evaluation of emerging shock | 96 | 96 | Factual
aggravation of heart dysfunction | 96 | 96 | Factual
echocardiogram showed decreased LV function | 96 | 96 | Factual
septal hypokinesia | 96 | 96 | Factual
ejection fraction 30% | 96 | 96 | Factual
dobutamine added | 96 | 120 | Factual
vasoactive drugs discontinued | 120 | 120 | Factual
afebrile | 120 | 120 | Factual
clinical symptoms improved | 120 | 120 | Factual
arterial pressure stable | 120 | 120 | Factual
no pathogenic agents detected | 120 | 120 | Factual
histopathological examination showed catarrhal appendicitis | 120 | 120 | Factual
D-dimer showed downward trend | 120 | 120 | Factual
troponemia resolved | 120 | 120 | Factual
inflammatory parameters normal | 120 | 120 | Factual
LV function improved | 120 | 120 | Factual
no aneurysms observed | 120 | 120 | Factual
discharged | 288 | 288 | Factual
follow-up outpatient visit | 336 | 336 | Factual
blood tests normalized | 336 | 336 | Factual
COV-2 IgG elevated | 336 | 336 | Factual
abdominal and cardiac ultrasounds normal | 336 | 336 | Factual
follow-up outpatient visits planned | 336 | 336 | Factual