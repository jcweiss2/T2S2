57 years old | 0
male | 0
Caucasian | 0
admitted to the hospital | 0
hypertension | -672
hepatitis C | -672
Crohn’s disease | -672
Prinzmetal angina | -672
recurrent chest pain | -168
single episode of fever | -168
general malaise | -168
diarrhea | -168
infliximab therapy | -336
azathioprine | -336
alcohol abuse | -672
tobacco abuse | -672
cocaine abuse | -10080
poultry farming | -672
exposure to animals | -672
substernal chest pain | -504
coronary angiography | -504
Prinzmetal angina diagnosis | -504
no need for coronary angioplasty | -504
recurred substernal chest pain | -24
presentation to rural hospital | -24
CT scan of the chest | -24
large pericardial effusion | -24
transfer to facility | -24
blood pressure 90/60 mmHg | 0
temperature 36.8 °C | 0
tachycardia | 0
respiratory rate 26 breaths per minute | 0
dehydration | 0
leukocytosis with left shift | 0
negative troponin level | 0
transthoracic echocardiogram | 0
cardiac tamponade physiology | 0
cardiothoracic consultation | 0
pericardial window | 0
drainage of 500 mL purulent fluid | 0
pericardial fluid grew nontyphoid Salmonella enterica | 0
stool specimen grew nontyphoid Salmonella enterica | 0
no growth on blood cultures | 0
vancomycin | 0
piperacillin/tazobactam | 0
ceftriaxone | 0
intensive care unit | 0
ten days of care | 240
transfer to general medical ward | 240
recurrence of fevers | 240
fevers up to 40 °C | 240
no hemodynamic instability | 240
comprehensive investigation for other causes of fever | 240
no change in therapy | 240
fever resolved | 480
last dose of infliximab | -336
completion of four weeks of ceftriaxone | 672
asymptomatic at eight-week follow-up | 1008