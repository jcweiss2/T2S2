44 years old | 0
female | 0
arterial hypertension | -672
dyslipidemia | -672
obesity | -672
aspirin | -672
losartan | -672
atorvastatin | -672
erythematous rash | -48
rash on thighs | -48
rash on armpits | -48
rash on inframammary fold | -48
rash progression to whole body | -24
application of dexamethasone | -24
use of tampons | -48
admitted to the hospital | 0
hypotensive | 0
low blood pressure | 0
high heart rate | 0
febrile | 0
somnolent | 0
morbilliform rash | 0
pustular lesions | 0
septic shock | 0
toxic shock syndrome | 0
DRESS | 0
AGEP | 0
broad spectrum antibiotics | 0
vancomycin | 0
piperacillin/tazobactam | 0
clindamycin | 0
vasopressor drugs | 0
norepinephrine | 0
vasopressin | 0
leukocytosis | 0
neutrophilia | 0
acute kidney failure | 0
elevated serum creatinine | 0
elevated blood urea nitrogen | 0
low estimated glomerular filtration rate | 0
elevated total bilirubin | 0
elevated serum transaminases | 0
metabolic acidosis | 0
hyperlactatemia | 0
parahiliar bilateral reticular infiltrates | 0
SARS-CoV-2 infection | 0
nasopharyngeal swab RT-PCR | 0
discontinuation of vancomycin | 24
daptomycin | 24
elevated creatine phosphokinase | 24
rhabdomyolysis | 24
skin biopsy | 24
diffuse spongiosis | 24
intradermic subcorneal micro pustules | 24
neutrophilic content | 24
reactive changes of microvascular endothelium | 24
fludrocortisone | 48
hydrocortisone | 48
meropenem | 48
local management of skin lesions | 48
hyperoxygenated fatty acids | 48
progressive improvement | 72
no longer required vasopressor agents | 120
extubated | 120
complete recovery of kidney function | 168
complete recovery of liver function | 168
lung images without COVID-19 pneumonia | 168
critical polyneuropathy | 168
proximal limb weakness | 168
physical rehabilitation | 168
discharged | 336