70 years old | 0
female | 0
presented to the emergency department | 0
constipation | -240
abdominal pain | -240
vomiting | -240
dehydration | 0
fever | 0
temperature of 37.8 centigrade | 0
pulse of 130/minute | 0
blood pressure of 100/70 mm Hg | 0
respiratory rate of 26/min | 0
BMI of 16 kg/m² | 0
history of asthma | 0
steroid inhalers | 0
bilateral rhonchi | 0
tense abdomen | 0
tender abdomen | 0
generalized guarding | 0
hyperdynamic bowel sounds | 0
inconclusive digital rectal examination | 0
white cell count of 16×10⁹/L | 0
erect abdomen x-ray with multiple scattered air fluid levels | 0
ultrasonography showing dilated small bowel loops | 0
normal peristaltic activity | 0
deteriorating condition | 0
acute peritonitis | 0
urgent laparotomy | 0
provisional diagnosis to surgery interval of 3 hours | 0
resuscitation | 0
blood pressure optimization | 0
electrolyte abnormalities optimization | 0
exploratory laparotomy | 0
strangulated obturator hernia | 0
ileum loop in hernia sac | 0
Meckel diverticulum in hernia sac | 0
perforation at base of Meckel diverticulum | 0
300 mL feculent matter removed | 0
dusky ileum | 0
ischemic ileum | 0
ileum resection | 0
hernia defect repair | 0
non-absorbable purse string sutures | 0
loop ileostomy creation | 0
abdomen cleansing with 6 liters saline | 0
retention sutures applied | 0
abdomen closure | 0
skin defect left open | 0
transfer to ICU | 0
ventilator support | 0
expired after 3 days in ICU | 72
multiple organ dysfunction | 72
overwhelming sepsis | 72
BMI of 16 kg/m² |6
