26 years old | 0
male | 0
abdominal pain | -24
night sweats | -24
fever | -24
intra-abdominal mass | -24
low-grade sarcoma | -24
mixed epithelioid and spindle cell morphology | -24
mucin 4-positive tumour | -24
EWSR1 gene rearrangement | -24
doxorubicin-ifosfamide chemotherapy | 0
stable disease | 24
disease progression | 96
cytoreductive surgery | 96
hyperthermic intraperitoneal chemotherapy | 96
cisplatin | 96
doxorubicin | 96
intravenous ifosfamide | 96
remission | 192
recurrence | 312
CRS | 312
HIPEC | 312
gemcitabine | 504
docetaxel | 504
disease progression | 504
symptomatic treatment | 504
COVID-19 | 624
enterocutaneous fistulas | 624
nil-by-mouth status | 624
parenteral nutrition | 624
sepsis | 624
intra-abdominal collections | 624
nivolumab | 624
no clinical response | 624
molecular tumour board | 720
next-generation sequencing | 720
ALK mutation | 720
crizotinib | 744
disease progression | 744
tumour size regression | 760
haematological toxicity | 776
fatigue | 776
reduced dose of crizotinib | 776
tumour response | 776
enterocutaneous fistulas improvement | 776