70 years old | 0
African-American | 0
male | 0
admitted to the hospital | 0
fever | 0
headaches | 0
chills | 0
nausea | 0
ESRD | -8760
non-insulin-dependent diabetes mellitus | -8760
hypertension | -8760
severe peripheral arterial disease | -8760
recurrent vascular access thrombosis | -8760
symptomatic bradyarrhythmia | -8760
AICD | -8760
aspirin | 0
calcium acetate | 0
carvedilol | 0
cinacalcet | 0
insulin | 0
warfarin | 0
gabapentin | 0
simvastatin | 0
esomeprazole | 0
temperature of 105 Fahrenheit | 0
blood pressure of 108/51 mm Hg | 0
heart rate of 114 beats per minute | 0
respiratory rate of 14 per minute | 0
oxygen saturation of 99% | 0
alert | 0
cooperative | 0
oriented | 0
no rash | 0
no finger clubbing | 0
lungs clear to auscultation | 0
no erythema | 0
no tenderness | 0
no fluctuation over the AICD site | 0
regular heart sounds | 0
no gallop rhythm | 0
audible grade 2/6 late diastolic murmur | 0
sodium of 135 mmol/L | 0
potassium of 4.8 mmol/L | 0
chloride of 96 mmol/L | 0
bicarbonate of 23 mmol/L | 0
blood urea nitrogen of 68 mg/dL | 0
creatinine of 11.12 mg/dL | 0
lactic acid of 1.7 mmol/L | 0
international normalized ratio 2.57 | 0
white blood cells of 10.8 k/mm3 | 0
hemoglobin 8.6 gm/dL | 0
hematocrit 25.5% | 0
platelets’ count of 79 k/mm3 | 0
empiric broad-spectrum antibiotics | 0
cefepime | 0
vancomycin | 0
CT scan of the head | 24
chest x-ray | 24
CSF examination | 24
blood cultures | 24
MRSA | 48
cuffed catheter tip culture | 48
negative | 48
transthoracic echocardiogram | 48
tricuspid valve mass | 48
trans-esophageal echocardiography | 72
tricuspid valve infectious endocarditis | 72
AICD pocket infection | 72
ampicillin | 72
vancomycin | 72
cefepime | 72
AICD removal | 96
tunneled catheter exchange | 96
new catheter | 96
fever persisted | 120
blood cultures positive for MRSA | 120
cuffed catheter exchange | 144
temporary non-cuffed catheter | 144
delirium | 168
deterioration of hemodynamic status | 168
intravenous fluids | 168
vasopressors’ support | 168
right femoral catheter removal | 192
peritoneal catheter insertion | 192
PD | 192
gradual escalation of PD exchanges | 216
improvement in clinical status | 240
resolution of fever | 240
intravenous daptomycin | 240
discharged to a long-term nursing facility | 432
long-term chronic manual ambulatory PD | 432