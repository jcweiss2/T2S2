60 years old | 0
female | 0
impaired consciousness | 0
atrial fibrillation | -672
dilated cardiomyopathy | -672
oral warfarin | -672
biventricular pacing implantable cardioverter defibrillator | -672
found lying at home | -1
transported to hospital | -1
JCS score II-10 | 0
GCS score 14 | 0
no clear neurological deficits | 0
hemorrhage in the third and fourth ventricles | 0
hemorrhage in bilateral lateral ventricles | 0
left dominance | 0
spot enhancement on the lateral wall of the anterior horn of the left lateral ventricle | 0
blood pressure control | 0
ventricular drainage not performed | 0
aneurysm at the distal site of the mLSA | 72
embolization | 72
endovascular treatment | 72
NBCA injection | 72
no signs of hemorrhagic complications | 72
no cerebral infarction | 72
sepsis triggered by pneumonia | 168
decrease in muscle strength | 168
disuse | 168
discharged | 432
modified Rankin Scale 1 | 432