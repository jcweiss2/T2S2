28 years old | 0
male | 0
thermal burn due to improper handling of a gasoline can | 0
superficial burns | 0
deep partial-thickness burns (grade IIA) | 0
deep partial-thickness burns (grade IIB) | 0
full-thickness burns (grade III) | 0
total body surface area lesions (approximately 80%) | 0
chest debridement | 0
abdominal debridement | 0
decompression incisions | 0
protective tracheal intubation | 0
suspicion of airway burns | 0
increased C-reactive protein (312.38 mg/L) | 0
moderately elevated procalcitonin (1.9 ng/ml) | 0
severe hypoproteinemia | 0
total protein (29.1 g/L) | 0
albumin (18 g/L) | 0
ABSI score (12 points) | 0
Baux score (108 points) | 0
R-Baux score (85 points) | 0
transferred to Clinical Hospital of Plastic, Reparatory, and Burn Surgery | 48
local conservative nonsurgical treatment for superficial burns | 48
lavage | 48
dressing with silver-containing products | 48
admission to Intensive Care Unit | 48
respiratory support using mechanical ventilation | 48
signs of aggressive burn-induced inflammatory reaction | 48
CRP (679 mg/L) | 48
albumin (25 g/L) | 48
presepsin (642 ng/L) | 48
serum iron (15 µg/dL) | 48
stabilized respiratory function | 48
no signs of inhalation injury | 48
oxygenation index | 48
ventilator parameters | 48
chest X-ray image | 48
extubation | 72
standard procedure for large mixed-type second-degree burns | 48
conservative local treatment methods | 48
removing devitalized tissue | 48
application of special topical antimicrobial agents | 48
superficial burns treated conservatively | 48
deep partial-thickness burns treated conservatively | 48
full-thickness burns excised and grafted | 48
expanded meshed autografts | 48
burn-protocol treatment | 0
proton-pump inhibitor (pantoprazole 40 mg) | 0
thromboprophylaxis with enoxaparin (40 mg per day) | 0
analgesics (paracetamol 4 g/day) | 0
morphine on request | 0
antioxidants (acetylcysteine) | 0
oligoelements | 0
enteral nutrition | 0
parenteral nutrition | 0
normal feeding | 0
Toronto formula estimation for caloric intake | 0
crystalloid solutions | 0
maintaining MAP >65 mmHg | 0
diuresis >0.5 ml/bw/h | 0
lactate <2 mmol/L | 0
ScVO2 >70% | 0
colonization of the wound with Pseudomonas aeruginosa | 192
increase in presepsin value to 1498 pg/ml | 192
antibiotic therapy with colistin | 192
antibiotic therapy with cefoperazone/sulbactam | 192
antibiotic therapy continued for 2 weeks | 192
swab cultures negative | 336
presepsin decreased to cut-off value for sepsis | 336
swab cultures sampled twice per week | 0
iron level tracked | 0
favorable evolution of intermediary burn injuries | 504
complete recovery | 504
transferred to burn unit | 504
stayed in burn unit for 3 weeks | 504
full-thickness burn excised and grafted | 840
expanded meshed autograft harvested from right forearm | 840
expanded meshed autograft harvested from anterior side of thigh | 840
second-degree lesions treated conservatively | 0
spontaneous epithelialization | 0
healing of second-degree lesions | 840
discharge | 1056
no vasopressor requirement | 0
no anemia | 0
no desaturation | 0
