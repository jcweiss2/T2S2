83 years old | 0
female | 0
accident involving wheelchair | 0
subcutaneous abscess on abdomen | -48
seen by family physician | -24
on way to see general surgeon | -24
flung from wheelchair | 0
fully immobilized and on backboard | 0
taken off backboard | 2
no complaints of pain other than left lower quadrant | 2
physical examination performed | 2
vital signs: blood pressure 124/59 | 2
vital signs: heart rate 107 | 2
vital signs: respiratory rate 18 | 2
vital signs: temperature 97.5°F | 2
vital signs: pulse oximetry 95% on room air | 2
lungs clear bilaterally | 2
cardiac auscultation normal | 2
abdomen bowel sounds in all 4 quadrants | 2
pain in left lower quadrant | 2
subcutaneous abscess 18 × 8-cm | 2
abscess fluctuant with central black necrotic skin | 2
oozing noted centrally | 2
Parkinson disease | 0
dementia | 0
husband became primary historian | 2
mass noticed in previous 2 days | -48
central black necrosis present since previous day | -24
increasing pain over past few days | -48
worsened pain with bowel movements | -48
history of gastroesophageal reflux | 0
history of hypertension | 0
history of hypothyroidism | 0
history of renal failure | 0
history of pulmonary hypertension | 0
history of diastolic heart failure | 0
recently hospitalized for acute diverticulitis with perforation | -168
treated medically for diverticulitis | -168
complete blood count ordered | 2
basic metabolic panel ordered | 2
urinalysis ordered | 2
abdominal computed tomography with IV contrast ordered | 2
surgical consult made | 2
white blood cell count 27.9 × 1,000/uL | 4
hemoglobin 9.4 g/dL | 4
hematocrit 27.6% | 4
platelet count 446 | 4
serum sodium 134 mmol/L | 4
potassium 3.4 mmol/L | 4
blood urea nitrogen 23 mg/dL | 4
creatinine 1.1 mg/dL | 4
urinalysis positive for nitrites | 4
microscopy showing 1+ leukocytes and 4+ bacteria | 4
CT revealed inflamed colon with fistulous tract | 4
necrotizing fasciitis diagnosed | 4
broad-spectrum antibiotics given | 6
IV fluids given | 6
presurgical laboratory tests performed | 6
admitted to intensive care unit | 6
surgical intervention performed | 12
debridement of abscess | 12
necrosis within subcutaneous fat | 12
opening at base of abscess | 12
pus from abdominal cavity | 12
sigmoid resection with placement of diverting colostomy | 12
wound vacuum placement | 12
wound site cultured | 12
Proteus mirabilis grown | 24
Escherichia coli grown | 24
E faecalis grown | 24
Bacillus fragilis grown | 24
coagulase-negative staphylococcus grown | 24
transferred to ICU on ventilatory support | 24
medical therapy for sepsis | 24
failure to wean from ventilatory support | 48
multiple bouts of fever secondary to sepsis | 48
underwent 3 other surgeries for abscess debridement | 72
transferred to long-term acute care hospital | 168