33 years old | 0
male | 0
admitted to the hospital | 0
diarrhea | -24
fever | -24
vomiting | -24
repeated belching | -6048
bloating | -6048
diarrhea for 7 years | -6048
blood tests | -6048
abdominal ultrasonography | -6048
computed tomography (CT) examinations | -6048
gastrointestinal endoscopy | -24
bowel preparation | -24
PEG | -24
gastroscopy | -24
colonoscopy | -24
hiatal hernia | -24
chronic nonatrophic gastritis | -24
erosions | -24
multiple polyps | -24
biopsy | -24
fundic gland polyps | -24
body temperature 39 °C | 0
blood pressure 114/65 mmHg | 0
heart rate 115 beats per min | 0
respiratory rate 18 breaths per min | 0
Plasma D-dimer 21800.00 μg/L | 0
brain natriuretic peptide (BNP) 7330.00 pg/mL | 0
white blood cells 35.07 × 10^9/L | 0
C-reactive protein 142.55 mg/dL | 0
procalcitonin 78.43 ng/mL | 0
lactic acid 3.3 mmol/L | 0
creatinine 391 μmol/L | 0
alanine aminotransferase 255 U/L | 0
aspartate aminotransferase 204 U/L | 0
total bile 72.3 μmol/L | 0
direct bile 41.1 μmol/L | 0
γ-glutamyltransferase 219 U/L | 0
abdominal CT examination | 0
lung CT | 0
inflammation in the lower lobe of the left lung | 0
symptomatic and supportive treatment | 0
stomach protection | 0
liver protection | 0
anti-infection | 0
levofloxacin | 0
omeprazole | 0
compound glycyrrhizin injection | 0
ademetionine 1,4-butanedisulfonate for injection | 0
elevated body temperature | 12
persistently high leukocyte index | 12
metabolic acidosis | 12
oxygenation maintained at 100% | 12
respiratory rate increased to 25 breaths per min | 12
heart rate 124 beats per min | 12
blood pressure 89/60 mmHg | 12
systemic inflammatory response | 12
septic shock | 12
acute renal insufficiency | 12
hepatic insufficiency | 12
multiple organ failure | 12
transferred to the intensive care unit (ICU) | 12
highest body temperature 40.1 °C | 24
anti-infection treatment with piperacillin sodium and tazobactam sodium | 24
body temperature dropped to 36.8 °C | 48
lactate level 1.0 | 48
white blood cell count dropped to 11.54 × 10^9/L | 48
transferred to the general ward | 48
discharged | 72
severe infection | 0
septic shock | 12
multiple organ failure | 12
follow-up | 4320