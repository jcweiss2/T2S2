72 years old | 0
male | 0
paroxysmal complete atrioventricular block | -132 
dual-chamber pacing and sensing system pacemaker implantation | -132 
box change | -36 
pacemaker box replacement | -36 
admitted to the hospital | 0
subacute endocarditis | 0
Streptococcus sanguinis bacteraemia | 0
Right atrium vegetation | 0
discovery of localized colon cancer | 0
discharged home | 24
developed acute cholangitis | 0
endoscopic retrograde cholangiopancreatography | 0
main bile duct lithiasis | 0
hilar bile duct stenosis | 0
improvement following intravenous antibiotics | 24
endoscopic stones extraction | 24
normal pacemaker function | 24
laparoscopic sigmoidectomy | 48
admitted in the intensive care unit | 96
biliary septic shock | 96
treated with vasopressors | 96
intravenous antibiotics | 96
endoscopic biliary drainage | 96
transferred to gastroenterology ward | 120
cholangitis recurrence | 120
discovery of complete ventricular lead rupture | 120
lead explantation postponed | 120
discharged home on a long-term antibiotic | 144
critically ill patient | 168
biliary sepsis recurrence | 168
decision not to replace the biliary drains | 168
antibiotic management alone | 168
lead explantation abandoned | 168
discharged home with a lifelong antibiotic | 168
patient died from biliary sepsis | 192
fever | -72
chills | -72
confusion | -72
valproic acid | -72
two strokes | -240 
cognitive impairment | -240 
right hemiparesis | -240 
blood samples demonstrated cholestasis | 0
blood cultures isolated penicillin-sensitive Streptococcus sanguinis | 0
serum alkalin phosphatase | 0
total bilirubin | 0
direct bilirubin | 0
alanine transaminase | 0
absolute neutrophil count | 0
C-reactive protein | 0
chest computed tomography | 0
multiple pulmonary embolisms | 0
transoesophageal echocardiography | 0
vegetation located on the intracardiac portion of the ventricular lead | 0
signs of biliary sepsis | 24
endoscopic retrograde cholangiopancreatography | 24
common bile duct lithiasis | 24
hilar bile duct stenosis | 24
intravenous antibiotics | 24
endoscopical stones extraction | 24
brush and forceps biopsies | 24
localized sigmoid cancer | 24
18Fluorodesoxyglucose positron emission tomography–CT | 24
sigmoidectomy | 48
endovascular lead explantation | 48
oral first-generation cephalosporin | 48
lead explantation postponed indefinitely | 120
discharged home on a long-term antibiotic | 120
critically ill patient | 168
biliary sepsis recurrence | 168
decision not to replace the biliary drains | 168
antibiotic management alone | 168
lead explantation abandoned | 168
discharged home with a lifelong antibiotic | 168
patient died from biliary sepsis | 192