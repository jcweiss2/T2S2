51 years old | 0
    indigenous woman | 0
    presented to a remote health service | 0
    back pain | 0
    radiating to the left flank | 0
    symptoms of dehydration | 0
    insulin dependent type two diabetes mellitus | 0
    medically managed ischaemic heart disease | 0
    hypertension | 0
    chronic lower back pain | 0
    treated with intra-muscular anti-inflammatories | 0
    discharged | 0
    acute exacerbation of lower back pain | 0
    represented five days later | -120
    vomiting | -120
    flank pain | -120
    confusion | -120
    transferred to a regional health service | -120
    blood pressure 76/53 mmHg | 0
    tachypnoeic at 55bpm | 0
    impaired consciousness | 0
    oliguria | 0
    non-ketotic high anion gap metabolic acidosis | 0
    pH 7.15 | 0
    lactate 10.1mmol/L | 0
    hyperglycaemia | 0
    blood glucose 23.5mmol/L | 0
    acute kidney injury | 0
    serum creatinine 348μmol/L | 0
    urinalysis demonstrated leukocytes | 0
    haemolysed blood | 0
    protein (300–500) | 0
    no nitrites | 0
    inflammatory markers elevated | 0
    white cell count 14x109 | 0
    CRP 156mg/L | 0
    hyponatraemic 126mmol/L | 0
    thrombocytopaenic 57x109 | 0
    septic shock | 0
    received broad-spectrum antibiotics | 0
    piperacillin-tazobactam | 0
    gentamicin | 0
    resuscitation | 0
    non-contrast computed tomography (CT) scan | 0
    marked oedema of the left kidney | 0
    hydronephrosis | 0
    extensive loculated and mottled areas of gas | 0
    trace perinephric gas | 0
    no fluid levels | 0
    no drainable collection | 0
    simple cyst of the superior pole | 0
    no gas internally | 0
    emphysematous pyelonephritis (EP) | 0
    admitted to the intensive care unit | 0
    vasopressor support | 0
    antibiotics | 0
    strict fluid balance | 0
    indwelling catheter | 0
    continuous veno-venous haemodialysis (CVVHD) | 0
    insulin infusion | 0
    urine culture for Klebsiella Pneumoniae | 0
    blood culture for Klebsiella Pneumoniae | 0
    antibiotic therapy narrowed | 0
    ceftriaxone | 0
    metronidazole | 0
    48-h of medical management | 48
    no clinical progression | 48
    8Fr nephrostomy tube placed | 48
    under CT guidance | 48
    further 72-h trial of non-operative management | 120
    nephrostomy drainage | 120
    organ support | 120
    cease CVVHD after 3 days | 72
    persisting confusion | 120
    high grade fevers | 120
    tachycardia | 120
    dependence on vasopressors | 120
    parenteral analgesia infusion | 120
    new anaemia Hb 82g/L | 120
    persisting inflammatory rise WCC 13.6x109 | 120
    thrombocytopaenia 114x109 | 120
    recurring deterioration in renal function Cr 142μmol/L | 120
    post CVVHD nadir Cr 71μmol/L | 72
    repeat imaging | 120
    no parenchymal improvement | 120
    high risk state | 120
    lack of drainable collections | 120
    worsening clinical status | 120
    ongoing refractory end organ dysfunction | 120
    decision for open nephrectomy | 120
    fibrous adhesions intraoperatively | 120
    subcapsular approach | 120
    post-operative recovery | 168
    intravenous antibiotics transitioned to oral after 4 days | 168
    discharged with creatinine 106μmol/L | 168
    
    