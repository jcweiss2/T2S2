40 years old | 0
male | 0
Japanese | 0
HIV-1 infection | -7776
high fever | 0
severe malaise | 0
headache | 0
generalized skin rash | 0
mild sinusitis | -720
symptomatic treatment | -720
admitted to the hospital | 0
fever | 0
shock status | 0
mildly altered consciousness | 0
neck stiffness | 0
diminished skin turgor | 0
no focal neurological deficits | 0
no visual disturbances | 0
leukocytosis | 0
elevated C-reactive protein | 0
hyperproteinemia | 0
acute renal dysfunction | 0
severe hyponatremia | 0
hyperkalemia | 0
moderate swelling of lymph nodes | 0
elevated total protein in CSF | 0
elevated IgG in CSF | 0
elevated leukocytes in CSF | 0
normal glucose level in CSF | 0
previous infection with human simplex virus 1 and 2 | -7776
previous infection with varicella-zoster virus | -7776
previous infection with hepatitis B virus | -7776
previous infection with cytomegalovirus | -7776
previous infection with Epstein–Barr virus | -7776
previous infection with syphilis | -7776
diagnosis of atypical generalized zoster | 0
high-dose acyclovir therapy | 0
rapid resolution | 24
electrolyte imbalance | 24
adrenal insufficiency | 24
comprehensive endocrinological workup | 24
panhypopituitarism | 24
head MRI scan | 48
inhomogeneous pituitary gland enlargement | 48
disappearance of T1 hyperintense signal | 48
sphenoid sinus mucosa thickening | 48
pituitary lesion with gadolinium ring enhancement | 48
high-intensity signals on diffusion-weighted imaging | 48
low-intensity signals on apparent diffusion coefficient imaging | 48
cefepime | 0
switch to ceftriaxone | 168
ceftriaxone | 168
improvement of lesions on follow-up MRI scans | 504
hydrocortisone and levothyroxine replacement | 168
plasma electrolytes normalized | 168
polyuria | 168
polydipsia | 168
desmopressin stimulation test | 168
hypotonic salt solution test | 168
diagnosis of masked diabetes insipidus | 168
desmopressin acetate | 168
no surgical drainage | 0
empirical medication improved clinical status | 0
intensive investigation regarding etiology of pituitary abscess | 0
blood and CSF cultures | 0
immunological tests for fungal infections | 0
polymerase chain reaction for mycobacteria and VZV | 0
no causative agent determined | 0
hormone replacement therapy | 0
2 years of follow-up | 17520
patient doing well | 17520