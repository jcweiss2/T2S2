50 years old | 0  
    male | 0  
    admitted to the ICU | 0  
    no spontaneous respiration | 0  
    pupils dilated and fixed at 7 mm | 0  
    no past history | 0  
    emergency decompressive craniectomy | -192  
    hematoma removal | -192  
    spontaneous intracerebral hemorrhage | -192  
    intraventricular hemorrhage | -192  
    no neurological recovery | -192  
    follow-up brain CT | -192  
    rebleeding | -192  
    second surgery | -192  
    transferred to our hospital for organ donation | -192  
    BP 75/50 mmHg | 0  
    HR 72 bpm | 0  
    SpO2 75% | 0  
    fluid administration | 0  
    continuous intravenous infusion of dopamine 15 µg/kg/min | 0  
    pressure control ventilation | 0  
    FiO2 1.0 | 0  
    PIP 26 cmH2O | 0  
    PEEP 10 cmH2O | 0  
    RR 20 breaths/min | 0  
    general edema | 0  
    large amount of pink frothy sputum | 0  
    rales bilaterally | 0  
    bilateral infiltration on chest X-ray | 0  
    concentric left ventricular hypertrophy | 0  
    preserved contractility | 0  
    no pulmonary arterial hypertension | 0  
    ABGA pH 7.310 | 0  
    PaCO2 40.5 mmHg | 0  
    PaO2 84.9 mmHg | 0  
    HCO3- 19.9 mEq/L | 0  
    BE -5.9 mEq/L | 0  
    SaO2 94.3% | 0  
    no heart failure | 0  
    no pneumonia | 0  
    no pulmonary embolism | 0  
    NPE | 0  
    hypoxemia | 0  
    SaO2 85.7% | 0  
    PaO2 66.7 mmHg | 0  
    SpO2 91-93% | 0  
    alveolar recruitment maneuvers | 0  
    CPAP 35-40 cmH2O | 0  
    BP monitoring | 0  
    RR 15-20 breaths/min | 0  
    PEEP 15 cmH2O | 0  
    SaO2 maintained at 96.3% or above | 0  
    PaO2 maintained at 93.4 mmHg or above | 0  
    endotracheal suction | 0  
    systolic pressure 90-120 mmHg | 0  
    diastolic pressure 50-80 mmHg | 0  
    HR 80-95 bpm | 0  
    central venous pressure 11-13 mmHg | 0  
    diabetes insipidus | 0  
    metabolic acidosis | 0  
    hyperglycemia | 0  
    hypernatremia | 0  
    fluid supplementation | 0  
    electrolyte correction | 0  
    sodium bicarbonate administration | 0  
    continuous intravenous insulin | 0  
    warm air blanket | 0  
    body temperature maintained at 36℃ or above | 0  
    crystalloid solution 6,280 ml | 0  
    colloid solution 80 ml | 0  
    urine output 3,840 ml | 0  
    nasogastric tube drainage 1,300 ml | 0  
    loss of brainstem reflexes | 0  
    two apnea tests | 0  
    transcranial Doppler | 0  
    electroencephalography | 0  
    brain death declared | 0  
    transferred to OR | 10.5  
    oxygen 12 L/min during transfer | 10.5  
    manual ventilation with resuscitation bag | 10.5  
    BP 120/70 mmHg | 10.5  
    HR 75 bpm | 10.5  
    SpO2 99% | 10.5  
    BP 87/55 mmHg | 10.5  
    HR 100 bpm | 10.5  
    SpO2 80% | 10.5  
    anesthesia machine connected | 10.5  
    no inhalational agent | 10.5  
    mechanical ventilation same settings as ICU | 10.5  
    SpO2 slowly rose | 10.5  
    alveolar recruitment maneuvers | 10.5  
    PEEP 15 cmH2O | 10.5  
    PIP 30 cmH2O | 10.5  
    SpO2 not above 91% | 10.5  
    ABGA pH 7.412 | 10.5  
    PaCO2 33.0 mmHg | 10.5  
    PaO2 62.3 mmHg | 10.5  
    HCO3. 20.5 mEq/L | 10.5  
    BE -3.6 mEq/L | 10.5  
    SaO2 90.8% | 10.5  
    dopamine 15 µg/kg/min | 10.5  
    epinephrine 0.05 µg/kg/min | 10.5  
    BP target achieved | 10.5  
    SpO2 did not rise further | 10.5  
    NO gas inhalation started | 10.75  
    NO infusion 20 ppm | 10.75  
    monitored NO2 concentration | 10.75  
    SpO2 rose to 99% | 10.75  
    ABGA pH 7.270 | 10.75  
    PaCO2 46.3 mmHg | 10.75  
    PaO2 328.7 mmHg | 10.75  
    HCO3. 20.8 mEq/L | 10.75  
    BE -6.0 mEq/L | 10.75  
    SaO2 99.5% | 10.75  
    hypoxemia improved | 10.75  
    NO administration continued | 10.75  
    SaO2 maintained at 98.4% or above | 10.75  
    PaO2 maintained at 132.4 mmHg or above | 10.75  
    supportive treatment continued | 10.75  
    endotracheal suctioning continued | 10.75  
    vecuronium administration | 10.75  
    crystalloid solution 2,380 ml | 10.75  
    colloid solution 500 ml | 10.75  
    red blood cells 4 units | 10.75  
    estimated blood loss 1,300 ml | 10.75  
    urine output 1,400 ml | 10.75  
    nasogastric tube drainage 340 ml | 10.75  
    cross-clamping of aorta | 13.25  
    BP suddenly decreased | 13.25  
    SpO2 suddenly decreased | 13.25  
    arrhythmia | 13.25  
    bradycardia | 13.25  
    cardiac arrest | 13.25  
    declared dead | 13.25  
    two kidneys retrieved | 13.25  
    organ transplantation successful | 13.25  
    