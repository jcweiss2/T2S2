28 years old | 0
male | 0
sickle cell trait | 0
history of previous intravenous drug use | 0
fever lasting nine days | -216
right-sided chest pain | -216
abdominal pain | -216
flank pain | -216
dysuria | -216
intermittent hematuria | -216
denied valvular heart disease | 0
denied congenital heart disease | 0
no prosthetic heart valves | 0
blood pressure 129/68 mmHg | 0
heart rate 129 beats per minute | 0
respiratory rate 19 breaths per minute | 0
temperature 39.4°C | 0
oxygen saturation 99% on room air | 0
clear chest auscultation | 0
no abnormal heart sounds | 0
severe abdominal tenderness | 0
guarding at right flank | 0
hypochondrium tenderness | 0
renal angle tenderness | 0
elevated white blood cells | 0
elevated c-reactive protein | 0
abnormal liver function tests | 0
urine dipstick analysis 3+ urobilinogen | 0
urine dipstick analysis 3+ erythrocytes | 0
diffuse bilateral nodular densities on chest radiograph | 0
poorly marginated nodules | 0
varying stages of cavitation | 0
normal sinus rhythm on electrocardiography | 0
acute abdominal pain | 0
ultrasound possible acalculous cholecystitis | 0
ill-defined mass near liver | 0
abdominal/pelvic CT with intravenous contrast | 0
CT indicated sealed bowel perforation | 0
CT indicated infection | 0
cryptogenic organizing pneumonia | 0
admitted pending repeat CT with oral contrast | 0
drowsy | 0
ill-looking | 0
tachypneic | 0
profuse sweating | 0
tachycardia | 0
hypotension | 0
IE strongly suspected | 0
pulmonary septic emboli on chest radiograph | 0
CT with oral contrast suggested pyelonephritis | 0
diagnosed with possible acute chest syndrome | 0
chest radiograph consistent with septic pulmonary emboli | 0
echocardiography confirmed tricuspid valve vegetation | 0
admitted to ICU | 0
treated with intravenous vancomycin | 0
treated with cefepime | 0
antibiotics switched to flucloxacillin | 0
blood cultures confirmed methicillin-sensitive Staphylococcus aureus | 0
blood cultures confirmed viridans group streptococci | 0
urine culture no growth | 0
CT re-evaluation showed renal infarction | 0
multiple cortical wedge-shaped areas of delayed striated contrast enhancement | 0
condition improved after 60 days | 1440
tests negative for HIV | 0
tests negative for hepatitis | 0
tests negative for thrombophilia | 0
discharged on day 61 | 1464
follow up with cardiology clinic | 1464
