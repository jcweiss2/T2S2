72 years old | 0  
    man | 0  
    dual-chamber pacing and sensing system pacemaker implantation for paroxysmal third-degree atrioventricular block | -113040  
    paroxysmal third-degree atrioventricular block | -113040  
    pacemaker box replacement due to battery end-of-life | -25920  
    battery end-of-life | -25920  
    admitted for subacute endocarditis | 0  
    Streptococcus sanguinis bacteraemia | 0  
    right atrium vegetation around one of the leads | 0  
    discovery of localized colon cancer on positron emission tomography–computed tomography (PET-CT) | 0  
    discharged home with long-term antibiotic therapy | 120  
    developed acute cholangitis | 0  
    endoscopic retrograde cholangiopancreatography showed main bile duct lithiasis | 0  
    hilar bile duct stenosis (biopsied) | 0  
    improvement following intravenous antibiotics | 0  
    endoscopic stones extraction | 0  
    normal pacemaker function in routine assessment | 240  
    laparoscopic sigmoidectomy for localized colon cancer | 408  
    admitted in the intensive care unit for biliary septic shock | -2640  
    treated with vasopressors | 0  
    intravenous (IV) antibiotics | 0  
    endoscopic biliary drainage | 0  
    transferred to gastroenterology ward once stabilized | 480  
    presented with cholangitis recurrence due to drains obstruction | 480  
    improved on IV antibiotics | 480  
    after biliary drain replacement | 480  
    discovery of complete ventricular lead rupture on chest X-ray | 960  
    PET-CT confirms persistent pacemaker leads and box infection | 960  
    lead explantation is postponed indefinitely | 960  
    discharged home on a long-term antibiotic | 960  
    critically ill patient following biliary sepsis recurrence | 1440  
    decision not to replace the biliary drains | 1440  
    antibiotic management alone | 1440  
    lead explantation is abandoned | 1440  
    discharged home with a lifelong antibiotic | 1440  
    patient died from biliary sepsis | 17520  
    chills | -2160  
    confusion | -2160  
    valproic acid for erroneously suspected epileptic seizures | -2160  
    two strokes (2000 and 2009) | -175200  
    phasic disorder | -175200  
    cognitive impairment | -175200  
    right hemiparesis | -175200  
    no past history of parenteral drug use | 0  
    hospital admission | 0  
    blood samples demonstrated cholestasis | 0  
    blood cultures isolated penicillin-sensitive Streptococcus sanguinis | 0  
    serum alkalin phosphatase reached 558 U/L | 0  
    total bilirubin was 2.3 mg/dL | 0  
    direct bilirubin at 1.6 mg/dL | 0  
    alanine transaminase 51 U/L | 0  
    absolute neutrophil count 23.840/mm3 | 0  
    C-reactive protein 89 mg/L | 0  
    chest computed tomography (CT) showed multiple pulmonary embolisms | 0  
    transoesophageal echocardiography revealed a 41 × 33 × 15 mm mobile vegetation located on the intracardiac portion of the ventricular lead | 0  
    developed signs of biliary sepsis | 0  
    endoscopic retrograde cholangiopancreatography revealed common bile duct lithiasis | 0  
    hilar bile duct stenosis | 0  
    intravenous antibiotics (Cefuroxime 1.500 mg/every 8 h (q8h) plus Metronidazole 500 mg/q8h) | 0  
    endoscopical stones extraction improved his condition | 0  
    brush and forceps biopsies were performed in search for a bile duct malignancy | 0  
    localized sigmoid cancer identified on 18Fluorodesoxyglucose (18F-FDG) positron emission tomography–CT (PET/CT) | 0  
    underwent sigmoidectomy the following month | 720  
    endovascular lead explantation was scheduled after rehabilitation | 720  
    prescribed an oral first-generation cephalosporin (cephalexin 500 mg b.i.d.) as prolonged antibiotic therapy whilst awaiting lead removal | 720  
    patient’s condition worsened | 1440  
    readmitted for recurrent cholangitis | 1440  
    repetitive antibiotic therapies | 1440  
    endoscopic biliary drainages | 1440  
    cholangiocarcinoma suspected | 1440  
    negative cytological and histological results | 1440  
    rest electrocardiogram (ECG) demonstrated sinus rhythm with normal AV delay | 1440  
    ventricular pacing spike with loss of ventricular capture | 1440  
    ventricular undersensing | 1440  
    chest X-ray revealed a complete intracardiac ventricular lead fracture | 1440  
    pacemaker interrogation reported ventricular undersensing | 1440  
    loss of capture | 1440  
    high impedance (>3000 ohms) | 1440  
    routine pacemaker assessment performed 4 months prior showed normal function | -2880  
    low rate of ventricular pacing (<1%) | -2880  
    gradual decrease in ventricular pacing impedance | -2880  
    another 18F-FDG PET/CT scan demonstrated increased uptake of 18F-FDG in both the intrathoracic and extrathoracic portions of the pacemaker | 1440  
    considering the extension of the infectious diseases | 1440  
    comorbidities of the patient (palliative approach for suspected cholangiocarcinoma, two strokes and cognitive impairment) | 1440  
    complete hardware removal was not a reasonable option | 1440  
    discharged home on lifelong antibiotic therapy (cephalexin) | 1440  
    patient became critically ill | 1440  
    transferred to a palliative care unit | 1440  
    passed away due to biliary sepsis | 17520  

    