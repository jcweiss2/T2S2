49 years old | 0
female | 0
esophageal squamous cell carcinoma | -672
neoadjuvant chemotherapy | -672
minimally invasive Ivor–Lewis esophagectomy | 0
inflammatory indexes increased | 72
CRP 178.2 ng/mL | 72
endoscopy | 96
CT scan | 96
large anastomotic leak | 96
anastomotic leak involving 75% of the anastomosis | 96
giant wound cavity in the pleural space of 8 cm in size | 96
fibrosis | 96
abundant necrotic tissue | 96
acute respiratory distress syndrome | 96
sepsis | 96
ventilatory support | 96
antibiotic therapy | 96
anastomotic dehiscence | 96
EVAC therapy | 96
Esosponge placement | 96
Esosponge in pleural space | 96
overtube | 96
14 treatment sessions | 96
treatment sessions over 35 days | 168-840
leak and cavity size improved | 168-840
development of healthy-appearing granulation tissue | 168-840
inflammatory indexes improved | 168-840
clinical conditions improved | 168-840
endoscopic findings | 168-840
CT scans | 168-840
no complications | 168-840
endoscopic evaluation | 840
cleaner and smaller cavity | 840
1 cm cavity | 840
two esophageal fully covered SEMS | 840
Taewoong Niti-S Beta Stent | 840
liquid diet | 840
SEMS placement | 840
SEMS kept for 3 weeks | 840-1008
endoscopy | 1008
esophagram | 1008
leak resolution | 1008
tiny persistent depression | 1008
no symptoms of recurrent fistula formation | 1512
SEMS removal | 1008