24 years old | 0
    female | 0
    26th week of first pregnancy | 0
    abdominal pain | -120
    abdominal distension | -120
    constipation | -120
    pain gradually increasing in severity | -120
    hypotension | 0
    tachycardia | 0
    tachypnea | 0
    asymmetrically distended abdomen | 0
    tenderness all over abdomen | 0
    empty rectum on digital examination | 0
    elevated white cell count (16,000/mm3) | 0
    normal urine analysis | 0
    distended bowel loop on ultrasound | 0
    moderate amount of free fluid in peritoneal cavity on ultrasound | 0
    single viable fetus confirmed | 0
    clinical diagnosis of intestinal obstruction | 0
    abdominal X-ray showing dilated large bowel with abnormal gas pattern | 0
    coffee bean appearance on X-ray | 0
    sigmoidoscopy confirmed twisted sigmoid colon | 0
    failure to negotiate obstruction | 0
    foetal distress (deceleration in heart rate) | 0
    emergency laparotomy | 0
    midline laparotomy | 0
    distended sigmoid loop with ischemic and gangrenous changes | 0
    necrosis due to twisted sigmoid mesocolon | 0
    posterior displacement of necrotic colon by pregnant uterus | 0
    lower segment caesarean section | 0
    male preterm infant (750 g) delivered | 0
    infant admitted to neonatal ICU | 0
    mechanical ventilation for lung immaturity | 0
    resection of gangrenous sigmoid colon | 0
    Hartmann’s procedure | 0
    end colostomy fashioned | 0
    closure of rectal stump below peritoneal reflection | 0
    uneventful post-operative course | 0
    discharged home on 9th post-operative day | 216
    infant discharged after 10 weeks in neonatal ICU | 0
    reversal of Hartmann’s procedure after 6 months | 0
    colo-rectal anastomosis | 0
