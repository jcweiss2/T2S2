62 years old | 0
male | 0
admitted to the hospital | 0
dental pain | -120
right buccal facial swelling | -120
attended general dental practitioner | -72
prescription for amoxicillin and metronidazole | -72
trismus | -24
voice changes | -24
dysphagia | -24
stroke | -2628
diet-controlled type 2 diabetes mellitus | 0
hypertension | 0
chronic alcohol abuse | 0
non-smoker | 0
trismus | 0
maximal mouth opening of 15 mm | 0
large right facial swelling | 0
tender to percussion | 0
firm collection | 0
NEWS of 0 | 0
Glasgow Coma Scale of 15 | 0
haemoglobin level of 119 g/L | 0
white cell count of 17.1×10^9/L | 0
neutrophil count of 9.5×10^9/L | 0
platelet count of 575×10^9/L | 0
urea and electrolytes normal | 0
CRP of 145 | 0
periapical radiolucencies on both the lower right second and third molars | 0
large collection in the deep peritonsillar and parapharyngeal spaces | 0
superficial component buccal to the mandible | 0
odontogenic parapharyngeal abscess | 0
intravenous co-amoxiclav | 0
dexamethasone | 0
urgent awake fibre-optic intubation | 0
examination under anaesthesia | 0
parapharyngeal swelling | 0
extension to the soft palate | 0
crossing the midline | 0
lower right second and third molar teeth extracted | 0
intraoral incision | 0
exploration of the tissue spaces | 0
copious pus | 0
intraoral drain | 0
recovered in intensive care | 48
extubated | 48
transferred to the head and neck ward | 48
breathing difficulties | 72
tired | 72
sweaty | 72
accessory muscles to breathe | 72
respiratory rate of 24 | 72
oxygen saturations of 82% | 72
improving to 96% on high flow oxygen | 72
breath sounds clear | 72
type 1 respiratory failure | 72
transferred to the surgical high dependency unit | 72
chest radiograph clear | 72
ECG clear | 72
CT pulmonary angiogram clear | 72
airway oedema | 72
regular chest physiotherapy | 72
effective, safe cough | 72
discharged | 120