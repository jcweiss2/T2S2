4 years old | 0
male | 0
presented to the emergency room | 0
fever | -72
abdominal pain | -72
neck pain | -72
trauma to the back of the skull | -168
grunting | 0
poor perfusion | 0
severe neck pain | 0
temperature 39 °C | 0
heart rate 200 per minute | 0
blood pressure 111/79 mmHg | 0
respiratory rate 40 per minute | 0
intravenous line insertion | 0
two boluses of intravenous fluid administered | 0
full septic work-up | 0
broad spectrum antibiotics started | 0
admitted to the pediatric intensive care unit | 0
progressive left neck pain | 0
neck swelling | 0
lateral neck radiograph taken | 0
slightly thickened prevertebral soft tissue | 0
computed tomography scan of the neck with contrast | 0
minimal fluid collection in the retropharyngeal space | 0
no definite abscess | 0
left jugular vein filling defect | 0
partial thrombosis of the left internal jugular vein | 0
brain venogram computed tomography confirmed thrombosis | 0
blood culture positive for Methicillin-sensitive Staphylococcus aureus | 0
repeated culture with same pathogen | 0
cerebrospinal fluid culture negative | 0
persistent growth of MSSA | 0
echocardiography done | 0
no vegetation | 0
no signs of infective endocarditis | 0
jugular vein thrombosis | 0
MSSA bacteremia/sepsis | 0
diagnosis of Lemierre syndrome | 0
new left-sided neck swelling | 0
imaging studies confirmed left vertebral artery aneurysm | 0
coiling of the aneurysm | 0
insertion of a peripherally inserted central catheter (PICC) line | 0
episodes of bradycardia | 0
ECG done | 0
Type I Brugada syndrome pattern | 0
follow up ECGs repeated | 0
abnormal ECG findings completely disappeared | 0
no family history of cardiac diseases | 0
no family history of sudden death | 0
genetic studies for Brugada syndrome negative | 0
SCN5A gene negative | 0
discharge from the hospital | 0
ECGs repeated after discharge | 0
normal ECGs | 0
no Brugada pattern | 0
follow-up with pediatric cardiology | 0
family counseled regarding Brugada syndrome | 0
precautions to treat any fever immediately | 0
precautions during swimming | 0
avoid over the counter medications | 0
no documented fever at time of Brugada pattern appearance | 0
Brugada syndrome unmasked after PICC line insertion | 0
