22 years old | 0
primigravida | 0
pregnancy | 0
hyperemesis gravidarum | 0
vaginal delivery | 0
male infant | 0
born at 40 6/7 weeks | 0
uncomplicated delivery | 0
no family history of inborn errors of metabolism | 0
newborn screen collected | 24
tachypnea | -72
discharged home | 96
poor oral intake | 96
difficulty establishing breastfeeding | 96
fever | 120
poor feeding | 120
dehydration | 120
admitted to intensive care unit | 120
rehydration | 125
sepsis evaluation | 125
newborn screen returned | 125
elevated C14:1 | 125
elevated C14:2 | 125
elevated C14 | 125
increased C14:1/C16 ratio | 125
VLCADD | 125
normal EKG | 125
normal echocardiogram | 125
infectious work-up completed | 125
antibiotic medication | 125
antiviral medication | 125
negative cultures | 125
negative testing | 125
normal glucose concentrations | 76
elevated creatine kinase | 76
rhabdomyolysis | 76
elevated BUN | 76
elevated creatinine | 76
renal dysfunction | 76
mildly elevated liver function tests | 76
aggressive hydration | 125
10% dextrose-containing fluids | 125
medical food low in long chain fat | 125
enriched with medium chain triglycerides | 125
total fluid intake at two times maintenance | 125
CK decline | 125
creatinine improvement | 125
labs improvement | 125
discharged | 456
initial plasma acylcarnitine concentrations | 125
decreased with treatment | 125
ACADVL mutations | 125
c.848T>C (p.Val243Ala) | 125
c.751A>G (p.Ser251Gly) | 125
normal growth | 0
normal development | 0
diet treatment | 0
C14:1 elevated | 0
l-Carnitine supplementation | 504
low plasma free carnitine concentrations | 504
hospitalizations | 0
illness | 0
poor oral intake requiring g-tube placement | 0
no further rhabdomyolysis | 0
transient elevations in CK | 0
recurrent rhabdomyolysis | 0
hypoglycemia | 0
fasting test | 0
difficulty establishing breastfeeding | 120
severity of disease | 120
elevated C14:1 on newborn screen | 24
confirmatory plasma acylcarnitine profile | 125
glucose administration | 125
supplementation with MCT | 125
resolved rhabdomyolysis | 125
normal reference ranges | 0
