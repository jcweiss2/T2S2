10 years old | 0
male | 0
admitted to the hospital | 0
pain in epigastrium | -72
hepatomegaly | -72
dull pain | -72
mild to moderate pain | -72
no radiation | -72
computed tomography scan abdomen | -24
cystic lesion of liver | -24
cystic lesion of kidney | -24
positive Anti-Echinococcus IgG antibody | -24
diagnosis of hydatid cyst of liver and kidney | -24
inhalational induction with sevoflurane | 0
administration of fentanyl | 0
administration of vecuronium | 0
trachea intubated | 0
injection of 10% PI | 0
heart rate increased | 1
hypercarbia | 1
hyperthermia | 1
administration of paracetamol | 1
infusion of normal saline | 1
arterial blood gas analysis | 1
metabolic acidosis | 1
acute renal failure | 1
decreased urine output | 1
administration of fluid bolus | 1
administration of frusemide | 1
improved urine output | 2
presumptive diagnosis of anaphylaxis | 2
administration of hydrocortisone | 2
administration of pheniramine maleate | 2
shifted to ICU | 2
investigations in ICU | 2
severe metabolic acidosis | 2
plan for haemodialysis | 2
tachycardia | 2
fluid responsive | 2
administration of Sterofundin | 2
administration of albumin | 2
administration of hydrocortisone | 2
bedside echocardiography | 3
good cardiac contractility | 3
under filled heart chambers | 3
inferior vena cava diameter | 3
collapsibility | 3
initiation of haemodialysis | 3
correction of acidosis | 6
settling of heart rate | 6
trachea extubated | 24
completion of dialysis | 24
tapering of hydrocortisone infusion | 24
stopping of hydrocortisone infusion | 24
discharge from ICU | 48
shifting to ward | 48