55 years old | 0
male | 0
non-smoker | 0
presented acutely | 0
fever | 0
joint pain | 0
cold | 0
painful extremities | 0
non-erosive rheumatoid arthritis | -52560
rheumatoid factor positive | -52560
anti-cyclic citrullinated peptide negative | -52560
methotrexate | -17520
limited cutaneous systemic sclerosis overlap syndrome | -17520
Raynaud’s phenomenon | -17520
sclerodactyly | -17520
telangiectasia | -17520
sicca symptoms | -17520
anti-nuclear antibodies positive | -17520
anti-RNP (U1RNP) specificity | -17520
cold digits | 0
small joint synovitis of the hands | 0
small joint synovitis of the feet | 0
raised white cell count | 0
neutrophil count 17.8×109/L | 0
C-reactive protein 301 mg/L | 0
chest x-ray | 0
urine dip | 0
empirical intravenous antibiotics | 0
oral corticosteroids | 0
prednisolone 20 mg od | 0
continuous prostaglandin analog infusion | 0
iloprost infusion | 0
body temperature spiked | 0
inflammatory markers rose further | 0
antibiotic therapy broadened | 0
transesophageal echocardiogram | 0
negative blood cultures | 0
computed tomography of chest | 0
computed tomography of abdomen | 0
computed tomography of pelvis | 0
necrosis of hands | 168
necrosis of feet | 168
therapeutic dose of low-molecular weight heparin | 168
clopidogrel | 168
iloprost infusion uptitrated | 168
deterioration in extremities | 168
magnetic resonance angiography | 168
intravenous methylprednisolone 500 mg | 168
C-reactive protein fell to 153 mg/L | 168
wet gangrene of lower limbs | 240
bilateral below-knee amputations | 240
prednisolone 60 mg daily | 240
intravenous immunoglobulin over 5 days | 240
demarcation of tissue gangrene | 240
no further progression of necrosis | 240
strong ulnar pulses | 240
strong radial pulses | 240
CRP fell rapidly | 240
antibiotics stopped | 240
mycophenolate mofetil initiated | 240
negative anti-centromere antibodies | 240
negative anti-Scl70 antibodies | 240
negative anti-neutrophil cytoplasmic antibody | 240
negative antiphospholipid antibodies | 240
negative cryoglobulins | 240
negative serology for hepatitis B | 240
negative serology for hepatitis C | 240
negative serology for HIV | 240
normal lipid profile | 240
examination by plastic surgeon | 240
advised amputation at both elbows | 240
conservative management | 240
dry gangrene | 240
await auto-amputation | 240
slow improvement in proximal areas of hands | 240
monthly IVIG | 240
weaning dose of prednisolone | 240
vasodilator therapy | 240
sildenafil | 240
mycophenolate mofetil uptitrated to 1g BD | 240
rivaroxaban | 240
discharged to rehabilitation | 2880
learned to use prostheses independently | 2880
fifth digits auto-amputated | 4320
limited surgical resection of necrotic digits | 12960
remains in remission | 12960
significant functional impairment | 12960
manages well | 12960
