52 years old | 0
female | 0
admitted to the emergency department | 0
diffuse myalgias predominantly in the lower limbs | -72
fever | -72
cough | -72
temperature of 35.9°C | 0
pulse oxygen saturation of 99% on room air | 0
heart rate of 62 per minute | 0
blood pressure of 127/89 mmHg | 0
diffuse muscle pain | 0
creatine kinase levels at 15000 IU/L | 0
SARS-CoV-2 RNA positive | 0
L452R mutation | 0
unremarkable renal function | 0
CT showing mild pulmonary infiltrates | 0
no pulmonary embolism | 0
hospitalized in the respiratory department | 0
admitted to the intensive care unit | 48
Glasgow score of 12/15 | 48
temperature of 40°C | 48
heart rate of 130 per minute | 48
hypotension at 70/30 mmHg | 48
anuria | 48
diffuse mottling | 48
no dyspnea | 48
treated with oxygen (15 L/min) | 48
intravenous saline | 48
bicarbonate 1.4% | 48
vasopressor support with norepinephrine | 48
intubated | 48
mechanically ventilated | 48
metabolic acidosis | 48
hyperkalemia | 48
anuria leading to renal replacement therapy | 48
hydrocortisone 50 mg/6 h | 48
antibiotics (amoxicillin/clavulanic acid) | 48
preventive anticoagulation with enoxaparin (4000 IU) | 48
continued hemodynamic deterioration | 48
cardiorespiratory arrest | 48
unsuccessful resuscitation after 45 minutes | 48
primary hypertension | 0
WBC 10.11 g/L | 0
lymphocytes 1.32 g/L | 0
CRP 37.8 mg/L | 0
D-dimer 2.50 μg/ml | 0
hypersensitive troponin T 962 ng/l | 0
creatinine 129 mmol/L | 0
eGFR 38 ml/min/1.73 m² | 0
urea 12.8 mmol/L | 0
K+ 6.4 mmol/L | 0
CPK 100557 IU/L | 0
myoglobin >30000 g/L | 0
AST 2394 U/L | 0
ALT 561.8 U/L | 0
COVID-19 viral load 310/ml | 0
negative pneumococcal/legionella antigenuria | 0
pH 7.43 | 0
PO2 98 mmHg | 0
PCO2 18 mmHg | 0
HCO3- 11.9 mmol/L | 0
lactate 6.7 | 0
pH 7.11 | 48
PO2 67 mmHg | 48
PCO2 34 mmHg | 48
HCO3; 10.8 mmol/L | 48
lactate 15.6 | 48
hypersensitive troponin T 2028 ng/l | 48
K+ 6.7 mmol/L | 48
CPK 101624 IU/L | 48
AST 1978 U/L | 48
ALT 517 U/L | 48
