43 years old | 0
    man | 0
    myelodysplastic syndrome with excess blasts-1 | 0
    scheduled for bone marrow transplantation | 0
    received 6 courses of treatment with azacytidine | -672
    Kawasaki disease | -960
    hypertension | -960
    hyperuricemia | -960
    angina pectoris | -960
    surgery for coronary artery lesions caused by Kawasaki disease | -960
    postoperative no functional cardiac abnormalities | -960
    no treatment for inactive Kawasaki disease | -960
    height 175 cm | 0
    weight 90 kg | 0
    does not smoke | 0
    denies alcohol use | 0
    denies illicit drug use | 0
    COVID-19 IgG/IgM combined antibody test negative | 0
    PICC inserted into the right upper arm | 0
    hematologist performed 30 PICC procedures | 0
    venous access achieved without difficulty | 0
    ultrasound-guided puncture | 0
    fluoroscopic wire/catheter guidance | 0
    hematologist wore surgical cap | 0
    surgical mask | 0
    sterile gown | 0
    sterile gloves | 0
    clean working space | 0
    day 4 | 96
    local redness observed at insertion site | 96
    hematologist removed the catheter | 96
    initiated broad-spectrum antimicrobial therapy with piperacillin/tazobactam | 96
    initiated teicoplanin | 96
    day 6 | 144
    fever up to 39.6°C | 144
    hematologist changed antimicrobials to meropenem | 144
    continued teicoplanin | 144
    initiated clindamycin | 144
    right upper arm swelled gradually | 144
    difficulty bending elbow | 144
    day 8 | 192
    fever 40.2°C | 192
    hematologist consulted orthopedic surgeon | 192
    antibacterial therapy had no effect | 192
    fever did not decrease | 192
    swelling worsened | 192
    orthopedic surgeon decided further antimicrobial therapy advisable | 192
    patient seemed to be doing well | 192
    less redness around insertion site | 192
    decided to continue conservative treatment for next 2 days | 192
    afternoon of day 10 | 240
    Glasgow Coma Scale E4V5M6 | 240
    temperature 39.1°C | 240
    blood pressure 79/43 mmHg | 240
    heart rate 90 beats/min | 240
    respiratory rate 16 breaths/min | 240
    oxygen saturation 100% | 240
    non-rebreather reservoir mask at 10 L/min oxygen | 240
    physical examination exacerbation of swelling and redness in right upper arm | 240
    no blistering | 240
    muscle pain | 240
    tenderness to palpation along right biceps brachii muscle | 240
    white blood cell count 10.4×103/μL with 94.0% neutrophils | 240
    hemoglobin 7.0 g/dL | 240
    platelet 18.8×104/μL | 240
    CRP 24.6 mg/dL | 240
    total protein 5.1 g/dL | 240
    albumin 2.6 g/dL | 240
    aspartate aminotransferase 18 U/L | 240
    alanine aminotransferase 15 U/L | 240
    total bilirubin 1.7 mg/dL | 240
    creatine kinase 281 U/L | 240
    blood urea nitrogen 39 mg/dL | 240
    creatinine 2.53 mg/dL | 240
    prothrombin time/international normalized ratio 1.61 | 240
    fibrinogen 699 mg/dL | 240
    fibrin and fibrinogen degradation products 15.1 μg/mL | 240
    D-dimer 9.6 μg/mL | 240
    procalcitonin 46.2 ng/mL | 240
    presepsin 1420 pg/mL | 240
    plain radiograph of upper arm showed no gas in soft tissue | 240
    fat-suppressed T2-weighted MRI showed diffuse heterogeneous high signal intensity in biceps brachii, brachialis, and triceps brachii muscles | 240
    suspected emergency necrotizing soft tissue infection | 240
    progression to septic shock | 240
    patient underwent urgent debridement surgery | 240
    administration of large fluid infusion | 240
    noradrenaline infusion | 240
    broad-spectrum antimicrobial agents with meropenem | 240
    initiated daptomycin | 240
    continued clindamycin | 240
    initiated posaconazole | 240
    no infectious findings between skin and subcutaneous tissue | 240
    brachial fascia severely swollen with evidence of internal pressure | 240
    incising brachial fascia | 240
    no obvious exudation of pus | 240
    more than half of biceps brachii and brachialis muscles poorly colored | 240
    scattered white spots on surface of muscles | 240
    muscles easily torn with finger | 240
    infectious myositis | 240
    myonecrosis | 240
    DVT of brachial vein observed | 240
    catheter insertion site confirmed | 240
    submitted muscle tissues and surrounding exudate for tissue culture | 240
    submitted muscle tissues for histopathological examination | 240
    excised infected or necrotic muscle | 240
    cleaned wound thoroughly | 240
    wound left open postoperatively | 240
    day 11 | 264
    evaluated extent of upper-extremity DVT with echo and enhanced computed tomography | 264
    no thrombosis in infra-clavicular and axillary veins | 264
    received intravenous heparin 10,000 units per day for 14 days | 264
    admitted to ICU postoperatively | 264
    vital signs stable on day 13 | 312
    culture tests negative | 312
    histopathological examination showed infectious myositis in biceps brachii and brachialis muscles | 312
    day 14 | 336
    rehabilitation of right upper extremity initiated | 336
    treated in ICU until day 16 | 384
    regular wound cleaning in ward | 384
    regular debridement in operation room | 384
    signs of infection disappeared on day 20 | 480
    aimed to improve edema and granulation with negative-pressure wound therapy | 480
    RENASYS TOUCH™ used for 3 weeks | 480
    shoe-lace technique using vessel tape for rapid wound closure | 480
    day 25 | 600
    changed antimicrobials and antifungals to oral tosufloxacin | 600
    changed to oral posaconazole | 600
    continued until day 40 | 960
    day 35 | 840
    CRP levels negative | 840
    day 52 | 1248
    wound closed spontaneously | 1248
    six months after PICC insertion | 4320
    range of motion of right elbow 100 degrees flexion | 4320
    range of motion of right elbow -30 degrees extension | 4320