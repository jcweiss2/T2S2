67 years old | 0
male | 0
admitted to the hospital | 0
obstructive jaundice | -672
anorexia | -672
weight loss | -672
biliary obstruction | -672
raised serum bilirubin | -672
raised serum aspartate aminotransferase | -672
raised serum alkaline phosphatase | -672
ultrasound scan | -24
CT scan | -24
intraluminal filling defect | -24
endoscopic retrograde cholangiopancreatography | -24
biliary stenting | -24
high-grade dysplastic cells | -24
no evidence of invasive malignancy | -24
provisional diagnosis of cholangiocarcinoma | -24
pylorus-preserving pancreatoduodenectomy | 0
Roux-en-Y reconstruction | 0
pancreatojejunostomy | 0
hepaticojejunostomy | 0
gastrojejunostomy | 0
histological examination | 24
high-grade biliary dysplasia | 24
cystic duct | 24
intrapancreatic segment of the common bile duct | 24
low-volume pancreatic leak | 48
sepsis | 48
haemoglobin | 48
white cell count | 48
neutrophil count | 48
platelet count | 48
bilirubin | 48
aspartate aminotransferase | 48
alanine aminotransferase | 48
alkaline phosphatase | 48
C-reactive protein | 48
pleural and peritoneal drain placement | 72
gastroparesis | 72
nasojejunal tube | 72
discharged | 168
haematemesis | 168
collapse | 168
haemodynamically unstable | 168
transfused with packed red blood cells | 168
transfused with platelets | 168
transfused with coagulation products | 168
angiogram | 168
gastro-duodenal artery stump haemorrhage | 168
covered stent | 168
bile leak | 192
retrievable covered stent | 192
percutaneous transhepatic cholangiography | 192
CT-guided drainage | 192
broad-spectrum antibiotics | 192
Enterococcus faecalis | 192
discharged | 336
jaundice | 8064
biliary sepsis | 8064
liver function tests | 8064
bilirubin | 8064
aspartate aminotransferase | 8064
alanine aminotransferase | 8064
alkaline phosphatase | 8064
C-reactive protein | 8064
CT scan | 8064
central soft tissue mass | 8064
liver lesions | 8064
metastatic disease | 8064
ultrasound-guided liver biopsy | 8064
antibiotics | 8064
percutaneous transhepatic cholangiogram | 8064
biliary drains | 8064
repeat CT | 8448
repeat biopsy | 8448
moderately differentiated adenocarcinoma | 8448
metastatic cholangiocarcinoma | 8448
re-assessment of pancreatico-duodenectomy specimen | 8448
no focus of invasive cancer | 8448
liver function tests | 8448
bilirubin | 8448
alanine aminotransferase | 8448
aspartate aminotransferase | 8448
alkaline phosphatase | 8448
gamma-glutamyl transferase | 8448
palliative care | 8448
died | 8512