39 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
height 155 cm | 0 | 0 | Factual
weight 44.5 kg | 0 | 0 | Factual
mild dyspnea | 0 | 0 | Factual
carinal resection | 0 | 0 | Factual
reconstruction | 0 | 0 | Factual
adenoid cystic carcinoma | 0 | 0 | Factual
chest computed tomography | -24 | -24 | Factual
bronchoscopy | -24 | -24 | Factual
left mainstem bronchus obstruction | -24 | 0 | Factual
carina obstruction | -24 | 0 | Factual
right mainstem bronchus obstruction | -24 | 0 | Factual
no underlying diseases | 0 | 0 | Factual
preoperative examinations normal | 0 | 0 | Factual
moderate obstructive pattern | 0 | 0 | Factual
forced expiratory volume | 0 | 0 | Factual
forced vital capacity | 0 | 0 | Factual
general anesthesia | 0 | 0 | Factual
propofol | 0 | 0 | Factual
remifentanil | 0 | 0 | Factual
rocuronium | 0 | 0 | Factual
tracheal intubation | 0 | 0 | Factual
right-sided double-lumen tube | 0 | 0 | Factual
right lateral position | 0 | 0 | Factual
left bronchi dissection | 0 | 20 | Factual
left vasculature dissection | 0 | 20 | Factual
thoracoscopic surgery | 0 | 20 | Factual
right OLV | 0 | 20 | Factual
arterial oxygen tension 462 mmHg | 20 | 20 | Factual
FIO2 1.0 | 20 | 20 | Factual
single-lumen endotracheal tube | 20 | 20 | Factual
bronchial blocker | 20 | 20 | Factual
left lateral position | 20 | 40 | Factual
right thoracotomy | 20 | 40 | Factual
left OLV | 20 | 40 | Factual
peak airway pressure 28 cmH2O | 40 | 40 | Factual
tidal volume 300 ml | 40 | 40 | Factual
PaO2 110 mmHg | 40 | 40 | Factual
FIO2 1.0 | 40 | 40 | Factual
carinal resection | 40 | 60 | Factual
LMB resection | 40 | 60 | Factual
sterile reinforced endotracheal tube | 40 | 60 | Factual
left OLV | 40 | 60 | Factual
airway pressure 35 cmH2O | 60 | 60 | Factual
oxygen saturation 70% | 60 | 60 | Factual
RMB resection | 60 | 80 | Factual
additional sterile endotracheal tube | 60 | 80 | Factual
differential bilateral lung ventilation | 60 | 80 | Factual
oxygen saturation 100% | 80 | 80 | Factual
carina removal | 80 | 100 | Factual
tracheobronchial anastomosis | 80 | 100 | Factual
no air leak | 100 | 100 | Factual
left lung removal | 100 | 120 | Factual
right hemithorax closure | 100 | 120 | Factual
non-dependent right OLV | 120 | 140 | Factual
oxygen saturation 80% | 140 | 140 | Factual
left pulmonary artery clamping | 140 | 140 | Factual
oxygen saturation 100% | 140 | 140 | Factual
left pulmonary artery ligation | 140 | 140 | Factual
right thoracotomy closure | 140 | 160 | Factual
left thoracotomy | 160 | 180 | Factual
left pneumonectomy | 160 | 180 | Factual
tracheal extubation | 180 | 180 | Factual
intensive care unit | 180 | 312 | Factual
discharge | 312 | 312 | Factual