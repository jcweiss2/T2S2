27 years old | 0
woman | 0
decompensated liver cirrhosis | 0
Model for End-Stage Liver Disease score of 30 | 0
primary biliary cholangitis | 0
autoimmune hepatitis overlap | 0
admitted to the intensive care unit | 0
septic shock | 0
acute kidney injury | 0
multidrug-resistant Escherichia coli urinary tract infection | 0
propranolol | 0
primary variceal prophylaxis | 0
chronic normocytic anemia | 0
baseline hemoglobin 8.5 mg/dL | 0
hematochezia | -1344
esophagogastroduodenoscopy | -1344
nonbleeding grade I esophageal varices | -1344
moderate portal hypertensive gastropathy | -1344
flexible sigmoidoscopy | -1344
mild nonbleeding internal hemorrhoids | -1344
no rectal varices | -1344
negative for spontaneous bacterial peritonitis | 0
hematochezia | 48
worsening anemia | 48
hemoglobin 5.7 mg/dL | 48
EGD | 48
severe portal hypertensive gastropathy | 48
4 nonbleeding grade III esophageal varices | 48
banded 4 times | 48
flexible sigmoidoscopy | 48
distal rectum with overlying clot | 48
oozing on water irrigation | 48
bleeding rectal varix | 48
placement of 1 band | 48
worsening anemia | 72
hemoglobin 6.7 mg/dL | 72
packed red blood cells | 72
fresh frozen plasma | 72
repeat flexible sigmoidoscopy | 72
large blood clot | 72
ulceration | 72
mild oozing | 72
previously seen rectal varix | 72
prior band dislodgement | 72
placement of 2 bands | 72
successful hemostasis | 72
persistent hematochezia | 192
hemoglobin drop | 192
hemoglobin 6.7 mg/dL | 192
packed red blood cells | 192
colonoscopy | 192
medium-sized bleeding rectal varix | 192
stigmata of prior banding | 192
overlying clot | 192
necrotic ulcer base | 192
hot snare with soft coagulation | 192
resection of protuberant part of clot | 192
resection of bands | 192
bleeding vessel at base | 192
placement of over-the-scope clip | 192
complete hemostasis | 192
no bleeding at end of procedure | 192
transferred to transplant center | 192
died from septic shock | 240
