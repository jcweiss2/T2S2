76 years old | 0
female | 0
admitted to the hospital | 0
fevers | -72
nonproductive cough | -72
dyspnea | -72
hypertension | -8760
hyperlipidemia | -8760
hypothyroidism | -8760
intubated | 0
respiratory distress | 0
hypoxic respiratory failure | 0
tachycardia | 0
diffusely decreased breath sounds | 0
crackles | 0
severe respiratory distress | 0
blood pressure 110/53 mm Hg | 0
pulse rate 124 beats/min | 0
respiratory rate 31 breaths/min | 0
oxygen saturation 79% | 0
temperature 102.3°F | 0
cardiovascular examination revealed tachycardia | 0
lung exam revealed diffusely decreased breath sounds and crackles | 0
potassium 2.2 mEQ/L | 0
creatinine 1.79 mg/dL | 0
C-reactive protein 23.10 mg/L | 0
interleukin-6 (IL-6) 781.46 mg/L | 0
lactate dehydrogenase 334 U/L | 0
ferritin 457 ng/mL | 0
procalcitonin 15.20 ng/mL | 0
prothrombin time 18.9 seconds | 0
fibrinogen >600 mg/dL | 0
white blood cell count 16.1 cells/L | 0
IgG 1622 mg/dL | 0
tested positive for SARS-CoV-2 | 0
troponin 0.03 ng/dL | 0
high-sensitivity troponin 503 ng/L | 48
proBNP 35,000 pg/mL | 48
chest radiograph showed diffuse bilateral pulmonary edema | 0
electrocardiogram showed no signs of ischemia | 0
normal sinus rhythm | 0
left ventricular (LV) hypertrophy | 0
QTc interval of 680 ms | 0
transthoracic echocardiogram (TTE) revealed a severely decreased LV systolic function | 24
segmental wall motion abnormalities | 24
akinesis of the distal segments of the left ventricle | 24
akinesis of the mid and distal portions of the right ventricle | 24
ejection fraction (EF) of 25%–30% | 24
vasopressor support with norepinephrine | 24
ARDSnet protocol | 24
treated with tocilizumab | 24
treated with intravenous immunoglobulin | 24
treated with ceftriaxone | 24
treated with cefdinir | 24
treated with cefepime | 24
treated with intravenous furosemide | 48
cardiac enzymes were found to be elevated | 48
repeat bedside TTE was performed | 48
LVEF of 20%–25% | 48
severe viral myocarditis | 48
transferred to a tertiary center | 72
complete 2D echocardiogram revealed an LVEF of 25%–30% | 72
wall motion abnormalities | 72
non-ST-elevation myocardial infarction | 72
treated with therapeutic enoxaparin | 72
LVEF recovered to 50% on TTE | 120
mildly reduced LV systolic function | 120
mid-septal and apical hypokinesis | 120
mildly reduced right ventricular function | 120
inflammatory markers greatly improved | 120
IL-6 continued to downtrend | 120
high-sensitivity troponin decreased | 120
discharged from tertiary center | 168
transferred back to intensive care unit | 168