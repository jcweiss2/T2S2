91 years old | 0
female | 0
admitted to the hospital | 0
febrile sensation | -48
general weakness | -48
hypertension | -672
dementia | -672
bevantolol | -672
donepezil | -672
risperidone | -672
ambulate | -672
communicate | -672
short-leg splint | -336
undisplaced fractures | -336
4th metatarsal bone | -336
5th metatarsal bone | -336
right foot | -336
watery diarrhea | -168
sputum | -48
abdominal CT scan | -24
fluid retention | -24
gas shadow | -24
right gluteal area | -24
greater trochanter | -24
femur | -24
sepsis | -24
soft tissue infection | -24
transferred to hospital | 0
intensive care | 0
systolic blood pressure | 0
diastolic blood pressure | 0
pulse rate | 0
respiratory rate | 0
body temperature | 0
physical examination | 0
skin necrosis | 0
fluctuation | 0
heat generation | 0
hip | 0
thigh | 0
white blood cell count | 0
neutrophils | 0
erythrocyte sedimentation rate | 0
C-reactive protein | 0
broad-spectrum antibiotics | 0
ceftriaxone | 0
clindamycin | 0
gas observed | 0
plain radiographs | 0
pelvis | 0
magnetic resonance imaging | 0
abscess formation | 0
right gluteus maximus | 0
gluteus medius | 0
left gluteus maximus | 0
air formation | 0
inflammatory lesions | 0
cystic shadows | 0
posterosuperior surface | 0
uterus | 0
bilateral NF | 0
hip joints | 0
fascia | 0
muscles | 0
surgery | 24
incisions | 24
debridements | 24
posterolateral approach | 24
right lateral position | 24
skin lesion | 24
thigh | 24
hip | 24
bacterial cultures | 24
abscess | 24
necrotic tissues | 24
gluteus medius | 24
greater trochanter | 24
femur | 24
deep muscles | 24
fascia | 24
subcutaneous tissues | 24
right hip joint puncture | 24
culture tests | 24
drainage catheter | 24
sutured | 24
gynecologist | 24
cystic lesions | 24
superior surface | 24
uterus | 24
transvaginal sonography | 24
puncture | 24
aspiration | 24
aspirated fluid | 24
non-inflammatory | 24
intensive care | 48
systolic blood pressure | 48
body temperature | 48
white blood cell count | 48
neutrophil | 48
erythrocyte sedimentation rate | 48
C-reactive protein | 48
Escherichia coli | 48
ciprofloxacin | 48
drainage catheter | 168
tip culture | 168
suture removal | 336
complications | 336
ambulation | 336
sepsis | 336
trauma | 336
operation | 336
infection | 336
pressure ulcer | 336
ischial areas | 336
management | 336
general symptoms | 336
high fever | 336
findings | 336
postoperative day 14 | 336
C-reactive protein | 336
body temperature | 336
antibiotic administration | 336
follow-up MRI | 336
abscess | 336
left greater trochanter | 336
gluteus medius | 336
incision | 360
debridement | 360
left aspect | 360
necrotic tissues | 360
wide posterolateral incision | 360
pus | 360
bacterial cultures | 360
drained serosanguinous fluid | 360
drainage catheter | 360
intensive care unit | 360
recovered | 360
bacteria | 360
culture tests | 360
body temperature | 360
ischial pressure ulcer | 360
wound dressing | 360
care | 360
ambulation | 504
wheelchair | 504
infection-related complications | 720
follow-up | 1440
patient conditions | 1440
systematic rehabilitation | 1440