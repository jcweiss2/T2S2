62 years old | 0
male | 0
COPD | 0
tobacco abuse | 0
former alcoholism | 0
hypertension | 0
bloating | -96
abdominal pain | -96
elevated liver function tests | -96
leukocytosis | -96
normocytic anemia | -96
lipase >4000 U/L | -96
lactate 1.7 mmol/L | -96
CRP 25.3 mg/dL | -96
troponin <0.012 ng/mL | -96
mass like density in the suprahilar region of the left upper lobe | -96
hepatomegaly | -96
diffuse, innumerable hypoattenuating nodules | -96
nodular enlargement of the adrenal glands | -96
periportal, peripancreatic and mild retroperitoneal lymphadenopathy | -96
bilateral lower extremity venous duplex scans | -96
abnormal liver parenchyma | -96
cholelithiasis | -96
liver biopsy | -48
CT chest with IV contrast | -48
MRI of the brain | -48
emphysema | -48
bulky left upper lobe tumor | -48
obstructed upper lobe bronchus | -48
encased main pulmonary artery and main-stem bronchus | -48
extensive mediastinal and supraclavicular lymphadenopathy | -48
chest wall invasion | -48
multiple metastatic lesions | -48
palliative radiation | -48
piperacillin/tazobactam | -48
port placement | -24
chemotherapy treatment | -24
carboplatin | -24
etoposide | -24
IV furosemide | -24
acute kidney injury | -12
worsening leukocytosis | -12
infectious disease consultation | -12
post-obstructive pneumonia | -12
lethargic | -12
hypotensive | -12
hypoxic respiratory failure | -12
arterial blood gas | -12
hypoxia | -12
septic shock | -12
tachycardic | -12
low dose Levophed | -12
colloid | -12
levofloxacin | -12
meropenem | -12
renal failure | -6
intubated | -6
high doses of norepinephrine | -6
vasopressin | -6
bronchoscopy | -6
sputum culture | -6
Enterobacter aerogenes | -6
blood cultures | -6
intermittent sinus tachycardia | -6
supraventricular tachycardia | -6
vasopressor requirement | -6
new heart rhythm | -6
echocardiogram | -6
troponins | -6
ECG | -6
fever | -6
type I Brugada wave | -6
heparin drip | -6
antiplatelet therapy | -6
type II NSTEMI | -6
hyper-dynamic left ventricle | -6
right heart chamber dilatation | -6
elevated right ventricular systolic pressure | -6
vasopressor requirement improved | 0
defervescence | 0
sinus tachycardia resolved | 0
repeat ECG | 0
resolution of Brugada wave | 0
extubated | 12
bilevel positive airway pressure | 12
nephrology evaluation | 12
dialysis | 12
anuric | 12
comfort care | 24
life saving measures ceased | 24
death | 24