57 years old | 0
female | 0
no pertinent family history | 0
hypertension | -672
amlodipine | -672
hyperlipidemia | -672
atorvastatin | -672
irritable bowel syndrome | -672
gastroesophageal reflux disease | -672
famotidine | -672
ankle injury | -12
right lateral ankle pain | -12
significant pain | -8
swelling on the lateral aspect | -8
presented to the ED | 0
physical exam of the right lower extremity | 0
swelling with a 2 cm round ecchymotic lesion | 0
limited range of motion secondary to pain | 0
intact pulses | 0
no other skin findings | 0
right leg and ankle x-ray | 0
lateral malleolar edema | 0
no acute osseous findings | 0
discharged home | 0
worsening swelling of her right lower extremity | 6
expansion of the ecchymotic lesion | 6
more painful | 6
shortness of breath | 6
emergency medical services contacted | 6
cardiac arrest | 6
hypoxic respiratory failure | 6
intubated in the field | 6
hypotension | 6
sinus tachycardia | 6
mechanically ventilated | 6
extensive hemorrhagic lesion | 6
bullous formation | 6
white blood cell count of 3.3 K/mm3 | 6
hemoglobin of 8.9 gm/dL | 6
mean corpuscular volume of 112.8 fL | 6
platelet count of 36 K/mm3 | 6
potassium 5.1 mmol/L | 6
carbon dioxide 11 mmol/L | 6
anion gap 33 mEq/L | 6
creatinine 2.9 mg/dL | 6
lactic acid 21.4 mmol/L | 6
total bilirubin 1.7 mg/dL | 6
aspartate transaminase 327 U/L | 6
alanine transaminase 164 U/L | 6
troponin of 0.110 ng/mL | 6
prothrombin time of 25.9 seconds | 6
international normalized ratio of 2.25 | 6
fibrinogen 318 mg/dL | 6
d-dimer 5200 ng/mL | 6
creatinine kinase levels of 3197 U/L | 6
metabolic acidosis | 6
pH 6.69 | 6
pCO2 69.1 mmHg | 6
HCO3 8.3 mmol/L | 6
clear lungs | 6
endotracheal tube in place | 6
small volume left inferior sylvian fissure subarachnoid hemorrhage | 6
no pulmonary embolism | 6
admitted to the intensive care unit | 6
septic shock | 6
intravenous fluids with 0.9% normal saline | 6
blood cultures obtained | 6
general surgery consulted | 6
empiric coverage with intravenous vancomycin | 6
meropenem | 6
clindamycin | 6
bedside fasciotomy of her right lower extremity | 12
bedside below the knee guillotine amputation | 12
tissue cultures obtained | 12
second set of blood cultures obtained | 12
continuous renal replacement therapy | 24
P. fluorescens and P. putida grew in blood cultures | 48
P. fluorescens and P. putida grew in tissue cultures | 48
expired due to multisystem organ failure | 48