23 years old | 0
female | 0
visited the emergency room | 0
abdominal pain | 0
nausea | 0
vomiting | 0
major depression | -936
bulimia nervosa | -936
frequent vomiting after episodes of binge eating | -936
numerous suicide attempts | -936
ate a very large quantity of food | -240
abdominal distension | -240
tenderness | -240
clear gastric distension on CT | -240
normal blood tests | -240
declined hospitalization | -240
re-visited the emergency room | -7
persistent abdominal pain | -7
mental confusion | -7
unconscious | -7
severe abdominal distension | -7
abdominal rigidity | -7
pale legs | -7
no abdominal auscultation sounds | -7
absent dorsalis pedis pulse | -7
shock | -7
blood pressure 60/40 mmHg | -7
heart rate 160 beats/min | -7
aspiration rate 22 times/minute | -7
temperature 36.4℃ | -7
metabolic acidosis | -7
electrolyte imbalance (Na+ 157 mM/L, K+ 6.2 mM/L, Cl"130 mM/L) | -7
severe hypoglycemia (15 mg/dl) | -7
acute renal failure (creatinine 2.84 mg/dl) | -7
sodium bicarbonate administration | -7
abdominal X-ray showing gastrointestinal tract filled with food | -7
abdominal CT showing dilated stomach, esophagus, duodenum | -7
mental state lethargic | -6
communication impossible | -6
decreased spontaneous respiration | -6
SpO2 88% | -6
endotracheal intubation | -6
Foley catheter insertion | -6
no urine output | -6
emergency hemodialysis preparation | -6
central venous catheter insertion | -6
radial artery conduit placement | -6
nasogastric tube insertion attempt | -6
abdominal CT follow-up showing food and twisted nasogastric tube | -6
no decompression via nasogastric tube | -6
mental confusion | -6
unstable vital signs | -6
decision for surgical decompression | -6
transferred to operation room | -6
crystalloid fluid administered (3,170 ml) | -6
no urine volume measured | -6
blood pressure 70/46 mmHg | 0
heart rate 128 beats/min | 0
crystalloid fluid administration | 0
norepinephrine infusion | 0
vasopressin infusion | 0
general anesthesia induction | 0
arterial blood gas analysis (pH 7.45, PaCO2 20.8 mmHg, etc.) | 0
erythrocytes prescribed | 0
furosemide injection | 0
rapid infusion system connected | 0
gastrotomy performed | 0
skin incision 10 cm | 0
drained 5,000 ml from stomach | 0
blood pressure 60/40 mmHg | 0
continuous gastric bleeding | 0
drained 6,000 ml into suction bottle | 0
arterial blood gas analysis (pH 6.75, PaCO2 46 mmHg, etc.) | 0
sodium bicarbonate administration | 0
insulin administration | 0
calcium chloride administration | 0
epinephrine injection | 0
continued gastric bleeding | 0
hemoglobin decrease | 0
additional erythrocytes prescribed | 0
fresh frozen plasma prescribed | 0
abdomen closed urgently | 0
transferred to ICU | 0
suturing completed | 0
no blood pressure measured | 0
flat radial artery waveforms | 0
no pulse detected | 0
pulseless electrical activity | 0
CPR initiated | 0
vasopressin injection | 0
abdominal closure during CPR | 0
no urine output | 0
operation duration 1 h 20 min | 0
anesthesia duration 1 h 50 min | 0
transfused 800 ml erythrocytes | 0
administered 6,200 ml crystalloid fluid | 0
drained 6,000 ml | 0
continued transfusion in ICU | 0
blood pressure unmeasurable | 0
nasogastric tube bleeding 1,000 ml | 0
abdominal bleeding continued | 0
DIC confirmed | 0
hemoglobin 1.8 g/dl | 0
heartbeat disappeared | 0
death declared | 0
