50 years old | 0
female | 0
admitted to the Emergency Department | 0
abdominal pain | -144
vomiting | -144
lactic acidosis | -144
thrombocytopenia | -144
aortic valve and mitral valve replacement | -1824
anemia | -728
chronic renal failure | -728
palpitation | -720
fever | -720
endocarditis | -720
methicillin-resistant Staphylococcus intermedius | -720
neoplasm around the mechanical aortic valve | -720
serum creatinine 331 µmol/L | -720
estimated glomerular filtration rate of 23 mL/min/1.73 m2 | -720
hemoglobin 78 g/L | -720
leukocytes 8.7×109/L | -720
polymorphonuclear neutrophils 7.57×109/L | -720
platelets 216×109/L | -720
LZD treatment | -720
warfarin treatment | -720
improved condition | -408
discharged from West China Hospital | -408
LZD treatment in a local hospital | -408
re-admitted to the ED | 0
LZD therapy | 0
drowsy | 600
dyspneic | 600
nausea | 600
vomiting | 600
persistent periumbilical pain | 600
tachypneic | 600
atrial fibrillation | 600
normotensive | 600
afebrile | 600
severe lactic acidosis | 624
severe thrombocytopenia | 624
transferred to the Emergency Intensive Care Unit | 624
hemodynamic support with norepinephrine | 624
mechanical ventilation | 624
continuous renal replacement therapy | 624
erythrocytes transfusion | 624
platelets transfusion | 624
shock | 720
multiple organ failure | 720
death | 816