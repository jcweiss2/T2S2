47 years old | 0
male | 0
admitted to the hospital | 0
chest pain | -27
shortness of breath | -27
dull pain in the left chest | -27
aggravated chest pain upon deep inhalation | -27
relieved by nitroglycerin | -26
reappearance of chest pain | -26
electrocardiogram | -18
troponin T examination | -18
normal electrocardiogram results | -18
normal troponin T results | -18
referred to the Department of Cardiology | -18
chest computed tomography (CT) | -18
inflammation of lower lobes in both lungs | -18
inflammation of inferior lingular segment of the left lung | -18
left pleural effusion | -18
ceftazidime treatment | -18
intravenously administered ceftazidime | -18
physical examination | -18
clear consciousness | -18
dulled left lower lung in percussion | -18
low left lung breath sounds | -18
no rale heard in both lungs | -18
transferred to the Department of Respiratory and Critical Care Medicine | -48
levofloxacin treatment | -48
intravenous injection of levofloxacin | -48
ultrasound-guided thoracentesis drainage | -72
examination of pleural effusion | -72
adenosine deaminase (ADA) of 50.3 U/L | -72
lactate dehydrogenase (LDH) of 2523 U/L | -72
protein level of 49.64 g/L | -72
no bacteria found in pleural fluid cytology | -72
no tumor cells found in pleural fluid cytology | -72
antibiotics regimen adjustment | -72
ceftazidime and moxifloxacin treatment | -72
rise in peak body temperature | -72
regimen readjusted to meropenem and moxifloxacin | -60
re-examination via chest CT | -56
double-under pneumonia | -56
increased pleural effusion | -56
C reactive protein examination | -52
erythrocyte sedimentation rate examination | -52
blood routine examination | -52
no obvious changes in examination results | -52
communication with the patient | -40
written informed consent form | -40
bronchoscopy | -40
alveolar lavage collection | -40
mNGS analysis | -40
no abnormalities in bronchoscopy results | -40
disappearance of fever | -40
mNGS results | -32
Gardnerella vaginalis infection | -32
Corynebacterium urealyticum infection | -32
negative sputum culture results | -32
negative blood culture results | -32
negative urine culture results | -32
discharged from hospital | 216
ornidazole treatment | 216
re-examination via chest CT | 216
pleural effusion in the left interlobular fissure | 216
reduction in pleural effusion | 216
follow-up | 504
physical examination | 504
no chest tightness | 504
no discomfort | 504
re-examination via chest CT | 504
absorption of inflammation in the right lower lobe | 504
reduction in pleural effusion | 504
Heart Stent Implantation | -10080
hypertension | -10080
smoking index of 500 | -10080
lobster Catering Company | -10080
dull pain in the left chest at 9 am | -27
shortness of breath after activity | -27
aggravated chest pain upon deep inhalation | -27
relieved by nitroglycerin | -26
reappearance of chest pain | -26
electrocardiogram at 7 pm | -18
troponin T examination at 7 pm | -18
normal electrocardiogram results at 7 pm | -18
normal troponin T results at 7 pm | -18
referred to the Department of Cardiology at 7 pm | -18
chest computed tomography (CT) at 7 pm | -18
inflammation of lower lobes in both lungs at 7 pm | -18
inflammation of inferior lingular segment of the left lung at 7 pm | -18
left pleural effusion at 7 pm | -18
ceftazidime treatment at 7 pm | -18
intravenously administered ceftazidime at 7 pm | -18
physical examination at 7 pm | -18
clear consciousness at 7 pm | -18
dulled left lower lung in percussion at 7 pm | -18
low left lung breath sounds at 7 pm | -18
no rale heard in both lungs at 7 pm | -18
transferred to the Department of Respiratory and Critical Care Medicine on October 7th | -48
levofloxacin treatment on October 7th | -48
intravenous injection of levofloxacin on October 7th | -48
ultrasound-guided thoracentesis drainage on October 9th | -72
examination of pleural effusion on October 9th | -72
adenosine deaminase (ADA) of 50.3 U/L on October 9th | -72
lactate dehydrogenase (LDH) of 2523 U/L on October 9th | -72
protein level of 49.64 g/L on October 9th | -72
no bacteria found in pleural fluid cytology on October 9th | -72
no tumor cells found in pleural fluid cytology on October 9th | -72
antibiotics regimen adjustment on October 10th | -72
ceftazidime and moxifloxacin treatment on October 10th | -72
rise in peak body temperature on October 10th | -72
regimen readjusted to meropenem and moxifloxacin on October 13th | -60
re-examination via chest CT on October 14th | -56
double-under pneumonia on October 14th | -56
increased pleural effusion on October 14th | -56
C reactive protein examination on October 15th | -52
erythrocyte sedimentation rate examination on October 15th | -52
blood routine examination on October 15th | -52
no obvious changes in examination results on October 15th | -52
communication with the patient on October 19th | -40
written informed consent form on October 19th | -40
bronchoscopy on October 19th | -40
alveolar lavage collection on October 19th | -40
mNGS analysis on October 19th | -40
no abnormalities in bronchoscopy results on October 19th | -40
disappearance of fever on October 19th | -40
mNGS results on October 21st | -32
Gardnerella vaginalis infection on October 21st | -32
Corynebacterium urealyticum infection on October 21st | -32
negative sputum culture results on October 21st | -32
negative blood culture results on October 21st | -32
negative urine culture results on October 21st | -32
discharged from hospital on October 23rd | 216
ornidazole treatment on October 23rd | 216
re-examination via chest CT on October 22nd | 216
pleural effusion in the left interlobular fissure on October 22nd | 216
reduction in pleural effusion on October 22nd | 216
follow-up on November 14th | 504
physical examination on November 14th | 504
no chest tightness on November 14th | 504
no discomfort on November 14th | 504
re-examination via chest CT on November 14th | 504
absorption of inflammation in the right lower lobe on November 14th | 504
reduction in pleural effusion on November 14th | 504
follow-up on February 6th | 1008
physical examination on February 6th | 1008
no chest tightness on February 6th | 1008
no discomfort on February 6th | 1008
re-examination via chest CT on February 6th | 1008
absorption of inflammation in the right lower lobe on February 6th | 1008
absorption of inflammation on the left on February 6th | 1008