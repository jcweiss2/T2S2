80 years old | 0
male | 0
admitted to the hospital | 0
urethral catheter replacement every 2 weeks | -336
urinary retention | -672
scrotal mass | -120
purulent discharge from left scrotal wall | -120
fever | -120
urethral catheter replacement | -24
pain on the left scrotum | -24
lump on the left scrotum | -24
referred to Hasan Sadikin Hospital | -24
blood pressure 90/60 mmHg | 0
heart rate 120 beats per minute | 0
respiratory rate 24 times per minute | 0
body temperature 37.5 °C | 0
lump in the left scrotum | 0
cystic on palpation | 0
pus coming out from the left scrotum | 0
purulent fluid in the urethral catheter tube | 0
scrotal ultrasound examination | 0
balloon catheter in the left scrotum | 0
hyperechoic lesion with an acoustic shadow in the posterior urethra | 0
kidney ureter bladder x-ray | 0
two radio opaque shadows in the pelvic area | 0
white blood cell count 19.790 WBC/mL | 0
hemoglobin of 7.8 g/dL | 0
serum BUN 103.14 mg/dL | 0
serum creatinine of 5.29 mg/dL | 0
serum lactate 2.1 | 0
blood glucose level of 114 mg/dL | 0
urinalysis showed >50/HPF red blood cells | 0
urinalysis showed >50/HPF white blood cells | 0
Fournier Gangrene Scoring Index (FGSI) was 18 points | 0
correction of fluid and electrolyte imbalance | 0
third generation of cephalosporin | 0
emergency necrotomy debridement | 12
retrograde urethrography | 12
contrast extravasation at the pendulare area | 12
open vesicolithotomy | 12
two stones from the bladder and urethra extracted | 12
bladder stone size was 45 × 20 × 15 mm | 12
urethral stone size was 20 × 18 × 12 mm | 12
cystostomy tube inserted | 12
incision drainage and necrotomy debridement of the scrotum | 12
5 cm defect on the urethral | 12
level of consciousness was 11 (E3M6V4) | 24
white cell count 16000 WBC/mL | 24
hemoglobin of 9.5g/dL | 24
serum BUN 67.2mg/dL | 24
serum creatinine decreased to 2.4 mg/dL | 24
shortness of breath | 48
hospital-acquired pneumonia | 48
intubated | 72
moved to the intensive care unit (ICU) | 72
respiratory problem worsened | 72
died due to respiratory failure | 96