22 years old | 0
female | 0
East Asian | 0
admitted to the hospital | 0
general malaise | -168
myalgia | -168
dyspnea | -168
fevers | -168
anorexia | -168
nasal discharge | -168
congestion | -168
abdominal pain | -168
vaginal pain | -168
dysuria | -168
cough | -168
sore throat | -168
throat pain | -168
hoarseness | -168
recent travel to Australia | -720
unprotected sex | -720
functionally independent | 0
smoked cigarettes | 0
alcohol use | 0
drug use | 0
sick contact | 0
afebrile | -24
tachycardic | -24
hypotensive | -24
oxygen requirement increased | -24
white blood cell count 6200/µL | -24
platelet count 23,000/µL | -24
creatinine 1.33 mg/dL | -24
alanine transaminase 36 U/L | -24
aspartate transaminase 59 U/L | -24
alkaline phosphatase 466 U/L | -24
total bilirubin 2.9 mg/dL | -24
serum lactic acid 4.9 mmol/L | -24
bilateral pleural effusions | -24
liver cystic lesions | -24
intrahepatic and extrahepatic bile duct dilatation | -24
mild splenomegaly | -24
right sided Bartholin gland cyst | -24
hepatic abscesses | -24
reactive gall bladder thickening | -24
Fusobacterium necrophorum in blood cultures | -24
meropenem | -24
transferred to hospital | -48
febrile | -48
tachycardic | -48
tachypneic | -48
high flow nasal cannula | -48
lung exam with crackles | -48
cardiac exam with tachycardia | -48
abdominal exam with mild right upper quadrant tenderness | -48
genitourinary exam with erythema and edema of labia | -48
no poor dentition or gingivitis | -48
white blood cell count 14,700/µL | -48
hemoglobin 11 g/dL | -48
platelet count 16,000/µL | -48
erythrocyte sedimentation rate 31 mm/h | -48
serum lactate dehydrogenase 323 U/L | -48
alkaline phosphatase 129 U/L | -48
c-reactive protein 17.05 mg/dL | -48
fibrinogen 349 mg/dL | -48
haptoglobin 59 mg/dL | -48
COVID-19 PCR negative | -48
HIV antibody screening negative | -48
urine gonorrhea and chlamydia PCR tests negative | -48
CT of neck with no evidence of abscess formation | -48
CT of chest with multiple nodular foci | -48
septic emboli | -48
multifocal pneumonia | -48
bilateral pleural effusion | -48
interval worsening of hepatic abscess burden | -48
piperacillin-tazobactam | -48
respiratory status improved | -42
diuresis | -42
transferred to general medicine ward | -42
nasal cannula | -42
ultrasound guided thoracentesis | -33
pleural fluid analysis | -33
exudative fluid | -33
fungal smear with no growth | -33
acid-fast stain negative | -33
gram stain with no organisms | -33
no aerobic or anaerobic bacterial growth | -33
repeat CT of chest, abdomen and pelvis | -31
bilateral multifocal pneumonia | -31
pleural effusions | -31
necrotizing pneumonia | -31
pulmonary abscess | -31
hepatic abscesses | -31
subcutaneous right perineal region fluid collection | -31
cardiothoracic surgery and gynecology consulted | -31
video-assisted thoracoscopic surgery (VATS) washout and decortication | -30
pleural rind acid fast staining negative | -30
biopsy with fibrinous and organizing pleuritis | -30
fibrinopurulent exudate | -30
cultures with no organisms | -30
pelvic examination | -30
right labial abscess | -30
incision and drainage | -30
clear serous fluid | -30
thick white caseous material | -30
gram stain with no organisms | -30
bacterial culture with Candida albicans | -30
contrasted CT of abdomen and pelvis | -25
nonocclusive thrombus in right common iliac vein | -25
internal iliac vein thrombus | -25
right distal external iliac vein nonocclusive thrombus | -25
transthoracic and transesophageal echocardiography | -25
no valvular vegetations | -25
no anticoagulation | -25
diagnosis of atypical Lemierre syndrome | -25
oxygen requirement decreased | -17
dyspnea decreased | -17
vulvar pain decreased | -17
intravenous ceftriaxone | -17
oral metronidazole | -17
discharged | 0
follow up appointment | 17
improvement of symptoms | 17
breathing improved | 17
vaginal pain improved | 17
appetite improved | 17
energy improved | 17
weight improved | 17
amoxicillin-clavulanate | 17