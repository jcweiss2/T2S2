69 years old | 0
male | 0
admitted to the hospital | 0
productive cough | -120
prescribed cold medicine | -120
fever | -24
chills | -24
breathlessness | -24
pain in the right chest wall | -24
visited emergency room | -24
farmer | 0
smoked for 25 years | 0
alert | 0
blood pressure 90/60 mmHg | 0
pulse rate 84/min | 0
body temperature 37.1℃ | 0
oxygen saturation 79% | 0
crackles in both lower lung fields | 0
arterial blood gas analysis | 0
pH 7.434 | 0
carbon dioxide partial pressure 34.9 mmHg | 0
oxygen partial pressure 41.0 mmHg | 0
bicarbonate 23.6 mmol/L | 0
oxygen saturation 78.3% | 0
white blood cell count 1,710/µL | 0
hemoglobin 14.6 g/dL | 0
hematocrit 45.1% | 0
platelet count 122,000/µL | 0
leucopenia | 0
no hematologic disease | 0
spontaneous recovery from leucopenia | 0
urea nitrogen 27 mg/dL | 0
creatinine 1.4 mg/dL | 0
total protein 5.8 g/dL | 0
albumin 3.5 g/dL | 0
aspartate aminotransferase 28 IU/L | 0
alanine aminotransferase 20 IU/L | 0
C-reactive protein 11.40 mg/dL | 0
prothrombin time 11.9 seconds | 0
activated partial thromboplastin time 34.7 seconds | 0
initial chest X-ray | 0
haziness in both lower lung fields | 0
endotracheal intubation | 0
transferred to ICU | 0
mechanical ventilator support | 0
ciprofloxacin | 0
piperacillin/tazobactam | 0
respiratory distress | 0
hypoxic | 48
septic shock | 48
inotropic agents | 48
pneumonia improved | 168
oxygen demand improved | 168
blood examination improved | 168
radiographic findings improved | 168
abdominal pain | 288
suprapubic catheter insertion | 288
abdominal computed tomography | 288
fluid in the proximal large intestine | 288
reduced contrast enhancement | 288
edema in the proximal large intestine | 288
exploratory laparotomy | 288
large fluid collection in the abdominal cavity | 288
necrosis of the colon | 288
subtotal colectomy | 288
ileostomy | 288
hypoxic damage of the bowel | 288
colonic infarction | 288
mucormycosis | 288
amphotericin B | 322
deteriorated | 816
died | 816