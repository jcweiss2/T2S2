45 years old | 0
    male | 0
    chronic smoker | 0
    chest pain | -2160
    progressively increasing respiratory distress | -2160
    blunt chest trauma | -2160
    two prior admissions in a local hospital | -2160
    high-resolution computed tomography (HRCT) showed bilateral hydropneumothorax | 0
    multiple rib fractures | 0
    shifted to intensive care unit (ICU) | 0
    signs of respiratory failure | 0
    bilateral chest tubes in situ | 0
    intermittent non-invasive ventilation (NIV) | 0
    antibiotics | 0
    adequate analgesia | 0
    supportive management | 0
    chest tubes removed | 24
    minimal fluid on ultrasound chest | 24
    dyspnoea persisted | 24
    repeat HRCT chest reported infective pathology (atypical pneumonia) | 24
    lesions in the apical segment of right upper lobe consistent with lymphangitis carcinomatosa | 24
    arterial blood gases reported persistently high pCO2 | 24
    mild hypoxia | 24
    acute exacerbation of COPD | 24
    type 2 respiratory failure | 24
    short course of oral steroid | 24
    20–30% improvement in dyspnoea | 72
    required NIV 3–4 hours/day | 72
    echocardiography done later | 72
    repeat contrast-enhanced computed tomography (CECT) lung done 2 weeks later | 336
    spiculated nodule in upper part of right lower lobe | 336
    multiple sclerotic lesions in vertebral body of D1 and sternum | 336
    lytic lesion in D11 (with pedicles) | 336
    ultrasound abdomen showed hepatomegaly | 336
    multiple spaceDoccupying lesions in both lobes of the liver | 336
    likely to be metastasis | 336
    fineDneedle aspiration cytology of space occupying lesion in liver reported adenocarcinoma metastasis | 336
    chemotherapy could not be started | 336
    poor general condition | 336
    expired after 10 days of diagnosis of occult primary malignancy | 456
    pulmonary lymphangitis carcinomatosa (PLC) | 336
    liver metastasis | 336
    ground glass appearance with septal thickening | 336
    peribronchovascular thickening | 336
    prominence of centrilobular interstitium | 336
    nodular thickening of interlobular septa | 336
    peribronchovascular interstitium | 336
    groundDglass appearance with septal thickening | 336
    lack of response to steroids within 2–4 weeks | 336
    rapid deterioration of dyspnoea | 336
    predominant disease in the lower lobes of the lungs | 336
    no conflicts of interest | 0
    nil financial support and sponsorship | 0
    