68 years old | 0
male | 0
obesity (body mass index: 34 kg/m2) | 0
admitted to intensive care unit (ICU) | 0
acute respiratory failure | 0
fever (38 °C) | 0
respiratory rate 30/min | 0
pulse 80/min | 0
blood pressure 102/68 mmHg | 0
low oxygen saturation (SpO2 85% on room air) | 0
SARS-CoV-2 negative | 0
Influenza A negative | 0
Influenza B negative | 0
Pneumococcal urinary antigen negative | 0
hemocultures negative | 0
endotracheal intubation | 24
mechanical ventilation | 24
progressive clinical worsening | 24
hypoxemia | 24
APACHE II Score 18 | 24
chest computed tomography (CT) scan bilateral infiltrates | 24
fibrosis | 24
areas of coalescence | 24
SARS-CoV-2 serological testing positive | 72
ventilator-associated bacterial pneumonia due to Acinetobacter baumanii | 216
multidrug resistant Acinetobacter baumanii | 216
metallo-beta-lactamase producing Acinetobacter baumanii | 216
colistin therapy | 216
tigecycline therapy | 216
catheter-related A. baumanii bacteraemia | 408
colistin therapy again | 408
tigecycline therapy again | 408
tracheal aspirate positive for Pseudomonas putida | 888
blood culture positive for Enterobacter cloacae | 888
