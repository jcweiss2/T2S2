28 years old | 0
    female | 0
    admitted to the hospital | 0
    fever | -168
    shortness of breath | -168
    spontaneous abortion | -168
    IVF-ET treatment | -1032
    obstruction in the fallopian tube | -1032
    pregnancy established | -1032
    vaginal bleeding | -216
    uterine clearance | -216
    feeling cold | -216
    chills | -216
    body temperature 38.7°C | -216
    occasional dry cough | -216
    dizziness | -216
    general fatigue | -216
    oral treatment with cefpodoxime proxetil | -216
    worsening shortness of breath | -48
    body temperature 38°C | -48
    occasional cough | -48
    chest CT revealing scattered ground-glass dense opacities | -24
    few nodular shadows in upper lobes | -24
    diagnosis of severe pneumonia | 0
    ARDS | 0
    septic shock | 0
    moderate anemia | 0
    anti-infective moxifloxacin therapy | 0
    fluid rehydration | 0
    noradrenaline administration | 0
    thymopetidum injection | 0
    vitamin C administration | 0
    double-lung pneumonia on chest X-ray | 0
    fiberoptic bronchoscopy | 0
    small yellow sputum scab | 0
    alveolar lavage fluid collected | 0
    body temperature 38°C | 24
    blood pressure 109/84 mmHg | 24
    oxygen concentration 80% | 24
    shortness of breath | 24
    sweating | 24
    sedation and analgesic treatments | 24
    PCT increased to 18.24 ng/mL | 24
    CRP 142.4 mg/L | 24
    anti-infection treatment with meropenem and linezolid | 72
    PCT 2.24 ng/mL | 96
    blood leukocyte count 4.49×10^9/L | 96
    neutrophils 82.2% | 96
    blood pressure 110/70 mmHg | 96
    heart rate 86 bpm | 96
    respiration rate 18 breaths per minute | 96
    SpO2 98% | 96
    ventilator settings reduced | 96
    arterial blood gas analysis | 96
    fever 38.4°C | 96
    CRP 90.5 mg/L | 96
    chest CT re-examination | 96
    multiple nodules in upper lobes | 96
    multiple patchy high-density shadows | 96
    mNGS test ordered | 96
    mNGS showed M. tuberculosis complex sequences | 96
    Xpert positive for M. tuberculosis | 96
    diagnosis of pulmonary TB | 96
    hematogenous disseminated pulmonary TB | 96
    discontinuation of moxifloxacin | 96
    discontinuation of meropenem | 96
    discontinuation of linezolid | 96
    quadruple anti-TB therapy initiated | 96
    chest radiograph showing extensive exudation | 168
    referral to TB hospital | 264
    M. tuberculosis culture positive | 264
    quadruple anti-TB therapy continued | 264
    ventilator assistance continued | 264
    death due to multiple organ failure | 720
    
    
<|eot_id|>
