70 years old | 0
male | 0
hypertension | 0
chronic obstructive pulmonary disease | 0
erythroderma | -1728
intense pruritus | -1728
refractory to topical corticosteroid therapy | -1728
refractory to oral corticosteroid therapy | -1728
shiny, bright red erythroderma | 0
bilateral axillary and inguinal lymph nodes were palpable | 0
basophilia of 14.1% | 0
elevated LDH | 0
parakeratosis | 0
dense lymphocytic infiltrate in the papillary dermis | 0
epidermotropism | 0
positive for CD2 | 0
positive for CD3 | 0
positive for CD4 | 0
positive for CD5 | 0
negative for CD7 | 0
negative for CD8 | 0
numerous enlarged lymph nodes in the cervical, axillary and inguinal regions | 0
Sézary cell count of 1031/mm3 | 0
axillary lymph node biopsy revealed paracortical infiltration due to Sézary syndrome | 0
Sézary syndrome diagnosis | 0
treatment with PUVA therapy | 0
treatment with interferon alpha | 0
treatment with bexarotene | 0
treatment with extracorporeal photopheresis | 0
disease progression | 0
enlarged lymph nodes | 0
uncontrollable pruritus | 0
LUC of 56.8% | 0
basophilia of 26% | 0
treatment with alemtuzumab | 0
cotrimoxazole prophylactic treatment | 0
famciclovir prophylactic treatment | 0
valganciclovir prophylactic treatment | 0
marked improvement | 72
80% erythroderma clearance | 72
pruritus cessation | 72
decrease in Sézary cell count to 0 | 72
severe neutropenia | 96
grade IV heart failure | 96
acute exacerbation of chronic obstructive pulmonary disease | 96
bronchospasm | 96
intensive care unit admission | 96
recovery with supportive treatment | 96
G-CSF therapy | 96
no signs of clinical or haematological disease activity | 624
treatment withdrawal | 96