51 years old | 0
male | 0
Caucasian | 0
admitted to the hospital | 0
hypertension | -672
severe COVID-19 | -168
acute respiratory distress syndrome | -168
mechanical ventilation | -168
ventilator-associated pneumonia | -168
carbapenem-resistant Acinetobacter baumannii | -168
ampicillin-sulbactam | -168
polymyxin B | -168
central line-related bloodstream infection | -168
carbapenem-resistant Pseudomonas aeruginosa | -168
meropenem | -168
sacral pressure injury | -168
critical illness polyneuropathy/myopathy | -168
discharged | -112
insidious pain in the lumbar region | -56
insidious pain in the right hip | -56
impairing ambulation | -56
referred to hospital | 0
severe pain on palpation | 0
severe pain on mobilization | 0
lumbar spine | 0
moderate pain in the right hip | 0
muscle strength normal | 0
reflexes normal | 0
sensitivity normal | 0
hemoglobin level 12.1 g/dL | 0
total leukocyte count 8700 cells/mm³ | 0
erythrocyte sedimentation rate 120 mm/hr | 0
C-reactive protein level 1.5 mg/dL | 0
computed tomography of the right hip | 0
periarticular calcifications | 0
heterotopic ossifications | 0
magnetic resonance imaging of the lumbar spine | 0
bone edema in the T12 and L1 vertebral bodies | 0
irregularity of the vertebral endplate | 0
psoas muscles involvement | 0
T12-L1 spondylodiscitis | 0
psoitis | 0
blood cultures negative | 0
CT-guided bone biopsy | 24
bacteria identification | 24
antimicrobial-susceptibility testing | 24
Pseudomonas aeruginosa | 24
sensitive to polymyxin B | 24
sensitive to ceftazidime-avibactam | 24
resistant to meropenem | 24
resistant to imipenem | 24
resistant to cefepime | 24
resistant to ceftazidime | 24
resistant to ciprofloxacin | 24
resistant to piperacillin-tazobactam | 24
resistant to tigecycline | 24
resistant to amikacin | 24
antimicrobial treatment initiated | 48
polymyxin B | 48
meropenem | 48
cutaneous rash | 72
switched to ceftazidime-avibactam | 72
dermatological lesions disappeared | 72
progressive improvement in inflammatory markers | 72
progressive improvement in pain | 72
progressive tolerance to rehabilitation exercises | 72
no adverse events | 72
antimicrobial treatment ended | 168
conservative treatment for heterotopic calcification | 168
nonsteroidal anti-inflammatory drugs | 168
physical therapy | 168
improvement of hip pain | 168
complete return to work | 336
asymptomatic | 336
inflammatory markers negative | 336
magnetic resonance imaging of the lumbar spine | 336
healing of the spondylodiscitis | 336
follow-up | 720