38 years old | 0
female | 0
type 2 diabetes mellitus | -8760
treated with sulfonylurea | -8760
abdominal pain | 0
polyuria | 0
polydipsia | 0
nausea | 0
vomiting | 0
blood pressure 93/53 mmHg | 0
pulse 119 beats/min | 0
respiratory rate 28 breaths/min | 0
oxygen saturation 99% | 0
temperature 97.8F | 0
Kussmaul breathing | 0
normal cardiopulmonary auscultation | 0
soft non-tender abdomen | 0
fully alert and oriented | 0
blood pH 6.98 | 0
serum bicarbonate 5mmol/L | 0
serum anion gap 22 | 0
serum glucose level 506mg/dL | 0
urinalysis positive for ketones | 0
urine pregnancy testing negative | 0
subtle prominence of the interstitial markings | 0
multiple ill-defined nodular opacities | 0
intravenous crystalloid | 0
insulin infusion | 0
blood cultures collected | 0
admitted to the intensive care unit | 0
progressively more hypoxemic | 2
dyspneic | 2
temperature rose to 104F | 2
level of consciousness declined to obtundation | 2
diffuse crackles | 2
endotracheally intubated | 2
hypoxemic respiratory failure | 2
volume assist-control ventilation | 2
diffuse bilateral opacities | 2
fraction of inspired oxygen 70% | 2
PaO2 59 mmHg | 2
PaO2/FiO2 ratio 84 | 2
lung-protective ventilation | 2
vancomycin | 2
piperacillin/tazobactam | 2
gram negative bacilli | 4
piperacillin/tazobactam switched to imipenem | 4
hemodynamics deteriorated | 6
high-dose norepinephrine infusion | 6
vasopressin | 6
FiO2 requirement rose to 100% | 72
PEEP increased to 15 cmH2O | 72
inhaled nitric oxide therapy | 72
oxygen saturation >90% | 72
pan-sensitive Klebsiella pneumoniae | 72
antibiotic coverage narrowed to ceftriaxone | 72
abdominal ultrasonography | 72
complex avascular hepatic mass-like lesion | 72
interventional radiology | 72
bedside placement of a drainage catheter | 72
pulseless electrical activity | 72
cardiopulmonary resuscitation | 72
resuscitative efforts aborted | 72
expired | 72
liver abscess | 72
extensive necrosis | 72
lung sections demonstrated diffuse abscess formation | 72
hyaline membranes | 72
diffuse alveolar damage | 72
invasive KLA syndrome | 72
ARDS | 2