27 years old | 0  
    male | 0  
    admitted to the hospital | 0  
    ulcerative colitis | -4032  
    primary sclerosing cholangitis | -4032  
    total abdominal colectomy | -4032  
    end-ileostomy | -4032  
    abdominal pain | 0  
    high ileostomy output | 0  
    9-kg weight loss over the last 7 days | -168  
    previous small bowel obstruction | -672  
    high ileostomy output in prior admissions | -672  
    prior medical management | -672  
    resolved within a few days | -672  
    home medications pantoprazole 40 mg | 0  
    ursodiol 300 mg twice daily | 0  
    lorazepam 0.5 mg as needed | 0  
    occasional alcohol consumption | 0  
    no smoking history | 0  
    no illicit drug use | 0  
    tachycardia (170 beats/min) | 0  
    afebrile | 0  
    blood pressure 103/74 mm Hg | 0  
    CT abdomen with intravenous contrast | 0  
    dilated loops of bowel | 0  
    white blood cell count 5.4 K/uL | 0  
    alanine aminotransferase 446 unit/L | 0  
    aspartate aminotransferase 268 unit/L | 0  
    alkaline phosphatase 1034 unit/L | 0  
    lactate 3.32 mmol/L | 0  
    admitted to colorectal surgery ward | 0  
    nil per os status | 0  
    resuscitated with 1900 mL IVF | 0  
    lactated Ringer's solution | 0  
    nasogastric tube placement | 0  
    decompression | 0  
    supportive care of small bowel obstruction | 0  
    no parenteral nutrition | 0  
    upper endoscopy | 0  
    chronic active ileitis | 0  
    medications metoprolol tartrate 25 mg twice daily | 0  
    hydromorphone 0.2 mg every 4 h | 0  
    ondansetron 4 mg every 6 h | 0  
    acetaminophen 1000 mg every 8 h | 0  
    pantoprazole 40 mg | 0  
    tachycardia persisted (150-180 beats/min) | 24  
    ostomy output >5 L/day | 24  
    aggressive IVF resuscitation (7272 mL LR) | 24  
    fever (39.7°C) | 72  
    tachypnea (32 breaths/min) | 72  
    tachycardia (128 beats/min) | 72  
    leukopenia (3.89 K/uL) | 72  
    mild agitation | 72  
    worsening abdominal pain | 72  
    increased ileostomy output | 72  
    suspected sepsis | 72  
    systemic inflammatory response syndrome criteria met | 72  
    upgraded to ICU | 72  
    IVF resuscitation (6982 mL LR) | 72  
    broad spectrum antibiotics piperacillin-tazobactam | 72  
    peripherally inserted central catheter removal | 72  
    metoprolol tartrate 12.5 mg | 72  
    no parenteral nutrition | 72  
    repeated CT scans | 72  
    small bowel obstruction up to stoma | 72  
    normal blood workup | 72  
    normal blood lactate levels | 72  
    negative urine culture | 72  
    negative blood culture | 72  
    negative Clostridium difficile toxin assay | 72  
    unremarkable echocardiogram | 72  
    sinus tachycardia on ECG | 72  
    thyroid function testing | 72  
    thyroid-stimulating hormone <0.02 ulU/mL | 72  
    triiodothyronine 13.0 pg/mL | 72  
    tetraiodothyronine 22.4 ug/dL | 72  
    normal parathyroid hormone 9.6 pg/mL | 72  
    hyperthyroidism diagnosis | 72  
    thyroid storm diagnosis | 72  
    antibiotics stopped | 72  
    Endocrinology consult | 72  
    esmolol infusion | 72  
    propylthiouracil 150 mg every 6 h | 72  
    cholestyramine 4 mg twice daily | 72  
    hydrocortisone 50 mg every 8 h | 72  
    continuous IVF hydration (150 mL/h LR) | 72  
    acetaminophen 1000 mg as needed | 72  
    elevated thyroid-stimulating immunoglobulins | 72  
    Graves' disease diagnosis | 72  
    ileostomy output decreased (5175 mL to 2150 mL) | 168  
    fevers resolved | 168  
    discharged home | 408  
    propranolol 30 mg twice daily | 408  
    propylthiouracil 200 mg twice daily | 408  
    prednisone 10 mg | 408  

