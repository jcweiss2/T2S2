42 years old | 0
woman | 0
relapsing-remitting multiple sclerosis (diagnosed) | -144000
McDonald criteria | -144000
methotrexate (treatment) | -17520
methotrexate discontinued | -17520
elevated liver enzymes | -17520
interferon beta 1-a (treatment) | -113520
interferon beta 1-a discontinued | -113520
disease activity | -113520
fingolimod (treatment) | -35040
muscle aches | -72
gait difficulty | -72
sensory disturbances | -72
weakness on the right side | -72
major depression disorder | 0
hypothyroidism | 0
recurrent urinary tract infection | 0
pulmonary embolism | 0
direct oral anticoagulation | 0
myasthenia gravis (diagnosed) | -43800
thymectomy | -43800
expanded disability status scale (EDSS) score | 0
positive Babinski sign on the right side | 0
MRI moderate disease burden in the brain | 0
right-sided cervical cord lesions | 0
lymphocyte count 842.4/μL | 0
symptoms started on March 1, 2020 | -144
symptoms gradually worsened over the next few days | -144
sought medical attention on March 5 | -96
outpatient MS clinic visit | -96
neurologic examination decreased sensation | -96
reduced muscle strength (4/5) | -96
brisk reflexes | -96
right positive Babinski sign | -96
EDSS 4 | -96
new relapse or recrudescence of old symptoms (pseudoexacerbation) | -96
admitted for relapse workup and treatment | -96
afebrile | 0
vital signs within normal limits | 0
C-reactive protein 76 mg/L | 0
erythrocyte sedimentation rate 46 mm | 0
suspected infectious etiology | 0
decrease in absolute lymphocyte count (601.6/μL) | 0
methylprednisolone IV 1,000 mg/d initiated | 0
chest X-ray ground glass opacity | 0
community-acquired pneumonia | 0
azithromycin 500 mg daily initiated | 0
allergy to fluoroquinolones | 0
dry cough | 48
dyspnea | 48
fever 38.7°C | 48
tachycardia 122 | 48
increased respiratory rate 30 | 48
blood pressure 100/70 mm Hg | 48
oxygen saturation 89% | 48
lymphocyte count 440.8/μL | 48
fingolimod discontinued | 48
ceftriaxone 1 g twice daily initiated | 48
oxygen via nasal cannula initiated | 48
chest CT performed | 48
ground glass opacities on CT | 48
suspected COVID-19 | 48
nasopharyngeal swab for PCR testing | 48
transferred to COVID ward | 48
hydroxychloroquine initiated | 48
oseltamivir initiated | 48
piperacillin/tazobactam initiated | 48
ceftriaxone discontinued | 48
azithromycin discontinued | 48
felt well on March 11 | 216
vital signs stabilized | 216
afebrile | 216
lymphocyte count 510.3/μL | 216
COVID-19 test positive | 216
all medications except hydroxychloroquine discontinued | 216
cough improved | 216
dyspnea improved | 216
neurologic symptoms improved | 216
discharged after 13-day admission | 312
glatiramer acetate initiated | 312
lymphocyte count 1,000.5/μL | 312
self-quarantined at home | 696
no respiratory symptoms | 696
no neurologic symptoms | 696
hemodynamic instability | 0
unclear neurologic symptoms etiology | 0
E.g., relapsing-remitting MS diagnosed | -144000 → should be -166440
relapsing-remitting multiple sclerosis (diagnosed) | -166440
McDonald criteria | -166440
muscle aches | -96
gait difficulty | -96
sensory disturbances | -96
weakness on the right side | -96
myasthenia gravis (diagnosed) | -210240
thymectomy | -210240
expanded disability status scale (EDSS) score | -4320
positive Babinski sign on the right side | -4320
MRI moderate disease burden in the brain | -4320
right-sided cervical cord lesions | -4320
lymphocyte count 842.4/μL | -4320
symptoms started on March 1, 2020 | -96
symptoms gradually worsened over the next few days | -96
sought medical attention on March 5 | 0
outpatient MS clinic visit | 0
neurologic examination decreased sensation | 0
reduced muscle strength (4/5) | 0
brisk reflexes | 0
right positive Babinski sign |
