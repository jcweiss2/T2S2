22 years old | 0
male | 0
admitted to the hospital | 0
one-day history of sudden onset fevers | -24
headache | -24
generalized myalgia | -24
several days of non-productive cough | -72
denied photophobia | 0
denied neck stiffness | 0
denied urinary symptoms | 0
denied bowel symptoms | 0
reported to be recently well before presentation | 0
Q fever | 0
febrile | 0
tachycardic | 0
no increased work of breathing | 0
chest clear on auscultation | 0
abdomen soft | 0
abdomen non-tender | 0
rest of examination unremarkable | 0
no localizing sign of infection | 0
deteriorated overnight | 0
progressive onset of severe epigastric pain | 0
vomiting | 0
persisting fevers | 0
generalized tenderness across the epigastrium | 0
developed septic shock | 0
urgently transferred to intensive care unit | 0
noradrenaline infusion commenced | 0
intravenous piperacillin-tazobactam commenced | 0
blood tests revealed ischaemic hepatitis | 0
acute kidney injury | 0
disseminated intravascular coagulopathy (DIC) | 0
screening for hepatitis B negative | 0
screening for hepatitis C negative | 0
screening for HIV negative | 0
lumbar puncture not performed | 0
abdominal ultrasound did not demonstrate any pathology | 0
contrast enhanced CT abdomen/pelvis did not demonstrate any pathology | 0
blood culture revealed N. meningitidis | 72
seven-day course of intravenous benzylpenicillin completed | 0
clinically improved | 240
discharged from hospital | 240
represented to hospital 4 days later | 384
mild intermittent left upper quadrant abdominal pain | 384
otherwise systemically well | 384
left upper quadrant tender on palpation | 384
remaining examination unremarkable | 384
haemodynamically stable | 384
spleen grossly abnormal on abdominal ultrasound | 384
significant fluid replacement of the normal splenic tissue | 384
splenic necrosis | 384
CT abdomen/pelvis reported extensive splenic necrosis | 384
associated abscess formation | 384
no normal splenic tissue on imaging | 384
associated vessels of normal appearance | 384
no evidence of thrombus | 384
excluded splenic artery aneurysm | 384
percutaneous drainage of the splenic abscess | 384
8 French percutaneous catheter inserted | 384
550 ml of thick altered blood drained | 384
no growth from collection | 384
recovered well from the procedure | 384
discharged 3 days later | 408
post-splenectomy vaccines | 408
antibiotics prophylaxis | 408
no free fluid inside the abdominal cavity | 384
no splenic artery aneurysm | 384
no residual enhancing splenic tissue | 384
