32 years old | 0
woman | 0
diagnosed with lymphangioleiomyomatosis | 0
placed on organ transplant waiting list | -4320
rapidly progressing respiratory insufficiency | -4320
multiple lymphangioleiomyomas in retroperitonium | 0
repeated spontaneous pneumothoraces | 0
required drainage | 0
transesophageal echocardiography performed | 0
low ejection fraction | 0
intubated | -3744
ventilated | -3744
respiratory failure | -3744
developed bronchopneumonia | -3744
multiresistant Pseudomonas aeruginosa | -3744
sepsis | -3744
disseminated intravascular coagulopathy | -3744
severe bleeding from nose | -3744
severe bleeding from hypopharynx | -3744
severe bleeding from lower respiratory tract | -3744
mechanical ventilation insufficient | -3744
venovenous ECMO commenced | -3744
bridge to urgent lung transplantation | -3744
donor found | -288
sequential bilateral lung transplant performed | -288
clamshell incision | -288
arteriovenous ECMO support | -288
cannulae from VV-ECMO left in place | -288
arterial cannula inserted into ascending aorta | -288
cannulation of vena jugularis interna dextra terminated | -288
donor lungs partially resected | -288
perioperative TEE | -288
severely hypokinetic right ventricle | -288
severely hypokinetic left ventricle | -288
large thrombus in left atrium | -288
diffuse bleeding | -288
coagulopathy | -288
10 L blood loss | -288
AV=ECMO left in place | -288
poor myocardial function | -288
sternotomy not closed | -288
arterial cannula remained in aorta | -288
severe pulmonary edema | 0
continuous leakage of edematous fluid from endotracheal tube | 0
tidal volumes 30-40 mL | 0
peak pressure 30 cm H2O | 0
positive end-expiratory pressure 10 cm H2O | 0
cardiovascular support with high-dose norepinephrine | 0
arterial blood gas results showed good oxygenation | 0
immunosuppression therapy commenced | 0
tacrolimus | 0
mycophenolate mofetil | 0
corticosteroids | 0
anticoagulation with heparin initiated | 0
target ACT 150-200 seconds | 0
TEE performed | 6
thrombi in left atrium | 6
thrombi in right atrium | 6
high risk of embolism | 6
crucial decision made | 6
thrombolysis initiated | 6
contraindicated in immediate postoperative period | 6
risk of massive embolism superior to bleeding risk | 6
primary thrombolysis with 25 mg alteplase | 6
alteplase given over 2 hours into pulmonary artery | 6
left atrial thrombus reduced | 8
second identical dose of alteplase given | 8
pulmonary edema resolved | 8
TEE showed no thrombi in left ventricle | 8
TEE showed no thrombi in pulmonary veins | 8
small thrombi remained in right atrium | 8
small thrombi remained in left atrium | 8
full dose thrombolytic agent given | 24
50 mg alteplase over 2 hours intravenously | 24
no further thrombi detected | 24
lung function improved | 168
radiological findings improved | 168
acute kidney injury | 168
continuous renal replacement therapy | 168
heart function improved | 192
lung function improved | 192
ECMO support stopped | 192
sternotomy closed | 192
resolution of P. aeruginosa infection | 192
weaning complicated by poor muscle strength | 192
rehabilitation complicated by poor muscle strength | 192
worsening lung function | 192
transbronchial biopsy performed | 192
tissue rejection A1-2 confirmed | 192
pulses of steroids | 192
loss of consciousness | 240
posterior reversible encephalopathy syndrome | 240
epileptic status | 240
antiepileptic medications prescribed | 240
stenosis of right main bronchus diagnosed | 2160
biodegradable stent implanted | 2160
pulmogenic sepsis | 4320
multiorgan failure | 4320
continuous renal replacement therapy needed | 4320
extubated | 4320
actively rehabilitated | 4320
discharged | 5040
good quality of life | 5040
no signs of stenosis of upper respiratory tract | 5040
stationary spirometric values | 5040
last FEV1 38% | 5040
