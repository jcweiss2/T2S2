42 years old | 0
Thai female | 0
motorcycle accident | 0
left knee pain | 0
drowsiness | 0
taken to emergency room | 0
ATLS examination | 0
life-threatening condition | 0
subdural hematoma | 0
right parietal lobe | 0
physical examination | 0
multiple shallow abrasion wounds | 0
left proximal tibia | 0
pain at lateral tibial plateau | 0
limited range of left knee motion | 0
anteroposterior radiographic images | 0
lateral radiographic images | 0
combined tibial plateau fracture | 0
tibial tubercle avulsion | 0
immobilized with long leg slab | 0
white blood cell count 19,490 /μL | 0
hematocrit 26.7% | 0
hemoglobin 8.6 g/dL | 0
polymorphonuclear neutrophils 85.5% | 0
lymphocytes 6.0% | 0
eosinophils 0.2% | 0
monocytes 8.2% | 0
platelets 336,000/μL | 0
afebrile | 0
admitted to intensive care unit | 0
close clinical observation | 0
no signs of wound infection | 0
regained full consciousness | 120
open reduction and internal fixation | 120
locking plate | 120
fracture site | 120
small amount of cloudy fluid | 120
gram stain | 120
culture | 120
Staphylococcus aureus | 120
intravenous ceftriaxone | 120
intravenous clindamycin | 120
fever | 168
redness around surgical wound | 168
investigated for sepsis | 168
chest radiograph no infiltration | 168
urine sample clear | 168
erythrocyte sedimentation rate >140 mm/h | 168
CRP >19.2 mg/dL | 168
irrigation and debridement | 192
necrotic tissue removed | 192
infected site copiously irrigated | 192
necrotic tissue culture Staphylococcus aureus | 192
hemoculture negative | 192
continued intravenous ceftriaxone | 192
continued intravenous clindamycin | 192
switched to oral Augmentin | 408
clinical condition improved | 408
complete course of Augmentin | 696
inflammatory markers disappeared | 696
able to walk without aid | 2880
plain radiograph showed union | 2880
4-month follow-up | 2880
