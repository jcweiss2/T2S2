33 years old | 0
    African American female | 0
    recurrent progressive metastatic squamous cell carcinoma cervical cancer | -672
    FIGO Stage IIB | -672
    external pelvic chemoradiation | -672
    chemotherapy weekly with cisplatin | -672
    intracavitary high-dose rate brachytherapy | -672
    recurrent disease in upper abdomen | -672
    recurrent disease in iliac bone | -672
    multiple admissions during prior cytotoxic chemotherapy | -672
    sepsis | -672
    pancreatitis | -672
    small bowel resection | -672
    permanent ostomy formation | -672
    single agent pembrolizumab | -672
    painful hyperpigmented maculopapular rash | -72
    blister-like lesions on lower back | -72
    blister-like lesions on feet | -72
    maculopapular rash evolved to forehead | -72
    maculopapular rash evolved to trunk | -72
    maculopapular rash evolved to thighs | -72
    painful blistering of lips | -72
    ocular involvement | -72
    biopsy confirmed SJS/TEN | -72
    apoptotic keratinocytes | -72
    lymphocytic infiltration involving dermis | -72
    transfer to University Burn Intensive Care Unit | 0
    IV antibiotic administration | 0
    complicated urosepsis | 0
    daptomycin | 0
    meropenem | 0
    started on pembrolizumab two weeks prior | -336
    moderate distress | 0
    15% BSA desquamative rash on buttocks | 0
    desquamative rash on sub mammary | 0
    desquamative rash on pressure areas | 0
    rash extending to upper extremities | 0
    rash extending to lower extremities | 0
    increasing odynophagia | 0
    worsening mouth ulcers | 0
    presumptive diagnosis of SJS/TEN due to meropenem | 0
    possible recent immunotherapy | 0
    meropenem held | 0
    pembrolizumab held | 0
    high-dose patient-controlled analgesics | 0
    Staphylococcus epidermidis sepsis | 0
    IV vancomycin 1500 mg every twelve hours | 0
    solumedrol 125 mg every 24 hours | 0
    improvement in cutaneous symptoms | 0
    dermatology consultation | 0
    ophthalmology consultation | 0
    burn consultation | 0
    gynecologic oncology consultation | 0
    wound care | 0
    prophylactic antibiotics | 0
    pain management | 0
    nutritional management | 0
    topical antibiotic ointment | 0
    cyclosporine 5 mg/kg/day twice a day | 0
    no ocular involvement | 0
    artificial tears 4–6 times per day | 0
    erythromycin ointment in both eyes | 0
    silverlon dressing | 0
    dampened 10-ply gauze | 0
    burn net | 0
    gauze changes daily | 0
    aggressive nutritional supplementation with protein | 0
    micronutrient supplementation with vitamin C | 0
    weekly nutrition labs | 0
    benign gynecology consultation | 0
    vulvovaginal involvement | 0
    intravaginal betamethasone therapy | 0
    estrogen therapy | 0
    gynecologic oncology consultation | 0
    pembrolizumab given four weeks prior | -672
    grade 4 immune-related dermatologic SJS/TEN-like reaction | 0
    cyclosporine discontinued | 0
    prednisone 1.5 mg/kg/day | 0
    symptom improvement | 24
    corticosteroid tapered to 1.25 mg/kg/day | 24
    discharge planned to inpatient rehab | 24
    insurance lapse | 24
    remained inpatient | 24
    extensive skin lesions | 24
    episode of fever | 48
    hypotension | 48
    empiric meropenem | 48
    empiric vancomycin | 48
    blood cultures grew Klebsiella | 48
    discharged to home | 72
    ciprofloxacin | 72
    remaining Prednisone steroid taper | 72