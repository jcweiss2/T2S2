44 years old|0
male|0
left flank pain| -120
abdominal pain| -120
painful ejaculation| -120
left flank pain radiating into left lower abdomen| -120
left flank pain radiating into left testicle| -120
achy to sharp pain| -120
nausea| -120
vomiting| -120
decreased appetite| -120
subjective fever| -120
chills| -120
utilization of prostate vibrator| -168
emergency department arrival|0
temperature 101.2 °F|0
blood pressure 92/54 mmHg|0
respiratory rate 21 breaths/min|0
weight 94.5 kg|0
SpO2 98%|0
distress due to pain|0
diaphoresis|0
ill appearance|0
dry oral mucosa|0
sinus tachycardia|0
no murmur|0
clear lungs bilaterally|0
left costovertebral angle tenderness|0
left upper abdominal tenderness|0
left lower abdominal tenderness|0
voluntary guarding|0
left inguinal canal tenderness|0
left epididymitis|0
no abscess|0
no cellulitis|0
no crepitus|0
sepsis protocol initiation|0
two peripheral IVs placed|0
urine cultures taken|0
blood cultures taken|0
laboratory evaluation started|0
fluid resuscitation with 30 mL/kg IV bolus|0
leukocytosis 18.2|0
neutrophil predominance|0
hemoglobin 11.6|0
platelet 220 bil/L|0
pre5-renal azotemia|0
BUN 27 mg/dL|0
creatinine 1.3 mg/dL|0
blood glucose 130|0
unremarkable hepatic function panel|0
lactic acid 3.2|0
lactic acid 1.5|0
urinalysis 2+ blood|0
+nitrites|0
3+ leukocyte esterase|0
>50 WBCs|0
3+ bacteria|0
25–50 RBCs|0
C-reactive protein 7.1|0
unremarkable laboratory evaluation|0
immunocompromised state due to HIV|0
high-risk sexual behavior|0
recent prostate manipulation|0
concern for acute bacterial prostatitis|0
ceftriaxone started|0
gentamicin started|0
ultrasound scrotum with Doppler|0
prominent epididymis with increased vascularity|0
small left hydrocele|0
scattered internal debris|0
no compromised arterial flow|0
no abscess formation|0
left hydrocele|0
CT abdomen/pelvis without contrast|0
left-sided peri-ureteral fat stranding|0
prominent left seminal vesicle|0
infiltrative fat stranding around left hemi-pelvis|0
multiple prominent pelvic lymph nodes up to 8.1 mm|0
prominent inguinal lymph nodes up to 6.5 mm|0
prostate size 5 cm|0
inflammatory changes within left hemi-pelvis|0
prominence of left seminal vesicle|0
prostatitis|0
peri-ureteral fat stranding reactive to prostatitis|0
hypotensive after fluid resuscitation|0
MAP <65|0
central venous catheter placement|0
inotropic medication initiation|0
intensive care unit admission|0
Escherichia coli in urine cultures|0
Escherichia coli in blood cultures|0
pansusceptible Escherichia coli|0
negative Chlamydia trachomatis|0
negative Neisseria gonorrhoeae|0
off inotropic medication by Day3|72
hemodynamically stable by Day3|72
tolerating regular diet by Day3|72
30 days antibiotics needed|72
discharged by Day4|96
cefuroxime at discharge|96
1-month follow-up|720
progressing well at follow-up|720
denies complaints at follow-up|720
