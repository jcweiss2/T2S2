15 years old | 0 | 0 
female | 0 | 0 
acute myelogenous leukemia | 0 | 0 
standard induction treatment | -672 | -336 
chemotherapy | -672 | -336 
pancytopenia | -336 | 0 
broad anti-infective treatment | -336 | 0 
ciprofloxacin | -336 | 0 
linezolid | -336 | 0 
meropenem | -336 | 0 
tobramycin | -336 | 0 
liposomal amphotericin | -336 | 0 
tachycardia | -24 | 0 
hypotension | -24 | 0 
lactic acidosis | -24 | 0 
admitted to the pediatric intensive care unit | 0 | 0 
severely impaired left ventricular ejection fraction | 0 | 0 
sinus tachycardia | 0 | 0 
incomplete right bundle branch block | 0 | 0 
elevated NT-proBNP | 0 | 0 
elevated high-sensitive troponin T | 0 | 0 
fluid therapy | 0 | 0 
noradrenaline | 0 | 0 
dobutamine | 0 | 0 
milrinone | 0 | 0 
deep sedation | 0 | 0 
mechanical ventilation | 0 | 0 
respiratory insufficiency | 0 | 0 
va-ECMO | 0 | 168 
cannulation of the left femoral artery and vein | 0 | 0 
arterial cannula | 0 | 0 
venous cannula | 0 | 0 
distal leg perfusion | 0 | 0 
sheath | 0 | 0 
Cardiohelp System | 0 | 168 
extracorporeal blood flow | 0 | 168 
mean arterial pressure | 0 | 168 
noradrenaline | 0 | 168 
vasopressin | 0 | 168 
levosimendan | 0 | 21 
hydrocortisone | 0 | 168 
continuous venovenous hemodiafiltration | 0 | 168 
anti-infective therapy | 0 | 168 
meropenem | 0 | 168 
ciprofloxacin | 0 | 168 
metronidazole | 0 | 168 
cotrimoxazole | 0 | 168 
liposomal amphotericin B | 0 | 168 
acyclovir | 0 | 168 
vancomycin | 0 | 168 
procalcitonin | 0 | 168 
C-reactive protein | 0 | 168 
decline of mean arterial blood pressure | 24 | 24 
increasing doses of vasopressors | 24 | 24 
decrease of LVEF | 24 | 24 
stop of levosimendan infusion | 24 | 24 
acute ischemic injury of the non-cannulated leg | 24 | 24 
dissection of the right femoral artery | 24 | 24 
insufficient blood inflow | 24 | 24 
Dacron conduit | 24 | 24 
second arterial cannula | 24 | 24 
Y-connector | 24 | 24 
enhancement of ECBF | 24 | 168 
maintenance of MAP | 24 | 168 
broad-complex tachycardia | 48 | 48 
esmolol | 48 | 48 
metoprolol | 48 | 48 
decrease of left ventricular function | 48 | 48 
aortic valve ceased to open | 48 | 48 
second venous cannula | 48 | 48 
percutaneous atrioseptostomy | 48 | 48 
left atrial venting | 48 | 168 
increase of ECBF | 48 | 168 
reduction of venous drainage pressures | 48 | 168 
cerebral oximetry | 48 | 168 
regional oxygen saturation | 48 | 168 
unfractionated heparin | 48 | 168 
peak of procalcitonin | 72 | 72 
peak of C-reactive protein | 72 | 72 
leukocytes | 72 | 72 
high-sensitive troponin T | 72 | 72 
creatine kinase MB | 72 | 72 
total creatine kinase | 72 | 72 
recovery of cardiac systolic function | 120 | 168 
removal of ECMO cannulas | 120 | 120 
removal of ECMO | 168 | 168 
recovery of LVEF | 168 | 168 
normal renal function | 168 | 168 
stop of CVVHDF | 168 | 168 
respirator weaning | 792 | 792 
allogenic stem cell transplantation | 1008 | 1008 
discharge to rehabilitation facility | 2160 | 2160 
severe critical illness | 2160 | 2160 
polyneuropathy | 2160 | 2160 
recovery of LVEF | 2160 | 2160 
ventricular dilatation | 2160 | 2160