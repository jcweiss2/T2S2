31 years old | 0
male | 0
black | 0
admitted to the ED | 0
complaining of open sores | 0
open sores covering his body | 0
cigarette burn to his left forearm | -336
sores began at the site of a cigarette burn | -336
sores spread diffusely over the body | -336
lesions were slightly tender to the touch | 0
review of systems was negative for a viral prodrome | 0
denied any fevers | 0
denied any chills | 0
denied any sweats | 0
denied any chest pain | 0
denied any shortness of breath | 0
no abdominal pain | 0
no nausea | 0
no vomiting | 0
no history of ill contacts | 0
no animal exposure | 0
no insect bites | 0
no recent travel | 0
denied intravenous drug use | 0
chronic use of tobacco | 0
chronic use of alcohol | 0
chronic use of marijuana | 0
not been taking any medications | 0
denied any known allergies | 0
denied any significant family history | 0
anxious | 0
avoided unnecessary movement | 0
temperature was 100.1°F | 0
heart rate was 145 beats per minute | 0
blood pressure 124/77 mm Hg | 0
respiratory rate 20 breaths per minute | 0
oxygen saturation 99% on room air | 0
heart tones were regularly tachycardic | 0
pulmonary exam was clear | 0
no edema of the extremities | 0
no lymphadenopathy | 0
no hepatosplenomegaly | 0
skin exam revealed diffuse regions of skin sloughing | 0
skin sloughing with necrosis | 0
mildly erythematous base along the dermis | 0
occasional small bullae | 0
occasional small vesicles | 0
over 50% of the patient’s total body surface area was involved | 0
back was involved | 0
abdomen was involved | 0
scrotum was involved | 0
perirectal area was involved | 0
forehead was spared | 0
scalp was spared | 0
no purulent discharge | 0
no pustules | 0
no purpura | 0
no ulcerations | 0
strong foul-smelling odor | 0
non-affected area of the patient’s skin easily sloughed | 0
oral mucosa was injected | 0
oral mucosa was sloughing | 0
conjunctivae were spared | 0
temperature increased to 101.7° F | 2
vancomycin was administered | 2
meropenem was administered | 2
blood cultures were sent | 2
received four liters intravenous normal saline | 2
morphine was administered | 2
white blood cell count of 12,000/mm | 2
lactic acid of 2.8 mmol/L | 2
serum bicarbonate 21 mmol/L | 2
serum glucose 140 mg/dL | 2
blood urea nitrogen 9 mg/dL | 2
creatinine 0.9 mg/dL | 2
anion gap 10 mmol/L | 2
severe sepsis developed | 24
blood cultures returned positive for oxacillin-sensitive Staphylococcal aureus | 24
steroids were administered | 24
intravenous immunoglobulin was administered | 24
multiple surgical debridement procedures | 48
skin biopsy revealed non-specific epidermal necrosis | 48
discharged home | 168
over-the-counter NSAID use | -168
admitted to the intensive care unit | 2
cared for in the Burn Care Unit | 24
septicemia | 24
secondary bacterial infection of the necrotic tissue | 24