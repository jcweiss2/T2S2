84 years old | 0
male | 0
emergency surgical consultation | 0
sudden lower abdominal discomfort | 0
lower abdominal pain | 0
chronic constipation | -87600
chronic heart failure | 0
atrial fibrillation | 0
generalized abdominal tenderness | 0
lower quadrants tenderness | 0
insignificant rebound tenderness | 0
hypogastric region tenderness | 0
loose bloody stool | 0
rectal perforation | 0
barium extravasation | 0
exploratory laparotomy | 24
midline incision | 24
no visible perforation in distal colon | 24
no visible perforation in sigmoid | 24
no visible perforation in upper rectum | 24
barium drops on posterior wall of peritoneum | 24
barium around sigmoid mesocolon | 24
barium around mesoileum | 24
barium penetration from retroperitoneum into intraperitoneal cavity | 24
extraction of barium drops | 24
massive irrigation | 24
peritoneal cavity lavage | 24
diverting ileostomy | 24
tissue sample taken from mesenteric tissue | 24
fat necrosis | 24
foreign-body reaction | 24
transfer to intensive care unit | 24
broad-spectrum intravenous antibiotics | 24
sepsis | 72
rigid proctoscopy | 72
massive inflammation on posterior wall of rectum | 72
blood clots on posterior wall of rectum | 72
open presacral drain | 72
generalized abdominal pain | 336
high fever | 336
abdominopelvic computed tomography scan | 336
hyperdense area in retroperitoneal space | 336
extension to psoas muscles | 336
second laparotomy | 336
barium dissemination up to inferior pole of kidneys | 336
mesentery covered by barium | 336
retroperitoneal tissues fragile and inflamed | 336
irrigation | 336
debridement of necrotic tissues | 336
two open corrugated drains | 336
fever disappeared | 504
regained appetite | 504
presacral drain removed | 504
abdominal drain removed | 504
oral diet | 504
discharged | 840
ileostomy closure | 2400
monthly visits | 2400
bimonthly visits | 2400
residual barium in retroperitoneal space | 17520
