36 years old | 0
male | 0
hypertension | -8760
systemic lupus erythematosus | -8760
coronary artery disease | -8760
seizure disorder | -8760
superior vena cava syndrome | -8760
end-stage renal disease | -8760
hemodialysis | -8760
dialysis catheter placements | -8760
sepsis | -720
disseminated intravascular coagulation | -720
bacteremia | -720
vancomycin-resistant Enterococcus | -720
extended-spectrum beta-lactamase–producing Klebsiella | -720
cefepime | -720
linezolid | -720
syncopal episode | -24
complete heart block | -24
junctional escape rhythm | -24
mildly sclerosed mitral and aortic valves | -24
mild-to-moderate mitral and tricuspid regurgitation | -24
normal LV function | -24
no regional wall motion abnormalities | -24
attempt to implant Micra leadless pacemaker | -12
vascular access unfeasible | -12
common iliac veins completely occluded | -12
superior vena cava chronically occluded | -12
transhepatic approach | -12
epicardial pacing | -12
surgical epicardial pacing | -6
left anterolateral minithoracotomy | -6
screw-in unipolar epicardial leads | -6
no capture | -6
frailty of the myocardium | -6
suture-on bipolar lead | -6
capturing in the operating room | -6
acceptable thresholds | -6
failure to capture | 0
WiSE-CRT system | 0
expedited plea to FDA | 0
institutional review board approval | 0
transmitter and battery implantations | 2
electrode insertion | 4
heparinization | 4
activated coagulation time | 4
retrograde access | 4
aortic valve | 4
lateral wall of the LV | 4
receiver electrode | 4
endocardiac pacing | 4
heparin reversal | 6
protamine | 6
arterial access closure | 6
Perclose ProGlide | 6
LV pacing | 6
appropriate capture | 6
sepsis | 336
intra-abdominal infection | 336
death | 336