31 years old | 0
female | 0
non-smoking | 0
Caucasian | 0
admitted to the hospital | 0
sudden-onset severe headache | -840
left arm numbness | -840
cranial computed tomography (CT) scan | -840
grade 2 SAH | -840
ruptured right middle cerebral artery aneurysm | -840
percutaneous endovascular coil embolization | -840
fever | -672
chills | -672
constant abdominal pain | -672
purulent uterine discharge | -672
sepsis | -672
septic shock | -672
transferred to the intensive care unit | -672
body temperature 38.3 °C | -672
invasive blood pressure 90/65 mmHg | -672
heart rate 135/min | -672
arterial oxygen saturation 82 % | -672
mild disorientation | -672
slower capillary refill | -672
coarse rales | -672
sequential organ failure assessment (SOFA) score 4 | -672
hemoglobin 6.8 g/dL | -672
d-dimers 4.58 μg/mL | -672
C-reactive protein 322 mg/L | -672
fibrinogen concentration 6.4 mL | -672
blood culture showed E. coli | -672
piperacillin/tazobactam | -672
vancomycin | -672
azithromycin | -672
chest radiography | -672
pulmonary nodules | -672
transvaginal ultrasound | -672
enlarged uterus | -672
complete loss of zonal anatomy | -672
abdominal magnetic resonance imaging (MRI) | -672
splenic metastatic lesion | -672
serum β-human chorionic gonadotrophin (β-hCG) 232,085 mUI/mL | -672
suction evacuation and curettage | -672
pathology report confirmed choriocarcinoma | -672
International Federation of Gynecology and Obstetrics (FIGO) modified WHO prognostic scoring system | -672
total score of 12 | -672
high risk of developing resistance to single-drug chemotherapy | -672
multiagent chemotherapy regimen | -24
low-dose etoposide | -24
cisplatin | -24
EMA/CO regimen | 0
etoposide | 0
methotrexate | 0
actinomycin D | 0
cyclophosphamide | 0
vincristine | 0
grade 3 neutropenia | 168
granulocyte colony stimulating factor (G-SCF) | 168
dose reduction of both etoposide and actinomycin D | 168
grade 2 alopecia | 168
grade 2 nausea | 168
dexamethasone | 168
ondansetron | 168
EP/EMA regimen | 336
grade 2 fatigue | 504
male condoms | 504
follow-up | 504
β-hCG levels plateaued | 504
restaging with MRI of the brain | 504
18F-fluorodeoxyglucose (FDG) positron emission tomography (PET)/CT scan | 504
decreased pulmonary nodules | 504
decreased uterine mass | 504
low standardized uptake value (SUV) | 504
revised FIGO score 7 | 504
therapeutic regimen changed | 504
normalization of β-hCG | 720
completion of three cycles | 720
disease-free for almost two years | 1008