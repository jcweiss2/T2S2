3 years old | 0
female | 0
Noonan syndrome | 0
heterozygous RIT1 mutation | 0
heart murmur | -12
HCM | -12
mid cavity left ventricular outflow tract obstruction | -12
severe right ventricular outflow tract obstruction | -12
dysplastic stenotic pulmonary valve | -12
surgical relief of LVOT obstruction | -10
myectomy | -10
relief of RVOT obstruction | -10
muscular resection | -10
transannular patch | -10
epicardial pacemaker | -10
post-operative complete heart block | -10
respiratory failure | -6
parainfluenza 3 infection | -6
bilateral pleural effusions | -6
pleural effusions drainage | -6
chylothorax | -6
low fat and high medium chain triglycerides diet | -6
octreotide infusion | -6
spontaneous bowel perforation | -5
terminal ileum resection | -5
stoma formation | -5
bacterial sepsis | -5
candida sepsis | -5
immunoglobulin replacements | -5
parenteral nutrition | -5
MCT diet | -3
discharged home | -3
reaccumulation of pleural effusions | 0
multiple chest drains | 0
pulmonary lymphangiectasia | 0
lymphatic dysplasia | 0
trametinib treatment | 0
severe eczema | 1
topical steroids | 1
stoma output increase | 1
parenteral nutrition | 1
reduction in left ventricular mass | 4
completion of 3-month trametinib course | 12
transition to enteral feeds | 12
discharged home | 12
no chylothorax recurrence | 20
stoma reversal | 20