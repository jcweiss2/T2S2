50 years old | 0
male | 0
admitted to the hospital | 0
fatigue | 0
mild splenomegaly | 0
pancytopenia | 0
poor reticulocyte response | 0
diagnosed with splenic marginal zone lymphoma | 0
splenic involvement | 0
bone marrow involvement | 0
remission | 0
relapse | -365
partial remission | -365
second line chemo-immunotherapy | -365
rituximab | -365
bendamustine | -365
supportive treatment | -365
intravenous immunoglobuline | -365
hypogammaglobulinemia | -365
second relapse | -120
third line chemo-immunotherapy | -120
rituximab-iphosphamide carboplatin and etoposide | -120
febrile neutropenia | -30
pneumonia | -30
bilateral ground-glass areas | -30
thorax computed tomography | -30
broad-spectrum antibiotherapy | -30
discharged | -14
admitted to the emergency room | 0
respiratory symptoms | 0
thoracic CT findings | 0
COVID-19 | 0
PCR result positive | 0
serum Na: 129 mmol/L | 0
CRP: 3.76 mg/dL | 0
D-dimer: 17.1 mg/L | 0
albumin: 3.4 g/dL | 0
sputum culture negative | 0
blood culture negative | 0
urine culture negative | 0
hydroxychloroquine | 0
oseltamivir | 0
favipiravir | 0
immune plasma therapy | 0
broad spectrum antibiotic treatments | 0
clinical condition partially improved | 30
PCR positivity continued | 30
hospitalized for 64 days | 64
PCR result negative | 60
discharged | 64
admitted to the emergency room again | 90
respiratory complaints | 90
fever | 90
consolidation | 90
ground-glass density | 90
thoracic CT | 90
PCR test positive | 90
serum Na: 135 mmol/L | 90
CRP: 12.7 mg/dL | 90
D-Dimer: 0.64 mg/L | 90
albumin: 3.2 g/dL | 90
Klebsiella pneumoniae | 90
sputum culture positive | 90
broad spectrum antibiotic treatments | 90
immune plasma therapy | 90
PCR negative | 95
radiological regression | 95
discharged | 106
monthly hematological intra venous immune globulin treatment | 106
admitted to the emergency room again | 120
diarrhea | 120
general condition disorder | 120
bilateral ground-glass areas | 120
CT scan | 120
PCR test positive | 120
serum Na: 130 mmol/L | 120
CRP: 7.59 mg/dL | 120
D-dimer: 0.52 mg/L | 120
albumin: 2.3 g/dL | 120
sputum culture negative | 120
blood culture negative | 120
urine culture negative | 120
metronidazole | 120
favipiravir | 120
prednol | 120
IVIG treatment | 120
COVID-19 PCR in stool positive | 125
high fever | 125
lobar pneumonia | 125
septic condition | 125
intensive care unit | 125
died | 161