25 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
housewife | 0 | 0 | Factual
given birth | -72 | -72 | Factual
baby girl | -72 | -72 | Factual
3.1-kg | -72 | -72 | Factual
37th week | -72 | -72 | Factual
first pregnancy | -72 | -72 | Factual
uncomplicated pregnancy | -72 | -72 | Factual
spontaneous vaginal delivery | -72 | -72 | Factual
episiotomy | -72 | -72 | Factual
severe pain | -24 | 0 | Factual
buttocks | -24 | 0 | Factual
shortness of breath | 0 | 0 | Factual
sudden onset | 0 | 0 | Factual
worsening pain | 0 | 0 | Factual
right thigh | 0 | 0 | Factual
drowsy | 0 | 0 | Factual
tachypneic | 0 | 0 | Factual
oxygen saturation | 0 | 0 | Factual
56% | 0 | 0 | Factual
high-flow oxygen supply | 0 | 0 | Factual
tachycardia | 0 | 0 | Factual
121 bpm | 0 | 0 | Factual
afebrile | 0 | 0 | Factual
36 °C | 0 | 0 | Factual
unrecordable blood pressure | 0 | 0 | Factual
hypotensive | 0 | 0 | Factual
56/30 mmHg | 0 | 0 | Factual
noradrenaline infusion | 0 | 0 | Factual
IV heparin | 0 | 0 | Factual
5000 units | 0 | 0 | Factual
IV amoxicillin-clavulanate | 0 | 0 | Factual
septicemic shock | 0 | 0 | Possible
pulmonary embolism | 0 | 0 | Possible
elective intubation | 0 | 0 | Factual
severe metabolic acidosis | 0 | 0 | Factual
lactic acidosis | 0 | 0 | Factual
worsening respiratory distress | 0 | 0 | Factual
120 mL/kg crystalloid | 0 | 0 | Factual
6 L | 0 | 0 | Factual
persistently hypotensive | 0 | 0 | Factual
adrenaline | 0 | 0 | Factual
vasopressin | 0 | 0 | Factual
dobutamine | 0 | 0 | Factual
grossly swollen right thigh | 0 | 0 | Factual
extensive blistering ecchymotic patches | 0 | 0 | Factual
right buttock | 0 | 0 | Factual
necrotizing fasciitis | 0 | 0 | Factual
septicemic shock | 0 | 0 | Factual
acute kidney injury | 0 | 0 | Factual
rhabdomyolysis | 0 | 0 | Factual
coagulopathy | 0 | 0 | Factual
thrombocytopenia | 0 | 0 | Factual
ischemic hepatitis | 0 | 0 | Factual
IV meropenem | 0 | 0 | Factual
IV clindamycin | 0 | 0 | Factual
IV vancomycin | 0 | 0 | Factual
high vaginal swab | 0 | 0 | Factual
culture and sensitivity | 0 | 0 | Factual
CT pulmonary angiography | 0 | 0 | Factual
small pulmonary embolism | 0 | 0 | Factual
bedside echocardiography | 0 | 0 | Factual
good contractility | 0 | 0 | Factual
heart chambers | 0 | 0 | Factual
not grossly dilated | 0 | 0 | Factual
intravenous immunoglobulin | 0 | 120 | Factual
toxin neutralization | 0 | 120 | Factual
5 days | 0 | 120 | Factual
continuous veno-venous hemofiltration | 0 | 0 | Factual
severe lactic acidosis | 0 | 0 | Factual
9.8-18 mmol/L | 0 | 0 | Factual
elevated creatinine kinase | 0 | 0 | Factual
29783 U/L | 0 | 0 | Factual
toxin removal | 0 | 0 | Factual
critical condition | 0 | 72 | Factual
4 inotropes | 0 | 72 | Factual
CVVH | 0 | 72 | Factual
skin lesion | 24 | 24 | Factual
bilateral upper and lower limbs | 24 | 24 | Factual
bluish discoloration | 24 | 24 | Factual
blistering | 24 | 24 | Factual
bilateral lower limbs | 24 | 24 | Factual
right lower abdomen | 24 | 24 | Factual
right upper limb | 24 | 24 | Factual
right elbow | 24 | 24 | Factual
Gram positive cocci | 24 | 24 | Factual
chains | 24 | 24 | Factual
S. pyogenes | 24 | 24 | Factual
group A beta hemolytic streptococcus | 24 | 24 | Factual
multidisciplinary discussion | 144 | 144 | Factual
day 6 | 144 | 144 | Factual
group A streptococcal toxic shock syndrome | 144 | 144 | Factual
necrotizing fasciitis | 144 | 144 | Factual
IV clindamycin | 144 | 168 | Factual
toxin suppression | 144 | 168 | Factual
IV crystalline penicillin G | 144 | 168 | Factual
every 4 hours | 144 | 168 | Factual
CVVH | 144 | 168 | Factual
toxin removal | 144 | 168 | Factual
surgical intervention | 144 | 168 | Factual
not feasible | 144 | 168 | Factual
skin biopsy | 144 | 168 | Factual
not performed | 144 | 168 | Factual
death | 168 | 168 | Factual
septic shock | 168 | 168 | Factual
tissue necrosis | 168 | 168 | Factual
toxic shock syndrome | 168 | 168 | Factual
S. pyogenes | 168 | 168 | Factual