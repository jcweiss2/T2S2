58 years old | 0
female | 0
metastatic melanoma | -504
nivolumab | -144
ipilimumab | -144
fever | -144
altered | 0
hypotensive | 0
tachycardic | 0
hypoxic | 0
peripheral edema | 0
elevated serum creatinine | 0
elevated alanine transaminase | 0
elevated aspartate transaminase | 0
elevated lactate | 0
elevated CRP | 0
mild leukocytosis | 0
pulmonary edema | 0
septic shock | 0
broad-spectrum antibiotics | 0
norepinephrine | 0
epinephrine | 0
vasopressin | 0
BiPAP | 0
methylprednisolone | 24
intubated | 24
tocilizumab | 48
IL-6 levels measured | 48
TNF-α levels measured | 48
etanercept | 72
symptoms improved | 96
extubated | 96
discharged | 168