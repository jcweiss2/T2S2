46 years old | 0
male | 0
HIV-positive | 0
admitted to the hospital | 0
shortness of breath | -144
cough | -144
pleuritic chest pain | -144
malaise | -144
diffuse joint pain | -144
intermittent fevers | -144
denies hemoptysis | -144
denies recent travel | -144
denies incarceration history | -144
denies homelessness | -144
worked as a farmer | -6720
coccidioidomycosis diagnosis | -336
fatigue | -336
fevers | -336
forearm lesions | -336
Coccidioides antibody IgG positive | -336
tachycardic | 0
tachypneic | 0
afebrile | 0
normotensive | 0
hypoxic | 0
coarse bilateral breath sounds | 0
labored breathing | 0
subcutaneous nodules | 0
no notable rashes | 0
no joint effusions | 0
no neurologic deficits | 0
cooperative | 0
alert | 0
oriented | 0
transitioned to non-invasive mechanical ventilation | 0
admitted to ICU | 0
acute hypoxemic respiratory failure | 0
severe sepsis | 0
CT scan of chest | 0
diffuse multifocal nodular consolidations | 0
ground glass opacities | 0
right upper lobe dense consolidations | 0
prominent mediastinal and hilar lymph nodes | 0
clear central airways | 0
no pulmonary embolism | 0
started on IV trimethoprim sulfamethoxazole | 0
started on IV cefepime | 0
started on oral fluconazole | 0
started on IV liposomal amphotericin B | 0
started on oral prednisone | 0
decompensated overnight | 12
required mechanical ventilation | 12
septic shock | 12
required norepinephrine | 12
blood cultures negative | 12
TB ruled out | 12
fungal studies negative for pneumocystis, cryptococcus, and toxoplasmosis | 12
coccidioidomycosis with titer levels of 1:64 in blood | 12
coccidioidomycosis with titer levels of 1:1 in CSF | 12
Infectious disease consulted | 12
antiretroviral therapy held | 12
declining mentation | 24
worsening respiratory status | 24
minimal response to proning | 24
intermittent severe metabolic acidosis | 24
renal failure | 24
improved with dialysis and bicarbonate drips | 24
CT scan of head | 24
corpus callosum mass | 24
features consistent with primary CNS lymphoma | 24
MRI of brain | 24
hemorrhagic mass | 24
surrounding edema | 24
high-grade glioma features | 24
echocardiogram | 24
right ventricular mobile mass | 24
started on IV flucytosine | 48
switched to IV fluconazole | 72
lack of clinical improvement | 120
decision to place on comfort care | 576
compassionately extubated | 576
expired | 576