70 years old | 0
    male | 0
    African-American | 0
    ESRD | 0
    IHD for 5 years | 0
    non-insulin-dependent diabetes mellitus | 0
    hypertension | 0
    severe peripheral arterial disease | 0
    recurrent vascular access thrombosis | 0
    symptomatic bradyarrhythmia | 0
    permanent implantable cardioverter-defibrillator (AICD) | 0
    upper half central veins significantly stenotic or occluded | 0
    right femoral last patent vein available for cannulation | 0
    home medications: aspirin | 0
    calcium acetate | 0
    carvedilol | 0
    cinacalcet | 0
    insulin | 0
    warfarin | 0
    gabapentin | 0
    simvastatin | 0
    esomeprazole | 0
    fever | -72
    headaches | -72
    chills | -72
    nausea | -72
    arrival to ED | 0
    temperature 105 Fahrenheit (40.50 Celsius) | 0
    blood pressure 108/51 mm Hg | 0
    heart rate 114 beats per minute | 0
    regular rhythm | 0
    respiratory rate 14 per minute | 0
    oxygen saturation 99% | 0
    alert | 0
    cooperative | 0
    oriented | 0
    no rash | 0
    no finger clubbing | 0
    lungs clear to auscultation | 0
    no erythema over AICD site | 0
    no tenderness over AICD site | 0
    no fluctuation over AICD site | 0
    cardiovascular exam: regular heart sounds | 0
    no gallop rhythm | 0
    grade 2/6 late diastolic murmur | 0
    right upper sternal border | 0
    no pericardial rub | 0
    no organomegaly | 0
    no peripheral edema | 0
    right femoral cuffed catheter minimal erythema | 0
    no warmth | 0
    no tenderness | 0
    no discharge over subcutaneous tunnel | 0
    no discharge over exit site | 0
    sodium 135 mmol/L | 0
    potassium 4.8 mmol/L | 0
    chloride 96 mmol/L | 0
    bicarbonate 23 mmol/L | 0
    blood urea nitrogen 68 mg/dL | 0
    creatinine 11.12 mg/dL | 0
    lactic acid 1.7 mmol/L | 0
    international normalized ratio 2.57 | 0
    white blood cells 10.8 k/mm3 | 0
    hemoglobin 8.6 gm/dL | 0
    hematocrit 25.5% | 0
    platelets 79 k/mm3 | 0
    empiric broad-spectrum antibiotics started | 0
    blood cultures sent | 0
    transfer to intensive care unit | 0
    CT scan of head unremarkable | 24
    chest x-ray unremarkable | 24
    CSF examination negative | 24
    blood cultures positive for MRSA | 24
    cuffed catheter tip culture negative | 24
    transthoracic echocardiogram echogenic tricuspid valve mass | 24
    trans-esophageal echocardiography confirmed tricuspid valve endocarditis | 24
    AICD pocket infection | 24
    antibiotics changed to ampicillin | 24
    vancomycin | 24
    cefepime | 24
    AICD removed | 24
    tunneled catheter exchanged over guidewire | 24
    new catheter at same femoral site | 24
    continued fever | 48
    blood cultures persistently positive for MRSA | 48
    exchange cuffed catheter with temporary non-cuffed catheter | 48
    frequent catheter changes every 48 hours | 48
    worsening delirium | 72
    deterioration of hemodynamic status | 72
    intravenous fluids started | 72
    vasopressors started | 72
    persistent metastatic infection | 96
    decision to remove right femoral catheter | 96
    transition to PD | 96
    peritoneal catheter inserted | 96
    PD plan gradual escalation of volume and frequency | 96
    well-tolerated PD | 96
    improvement in clinical status | 96
    mental improvement | 96
    hemodynamic improvement | 96
    resolution of fever | 96
    plasma biochemistry improvement | 96
    uremic status improvement | 96
    intravenous daptomycin continued for 6 weeks | 96
    discharged to long-term nursing facility | 240
    chronic manual ambulatory PD | 240
    blood cultures positive on days 1-11 | 24
    blood cultures negative on days 5, 12-21 | 168
    catheter tip culture negative on days 12 and 17 | 168
    initiation of peritoneal dialysis | 96
    