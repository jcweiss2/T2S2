23 years old | 0
female | 0
admitted to the hospital | 0
painful and swollen right breast | -12
breast pruritus | -72
dizziness | -12
nausea | -12
vomiting | -12
obesity | 0
polycystic ovarian syndrome | 0
non-smoker | 0
social alcohol consumption | 0
discoloured breast | 0
offensive nipple discharge | 0
grossly swollen breast | 0
tender breast | 0
discolouration | 0
erythema | 0
bullae | 0
severe sepsis | 0
end organ dysfunction | 0
increased white cell count | 0
neutrophilia | 0
increased C-reactive protein | 0
metabolic acidosis | 0
elevated lactate | 0
elevated creatinine | 0
reduced estimated glomerular filtration rate | 0
elevated international normalised ratio | 0
elevated activated partial thromboplastin time | 0
intravenous crystalloid resuscitation | 0
inotropic support | 0
metaraminol administration | 0
adrenaline administration | 0
noradrenaline infusion | 0
vasopressin infusion | 0
meropenem administration | 0
clindamycin administration | 0
vancomycin administration | 0
emergency right mastectomy | 3
debridement of necrotic tissue | 3
pectoralis major fascia debridement | 3
fresh frozen plasma administration | 3
vacuum assisted closure dressing | 3
intensive care unit admission | 3
continuous renal replacement therapy | 3
troponin-I rise | 12
ST elevation | 12
myocardial ischaemia | 12
aspirin administration | 12
heparin infusion | 12
noradrenaline infusion weaning | 6
noradrenaline infusion cessation | 48
continuous renal replacement therapy cessation | 12
extubation | 192
wound debridements | 24
VAC applications | 24
tissue culture positive for streptococcus pyogenes | 120
antibiotic therapy change to benzylpenicillin | 120
inflammatory markers improvement | 120
afebrile | 120
oral amoxicillin | 120
electrocardiogram | 120
transthoracic echocardiogram | 120
ejection fraction | 120
septal and inferior wall motion abnormality | 120
mild hypokinesis | 120
CT coronary angiograms | 384
ICU discharge | 288
ward transfer | 288
plastic surgery service transfer | 384
skin grafting | 384
discharge | 384