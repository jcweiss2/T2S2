50 years old | 0
female | 0
admitted to the hospital | 0
fever | -168
abdominal pain | -168
loose stools | -168
dry cough | -336
history of vomiting | -672
history of dyspnoea | -672
history of sputum production | -672
history of haemoptysis | -672
history of obstructive airway disease | -672
history of antitubercular treatment | -672
type 2 diabetes mellitus | -0
hypertension | -0
hypothyroidism | -0
thyroid surgery | -6480
surgical site infection | -6468
involvement of trachea | -6468
on and off dry cough | -2880
treated symptomatically | -2880
cough suppressants | -2880
antibiotics | -2880
symptoms used to recur | -2880
moderately built woman | 0
weight of 62 kg | 0
afebrile | 0
blood pressure of 80/50 mmHg | 0
pulse rate of 110/min | 0
SpO2 of 94 % on room air | 0
surgical scar of thyroid surgery | 0
no pallor | 0
no icterus | 0
no cyanosis | 0
no clubbing | 0
no pedal oedema | 0
no lymphadenopathy | 0
dehydrated | 0
peripheries were cool | 0
peripheral pulses were not well palpable | 0
gastrointestinal system examination was unremarkable | 0
upper respiratory tract examination was normal | 0
scattered coarse crackles at bilateral lung bases | 0
total count: 15,500 | 0
haemoglobin: 11.2 | 0
platelets: 231,000 | 0
C-reactive protein: 31.3 | 0
serum creatinine: 1.9 | 0
sodium: 133 | 0
potassium: 3.0 | 0
aspartate aminotransferase: 663 | 0
alanine transaminase: 317 | 0
sensitive thyroid-stimulating hormone: 0.69 | 0
chest radiograph: Normal | 0
high-resolution computed tomography (HRCT) of the thorax with dynamic tracheal imaging: Normal tracheal appearance seen during inspiration | 0
high-resolution computed tomography (HRCT) of the thorax with dynamic tracheal imaging: A typical crescentric tracheal appearance with >50% narrowing of lumen s/o TM seen during expiration | 0
centrilobular emphysematous cyst in anterior segment of right lower lobe | 0
diagnosis of acute gastroenteritis | 0
diagnosis of sepsis | 0
diagnosis of prerenal acute kidney injury | 0
diagnosis of upper respiratory infection | 0
elevated inflammatory markers | 0
growth of Escherichia coli in blood culture | 0
treated in Intensive Care Unit (ICU) | 0
appropriate antibiotics | 0
tracheal pathology suspected | 0
diagnosis of TM | 24
bronchoscopy | 24
tracheoplasty | 24
stenting | 24
conservative treatment with cough suppressant | 24
influenza vaccination | 24
discharged | 168