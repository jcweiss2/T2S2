74 years old | 0
male | 0
hypertension | 0
insulin-dependent diabetes mellitus type 2 | 0
diabetic retinopathy | 0
admitted to the hospital | 0
weight loss | -672
iron deficiency anemia | -672
tumor in the colon ascendens | -672
liver metastases | -672
right hemicolectomy | -672
low-grade pT3cN0 adenocarcinoma | -672
absence of metastases in 24 excised lymph nodes | -672
lymphovascular growth | -672
no vascular or perineural growth | -672
activated BRAF mutation | -672
loss of expression of MLH1 and PMS2 | -672
mismatch repair-deficient (MMR-D)/microsatellite-instable (MSI) tumor | -672
initiated therapy with pembrolizumab | 0
symptoms of a cold | 168
leukocytosis | 168
slight increase in C-reactive protein | 168
dry coughing | 528
no fever | 528
increase in AST and ALT | 528
ICI-induced hepatitis grade 2 | 528
initiated prednisolone therapy | 528
second dose of pembrolizumab not given | 528
dyspnea | 696
myocardial infarction suspected | 696
elevation of troponin T | 696
septal hypokinesia | 696
somnolence | 720
difficulty walking | 720
dysarthria | 720
hoarseness | 720
pain in neck and right leg | 720
difficulty raising right leg | 720
dose of prednisolone increased | 720
computed tomography did not show signs of stroke | 720
increased creatine kinase and myoglobin levels | 720
ICI-induced myositis suspected | 720
gradual decrease in creatinine levels | 720
antibodies against acetylcholine receptor and titin present | 720
albumin present in cerebrospinal fluid | 720
myasthenia gravis (MG) | 720
unable to sit up | 1008
severe dysarthria and dysphagia | 1008
absent reflexes | 1008
transferred to intensive care unit | 1008
intubated | 1104
given methylprednisolone | 1104
given intravenous immunoglobulins | 1104
given infliximab | 1104
felt better | 1128
better muscle strength in hands | 1128
developed carbon dioxide retention | 1164
needed noninvasive ventilation | 1164
developed sinus bradycardia | 1164
died | 1164
autopsy showed significant stenosis of right coronary artery | 1164
no fibrosis or signs of recent myocardial infarction | 1164
tongue softened | 1164
no surgical complication after hemicolectomy | 1164
metastasis in right liver lobe | 1164
pronounced inflammatory infiltration of lymphocytes | 1164
fibrosis consistent with myositis | 1164
fibrosis in heart consistent with myocardial infarction | 1164
inflammatory infiltrate in heart | 1164
hepatocellular cancer (HCC) | 1164
HCC positive for hepatocytes | 1164
HCC negative for glypican, CDX2, CK20 and CK7 | 1164
fibrosis stage 2-3 in liver | 1164
cause of death determined as respiratory insufficiency | 1164
due to polymyositis | 1164