33 years old | 0
female | 0
injection drug use | 0
untreated chronic hepatitis C infection | 0
fever | -72
pruritic lesion | -72
erythematous | -72
warm | -72
tender | -72
right-sided periorbital edema | -72
febrile | -72
white blood cell count 17.0 × 106 cells/L | -72
neutrophils 80.3% | -72
preseptal cellulitis | -72
IV vancomycin | -72
IV ceftriaxone | -72
discharged herself | -48
methicillin-resistant Staphylococcus aureus | -48
headache | -336
facial pain | -336
shortness of breath | -336
pain everywhere | -336
transferred to our facility | -336
alert | 0
oriented only to self | 0
blood pressure 137/79 mmHg | 0
heart rate 82 beats per minute | 0
temperature 37.6°C | 0
respiratory rate 26 breaths per minute | 0
oxygen saturation 97% | 0
bilateral severe eyelid edema | 0
chemosis | 0
right-sided peripheral facial droop | 0
no nuchal rigidity | 0
cardiac findings normal | 0
pulmonary exam revealed diffuse rhonchi | 0
WBC 31.3 × 106 cells/L | 0
C-reactive protein 409.9 mg/L | 0
erythrocyte sedimentation rate 97 mm/h | 0
peripheral blood cultures grew MRSA | 0
urine drug screen positive for opiates | 0
urine drug screen positive for cocaine | 0
CT of the head without contrast | 0
CT perfusion | 0
CT angiogram of the head and neck | 0
CT of the face with contrast | 0
MRI with and without contrast | 0
bilateral facial, preseptal, and postseptal cellulitis | 0
septic thrombophlebitis in multiple bilateral facial veins | 0
thrombosis in the bilateral cavernous sinuses | 0
thrombosis in multiple dural sinuses | 0
thrombosis in bilateral IJVs | 0
internal carotid artery stenosis | 0
endarteritis | 0
infarcts involving the right lateral hemipons | 0
infarcts involving bilateral cerebral hemispheres | 0
CT of the chest with contrast | 0
septic emboli | 0
transthoracic echocardiogram | 0
no valvular vegetations | 0
IV vancomycin | 0
heparin | 0
worsening of ventriculitis | 24
ACA/MCA watershed infarcts | 24
neurosurgery to place a stent in her right ICA | 48
lumbar puncture | 48
cerebrospinal fluid culture grew MRSA | 48
IV daptomycin | 72
goals-of-care discussion | 168
comfort care initiated | 168
transfer to hospice | 168
died | 504