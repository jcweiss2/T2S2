45 years old | 0
    male | 0
    swelling in the right lower limb | -120
    tenderness in the right lower limb | -120
    leukocytosis | -120
    necrotizing fasciitis | -120
    septic shock | 0
    right internal jugular venous central line placed | 0
    initial volume resuscitation | 0
    treatment with antibiotics | 0
    extensive debridement | 0
    intubated | 0
    mechanical ventilation | 0
    inotropic support | 0
    transferred to ICU | 0
    bedside ultrasonography | 0
    intraluminal hyperechoic shadow | 0
    X-ray ordered | 0
    confirmation of guidewire position | 0
    ultrasound examination of central venous line | 0
    guidewire in external part | 0
    left femoral central catheter inserted | 0
    inotropic infusion pump shifted to femoral line | 0
    right internal jugular line clamped | 0
    removal of guidewire | 24
    repeat bedside ultrasound documenting removal | 24