39 years old | 0
African-American | 0
male | 0
admitted from a nursing home | 0
weakness | 0
decreased appetite | 0
admitted to medical Intensive Care Unit | 0
suspected sepsis of unknown origin | 0
started empirically on vancomycin | 0
started empirically on meropenem | 0
urine cultures grew >100,000 CFU/mL of Candida glabrata | 0
chronic indwelling Foley catheter | 0
urinary retention | 0
stabilized | 144
transferred to general medical floor | 144
further management of sepsis | 144
subsequent workup on days 10–13 | 240-312
osteomyelitis | 240-312
Stage IV sacral decubitus ulcer | 240-312
exposed bone | 240-312
negative blood cultures | 240-312
urine cultures remained positive | 672
urine cultures yielded 15,000 CFU/mL of Candida albicans | 672
treated for osteomyelitis for 45 days | 0
combination therapy with vancomycin | 0
various Gram-negative therapies | 0
meropenem | 0
ertapenem | 0
ceftazidime | 0
workup for failure to thrive | 48
body mass index 14.7 kg/m² | 48
percutaneous endoscopic gastrostomy tube placement | 288
elevated alkaline phosphatase | 0
elevated aspartate aminotransferase | 0
elevated alanine aminotransferase | 0
failure to thrive | 0
poor nutritional status | 0
extremely brittle diabetes | 0
multiple hypoglycemic episodes | 0
corrected with 50% dextrose boluses | 0
started on insulin glargine 2 units every evening | 0
large fluctuations in blood sugars | 0
blood sugars ranging from 18 to 460 mg/dL | 0
average blood sugar 233 mg/dL | 0
switched to NPH insulin on day 51 | 1224
NPH insulin 2 units twice daily | 1224
avoid hypoglycemia | 1224
blood sugars drop to <50 mg/dL when not allowed to eat or drink | 0
required 5% dextrose infusion | 0
glycemic goals: avoid hypoglycemia | 0
glycemic goals: avoid diabetic ketoacidosis | 0
continued leukocytosis | 0
blood cultures drawn on day 34 | 816
urine cultures drawn on day 34 | 816
abdominal CT scan on day 36 | 864
right-sided pyelonephritis | 864
left-sided hydronephrosis | 864
left-sided hydroureter | 864
expanded antimicrobial therapy to include micafungin | 864
urology consulted on day 37 | 888
repeat abdominal CT scan on day 38 | 912
pyelonephritis in both kidneys | 912
filling defects (left > right) | 912
mild debris along bladder base | 912
fungus balls/mycetomas | 912
urine cultures on day 40 | 960
Candida glabrata | 960
Candida albicans | 960
fluconazole MIC 8 for C. glabrata | 960
caspofungin MIC 0.5 mg/L for C. glabrata | 960
fluconazole MIC 4 mg/L for C. albicans | 960
caspofungin MIC ≤0.25 mg/L for C. albicans | 960
blood cultures on day 40 | 960
fluconazole MIC 2 mg/L | 960
switched from micafungin to high-dose fluconazole | 960
urology recommended drainage of fungal balls | 960
irrigation with AmBd via bilateral nephrostomy tubes | 960
nephrostomy tube placed in left kidney on day 45 | 1080
drain fungal ball | 1080
preparation for AmBd irrigation | 1080
6 days of systemic antifungal therapy | 1080-1344
blood cultures cleared | 1344
renal ultrasound on day 54 | 1296
continued presence of fungal balls | 1296
lack of improvement in renal impairment | 1296
estimated glomerular filtration rate 10-30 mL/min/1.73 m² | 1296
comparable to pre-nephrostomy tube placement | 1296
required intermittent hemodialysis on day 56 | 1344
attempted placement of right nephrostomy tube on day 59 | 1416
placement failed | 1416
decision to discontinue fluconazole | 1416
initiated systemic AmBd at 0.7 mg/kg/day | 1416
treat renal fungal balls | 1416
LFTs significantly worsened on day 61 | 1464
Naranjo score 5 | 1464
LFTs returned near baseline | 1464
amphotericin B as culprit of acute liver injury | 1464
patient changed code status to DNR | 0
condition continued to decline | 0
daughter stopped 5% dextrose infusion | 0
patient expired | 1584
