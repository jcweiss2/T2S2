50 years old | 0
male | 0
presented with chest pain | 0
presented with shortness of breath | 0
chest computed tomography showed pulmonary emboli | -144
hospital day 6 | -144
transferred to intensive care unit | -144
intubated for severe respiratory distress | -144
hospital day 7 | -168
repeat CT showed progressive necrosis | -168
underwent thoracotomy with partial decortication | -168
underwent right thoracoscopy | -168
3 chest tubes placed | -168
started on empiric piperacillin-tazobactam | -168
started on intravenous vancomycin | -168
hospital day 9 | -216
bronchoalveolar lavage | -216
hospital day 12 | -288
meropenem-susceptible A. baumannii positive | -288
antibiotics switched to extended infusion meropenem | -288
underwent another thoracotomy | -288
underwent RLL resection | -288
underwent complete decortication | -288
pathology demonstrated acute fibrinopurulent exudate | -288
resected RLL demonstrated extensive abscess | -288
resected RLL demonstrated necrosis | -288
resected RLL demonstrated hemorrhage | -288
hospital day 18 | -432
pleural tissue culture demonstrated XDR A. baumannii | -432
intermediate susceptibility to colistin | -432
tigecycline MIC 2 mg/L | -432
switched from meropenem to tigecycline | -456
hospital day 19 | -456
hospital day 26 | -624
required vasoactive agents | -624
CT chest demonstrated RLL pyopneumothorax | -624
switched tigecycline to colistin | -624
switched to meropenem | -624
hospital day 28 | -672
underwent bronchoscopy | -672
identified right bronchopleural fistula | -672
acute tubular necrosis | -672
serum creatinine increased 7-fold | -672
hospital day 23 | -552
chest tube fluid culture | -552
hospital day 29 | -696
cefiderocol susceptible | -696
eravacycline susceptible | -696
switched colistin and meropenem to cefiderocol | -696
hospital day 40 | -960
bronchial washings culture | -960
hospital day 45 | -1080
XDR A. baumannii positive | -1080
cefiderocol-resistant | -1080
hospital day 49 | -1176
switched cefiderocol to eravacycline | -1176
hospital day 54 | -1296
febrile | -1296
tachycardic | -1296
increased chest tube output | -1296
eravacycline MIC increased to 1 mg/L | -1296
discontinued eravacycline | -1296
initiated combination therapy with cefiderocol | -1296
initiated combination therapy with tigecycline | -1296
hospital day 62 | -1488
started sulbactam-durlobactam | -1488
started meropenem | -1488
hospital day 75 | -1800
chest tube output resolved | -1800
completed 3 weeks of antibiotic therapy | -1800
antibiotics discontinued | -1800
cleared for discharge | -1824
followed up with infectious diseases | 0
at prehospital baseline | 672
