37 years old | 0
rheumatic mitral stenosis | 0
mild aortic insufficiency | 0
pulmonary hypertension | 0
referred to surgical treatment | -48000
heart failure | -33600
signs of endocarditis | -33600
sepsis with excessive organ failure | -33600
urgent surgery | -33600
implantation of mechanical mitral valve | -33600
minor commissurotomy of aortic valve cusps | -33600
double valve re-endocarditis | -4032
affecting prosthetic mitral valve | -4032
affecting native aortic valve | -4032
urgent surgery | -4032
implantation of biological mitral valve | -4032
St. Jude Medical Epic, size 27 mm | -4032
due to aortic root abscess | -4032
full root implantation of Medtronic Freestyle stentless bioprosthesis | -4032
MFB size 23 mm | -4032
reimplantation of coronary ostia | -4032
preoperative coronary angiography | -4032
normal coronary arteries | -4032
without stenosis | -4032
diagnosed with non-ST-elevation myocardial infarction | -432
preoperative computed tomography | -432
coronary angiography | -432
90% ostial stenosis of left main coronary artery | -432
90% ostial stenosis of right coronary artery | -432
emergent re-reoperation | -432
coronary artery bypass grafting of left anterior descending branch | -432
coronary artery bypass grafting of right coronary artery | -432
intraoperative findings | -432
endoluminar glass-like pseudointimal membranes | -432
covering distal anastomosis of MFB | -432
covering both coronary ostiae | -432
admission to Rigshospitalet | 0
complex mechanical mitral valve endocarditis | 0
native aortic valve endocarditis | 0
aortic root abscess | 0
medical history | 0
heart failure after rheumatic fever | 0
mitral stenosis | 0
mitral valve replacement | 0
minor commissurotomy of fused aortic valve cusps | 0
otherwise healthy | 0
no risk factors for coronary artery disease | 0
preoperative coronary angiography | 0
normal | 0
emergently operated | 0
implantation of biological mitral valve | 0
St. Jude Medical Epic, size 27 mm | 0
full root FB in aortic position | 0
FB chosen due to tissue quality | 0
irregularity of revised root | 0
presence of rigid biological mitral valve prosthesis | 0
homograft not available | 0
reimplantation of coronary ostia | 0
button technique | 0
orientation of porcine coronary ostia | 0
left coronary artery reimplanted in left porcine ostium | 0
right coronary artery reimplanted higher and further to the right | 0
to avoid kinking or stretching of the coronary | 0
discharged after 6 weeks | 504
targeted intravenous antibiotic therapy | 504
atrial fibrillation | 504
newly diagnosed diabetes mellitus type 2 | 504
prescribed warfarin | 504
target international normalized ratio 2-3 | 504
enalapril 2.5 mg | 504
metformin 1000 mg | 504
metoprolol 50 mg | 504
follow-up transoesophageal echocardiography | 504
41 days postoperatively | 504
well-functioning FB valve in aortic position | 504
presented with chest oppression | 4032
pain in left arm | 4032
pain in hand | 4032
shortness of breath | 4032
physical examination | 4032
discrete heart murmur | 4032
irregular rhythm | 4032
lung auscultation | 4032
normal vesicular breath sounds | 4032
extremities without edema | 4032
general condition good | 4032
further physical examination normal | 4032
electrocardiogram | 4032
atrial fibrillation | 4032
new ST depressions | 4032
T-wave inversions in I | 4032
T-wave inversions in II | 4032
T-wave inversions in V5 | 4032
T-wave inversions in V6 | 4032
ST elevation in aVR | 4032
Troponin T samples | 4032
increasing concentration | 4032
maximum 196 ng/L | 4032
contrast-enhanced cardiac computed tomography | 4032
significant left coronary ostial stenosis | 4032
significant right coronary ostial stenosis | 4032
no sign of atherosclerosis | 4032
preoperative coronary angiography | 4032
90% stenosis in both ostia | 4032
otherwise normal coronary arteries | 4032
preoperative transthoracic echocardiogram | 4032
left ventricular ejection fraction 50% | 4032
excellent prosthetic aortic valve function | 4032
excellent prosthetic mitral valve function | 4032
not suitable for percutaneous coronary intervention | 4032
underwent emergent reoperation | 4032
aim to replace FB | 4032
aim to perform revascularization | 4032
intraoperative findings | 4032
partial opening of distal anastomosis | 4032
pseudointimal glass-like membranes | 4032
covered distal anastomosis | 4032
covered both coronary ostia | 4032
high-grade stenoses | 4032
membranal tissue brittle | 4032
not invading FB tissue | 4032
peeled off in strips | 4032
pseudointimal membranes extended from anastomotic sites | 4032
into both coronary arteries | 4032
surgical detachment of membrane tissue | 4032
radical in proximal parts | 4032
replacement of FB considered | 4032
risk of dissection | 4032
coronary occlusion by remaining membrane tissue | 4032
PCI could dislodge membrane | 4032
cause occlusion | 4032
tissue sample of pseudointimal membrane | 4032
coronary artery bypass grafting | 4032
separate venous grafts | 4032
left anterior descending artery | 4032
right coronary artery | 4032
recovery uneventful | 4032
epigastric fascial rupture | 4032
smaller procedure | 4032
acetylsalicylic acid 75 mg | 4032
previous medication | 4032
metoprolol reduced to 25 mg | 4032
histological examination | 4032
fibro-intimal thickening | 4032
inflamed granulation tissue | 4032
no sign of acute inflammation | 4032
no calcifications | 4032
no foreign bodies | 4032
no amyloidosis | 4032
follow-up cardiac CT | 4320
transthoracic echocardiography | 4320
complaints of chest pains | 4320
small pseudoaneurysm | 4320
2.3 mL | 4320
arising from partial rupture | 4320
distal anastomosis between FB and aorta | 4320
conservative, non-surgical strategy | 4320
repeat follow-up cardiac CT | 4320
3 months later | 4320
reduction of pseudoaneurysm to 1.4 mL | 4320
during follow-up | 10824
suffered exercise-induced chest pains | 10824
myocardial perfusion scintigraphy | 10824
exercise-induced myocardial ischemia | 10824
6-8% | 10824
due to previous myocardial infarction | 10824
coronary angiography | 10824
complete revascularization | 10824
transthoracic echo | 10824
mild-moderate stenosis of FB valve | 10824
well-functioning biological mitral valve | 10824
