43 years old | 0
female | 0
admitted to the hospital | 0
fever | -336
lower abdominal pain | -336
foul-smelling discharge | -336
perianal region | -336
necrotic tissue | 0
foul-smelling thin pus | 0
surgery | 0
debridement | 0
abscess | 0
laparotomy | 48
thick abscess | 48
necrotic rectus muscle | 48
abscess drainage | 48
debridement | 48
abdomen left open | 48
Bogota bag | 48
antibiotics changed | 48
relaparotomy | 96
no disease progression | 96
ICU | 96
antibiotics | 96
reconstruction | 840
sub-umbilical fascia defect | 840
non-vascularized bilateral tensor fascia-lata graft | 840
abdomen closed | 840
secondary closure of perianal wound | 840
follow-up visit | 2160
computed tomography scan | 2160
normal anterior abdominal fascia | 2160
discharged | 2160