80 years old | 0
male | 0
admitted to the hospital | 0
COVID-19 | -168
intubated | -168
prone positioning | -168
moderately responsive | -168
transferred to ICU | -9
ARDS | -9
MOF | -9
oliguria | -9
septic shock | -9
hepatic dysfunction | -9
mixed acidosis | -9
SOFA-Score 13 | -9
noradrenalin 0.35 µg/kg/h | -9
ECMO not initiated | -9
ADVOS treatment started | 0
renal replacement therapy | 0
mixed acidosis | 0
hepatic failure | 0
blood flow 100–300 mL/min | 0
dialysate flow 160–320 mL/min | 0
dialysate pH 7.6–9.0 | 0
atrial fibrillation | 24
digitoxin administered | 24
ultrafiltration performed | 24
hemodynamic parameters improved | 48
vasopressor requirement reduced | 48
pH-normalization | 48
system clotting | 48
dialysis circuit renewed | 48
CO2 removal | 48
acid-base balance controlled | 48
infections detected | 95
Klebsiella oxytoca | 95
Aspergillus-antigen-testing positive | 95
anti-microbial systemic therapy | 95
hemoptysis | 95
cardiac arrest | 160
death | 160
autopsy not performed | 160