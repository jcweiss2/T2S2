62 years old | 0
male | 0
diabetes mellitus | -4320
hypertension | -4320
abdominal pain | -4320
palpable pulsatile epigastric mass | -4320
bilateral total hip replacements | -4320
infected hip replacements | -4320
levofloxacin | -4320
teicoplanin | -4320
vancomycin | -4320
implant removal | -4320
joint spacers implanted | -4320
blood cultures demonstrated MRSA | -4320
tissue cultures demonstrated proteus mirabilis | -4320
fever persisted | -4320
CT demonstrated septic spleen | -4320
splenectomy performed | -4320
recurrent sepsis | -1440
white blood count of 12,000/mm3 | -1440
CT angiography revealed paravisceral aortic pseudoaneurysm | -1440
transferred to tertiary care center | -1440
written consent obtained | -1440
attempted covered stent placement | -1440
midline laparotomy | 0
exposed paravisceral aorta | 0
exposed infrarenal aorta | 0
divided crura of diaphragm | 0
clamped aorta proximal to CA | 0
clamped aorta below renal arteries | 0
opened pseudoaneurysm | 0
removed infected tissues | 0
removed necrotic aortic wall | 0
reconstruction of CA not feasible | 0
ligated distal CA | 0
excised pseudoaneurysm | 0
repaired aorta with cryopreserved allograft | 0
aortic cross clamp time 34 min | 0
postoperative intensive care stay | 48
blood cultures confirmed MRSA | 48
tissue culture from aortic wall negative | 48
dismissed to rehabilitation facility | 168
meropenem | 168
free of infection at 1-year follow-up | 8760
control CTA showed patent SMA | 8760
control CTA showed patent renal arteries | 8760
control CTA showed no pseudoaneurysm | 8760
no symptoms of infection | 8760
