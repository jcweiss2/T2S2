28 years old | 0
male | 0
admitted to the hospital | 0
hepatomegaly | 0
splenomegaly | 0
leukopenia | 0
thrombocytopenia | 0
Gilbert’s syndrome | -672
fever | -72
recurrent episodes of fever | -72
abdominal pain | -72
enlarged spleen | 0
enlarged liver | 0
leukopenia with neutropenia | 0
thrombocytopenia | 0
elevated activity of aminotransferases | 0
increased total bilirubin level | 0
viral studies excluded HIV | 0
viral studies excluded HCV | 0
viral studies excluded HBV | 0
abdominal ultrasonography | 0
bone marrow smear evaluation | 0
multiparameter flow cytometric analysis | 0
bone marrow cytogenetic study | 0
positron emission tomography | 24
PET-CT examination | 24
fever | 72
persistent dry cough | 72
urine culture revealed Escherichia coli | 72
Chlamydophila pneumoniae antigen | 72
increased lactate dehydrogenase activity | 72
another bone marrow examination | 72
normal cytomorphology | 72
normal immunophenotype | 72
no ring sideroblasts | 72
paroxysmal nocturnal hemoglobinuria excluded | 72
CMV infection excluded | 72
EBV infection excluded | 72
parvovirus B19 infection excluded | 72
beta-glucocerebrosidase normal | 72
ceruloplasmin activity normal | 72
chest X-ray normal | 72
treated with levofloxacin | 72
treated with filgrastim | 72
recovered from fever | 96
leukocyte count increased | 96
recurrence of fever | 120
worsening of neutropenia | 120
filgrastim and prophylactic antibiotic therapy restarted | 120
steroid therapy initiated | 120
clinical improvement | 144
fever subsided | 144
leukocyte count increased | 144
additional tests excluded ANA | 144
additional tests excluded ANCA | 144
additional tests excluded anti-hepatic antibodies | 144
additional tests excluded anti-cardiolipin antibodies | 144
additional tests excluded anti-beta2-microglobulin antibodies | 144
liver biopsy | 168
elevated activity of aminotransferases | 168
concentration of bilirubin | 168
enlargement of liver and spleen | 168
histopathological examination of liver biopsy | 168
no clinically important abnormalities | 168
fever recurred | 168
empirical antibiotic therapy started | 168
doses of steroids escalated | 168
fever did not resolve | 168
transferred to Department of Hematology | 192
severe abdominal pain | 192
enlarged spleen and liver | 192
abdominal USG | 192
free fluid in abdominal cavity | 192
rapid drop in hemoglobin concentration | 192
abdominal CT | 192
enlargement of liver | 192
enlargement of spleen | 192
subcapsular rupture | 192
retroperitoneal enlarged lymph nodes | 192
transferred to Surgery Department | 216
splenectomy | 216
enlarged lymph nodes collected | 216
transferred to Intensive Care Unit | 216
numerous transfusions | 216
erythrocytes and platelets concentrates | 216
fresh frozen plasma | 216
recombinant factor VIIa | 216
hematoma in spleen extraction site | 216
another laparotomy | 216
aspiration biopsy | 216
numerous hemophagocytes | 216
significant increase in ferritinemia | 216
met 5 of 8 HLH 04 criteria | 216
treated with dexamethasone | 216
treated with etoposide | 216
treated with cyclosporine A | 216
condition deteriorated rapidly | 240
multiple-organ failure | 240
respiratory failure | 240
septic shock | 240
liver failure | 240
cerebral hemorrhage | 240
died | 240
histopathological assessment of retroperitoneal lymph nodes | 240
peripheral T-cell lymphoma | 240