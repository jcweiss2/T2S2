27 years old | 0
male | 0
admitted to the hospital | 0
fever | -336
fatigue | -336
unconsciousness | -24
recurrent fever | -336
highest documented temperature 40.0°C | -336
bilateral lung infection | -336
WBC count 14.63 × 10^9/L | -336
RBC count 3.35 × 10^12/L | -336
hemoglobin 107.00 g/L | -336
platelet count 98 × 10^9/L | -336
CRP 47.63 mg/L | -336
moxifloxacin 0.4 g daily | -336
chest CT showed bilateral pneumonia | -336
intubated | 0
mechanical ventilation | 0
norepinephrine infusion | 0
shallow breathing | 0
moist crackles | 0
anoxia | 0
hyperventilation | 0
low partial pressures of oxygen | 0
low pH | 0
transcutaneous oxygen saturation 75% | 0
WBC count 34.45 × 10^9/L | 0
CRP concentration 80.78 mg/L | 0
hemoglobin 90.00 g/L | 0
platelet count 80.78 × 10^9/L | 0
RBC count 3.36 × 10^12/L | 0
mean corpuscular volume 120.1 fL | 0
mean corpuscular hemoglobin 40.8 pg | 0
erythrocyte sedimentation rate 106 mm/h | 0
ferritin > 1500.00 ng/mL | 0
severe pneumonia | 0
respiratory failure | 0
septic shock | 0
anemia | 0
thrombocytopenia | 0
trisomy 8 | 0
vancomycin 1 g 12 hly | 0
imipenem 0.5 g 6 hly | 0
ambroxol | 0
omeprazole | 0
enteral nutrition | 0
vancomycin discontinued | 72
fluconazole 0.4 g daily | 120
methylprednisolone 500 mg daily | 120
imipenem discontinued | 216
piperacillin–tazobactam 4.5 g 8 hly | 216
methylprednisolone dose reduced to 250 mg daily | 216
extubated | 288
methylprednisolone dose reduced to 120 mg daily | 312
methylprednisolone dose reduced to 60 mg daily | 336
transferred to Department of Respiratory Medicine | 408
discharged | 432
Epstein–Barr virus detected | 0
Mycobacterium kansasii detected | 0
Cordyceps portugal detected | 48
bone marrow examination showed erythroid deficiency | 48
bone marrow examination showed grain maturation disorder | 48
chromosome analysis showed trisomy 8 | 48
Candida Portugal detected | 48
blood cultures performed | 48
informed consent obtained | -336
informed written consent obtained | 0