68 years old | 0
male | 0
admitted to the Emergency Department | 0
chest pain | -2
vomiting | -2
hypertension | -Infinity
hyperuricemia | -Infinity
Mallory-Weiss syndrome | -Infinity
arterial blood pressure 144/78 mmHg | 0
cardiac frequency 108/min | 0
peripheral oxygen saturation 90% | 0
temperature 37.7°C | 0
decreased respiratory sounds in both inferior pulmonary areas | 0
no changes on abdominal examination | 0
pH 7.45 | 0
pO2 57.2 mmHg | 0
pCO2 36.2 mmHg | 0
HCO3–36.4 mEq/L | 0
O2 saturation 90.4% | 0
pulmonary opacity on the left | 0
white blood cell count 10.200/mm3 | 0
normal electrocardiography | 0
normal high sensitivity troponin I | 0
admitted to the Internal Medicine Department | 0
presumptive diagnosis of pneumonia | 0
intravenous antibiotic | 0
oxygen | 0
severe chest pain | 48
respiratory distress | 48
type 1 respiratory failure | 48
increased white blood cell count | 48
increased c-reactive protein | 48
increased d-dimer | 48
chest computed tomographic angiography | 48
important pneumomediastinum | 48
hydropneumothorax on the left chest | 48
destruction of the lower esophagus | 48
spontaneous rupture of the esophagus | 48
emergent transhiatal esophagectomy | 48
primary anastomosis | 48
left thoracic drainage | 48
esophageal perforation | 48
no peritonitis | 48
pleural effusion | 48
nasojejunal tube | 48
transfered to the intensive care unit | 48
stayed in intensive care unit for 8 days | 48
oral swallow X-ray revealed no anastomotic leak | 48
clear liquid diet started | 144
discharged home | 504
oral contrast esophagogram 1 month after discharge | 672
no anastomotic leak | 672
no stenosis | 672
asymptomatic one year later | 8760
