82 years old | 0
female | 0
admitted to the emergency department | 0
cognitive regression | 0
deterioration | 0
decreased oral intake | 0
fever | -168
hypertension | 0
chronic atrial fibrillation | 0
bilateral salpingo-oophorectomy | 0
total abdominal hysterectomy | 0
clavicle fracture | -70080
bed-dependent state | -26208
GCS was 8 | 0
SaO2 was 92–95% | 0
ABP was 90/60 mmHg | 0
pulse was 120–136 bpm | 0
respiratory rate was 25–35/min | 0
ED transthoracic echocardiogram findings normal | 0
CT no active consolidation | 0
CT no pulmonary thromboembolism | 0
colonic loops distended | 0
no urgent surgery needed | 0
sepsis not ruled out | 0
breathing pattern deteriorated | 0
intubated | 0
vasopressor support | 0
admitted to ICU | 0
perianal abscess | 0
perianal fistula | 0
abscess drained | 0
mechanical ventilatory support | 0
laboratory assays stabilized | 0
sedation with dexmedetomidine/propofol | 0
analgesia with fentanyl/morphine | 0
ventilatory weaning failed | 672
daily sedation/analgesia intervals | 672
spontaneous breathing trials | 672
tracheostomy considered | 672
short thyromental distance | 672
short neck | 672
limited neck extension | 672
ENT evaluation | 672
OST performed | 672
no intraoperative complications | 672
no early post-operative complications | 672
enteral feeding remnants in tracheostomy | 48
pulsative air filling in nasogastric bag | 48
bedside bronchoscopy performed | 48
trachea and esophagus joined | 48
single passage lumen | 48
tracheal laceration | 48
fistulation | 48
contrast-enhanced CT verification | 48
wide communication of trachea and esophagus | 48
tube jejunostomy performed | 72
air filling into GIS ongoing | 72
reconstructive surgery concluded | 72
SBt inserted | 120
gastric balloon inflated | 120
esophagus balloon inflated | 120
SBt position confirmed | 120
SBt adaptation improved | 120
air leak prevented | 120
GIS reflux prevented | 120
ED transthoracic echocardiogram findings normal |' 0
