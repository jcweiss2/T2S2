40 years old| 0
    man | 0
    arrived as a patient with priority 1 trauma | 0
    gunshots to the chest | 0
    gunshots to the abdomen | 0
    gunshots to the pelvis | 0
    resuscitative thoracotomy | 0
    emergent exploratory laparotomy | 0
    splenectomy | 0
    direct repair of enterotomies | 0
    gastrotomy | 0
    traumatic IVC injury | 0
    abdominal packing | 0
    temporary abdominal closure | 0
    mass transfusion protocol | 0
    transfer to surgical trauma intensive care unit | 0
    continued resuscitation | 0
    high sanguineous output from abdominal wound | 0
    hemodynamic instability at 7:12 am | 0
    noticeable hemoperitoneum | 0
    increasing drain output | 0
    fluid balance within first 12 hours of admission | 0
    transfusion totals within first 12 hours of admission | 0
    hemoglobin levels | 0
    Abtheraa loss | 0
    intraoperative fluid loss | 0
    total administered fluid | 0
    total loss fluid | 0
    transfusion total | 0
    packed red blood cells transfusion | 0
    vascular surgery consultation | 0
    multidisciplinary team meeting | 0
    decision for IVC venogram | 0
    activation of semihybrid circulatory dynamics laboratory | 0
    continued massive transfusion protocol | 0
    hemodynamics supported with vasopressors | 0
    ultrasound-guided access of right femoral vein | 0
    8F sheath placement | 0
    IVC venogram | 0
    power injector through 5F Omni flush catheter | 0
    no apparent blush within retrohepatic IVC | 0
    retraction of catheter | 0
    imaging series with undiluted contrast | 0
    substantial blush within suprarenal IVC | 0
    angiographic sizing of IVC | 0
    IVUS probe advancement | 0
    measurements at proximal and distal IVC injury sites | 0
    decision to use Gore TAG 28.5-mm × 3.3-cm endograft cuff | 0
    table locked and screen marked | 0
    20F Gore DrySeal sheath exchange | 0
    deployment of endograft | 0
    completion venogram | 0
    tilting of first cuff | 0
    incomplete seal | 0
    continued blush | 0
    visualization of renal veins | 0
    deployment of second Gore TAG endograft cuff | 0
    complete seal | 0
    resolution of blush | 0
    access site closure | 0
    monofilament figure-of-eight cutaneous stitch | 0
    direct pressure for 10 minutes | 0
    hemostasis | 0
    coagulation panel ordered | 0
    return to trauma intensive care unit | 0
    hemodynamic stability overnight | 0
    return to operating room for abdominal washout | 24
    total operative case time 53 minutes | 24
    follow-up computed tomography scan | 336
    no stent graft migration | 336
    no extravasation around stent graft | 336
    discharge home | 168
    advised 30-day follow-up | 168
    prescription for daily 75 mg clopidogrel | 168
    prescription for 81 mg aspirin | 168
    plans for continuing clopidogrel for 6 months | 168
    long-term broad-spectrum antibiotics | 168
    no clinical signs of infection | 168
  