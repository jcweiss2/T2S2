55 years old | 0
female | 0
smoker | 0
chronic obstructive pulmonary disease | 0
diabetes | 0
presented to the emergency department | 0
worsening dyspnea | 0
respiratory distress | 0
tachypnea | 0
tachycardia | 0
wheezing | 0
decreased breath sounds in the left upper lung field | 0
chest radiography showed left upper lung airspace disease | 0
pneumonia | 0
acute respiratory failure | 0
admitted to the intensive care unit | 0
intravenous antibiotics | 0
fluid resuscitation | 0
noninvasive ventilatory support | 0
right upper quadrant pain | 0
high alkaline phosphate level | 0
abdominal ultrasonography conducted | 0
enlarged liver | 0
multiple liver masses | 0
condition stabilized | 0
chest computed tomography | 0
abdomen computed tomography | 0
7 cm mass in the left upper lung lobe | 0
obstructive pneumonitis | 0
bilateral mediastinal lymphadenopathy | 0
left hilar lymphadenopathy | 0
axillary lymphadenopathy | 0
supraclavicular lymphadenopathy | 0
multiple liver metastases | 0
histopathologic examination of liver biopsy specimen | 0
high grade small cell neuroendocrine cancer | 0
magnetic resonance imaging of the brain yielded normal findings | 0
extensive stage small cell lung cancer | 0
hospital day 4 | 96
oliguria detected | 96
elevated creatinine | 96
elevated potassium | 96
sepsis associated acute kidney injury | 96
increasing potassium levels | 96
maximum potassium 5.6 mEq/L | 96
increasing phosphorus levels | 96
maximum phosphorus 8.4 mg/dL | 96
increasing uric acid levels | 96
maximum uric acid 11.3 mg/dL | 96
spontaneous tumor lysis syndrome diagnosed | 96
aggressive treatment | 96
fluid resuscitation | 96
phosphate binders | 96
allopurinol | 96
rasburicase | 96
renal function deterioration | 96
creatinine increased from 0.5 mg/dL upon admission to 7.9 mg/dL over 6 days | 96
oncology consultation | 96
nephrology consultation | 96
daily hemolysis | 96
first cycle of palliative chemotherapy with cisplatin | 96
palliative chemotherapy with etoposide | 96
no major complications | 96
poor renal recovery | 96
dialysis dependent | 96
