unconscious state | 0
history of hypertension | 0
history of ischaemic heart disease | 0
history of peripheral vascular disease | 0
stroke | 0
head computed tomographic scan | 0
inotropic support | -48
septic shock | 48
elevated levels of inflammatory markers | 48
erythrocyte sedimentation rate, 70 mm/h | 48
C-reactive protein, 78 mg/L | 48
blood obtained | 48
yeast in both aerobic and anaerobic BacT/ALERT culture bottles | 48
caspofungin administered | 48
death | 72
identification as C. parapsilosis by the VITEK 2 yeast identification system | 72
turquoise blue colonies on CHROMagar Candida | 96
long ellipsoidal-shaped ascospores on acetate ascospore agar | 168
DNA sequence data comparisons | 168
hospitalization for lower limb ischaemia due to peripheral vascular disease | -336
discharge from hospital | -336
inoculation of the yeast from the skin | -48
translocation from the gastrointestinal tract | -48
antibiotics not administered | 0
no central lines emplaced | 0 
no shortness of breath | 0
denies chest pain | 0