63 years old | 0
male | 0
admitted to the hospital | 0
abdominal pain | -24
fever | -24
recurrent abdominal adhesions | -8760
multiple surgeries | -8760
Abcarian stoma | -8760
mucus fistula | -8760
body temperature 36.8°C | 0
blood pressure 109/54 mmHg | 0
pulse rate 109 beats/min | 0
respiratory rate 18 breaths/min | 0
coarse breathing sound | 0
regular heartbeats | 0
no audible murmur | 0
abdomen soft | 0
tenderness in the right upper quadrant | 0
positive murphy signs | 0
no palpable mass | 0
no hepatosplenomegaly | 0
mild anemia | 0
hemoglobin level 10.6g/dl | 0
neutrophilic leuocytosis | 0
white blood cell count 28,000/ml | 0
C-reactive protein level 100 mg/L | 0
troponin I level 48 ng/L | 0
renal function deranged | 0
creatinine level 176 umol/L | 0
urea 19 mmol/L | 0
normal electrolytes | 0
normal liver function tests | 0
normal serology | 0
normal urinalysis | 0
unremarkable chest X-ray | 0
thick gallbladder wall | 0
pericholecystic fluid | 0
sludge | 0
cholelithiasis | 0
sepsis secondary to acute cholecystitis | 0
antibiotics | 0
supportive measures | 0
highly febrile | 24
hypotensive | 24
inotropic support | 24
retrosternal chest pain | 48
profuse sweating | 48
ST-segment elevation on leads V2–V4 | 48
troponin-T level 781 ng/L | 48
anterior wall ST-segment elevation myocardial infarction | 48
emergent coronary angiography | 48
nonobstructive CAD | 48
dilated left ventricular cavity | 48
extensive apical dyskinesis | 48
relative preservation of the basal to midseptal and basal-lateral wall contraction | 48
estimated left ejection fraction 25% | 48
sepsis-induced TCM | 48
recovered | 240
discharged from the hospital | 240
repeated echocardiogram | 672
complete resolution of left ventricular systolic function | 672
estimated ejection fraction >55% | 672