85 years old | 0
male | 0
lived in a rural area | 0
no previous history of comorbidities | 0
dog bite on right arm | -360
fever | -48
aggressive behavior | -120
mental confusion | -120
psychomotor agitation | -120
impaired consciousness | -120
healing wound 3x2 cm on posterior right arm | 0
no signs of cutaneous or soft tissue infection | 0
nuchal rigidity | 0
Brudzinski’s sign | 0
leukocytosis (15,000/mm3) | 0
low platelet count (9,000/mm3) | 0
elevated C-reactive protein (187.7 mg/L) |E0
normal liver function tests | 0
normal renal function tests | 0
normal glycosylated hemoglobin level | 0
negative anti-HIV 1/2 Western blot | 0
negative blood cultures | 0
positive RT-PCR for SARS-CoV-2 | 0
diagnosis of COVID-19 | 0
normal cranial computed tomography | 0
cerebrospinal fluid (CSF) analysis performed | 0
CSF glucose 9 mg/dL | 0
CSF protein 171.3 mg/dL | 0
CSF white blood cell count 727 cells/mm3 | 0
CSF polymorphonucleocytes 89% | 0
CSF Gram stain with gram-negative bacilli | 0
CSF culture with translucent colonies on chocolate agar | 0
identification of C. canimorsus via MALDI-TOF | 0
no clinical improvement with ceftriaxone | 120
treatment switched to meropenem | 120
admission to ICU | 0
loss of consciousness | 0
no orotracheal intubation | 0
discharge from ICU | 120
discharged after 14-day meropenem | 336
full clinical resolution of symptoms | 336
no sequelae at six-month follow-up | 4320
no skin rash | 0
no purpura | 0
severe disease based on sepsis criteria | 0
central nervous system involvement | 0
no respiratory symptoms | 0
asymptomatic COVID-19 | 0
Gamma (P.1) variant | 0
CSF Gram stain of C. canimorsus | 0
CSF culture colonies after 48h incubation | 0
negative growth on MacConkey agar | 0
negative growth without CO2 | 0
Vitek®2 GN ID card low discrimination | 0
MALDI-TOF confirmation 99.9% confidence | 0
prompt clinical response to meropenem | 120
ICU stay 5 days | 120
treatment with meropenem for 14 days | 336
coinfection with SARS-CoV-2 | 0
immunocompetent patient | 0
rare case of C. canimorsus meningitis | 0
molecular diagnosis via MALDI-TOF | 0
