10 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
pre-term | 0 | 0 | Factual
gestational age of 33 weeks and 2 days | 0 | 0 | Factual
developmental delays in growth | 0 | 0 | Factual
developmental delays in motor function | 0 | 0 | Factual
short stature | -2190 | -2190 | Factual
Russell–Silver syndrome | -2190 | -2190 | Factual
proteinuria | -2190 | -2190 | Factual
hypoalbuminemia | -2190 | -2190 | Factual
nephrotic syndrome | -2190 | -2190 | Factual
high-dose steroid | -2190 | -1680 | Factual
calcineurin inhibitor | -2190 | -1680 | Factual
renal function deterioration | -1680 | -1680 | Factual
right renal vein thrombosis | -1095 | -1095 | Factual
pulmonary embolism | -1095 | -1095 | Factual
anticoagulants | -1095 | -730 | Factual
persistent pulmonary hypertension | -730 | 0 | Factual
sildenafil | -730 | 0 | Factual
living donor kidney transplantation | 0 | 0 | Factual
immunosuppression | 0 | 215 | Factual
prednisolone | 0 | 215 | Factual
mycophenolate mofetil (MMF) | 0 | 70 | Factual
tacrolimus | 0 | 215 | Factual
discontinued MMF | 70 | 70 | Factual
steroid tapered | 70 | 135 | Factual
pneumocystis pneumonia | 90 | 104 | Factual
mechanical ventilation | 90 | 104 | Factual
intravenous sulfamethoxazole/trimethoprim | 90 | 104 | Factual
steroid increased | 135 | 135 | Factual
dysuria | 135 | 215 | Factual
gross hematuria | 135 | 215 | Factual
blood urea nitrogen (BUN) 24 mg/dL | 135 | 135 | Factual
creatinine (Cr) 0.56 mg/dL | 135 | 135 | Factual
C-reactive protein (CRP) 0.42 mg/dL | 135 | 135 | Factual
urinalysis | 135 | 135 | Factual
red blood cell (RBC) count > 100/high power fields (HPF) | 135 | 215 | Factual
white blood cell (WBC) count > 100/HPF | 135 | 142 | Factual
urine culture for bacteria negative | 135 | 135 | Factual
urine BK virus negative | 135 | 135 | Factual
urine John Cunningham (JC) virus polymerase chain reaction (PCR) positive | 135 | 135 | Factual
urine adenovirus culture positive | 135 | 135 | Factual
hemorrhagic cystitis | 135 | 215 | Factual
hydration | 135 | 215 | Factual
pain control | 135 | 215 | Factual
fever | 159 | 215 | Factual
general weakness | 159 | 215 | Factual
chest tightness | 159 | 215 | Factual
mild cough | 159 | 215 | Factual
BUN 175 mg/dL | 159 | 159 | Factual
Cr 8.29 mg/dL | 159 | 159 | Factual
CRP 30.23 mg/dL | 159 | 159 | Factual
emergent hemodialysis | 159 | 215 | Factual
piperacillin/tazobactam | 159 | 215 | Factual
sputum culture negative | 159 | 159 | Factual
blood culture negative | 159 | 159 | Factual
urine culture negative | 159 | 159 | Factual
adenovirus real-time PCR of sputum positive | 159 | 159 | Factual
blood cytomegalovirus (CMV) antigen positive | 159 | 159 | Factual
disseminated adenovirus infection | 159 | 215 | Factual
immunosuppression reduction | 159 | 215 | Factual
ganciclovir | 159 | 215 | Factual
renal allograft biopsy | 159 | 159 | Factual
diffuse necrotizing granulomatous tubulointerstitial nephritis | 159 | 159 | Factual
infectious tubulointerstitial nephritis | 159 | 159 | Factual
JC virus PCR positive | 159 | 159 | Factual
serum CMV PCR positive | 159 | 159 | Factual
coinfection | 159 | 215 | Factual
cidofovir | 167 | 215 | Factual
nephrotoxicity | 167 | 215 | Factual
granulocyte colony-stimulating factor | 167 | 215 | Factual
immunoglobulin | 167 | 215 | Factual
transfusion | 167 | 215 | Factual
hemodialysis | 167 | 215 | Factual
anemia | 190 | 215 | Factual
leukopenia | 190 | 215 | Factual
thrombocytopenia | 190 | 215 | Factual
bone marrow suppression | 190 | 215 | Factual
generalized tonic-clonic seizure | 200 | 200 | Factual
vancomycin | 200 | 215 | Factual
meropenem | 200 | 215 | Factual
acyclovir | 200 | 215 | Factual
mechanical ventilation | 200 | 215 | Factual
continuous renal replacement therapy | 200 | 215 | Factual
death | 215 | 215 | Factual