54 years old | 0
female | 0
rheumatoid arthritis | 0
uncontrolled diabetes mellitus type II | 0
neuropathy | 0
hypothyroidism | 0
admitted to the hospital | 0
acute idiopathic necrotizing pancreatitis | -48
sepsis from an infected pseudocyst | -48
pressor support | -48
acute respiratory distress syndrome | -48
acute kidney injury | -48
deep vein thrombosis | -48
pulmonary embolism | -48
anticoagulation | -48
retroperitoneal drainage catheter | -24
abscess | -24
transfer to the tertiary care referral center | 0
admitted to the surgical intensive care unit | 0
anticoagulation therapy continued | 0
progressive abdominal pain | 24
low drain output | 24
imaging demonstrated appropriate drain position | 24
tissue-plasminogen activator (t-PA) injection | 24
fresh blood in the drainage catheter | 48
hypotensive | 48
decreased hemoglobin | 48
resuscitation | 48
crystalloid solution | 48
blood transfusions | 48
unenhanced CT of the abdomen and pelvis | 48
heterogeneously hyperdense subcapsular and perihepatic collections | 48
contrast-enhanced multiphase CT of the abdomen and pelvis | 48
active hemorrhage in the gallbladder fossa | 48
percutaneous endovascular embolization of the cystic artery | 72
gelatin foam | 72
detachable coil | 72
transfusion of packed red blood cells | 72
fresh frozen plasma | 72
albumin | 72
blood pressure stabilized | 72
hemoglobin stabilized | 72
anticoagulation not restarted | 72
serum transaminases increased | 120
alkaline phosphatase increased | 120
bilirubin increased | 120
hemoglobin decreased | 120
follow-up contrast-enhanced multiphase CT of the abdomen and pelvis | 120
increased size of the hepatic subcapsular hematoma | 120
hepatic ischemia | 120
liver enzymes worsened | 120
hepatic angiography | 144
punctate areas of contrast blush | 144
bleeding along the liver edge | 144
no embolization | 144
blood products and crystalloid resuscitation | 144
laboratory indicators worsened | 144
surgical evaluation | 168
laparoscopy | 168
extensive inflammatory adhesions | 168
large organized hematoma | 168
diffuse oozing from the liver parenchyma | 168
right subcostal incision | 168
evacuation of the large hepatic subcapsular hematoma | 168
numerous packs placed along the right hepatic edge | 168
hemostasis achieved | 168
subhepatic hematoma evacuated | 168
cholecystectomy | 168
retroperitoneal necrosectomy | 168
feeding jejunostomy tube placed | 168
primary closure of the surgical incision | 168
repeat laboratories drawn | 172
marked improvements in alkaline phosphatase | 172
ALT | 172
AST | 172
bilirubin | 172
no further bleeding events | 240
liver enzymes remained stable | 240
follow-up imaging | 768
persistent areas of infarction of large portions of the right hepatic lobe | 768
infarctions persisted on 5-month follow-up imaging | 4320