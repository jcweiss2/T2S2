69 years old | 0
female | 0
stabbed herself in the abdomen | -1
admitted to emergency department | 0
blood pressure could not be measured | 0
pulseless electrical activity | 0
body temperature 35.0 °C | 0
oxygen saturation 99 % | 0
Glasgow Coma Scale score 3 | 0
agonal respiration | 0
wound on upper abdomen | 0
intra-abdominal fluid collection | 0
emergency thoracotomy | 1
aortic cross-clamping | 1
open cardiac massage | 1
epinephrine administration | 1
temporary return of spontaneous circulation | 1
hemodynamically unstable | 1
laparotomy | 2
injuries to common hepatic and splenic arteries | 2
injuries to pancreas, spleen, and liver | 2
ligation of injured arteries | 2
distal pancreatectomy | 2
splenectomy | 2
liver sutured | 2
norepinephrine administration | 2
second-look surgery | 24
no active bleeding | 24
no ischemic change | 24
abdominal wall closure | 72
enhanced CT scan | 96
disruption of celiac artery | 96
gastroduodenal artery arising from superior mesenteric artery | 96
gastroscopy | 216
patchy mucosal necrosis | 216
conservative treatment | 216
fever 39 °C | 552
pain in stomach | 552
white blood cell count 34,000/mm3 | 552
C reactive protein 13.4 mg/dL | 552
CT scan | 552
air in gastric wall | 552
intra-abdominal free air | 552
gastric necrosis | 552
emergency surgery | 552
total gastrectomy | 552
Roux-en-Y reconstruction | 552
histological findings of stomach | 552
diffuse necrotic changes | 552
inflammatory cell infiltrations | 552
no invasive fungal infection | 552
leakage on duodenal stump | 696
continuous tube drainage | 696
sepsis | 720
multidrug-resistant Pseudomonas aeruginosa infection | 720
disseminated intravascular coagulation | 720
death | 1680