26 years old | 0
male | 0
admitted to the hospital | 0
height: 180 cm | 0
weight: 74 kg | 0
kidney transplant | -18960
end-stage kidney disease | -28800
immunosuppression | 0
mycofenolate sodium | 0
methylprednisolone | 0
estimated glomerular filtration rate (eGFR) 35.9 mL/min/1.73 m2 | 0
proteinuria 117 mg/d | 0
chronic kidney transplant disease stage 3bA1 | 0
status post vascular rejection | -18960
chronic calcineurin-inhibitor toxicity | -18960
new-onset headache | 0
blurred vision | 0
cranial CT- and MRI scans | 0
several contrast-enhancing intracerebral lesions | 0
perifocal edema | 0
methylprednisolone therapy stopped | 0
dexamethasone administered | 0
brain edema | 0
transmitted to the university department of Nephrology | 24
transmitted to the department of Neurosurgery | 48
brain biopsy | 72
diagnosis of cerebral PTLD | 72
diffuse large B-cell lymphoma | 72
positive for Ebstein-Barr virus | 72
initial chemotherapy regime | 120
high-dose cytarabin | 120
Rituximab | 120
MRI scan confirmed complete remission of PTLD | 240
impairment of the transplant function aggravated | 240
eGFR 25.4 mL/min/1.73 m2 | 240
cytomegalovirus (CMV) reactivated | 480
pneumocystis jirovecii pneumonia | 480
chemotherapy changed to Rituximab | 480
antiviral and antibiotic therapy | 480
dose of mycofenolate sodium tapered | 480
generalized seizure | 720
cerebral MRI scan demonstrated the recurrence of PTLD | 720
HDMTX therapy | 720
Leukovorine | 720
Rituximab | 720
vigorous hydration | 720
HFHD | 744
dialysis procedures started | 744
MTX-level measurements | 744
nadir of leucocytes | 840
severe CMV- and E.coli pneumonia | 936
sepsis | 936
acute kidney transplant failure | 936
transmission to an intensive care unit | 936
invasive ventilation | 936
sepsis managed | 1008
follow up cerebral MRI scan | 1104
small regredience of PTLD | 1104
cerebral radiation | 1104
no relevant response of the disease | 1176
discharged | 1200