64 years old | 0
female | 0
hypertension | 0
hypothyroidism | 0
tobacco use disorder | 0
takotsubo cardiomyopathy | 0
recovered ejection fraction | 0
stroke | 0
acute abdominal pain | 0
nausea | -48
vomiting | -48
dry mucous membranes | 0
periumbilical abdominal tenderness | 0
no peritoneal signs | 0
temperature 36.4 °C | 0
blood pressure 65/34 mmHg | 0
heart rate 78 bpm | 0
oxygen saturation 96% | 0
hemoglobin 12.0 g/dL | 0
white blood cell count 19,890 μL | 0
lactic acid level 3.4 mmol/L | 0
creatinine 2.65 mg/dL | 0
BUN 36 mg/dL | 0
CO2 22mEq/L | 0
voluminous non-bloody diarrhea | 0
CT abdomen and pelvis without contrast | 0
generalized colonic thickening | 0
no obvious transition point | 0
moderate fluid distension | 0
ascending colon distension | 0
transverse colon distension | 0
splenic flexure distension | 0
concern for stricture proximal descending colon | 0
stool Clostridium Difficile toxin negative | 0
fecal occult blood test positive | 0
septic shock diagnosis | 0
infectious colitis | 0
blood cultures pending | 0
fluid resuscitation | 0
piperacillin-tazobactam | 0
ICU admission | 0
vasopressor support | 0
colorectal surgery consultation | 0
gastroenterology consultation | 0
hemodynamic stability | 0
colonoscopy deferred | 0
second day hospitalization | 48
renal function improved | 48
repeat CT abdomen and pelvis with IV contrast | 48
pancolonic thickening | 48
left side more marked involvement | 48
fecal calprotectin 1190 μg/mg | 48
fecal lactoferrin positive | 48
normal stool culture | 48
blood cultures gram variable rods | 48
erythrocyte sedimentation rate 105 mm/h | 48
C-reactive protein 24 mg/dL | 48
D-dimer >20 μg/mlFEU | 48
third day hospitalization | 72
downgraded to general medical floor | 72
colonoscopy performed | 72
scattered severe mucosal changes | 72
altered vascularity | 72
congestion | 72
friability | 72
granularity | 72
mucus | 72
deep ulcerations | 72
ascending colon involvement | 72
transverse colon involvement | 72
descending colon involvement | 72
sigmoid colon involvement | 72
severe ischemic colitis | 72
endoscopic biopsies | 72
pancolonic mucosal ulcerations | 72
transverse colon most severe | 72
descending colon most severe | 72
rectal sparing | 72
Cytomegalovirus immunostaining negative | 72
MRI angiography | 72
no high grade stenosis celiac artery | 72
no high grade stenosis superior mesenteric artery | 72
no high grade stenosis inferior mesenteric artery | 72
diarrhea resolved | 168
abdominal pain continued | 168
nausea continued | 168
vomiting continued | 168
seventh day hospitalization | 168
blood cultures positive Fusobacterium Necrophorum | 168
piperacillin-tazobactam continued | 168
colorectal surgery consultation against surgery | 168
total colectomy deferral | 168
ileostomy deferral | 168
discharge three weeks after admission | 504
bowel movements normalizing | 504
tolerating low residue diet | 504
readmitted one week after discharge | 672
recurrent bloody diarrhea | 672
vancomycin-resistant Enterococcus bacteremia | 672
stabilized | 672
discharged with gastroenterology follow-up | 672
returned to hospital | 672
abdominal pain | 672
voluminous diarrhea | 672
severe anemia | 672
repeat CT angiogram abdomen and pelvis | 672
persistent diffuse colonic thickening | 672
no pneumatosis | 672
no vascular occlusion | 672
antineutrophil cytoplasmic antibodies negative | 672
persistent ischemic bowel disease | 672
surgical consultation deferred | 672
monitoring for symptom improvement | 672
colonoscopy plan after discharge | 672
repeat colonoscopy four months after initial presentation | 2880
deep ulcerations | 2880
serpentine ulcerations | 2880
continuous pattern | 2880
circumferential pattern | 2880
transverse colon involvement | 2880
sigmoid colon involvement | 2880
rectal sparing | 2880
IBD diagnosis | 2880
steroids prescribed | 2880
biologic therapy plan | 2880
died a few months later | N/A
no autopsy | N/A
