60 years old | 0
male | 0
admitted to the hospital | 0
syncope | 0
received second dose of BNT162b2 COVID-19 vaccine | -48
first vaccination administered | -504
fever of 38°C | -24
malaise | -24
decreased urine output | 0
right leg edema | 0
nausea | 0
dizziness | 0
dyspnea on exertion | 0
lost consciousness | 0
taken to emergency department | 0
awake and alert | 0
blood pressure 97/50 mmHg | 0
pulse rate 114/min | 0
body temperature 36.0°C |$0
respiratory rate 12 breaths/min | 0
percutaneous oxygen saturation 97% | 0
generalized pitting edema in legs | 0
elevated white blood cell count (12,000 /μL) | 0
hemoglobin 22.2/dL | 0
serum creatinine 1.51 mg/dL | 0
no proteinuria | 0
no hematuria | 0
no urinary casts | 0
normal chest radiography | 0
normal electrocardiography | 0
admitted to intensive care unit | 0
aggressive fluid therapy | 0
urine output increased (6,000 mL/day) | 24
blood pressure stabilized | 24
hemoconcentration improved | 24
hospitalized for 5 days | 0
discharged | 120
previous episodes: first episode 12 years ago | -105216
common cold-like symptoms | -105216
nausea and vomiting | -105216
pain and swelling in lower extremities | -105216
oliguria | -105216
hypotension | -105216
hemoconcentration | -105216
hospitalized for 36 days | -105216
fluid therapy | -105216
antimicrobial therapy | -105216
diagnosed with sepsis of unknown origin | -105216
second episode 4 years after first | -87696
preceded by cold-like symptoms | -87696
nausea | -87696
oliguria | -87696
swelling in lower extremities | -87696
discharged within 4 days | -87696
diagnosed with acute renal failure of unknown origin | -87696
third episode 5 years after second | -63120
left leg swelling | -63120
decrease in urine output | -63120
generalized body edema | -63120
nausea | -63120
dizziness | -63120
dyspnea on exertion | -63120
hypotension | -63120
laboratory data: inflammatory response | -63120
hemoconcentration | -63120
kidney dysfunction | -63120
admitted to intensive care unit | -63120
aggressive fluid therapy | -63120
urine output increased | -63120
blood pressure stabilized | -63120
hemoconcentration improved | -63120
hospitalized for 9 days | -63120
discharged | -63120
IgG-κ-type M-proteinemia | -63120
small JAK2 mutations | -63120
diagnosed with SCLS | -63120
fourth episode after COVID-19 vaccine | 0
highly sensitive Troponin I low | 0
brain natriuretic peptide low | 0
soluble interleukin-2 receptor not elevated | 0
C4 normal | 0
C1 elastase inhibitors normal | 0
negative blood culture | 0
negative anti-streptolysin O antibody | 0
negative antinuclear antibody | 0
negative anti-glomerular basement membrane antibody | 0
negative antineutrophil cytoplasmic antibody | 0
negative rheumatoid factor | 0
diagnosed with fourth attack of SCLS | 0
started oral terbutaline and theophylline prophylaxis | 0
no further SCLS episodes for 1 year | 0
no Conflict of Interest (COI) | 0
