63 years old | 0
female | 0
chronic hepatitis B-related cirrhosis | -87600
Child-Pugh class A status | -87600
undetectable HBV DNA | -87600
normal ALT levels | -87600
type II diabetic mellitus | -87600
hypertension | -87600
hepatocellular carcinoma | -17520
AJCC/TNM stage II | -17520
BCLC stage B | -17520
transarterial chemoembolization | -17520
contrast-enhanced CT | -876
two tumors at segment 5 | -876
two new poorly enhanced nodules in segments 2 and 8 | -876
no extrahepatic metastasis | -876
no major vascular invasion | -876
radiofrequency ablation | 0
ultrasound-guided RFA | 0
general anesthesia | 0
acute onset of fever | 6
chills | 6
dyspnea | 6
abdominal pain | 6
body temperature 39.6°C | 6
heart rate 130 beats per min | 6
blood pressure 90/46 mmHg | 6
WBC 24,600/μL | 6
neutrophil predominant 85% | 6
hyperlactatemia 65.4 mg/dL | 6
CRP 51 mg/L | 6
AST 239 U/L | 6
ALT 80 U/L | 6
total bilirubin 1.1 mg/dL | 6
albumin 3.5 g/dL | 6
INR 1.82 | 6
Cr 1.48 mg/dL | 6
ammonia 255 μg/dL | 6
abdominal ultrasound | 6
hyperechoic change with air formation | 6
contrast-enhanced CT | 6
necrotic changes with air component | 6
intra-tumoral abscess formation | 6
septic shock | 6
transferred to intensive care unit | 6
oxygen supplement | 6
aggressive fluid resuscitation | 6
empirical antibiotic with Flomoxef | 6
ultrasound-guided aspiration | 6
pus discharge | 6
packed red blood cell transfusion | 6
fresh frozen plasma transfusion | 6
liver abscess culture Clostridium perfringens | 72
blood culture Clostridium perfringens | 72
susceptible to Flomoxef | 72
sessions of ultrasound-guided aspiration | 72
antibiotic course completed | 720
infection under control | 720
discharged | 720
complete ablation of treated tumors | 720
no local tumor recurrence | 720
