52 years old | 0
    female | 0
    visited emergency room | 0
    abdominal pain | -48
    nausea | -48
    vomiting | -48
    increased ALT | -840
    alanine aminotransferase (ALT) 320 U/mL | -840
    health screening test | -840
    anti-nuclear antibody 1:1280 | -840
    anti-mitochondrial antibody positive | -840
    immunoglobulin G 1577 mg/dL | -840
    coarse liver surface | -840
    chronic liver disease | -840
    liver biopsy | -840
    overlap syndrome | -840
    autoimmune hepatitis | -840
    ursodeoxycholic acid | -840
    prednisolone 40 mg daily | -840
    ursodeoxycholic acid maintained | -840
    prednisolone reduced by 10 mg every week | -840
    prednisolone reduced to 5 mg | -144
    azathioprine 50 mg | -144
    mild heartburn | -48
    abdominal pain worsened | -24
    nausea increased | -24
    vomiting increased | -24
    diarrhea | -24
    blood pressure 130/80 mmHg | 0
    fever 37.6°C | 0
    tachycardia 110 beats/min | 0
    tachypnea 30 breaths/min | 0
    abdominal tenderness epigastric to left upper quadrant | 0
    abdomen slightly hard | 0
    no rebound tenderness | 0
    white blood cells reduced 700/µL | 0
    platelets reduced 61000/µL | 0
    neutrophil 5% | 0
    C-reactive protein 14.35 mg/dL | 0
    systemic infection suspected | 0
    aspartate aminotransferase 347 U/L | 0
    ALT 52 U/L | 0
    gamma glutamyl transferase 458 U/L | 0
    prothrombin time INR 1.2 | 0
    CT layered wall thickening stomach fundus and upper body | 0
    CT air in stomach wall | 0
    CT decreased mucosal enhancement | 0
    necrotizing gastritis | 0
    septic shock | 0
    blood pressure decreased <80 mmHg | 0.5
    transferred to ICU | 0.5
    intravenous hydration | 0.5
    antibiotic treatment | 0.5
    blood pressure increased 127/95 mmHg | 2
    inotropics norepinephrine | 2
    fluid treatment | 2
    heart rate slowed | 3
    echocardiography | 3
    stress-induced cardiomyopathy | 3
    ejection fraction <10% | 3
    extracorporeal membrane oxygenation preparation | 3
    sudden cardiac arrest | 3.5
    pulseless electrical activity | 3.5
    cardiopulmonary resuscitation | 3.5
    extracorporeal membrane oxygenation applied | 3.5
    death | 4
    