41 years old | 0
male | 0
originally from West Africa | 0
questionable history of ventriculoseptal defect | 0
presented with worsening exertional dyspnea | -6*168
presented with palpitations | -6*168
presented with loss of appetite | -6*168
presented with lower extremity edema | -6*168
presented with 30 pounds weight loss over 6 weeks | -6*168
temperature 98.8°F | 0
blood pressure 104/50 mm Hg | 0
heart rate 120/min | 0
respiratory rate 18/min | 0
oxygen saturation 98% on room air | 0
chronically ill cachexic male | 0
BMI 21 kg/m2 | 0
jugular venous distension | 0
bilateral rales | 0
tachycardia | 0
RV heave | 0
4/6 pan-systolic murmur | 0
palpable thrill throughout the precordium | 0
blood cultures obtained for suspected endocarditis | 0
empiric intravenous antibiotics started | 0
initial transthoracic echocardiogram | 0
subsequent transesophageal echocardiogram demonstrated large mass attached to aortic valve leaflet | 0
severe aortic regurgitation with holodiastolic flow reversal in the aorta | 0
mass attached to flail anterior mitral valve leaflet resulting in severe mitral regurgitation | 0
mass attached to pulmonic valve | 0
significant pulmonic regurgitation | 0
severe pulmonary hypertension with Pulmonary Artery Systolic Pressure 65 mm Hg | 0
dilatation of the aortic root | 0
fistula between aortic sinus and RV outflow tract | 0
blood culture revealed gram-positive cocci identified as Abiotrophia species | 24
transferred to tertiary care center | 24
underwent right heart catheterization demonstrating elevated filling pressures | 24
low cardiac index | 24
shunt fraction 2.1 | 24
emergent surgery revealed aortic root abscess | 24
underwent prophylactic grafting of left anterior descending coronary artery | 24
prophylactic grafting of obtuse marginal artery | 24
bio-prosthetic pulmonary valve replacement | 24
bio-prosthetic mitral valve replacement | 24
closure of congenital VSD | 24
closure of aorto-RV fistula using bovine pericardial patches | 24
aortic root replacement with porcine root prosthesis | 24
post-operative atrial fibrillation | 24
started on amiodarone therapy | 24
intravenous penicillin | 24
gentamycin during hospitalization | 24
transesophageal echocardiogram post intervention showed mild left ventricular dysfunction | 24
ejection fraction 45% | 24
competent bio-prosthetic valves | 24
repeat blood cultures remained negative | 24
discharged on intravenous vancomycin via peripherally inserted central catheter | 24
