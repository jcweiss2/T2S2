37 years old | 0
female | 0
Graves' disease | -1095
methimazole 120 mg/day | -1095
discontinued methimazole | -780
hyperthyroidism symptoms | -24
palpitations | -24
sweating | -24
easy fatigue | -24
propylthiouracil 900 mg/day | -24
switched to methimazole 90 mg/day | -12
high free thyroxine (FT4) levels | -12
methimazole increased to 120 mg/day | -12
pregnancy confirmed | -4
methimazole 120 mg/day | -4
FT4 level 8.8 ng/L | -4
did not visit hospital | -4
visited hospital at 12 weeks pregnant | 0
FT4 level 0.11 ng/L | 0
methimazole reduced to 60 mg/day | 0
levothyroxine (LT4) 50 µg/day | 0
methimazole reduced to 40 mg/day | 16
methimazole reduced to 20 mg/day | 20
ultrasound detected gastroschisis | 28
referred to RSCM | 28
ultrasound confirmed gastroschisis | 33
cesarean section | 36
Bogota bag placement | 36
baby died of septic shock | 56
gastroschisis | 28
restricted fetal growth | 33
nuchal cord | 33
DRESS syndrome | -672 
fever | -72 
rash | -72 
acne | -672 
minocycline | -672 
increased WBC count | 0 
eosinophilia | 0 
systemic involvement | 0 
diffuse erythematous or maculopapular eruption | 0 
pruritis | 0 
discharged | 24