26 years old | 0
female | 0
admitted to the hospital | 0
jaundice | -120
intermittent epigastric pain | -120
weight loss | -120
pruritus | -120
tea-colored urine | -120
obstructive jaundice | -120
choledocholithiasis | -120
icteric sclerae | 0
soft abdomen | 0
nondistended abdomen | 0
nontender abdomen | 0
generalized jaundice | 0
intrahepatic ductal dilatation | 0
bile duct sludges | 0
hepatobiliary tuberculosis | 0
ERCP | 0
cannulation | 0
cholangiogram | 0
common hepatic duct stricture | 0
dilation of CHD stricture | 0
partial sphincterotomy | 0
biliary stent insertion | 0
TB-PCR testing | 0
abdominal pain | 24
fever | 48
tachycardia | 48
epigastric tenderness | 48
post-ERCP pancreatitis | 48
elevated amylase level | 48
normal lipase level | 48
hypotension | 72
generalized abdominal pain | 72
abdominal distension | 72
direct tenderness | 72
rebound tenderness | 72
elevated WBC count | 72
prothrombin time elevation | 72
PT-INR elevation | 72
activated partial thromboplastin time elevation | 72
broad-spectrum antibiotics | 72
Vitamin K infusion | 72
FFP transfusion | 72
norepinephrine | 72
exploratory laparotomy | 96
duodenal perforation | 96
biliary stent migration | 96
peritonitis | 96
duodenorrhaphy | 96
primary repair | 96
peritoneal lavage | 96
tube jejunostomy | 96
persistent hypotension | 120
supraventricular tachycardia | 120
death | 120