15 years old | 0
male | 0
Saudi Arabian | 0
admitted to the emergency department | 0
vomiting | -72
headache | -72
hemoptysis | -72
shortness of breath | -72
no past medical illness | 0
referred from a secondary care hospital | -24
intubated | -24
decreased oxygen saturation | -24
initial diagnosis of meningitis | -24
initial diagnosis of acute respiratory distress syndrome | -24
physical examination | 0
intubated | 0
SpO2 100% | 0
temperature 37.2°C | 0
heart rate 132 bpm | 0
blood pressure 135/95 mmHg | 0
crepitus at both upper regions of the chest | 0
abdominal examination did not reveal any clinical abnormality | 0
cardiovascular examination did not reveal any clinical abnormality | 0
laboratory findings of blood count were not significant | 0
neck and chest contrast-enhanced CT | 0
large pre-vertebral collection of abscess | 0
abscess in the retropharyngeal space | 0
extension into the posterior mediastinum | 0
low attenuation density with peripheral rim enhancement | 0
mass effect on adjacent structures | 0
anterior displacement of the pharynx | 0
anterior displacement of the oesophagus | 0
anterior displacement of the trachea | 0
conservative management | 0
no improvement of his condition | 24
surgical intervention | 24
cervical approach | 24
longitudinal incision | 24
drainage of pus | 24
about 200 cc of pus was drained | 24
improvements in his condition | 48
C/S of the swab showed Ochrobactrum anthropi | 48
sensitive to imipenem | 48
sensitive to cefepime | 48
sensitive to amikacin | 48
sensitive to gentamicin | 48
sensitive to ciprofloxacin | 48
extubated | 48
recovered well | 48
discharged | 192
no complications | 192
follow-up | 384
well at a 2-month follow-up | 384