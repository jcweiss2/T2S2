4-year-old | 0
    boy | 0
    presented to the institution | 0
    headaches | -48
    vomiting | -48
    tonic-clonic seizure | -48
    subacute hydrocephalus | 0
    tested positive for COVID-19 | 0
    asymptomatic | 0
    external ventricular drain placed | 0
    awake | 0
    alert | 0
    stable neurological examination | 0
    postprocedural CT demonstrated satisfactory catheter placement | 0
    interval reduction in ventriculomegaly | 0
    MRI demonstrated membrane obstructing right foramen of Monro | 0
    congenital malformation | 0
    hydrocephalus | 0
    magnetic resonance venography | 24
    cervical spine MRI | 24
    new left-sided hemiparesis | 72
    repeat MRI | 72
    MRA of the brain | 72
    new diffusion restriction indicative of infarctions | 72
    both hemispheres | 72
    thalami | 72
    basal ganglia | 72
    MRA showed focal narrowing and irregularity | 72
    distal left carotid artery | 72
    left M1 and M2 | 72
    right postbifurcation M1 segments | 72
    right A1 segment | 72
    left P2 | 72
    right P1 segments | 72
    concerning for vasculitis or vasospasm | 72
    stroke workup initiated | 72
    echocardiography confirmed normal heart | 72
    no evidence of emboli | 72
    coagulopathy workup | 72
    D-dimer levels normal | 72
    protein S level mildly low | 72
    homozygous 4G/4G for PAI-1 gene | 72
    CSF infectious studies ordered | 72
    varicella zoster virus | 72
    herpes simplex viruses 1, 2, 6 | 72
    Haemophilus influenzae | 72
    Neisseria meningitidis | 72
    CSF PCR tests negative | 72
    CSF cultures sterile | 72
    SARS-CoV-2 IgG antibodies positive | 72
    SARS-CoV-2 PCR positive on four serum samples | 72
    no fever | 0
    no respiratory symptoms | 0
    CSF negative for SARS-CoV-2 | 72
    elevated levels of proinflammatory cytokines | 72
    IL-6 elevated | 72
    IL-8 elevated | 72
    empirical treatment with steroids initiated | 72
    no additional infarcts after treatment | 72
    intracranial pressure monitoring with EVD | 72
    patent external CSF diversion | 72
    treatment for provoked vasculitis | 72
    ventricular endoscopy | 168
    membranous obstruction at right foramen of Monro | 168
    septum pellucidotomy performed | 168
    CSF flow normalization | 168
    no surgical complications | 168
    external CSF drainage continued | 168
    drain weaned and removed | 168
    surveillance MRI/MRA confirmed resolution of vascular findings | 168
    no further infarcts | 168