28 years old | 0
male | 0
Caucasian | 0
police officer | 0
admitted to the hospital | 0
fever | -168
acute diarrhea | -168
poor oral intake | -168
hemophagocytic lymphohistiocytosis (HLH) | -672
fever | -672
pancytopenia | -672
splenomegaly | -672
bone marrow (BM) biopsy | -672
Epstein–Barr virus (EBV) titers | -672
dexamethasone | -672
intravenous (IV) immunoglobulin | -672
etoposide | -672
cyclosporine | -672
surveillance imaging studies | -672
computerized tomography chest | -672
abdomen | -672
pelvis | -672
positron emission tomography scan | -672
no evidence of malignancy | -672
good response to therapy | -672
febrile neutropenia | -24
IV vancomycin | -24
cefepime | -24
transferred to hospital | -24
temperature 38.5°C | 0
blood pressure 116/60 mmHg | 0
heart rate 80 beats/min | 0
weight 120 kg | 0
2-cm left cervical lymph node | 0
serum creatinine 2.6 mg/dL | 0
arterial blood gas (ABG) | 0
pH 7.23 | 0
pCO2 24 mmHg | 0
pO2 101 mmHg | 0
HCO3 10 mmol/L | 0
anion gap metabolic acidosis | 0
respiratory compensation | 0
urinalysis | 0
granular casts | 0
renal epithelial cells | 0
acute tubular necrosis | 0
cervical lymph node biopsy | 0
repeat BM biopsy | 0
peripheral T-cell lymphoma | 0
stool positive for Clostridium difficile | 0
diagnosis of peripheral T-cell lymphoma | 0
relapsing HLH | 0
C. difficile colitis | 0
acute kidney injury | 0
lactic acidosis | 0
treated with oral vancomycin | 0
dexamethasone | 0
etoposide | 0
basiliximab | 0
cyclosporin | 0
alemtuzumab | 0
nitrogen mustard | 0
rituximab | 0
septic shock | 48
multiorgan system failure | 48
vasopressors | 48
continuous venovenous hemofiltration (CVVH) | 48
replacement fluid rate 3.6 L/h | 48
anticoagulant citrate dextrose solution A | 48
hyperkalemia | 56
acid–base status | 56
hemofiltration rate increased to 7 L/h | 56
high bicarbonate replacement fluid | 56
low-potassium replacement fluid | 56
persistent hyperkalemia | 64
severe lactic acidosis | 64
intermittent hemodialysis (IHD) | 64
CVVHD | 64
volume overload | 64
hypoxemia | 64
CVVHD with dialysate rate of 7 L/h | 72
CVVH with replacement fluid at 5 L/h | 72
two machines | 72
volume status stabilized | 144
hemodynamics stabilized | 144
decreasing requirements for vasopressors | 144
improved serum lactate level | 144
CVVHD stopped | 144
CVVH continued | 144
hemofiltration rate of 5 L/h | 144
one machine | 144
plasma lactate level continued to decrease | 168
lactate clearance evaluation | 168
lactate concentrations in samples of plasma and effluent | 168
calculated lactate clearance | 168
79 mL/min | 168
0.56 mmol/min | 168
effluent fluid lactate | 168
6.2 mmol/L | 168
CVVH output | 168
91 mL/min | 168
plasma lactate | 168
7.1 mmol/L | 168
lactate clearance calculated | 168
plasma lactatefilter | 168
6.2 mmol/L | 168
total CVVH replacement fluid rate reduced to 3.6 L/h | 192
plasma lactic acid level continued to decrease | 192
5.6 mmol/L | 192
improvement in metabolic acidosis | 192
ABG | 192
pH of 7.35 | 192
pCO2 of 35 mmHg | 192
HCO3 of 18 mmol/L | 192
weaned off of vasopressors | 192
improvement in mental status | 192
massive lower gastrointestinal bleeding | 216
severe thrombocytopenia | 216
ischemic colitis | 216
palliative treatment | 216
passed away | 576