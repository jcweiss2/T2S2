21 years old | 0
woman | 0
Caucasian | 0
admitted to the hospital | 0
altered mental status | 0
lethargic | 0
plasma glucose 20 mg/dl | 0
hospitalized | 0
dextrose infusion | 0
10% dextrose in water | 0
hypoglycemic | 0
capillary glucose 50-60 mg/dl | 0
transferred to our facility | 0
suspicion of insulinoma | 0
medical records revealed treatment for hypoglycemia as a neonate | -20160
repeated episodes of seizures | -4032
syncope | -4032
dizziness | -4032
headaches | -4032
palpitations | -4032
sweating | -4032
symptoms since birth | -20160
intermittent symptoms | -20160
varying severity | -20160
seizure-free | -20160
without syncopal episodes | -20160
syncopal episode at age 17 | -20160
inpatient hypoglycemia evaluation | -20160
blood glucose 47 mg/dl after 2 h fasting | -20160
proinsulin levels 10.4 to 84.1 pmol/l | -20160
C-peptide level 3.1 ng/ml | -20160
negative insulin antibodies | -20160
negative sulfonylurea screen | -20160
MRI abdomen showed no insulinoma | -20160
genetic studies revealed Val452 Leu activating mutation of GCK gene | -20160
treated with diazoxide | -20160
discharged home on oral diazoxide 250 mg daily | -20160
discontinued diazoxide due to hirsutism and fluid retention | -20160
current admission | 0
treated with dextrose boluses | 0
blood glucose level remained low | 0
continuous infusion of 5% dextrose | 0
transfer to intensive care unit | 0
fasting blood glucose low | 0
postprandial blood glucose low | 0
review of medication list showed no implicating drugs | 0
no additional work-up | 0
placed on octreotide 200 µg subcutaneously twice daily | 0
diazoxide suspension 100 mg three times a day | 0
consultation with pediatric endocrinologist | 0
neuroglycopenic symptoms of hypoglycemia improved | 0
hypoglycemia improved with capillary glucose 55-110 mg/dl | 0
discharged | 24
emphasized compliance with treatment | 24
follow-up with endocrinologist | 24
congenital hyperinsulinism (CHI) | -20160
activating mutation of GCK gene | -20160
rare genetic cause | -20160
recurrent hypoglycemia | -20160
persistent hypoglycemia | -20160
insulinoma ruled out | -20160
negative MRI abdomen | -20160
negative autoimmune work-up | -20160
negative drug screen | -20160
negative fasting studies | -20160
negative pancreatic arterial calcium stimulation test (SPACI) | -20160
non-insulinoma pancreatogenous hypoglycemia syndrome (NIPHS) | -20160
effective treatment with diazoxide and octreotide | -20160
transition to adulthood care | -20160
coordination with pediatric endocrinologist | 0
improved hypoglycemia | 24
discharge with improved glucose levels | 24
emphasized treatment compliance | 24
emphasized follow-up | 24
rare genetic diagnosis | -20160
congenital GCK mutation | -20160
de novo mutation considered | 0
family history of hypoglycemia | -20160
lifelong low plasma glucose | -20160
increased BMI | -20160
positive response to octreotide | 0
transition of care importance | 0
rare disease management | 0
cost-effective patient information dissemination | 0
conflict of interest | 0
no funding or benefits | 0
