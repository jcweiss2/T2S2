70 years old | 0 | 0 
male | 0 | 0 
emergency esophageal diversion | -720 | -720 
injury to the cervical esophagus | -720 | -720 
spinal surgery | -720 | -720 
gastric pull-up procedure | -504 | -504 
postoperative anastomotic leakage | -504 | -504 
endoscopy | -504 | -504 
esophageal stent | -504 | -168 
discharged | -168 | -168 
local cervical infection | -168 | -168 
sepsis | -168 | -168 
transfer to tertiary university hospital | -168 | -168 
arterial hypertonus | 0 | 0 
non-active smoking status | 0 | 0 
ischemic stroke | 0 | 0 
incomplete senso-motoric hemiparesis | 0 | 0 
thyroidectomy | 0 | 0 
open prostatectomy | 0 | 0 
prostate cancer | 0 | 0 
malnutrition | 0 | 0 
systemic inflammation | 0 | 0 
jugular and cervical phlegmon | 0 | 0 
hemoglobin level of 6.7 g/dL | 0 | 0 
white blood cell count of 6400 cells/μL | 0 | 0 
platelet count of 210 × 10^3/μL | 0 | 0 
creatinine level of 0.76 mg/dL | 0 | 0 
unremarkable liver and cholestasis parameters | 0 | 0 
albumin level of 2.8 g/dL | 0 | 0 
chest computed tomography scan | 0 | 0 
endoscopy | 0 | 0 
dislodged esophageal stent | 0 | 0 
esophageal perforation | 0 | 0 
infected cavity | 0 | 0 
esophageal stenosis | 0 | 0 
stent removal | 0 | 0 
endoscopic vacuum therapy | 24 | 168 
EsoSponge system | 24 | 168 
jugular and cervical phlegmon resolved | 168 | 168 
repeated endoscopic balloon dilatation | 168 | 168 
subtotal esophageal resection | 168 | 168 
reconstruction using a free-jejunal graft interposition | 168 | 168 
CT angiography | 168 | 168 
partial sternotomy | 168 | 168 
laparotomy | 168 | 168 
jejunal segment harvested | 168 | 168 
left carotid artery and left jugular vein used as recipient vessels | 168 | 168 
graft implanted in an isoperistaltic position | 168 | 168 
cervical anastomosis performed in an end-to-end fashion | 168 | 168 
upper mediastinal gastro-jejunostomy performed in a side-to-side fashion | 168 | 168 
upper sternum resected | 168 | 168 
soft tissue defect covered with a sternocleidomastoid muscle flap | 168 | 168 
abdominal reconstruction achieved by an end-to-end jejunojejunostomy | 168 | 168 
postoperative course uneventful | 168 | 336 
oral alimentation reestablished | 168 | 336 
daily speech therapy | 168 | 336 
anastomotic healing confirmed radiologically and endoscopically | 336 | 336 
patient transferred to a rehabilitation clinic | 336 | 336 
esophagectomy with diversion and later reconstruction | 0 | 0 
anastomotic complications following gastric pull-up procedures | 0 | 0 
endoscopic management of leaks, fistulas and stenosis | 0 | 0 
esophageal reconstruction with a free jejunal graft | 168 | 168 
salvage option after failed gastric pull-up | 168 | 168 
complication rate in excess of 70% | 0 | 0 
free jejunal grafts | 168 | 168 
transient ischemia | 168 | 168 
advanced microsurgical skills for swift revascularization | 168 | 168 
challenging surgical site environment | 168 | 168 
multidisciplinary approach | 0 | 336 
interventional endoscopists and surgeons | 0 | 336 
successful salvage management | 336 | 336 
restoration and reconstruction of the esophagus | 336 | 336 
patients with chronic postoperative fistulas or stenoses of the esophagus | 0 | 0 
specialized centers | 0 | 0 
written consent for publication | 0 | 0 
CARE Checklist (2016) | 0 | 0 
manuscript source | 0 | 0 
peer-review started | 0 | 0 
first decision | 0 | 0 
article in press | 0 | 0 
specialty type | 0 | 0 
country/territory of origin | 0 | 0 
peer-review report’s scientific quality classification | 0 | 0 
P-Reviewer | 0 | 0 
S-Editor | 0 | 0 
L-Editor | 0 | 0 
P-Editor | 0 | 0