53 years old | 0
female | 0
admitted to hospital | 0
dizziness | -168
shortness of breath | -168
increasing chest pressure | -168
urinary tract infection | -168
sulfamethoxazole-trimethoprim | -168
ceftriaxone | -168
ciprofloxacin | -168
lethargy | 0
temperature 36.7°C | 0
blood pressure 104/88 mmHg | 0
heart rate 175 beats per minute | 0
respiratory rate 21 breaths per minute | 0
oxygen saturation 98% | 0
atrial fibrillation | 0
rapid ventricular rate | 0
brain natriuretic peptide elevated | 0
troponin I value 0.1 ng/mL | 0
heparin infusion | 0
diltiazem infusion | 0
lactic acidosis | 0
acute kidney injury | 0
thrombocytopenia | 0
thickened and restricted mitral valve | 0
large vegetation on posterior leaflet | 0
partial flail | 0
severe regurgitation | 0
aortic valve thickened | 0
perforation of non-coronary cusp | 0
ejection fraction normal | 0
right ventricular systolic pressure elevated | 0
right ventricular overload | 0
empiric vancomycin | 0
piperacillin/tazobactam | 0
ampicillin | 24
gentamycin | 24
severe thrombocytopenia | 24
bacteremia | 24
acute heart failure | 168
emergent intubation | 168
mechanical ventilation | 168
ampicillin/sulbactam | 168
daptomycin | 168
septic embolization to left lower limb | 168
critical ischemia | 168
splenic infarcts | 168
left lower extremity thrombectomy | 168
four-compartment fasciotomy | 168
surgical replacement of mitral and aortic valves | 168
intraoperative transesophageal echocardiogram | 168
enlarged left atrium | 168
thrombi in left and right atrial appendages | 168
aortic valve thinned | 168
severe aortic insufficiency | 168
posterior leaflet of mitral valve eroded | 168
micro-abscesses in posterior annulus | 168
nodular extension up endocardium | 168
inhaled epoprostenol | 168
elevated pulmonary artery pressures | 168
postoperative course uncomplicated | 240
blood culture pathogen identification | 240
Abiotrophia defectiva | 240
Gram-positive bacilli | 240
discharged from intensive care unit | 336
broad spectrum antibiotics | 336
total 6 weeks antibiotics | 504
urinary tract infection caused by Abiotrophia defectiva | -672
hematogenous spread | 0
cardiogenic shock | 0
septic shock | 0
open heart surgery | 168
complex anesthesia management | 168
uncomplicated postoperative course | 240