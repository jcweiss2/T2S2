63 years old | 0
male | 0
admitted to the hospital | 0
dyspnea | -3
central chest pain | -3
chest pain radiated into back | -3
workup for acute coronary syndrome | 0
pulse 94 per minute | 0
BP 135/72 mm Hg | 0
SaO2 97% on air | 0
temperature 37°C | 0
no history of alcohol ingestion | 0
no cardiovascular diseases | 0
no abdominal diseases | 0
no surgical emphysema in supraclavicular fossae | 0
physical examination revealed an acutely ill man | 72
temperature rose to 39 °C | 72
right lower chest region was dull to percussion | 72
decreased breath sound | 72
Chest X-ray demonstrated right pleural effusion | 72
no evidence of pneumomediastinum | 72
no subcutaneous emphysema | 72
diagnostic pleural fluid aspiration | 72
exudates | 72
gram stain negative | 72
culture negative | 72
CT scan demonstrated right sided pneumothorax | 72
extended right sided pleural effusion | 72
small amount of air in mediastinum | 72
hemoglobin concentration 11.5 gm/dl | 72
hematocrit 35.4% | 72
white-cell count 17500/ml | 72
85% neutrophils | 72
platelet count 145,000/ml | 72
serum electrolytes normal | 72
urea nitrogen level 30 mg per deciliter | 72
creatinine level 2.1 mg per deciliter | 72
liver function tests normal | 72
treated with antibiotics | 72
tube thoracostomy | 72
right closed thoracotomy | 72
water-seal drainage | 72
removal of 1500 ml of fluid | 72
treated with ceftriaxone | 72
treated with clindamycin | 72
imipenem added to treatment | 120
vancomycin added to treatment | 120
clinical deterioration | 120
increased respiratory distress | 120
discomfort | 120
fever | 120
delay in chest expansion | 120
chest pain | 120
suspicion of esophageal perforation | 120
underwent right thoracotomy | 120
repair of linear longitudinal tear | 120
marked mediastinal and pleural inflammation | 120
open thoracotomy | 120
surgical repair of esophageal perforation | 120
thoracic window | 120
intravenous vasopressors | 120
mechanical ventilation | 168
respiratory failure | 168
acute kidney failure | 168
pleural empyema | 168
re-operation | 168
died | 408