49 years old | 0
woman | 0
admitted to the emergency department | 0
Glasgow Coma Scale 7/15 | 0
right-sided anisocoria | 0
pupils reactive to light | 0
intubated | 0
thunderclap headache | -24
neck pain | -24
loss of consciousness | -24
computed tomography of the brain | 0
right occipital intracerebral hematoma | 0
subarachnoid hemorrhage Fischer Grade scale IV | 0
brain computed tomography angiography | 0
right 6-mm distal PCA saccular aneurysm | 0
parieto!-occipital artery | 0
splenial artery | 0
emergently operated | 0
right posterior occipital interhemispheric approach | 0
hematoma evacuation | 0
aneurysm clipping | 0
transferred to the intensive care unit | 0
extubated | 72
significant neurological recovery | 72
died | 192
acute respiratory distress syndrome | 192
septic shock | 192
