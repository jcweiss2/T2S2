74 years old | 0
male | 0
end-stage renal disease | 0
admitted to hospital | 0
syncope | -24
returned from cottage | -24
fever | 24
tachycardia | 24
confused | 24
no nuchal rigidity | 24
no jaundice | 24
no cardiorespiratory abnormalities | 24
no lymphadenopathy | 24
no hepatosplenomegaly | 24
no abdominal tenderness | 24
mild anemia | 24
elevation in aspartate transaminase | 24
normal computed tomography scans | 24
working diagnosis of sepsis | 24
started on intravenous piperacillin–tazobactam | 24
started on intravenous vancomycin | 24
high-grade fevers | 48
decreasing level of consciousness | 48
hypotensive | 48
transferred to intensive care unit | 48
intubation | 48
changed anti-infective drugs | 48
started on intravenous acyclovir | 48
started on intravenous ampicillin | 48
started on intravenous ceftriaxone | 48
anemia | 120
thrombocytopenia | 120
transaminitis | 120
hyperferritinemia | 120
suspected hemophagocytic lymphohistiocytosis | 120
normal magnetic resonance imaging of brain | 120
tick discovered on left calf | 120
Ixodes scapularis tick | 120
morulae within granulocytes | 120
started on oral doxycycline | 120
bone marrow aspiration and biopsy | 144
hemophagocytosis | 144
pursued broad infectious work-up | 144
negative blood cultures | 144
negative urine culture | 144
negative serological testing | 144
negative polymerase chain reaction tests | 144
positive serology for Anaplasma phagocytophilum | 168
positive serology for Borrelia burgdorferi | 168
positive serology for Powassan virus | 168
diagnosed with human granulocytic anaplasmosis | 168
diagnosed with hemophagocytic lymphohistiocytosis | 168
diagnosed with Lyme disease | 168
diagnosed with Powassan virus | 168
completed 10-day course of doxycycline | 240
completed 3-week course of ceftriaxone | 240
discharged from hospital | 1320
follow-up 3 months after presentation | 2160
clinically well | 2160
complete resolution of hematologic derangements | 2160