55 years old | 0
woman | 0
admitted to the hospital | 0
abdominal distress | 0
medical history of two kidney transplantations | -6720
IgA nephropathy | -6720
first allograft lost due to chronic allograft rejection | -6720
current allograft functioning with estimated glomerular filtration rate of approximately 60 ml/min per 1.73 m² | 0
computed tomographic scan revealed free intra-abdominal air | 0
sigma perforation (sigma diverticulitis type 2c2) | 0
sigma resection | 0
protective ileostomy | 0
required two more surgical interventions | 24
burst abdomen | 24
presumed peritonitis | 24
initial blood cultures positive with Alistipes onderdonkii | 0
intraoperative cultures grew Klebsiella oxytoca (3-multidrug-resistant gram-negative bacteria pattern) | 0
developed fever | 72
respiratory insufficiency | 72
signs of hemodynamic compromise | 72
switched to mechanical ventilation | 72
norepinephrine required to maintain mean arterial pressure above 60 mm Hg | 72
antibiotic therapy intensified | 72
administered vitamin C 1.5 g i.v. 4 times a day for 4 sequential days (1 dose missed, total dose 22.5 g) | 72
administered vitamin B1 200 mg i.v. 3 times a day for 3 sequential days | 72
urine output progressively declined | 96
plasma creatinine increased | 96
no obvious nephrotoxic medications administered | 96
immunosuppression included tacrolimus | 0
immunosuppression included mycophenolate | 0
immunosuppression included corticosteroids | 0
tacrolimus with fluctuating trough level concentrations (range 2.4–19.3 ng/ml) | 0
urinalysis revealed tubular proteinuria of 750 mg alpha-1-microglobulin per g creatinine | 96
albumin 180 mg per g creatinine | 96
urine microscopy could not detect erythrocytes | 96
urine microscopy could not detect leukocytes | 96
urine microscopy could not detect casts | 96
sonography excluded obstructive uropathy | 96
vascular resistance indices of the kidney allograft within normal range (0.66–0.78) | 96
continuous renal replacement therapy (citrate-based) initiated | 168
acute tubular damage in the context of sepsis | 168
allograft rejection considered unlikely | 168
current kidney allograft a complete HLA match organ | 168
patient had received one kidney allograft in the past | -6720
HLA-sensitized | -6720
performed kidney allograft biopsy | 168
kidney biopsy yielded 8 glomeruli | 168
histologic finding showed severe signs of acute tubular epithelial injury | 168
multifocal intratubular calcium oxalate depositions | 168
one glomerulus globally sclerosed | 168
discrete glomerulitis | 168
moderate peritubular capillaritis (C4d negative) | 168
no double contours of the glomerular basement membranes | 168
no significant mesangial hypercellularity | 168
no significant endocapillary hypercellularity | 168
no crescents | 168
interstitium showed discrete lymphoplasmacellular infiltrates | 168
mild tubulitis (corresponding to borderline changes) | 168
SV40 staining negative | 168
interstitial fibrosis and tubular atrophy amounted to 15% | 168
test for donor-specific antibodies negative | 168
leukocyte count 17,460/µl | 168
hemoglobin concentration 7.2 g/dl | 168
thrombocyte count 443,000/µl | 168
sodium 142 mmol/l | 168
potassium 4.1 mmol/l | 168
calcium, total 2.3 mmol/l | 168
creatinine 0.7 mg/dl | 168
urea 14 mg/dl | 168
procalcitonin 30.0 ng/ml | 168
LDH 186 U/l | 168
tacrolimus trough level 13.0 ng/ml | 168
urine protein ++ | 168
urine hemoglobin negative | 168
urine leukocytes negative | 168
urine protein-creatinine ratio 583 mg/g | 168
urine albumin-creatinine ratio 179 mg/g | 168
urine alpha 1-microglobulin–creatinine ratio 746 mg/g | 168
acute tubular injury | 168
oxalate nephropathy secondary to vitamin C administration | 168
discontinued vitamin C | 168
continued citrate-based continuous renal replacement therapy | 168
urinary output restored | 240
continuous renal replacement therapy terminated | 240
second episode of acute kidney injury | 240
kidney allograft function recovered | 336
estimated glomerular filtration rate approximately 45–50 ml/min per 1.73 m² at 1-year follow-up | 8760
