61 years old | 0
female | 0
type 2 diabetes mellitus | 0
chronic obstructive airway disease | 0
admitted to the hospital | 0
severe community-acquired pneumonia | 0
acute renal failure | 0
renal failure attributed to acute tubular necrosis | 0
sepsis | 0
hypotension | 0
no red cells or casts in urine | 0
renal function remained stable | 0
renal function worsened | 0
fluid overload | 0
haemodialysis | 0
renal function improved | 0
discharged home | 45
readmitted to the intensive care unit | 48
acute pulmonary oedema | 48
skin rash | 48
pulmonary hypertension | 48
splenomegaly | 48
hepatomegaly | 48
bilateral pleural effusion | 48
vasculitis | 48
dysmorphic red cells in urine | 48
proteinuria | 48
hypoalbuminaemia | 48
low complement levels | 48
positive serology for mixed cryoglobulinaemia | 48
renal ultrasound showed normal sized kidneys | 48
renal ultrasound showed normal echotexture | 48
rheumatoid factor weakly positive | 48
HCV RNA negative | 48
autoimmune screens negative | 48
renal biopsy | 48
diffuse mesangiocapillary glomerulonephritis | 48
hyaline capillary thrombi | 48
focal mild endarteritis | 48
cryoglobulinaemic vasculitis | 48
plasma exchange | 48
haemodialysis | 48
prednisolone | 48
cyclophosphamide | 48
good initial response | 72
decrease in cryoglobulin levels | 72
symptomatic improvement | 72
cyclophosphamide discontinued | 72
thrombocytopenia | 72
discharged on prednisolone | 72
renal function normal on discharge | 72
symptomatic again | 86
rash | 86
serum cryoglobulins positive | 86
complements low | 86
worsening proteinuria | 86
fluid retention | 86
urea level high | 86
creatinine level low | 86
plasmapheresis | 86
cyclophosphamide recommenced | 86
discharged from hospital | 98
serum cryoglobulin negative | 98
fluid overload | 110
pneumonia | 110
cyclophosphamide ceased | 110
thrombocytopenia | 110
sepsis | 110
herpes zoster | 110
haemodialysis | 110
plasmapheresis | 110
paraproteinaemia | 110
monoclonal IgM kappa | 110
Bence Jones protein negative | 110
skeletal survey normal | 110
light chains in serum negative | 110
bone marrow biopsy | 110
low-grade lymphoma | 110
CD20 expression on B cells | 110
rituximab | 110
dramatic improvements in symptoms | 117
absence of cryoglobulins | 117
normal complement levels | 117
discharged home | 117
renal function improved | 210
dialysis independent | 210
cryoglobulin titres negative | 840
serum complements normal | 840
prednisolone 5 mg daily | 840
no side effects | 840
no infections | 840