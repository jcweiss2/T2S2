37 years old | 0
male | 0
admitted to the hospital | 0
severe epigastric pain | -72
progressive lower limbs paresis | -72
alcohol-related acute pancreatitis | -672
heart rate 70 beats/minute | 0
blood pressure 126/76 mmHg | 0
saturation 99% at FiO2=0.21 | 0
body temperature 38°C | 0
bruising around the umbilicus | 0
abdominal wall tender to palpation | 0
absent deep tendon reflexes | 0
weakened middle and lower cutaneous reflexes | 0
attenuation of all kinds of sensation below the umbilicus | 0
complete loss of sensation below the knees | 0
increased amylase level | 0
leukocytosis | 0
giant pancreatic pseudocyst | 0
impaired contrast enhancement of the left kidney | 0
small subcapsular ischemic foci in both kidneys | 0
central hyper-intense signal on T2-weighted images in the thickened medullary cone | 0
medullary infarction | 0
prophylactic dose of low-molecular-weight heparin | 0
empiric antimicrobial therapy | 0
mild anemia | 12
thrombocytopenia | 12
general condition deteriorated | 48
acute renal failure | 48
acute liver failure | 48
complete paraplegia | 48
anemia | 48
thrombocytopenia | 48
decreased fibrinogen | 48
increased D-dimers | 48
international normalized ratio | 48
prolonged activated partial thromboplastin time | 48
hyperdense content in the pancreatic cysts | 48
fresh frozen plasma and packed red blood cells administered | 48
hypotensive | 72
septic shock | 72
emergency laparotomy | 72
omentum and cholecystectomy | 72
external drainage of pancreatic cyst | 72
multifocal coagulative necrosis of mucosa | 72
active inflammatory infiltrate | 72
small vessels with fresh thrombosis | 72
ischemic foci in the liver and spleen | 168
necrotic tissue in the pancreatic head and body | 168
relaparotomy | 168
pancreatic necrosectomy | 168
lesser sac and rectovesical pouch drainage | 168
mixed pancreatobiliary fistula | 168
total parenteral nutrition | 168
somatostatin | 168
hemodiafiltration | 168
hemodialysis | 168
red cell concentrate transfusion | 168
platelets count normalized | 216
hemoglobin level normalized | 288
transferred from the ICU to the surgical ward | 312
follow up MRI | 504
persistent hyperintense signal on T2-weighted images | 504
atrial fibrillation | 624
cardiac arrest | 624
endoscopic retrograde cholangiopancreatography | 624
stents introduced to the common bile duct and Wirsung duct | 960
discharged from the hospital | 1368
lower-limb muscle atrophy | 8760
contractures in the talocrural regions | 8760
no deep tendon reflexes | 8760
no middle and lower cutaneous reflexes | 8760
no sensation below the knees | 8760
moderate flexion and extension in the hips | 8760
urinary retention | 8760
erectile dysfunction | 8760
severe atrophy of the medullary cone | 10800
central gliosis | 10800