54 years old| 0
    woman| 0
    type 2 diabetes mellitus| 0
    brought into emergency department| 0
    acute onset of shortness of breath| -24
    drowsiness| -24
    stopped metformin| -8760
    stopped subcutaneous insulin| -8760
    lifestyle modifications| -8760
    regular exercise| -8760
    modified diet comprising mostly fruits and salads| -8760
    intermittent fasting from 09:00 to 21:00 daily| -8760
    started taking traditional Chinese medications| -8760
    fish oil| -8760
    black garlic| -8760
    lingzhi| -8760
    polydipsia| -4320
    back aches| -4320
    thigh aches| -4320
    intentional weight loss of 27%| -4320
    atrophy of leg muscles| -4320
    slow gait| -4320
    difficulty climbing stairs| -4320
    dehydrated| 0
    drowsy| 0
    Glasgow Coma Scale of 6| 0
    sinus tachycardia| 0
    tachypnoea| 0
    heart rate of 125| 0
    respiratory rate of 28| 0
    blood pressure of 157/113| 0
    afebrile| 0
    saturating well on room air| 0
    cachexic| 0
    malnourished| 0
    equal pupils| 0
    reactive pupils| 0
    no pink skin| 0
    no bright red lips| 0
    no signs of pancreatitis| 0
    blood samples lipaemic| 0
    strawberry pink blood| 0
    high anion gap metabolic acidosis| 0
    lactic acidosis| 0
    ketosis| 0
    serum ketones 16.47 mmol/L| 0
    lactate 3.47 mmol/L| 0
    inadequate respiratory compensation| 0
    hyperkalaemia| 0
    hypokalaemia| 0
    HAGMA| 0
    anion gap 44.0| 0
    delta gap 1.6| 0
    normokalaemia| 0
    serum glucose 31.5 mmol/L| 0
    urea 7.2 mmol/L| 0
    serum osmolality 312 mOsm/kg| 0
    severe hyperlipidaemia| 0
    hypertriglyceridaemia| 0
    total serum cholesterol 47.07 mmol/L| 0
    serum triglycerides 267.66 mmol/L| 0
    high-density lipoprotein 0.28 mmol/L| 0
    low-density lipoprotein 3.85 mmol/L| 0
    no significant biochemical evidence of pancreatitis| 0
    glycated haemoglobin 8.2%| 0
    normal serum troponin| 0
    normal liver function tests| 0
    normal thyroid function tests| 0
    normal creatine kinase| 0
    normal paracetamol levels| 0
    normal salicylate levels| 0
    normal carboxyhaemoglobin| 0
    normal calcium| 0
    normal magnesium| 0
    normal phosphate levels| 0
    urine positive for glucose 4+| 0
    urine positive for ketones 4+| 0
    urine positive for proteins 4+| 0
    ECG sinus tachycardia| 0
    ECG no signs of hyperkalaemia| 0
    ECG no signs of hypokalaemia| 0
    normal chest X-ray| 0
    normal abdominal X-ray| 0
    normal CT brain imaging| 0
    diagnosed with severe DKA| 0
    severe hypertriglyceridaemia| 0
    intubated for airway protection| 0
    fluid resuscitation| 0
    intravenous insulin| 0
    admitted to ICU| 24
    resuscitated with 7 L fluids| 24
    started on intravenous meropenem| 24
    continuous insulin infusion| 24
    lactic acidosis resolved| 48
    ketoacidosis resolved over 3 days| 72
    weaned off intravenous insulin on day 4| 96
    subcutaneous insulin started| 96
    extubated| 96
    transferred out of ICU| 96
    started on statins| 96
    started on fibrates| 96
    HT improved| 96
    hypercholesterolaemia improved| 96
    blood cultures positive for E. coli| 96
    urine cultures negative| 96
    normal CXR| 96
    normal contrasted CT abdomen and pelvis| 96
    referred to endocrinology| 96
    referred to renal medicine| 96
    insulin titration| 96
    chronic outpatient follow-up| 96
    reviewed by hospital dietician| 96
    occupational therapists consulted| 96
    physiotherapists consulted| 96
    rehabilitation| 96
    muscle recovery| 96
    educated on medication compliance| 96
    DKA improved| 408
    hypertriglyceridaemia improved| 408
    discharged on day 18| 432
    total serum cholesterol downtrended to 11.69 mmol/L| 432
    triglycerides downtrended to 0.78 mmol/L| 432
    asymptomatic at follow-up| 672
    compliant to insulin| 672
    compliant to diabetes medications| 672
    normal total serum cholesterol at 1 month| 672
    normal triglycerides at 1 month| 672
    random urine protein <0.04 mg/dL| 672
    UFEME negative for glucose| 672
    UFEME negative for ketones| 672
    no neuropathy| 672
    no retinopathy| 672
    routine outpatient follow-up| 672
