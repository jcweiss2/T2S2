75 years old | 0
male | 0
Caucasian | 0
admitted to the hospital | 0
history of UC | -155520
clinical remission | -116640
recurrent flares | -29120
maintenance therapy with 5-aminosalicylates | -29120
repeated courses of steroids | -29120
commenced on prednisolone | -8760
6-mercaptopurine | -8760
incessant nausea | -8760
abdominal pain | -8760
continued to take prednisolone | -5040
severe life-threatening flare | -168
intravenous steroids | -168
hydrocortisone | -168
rescue therapy with infliximab | -168
discharged home | 336
second dose of infliximab | 504
abdominal pain | 1008
collapse | 1008
hypotensive | 1008
tachycardic | 1008
febrile | 1008
hypoxic | 1008
oxygen saturations of 91% | 1008
tenderness in the right iliac fossa | 1008
haemoglobin of 8.6 g/dL | 1008
normal white cell count | 1008
raised CRP of 193 mg/L | 1008
bilateral lower zone consolidation | 1008
severe chest sepsis | 1008
on-going colitis | 1008
co-amoxiclavulanic acid | 1008
gentamicin | 1008
signs of meningism | 1068
cerebrospinal fluid Gram stain showed Gram-positive rods | 1068
meropenem | 1068
rifampicin | 1068
blood and CSF cultures grew Listeria species | 1128
Listeria monocytogenes | 1128
reduction in Glasgow coma scale | 1208
computed tomography scan of brain | 1208
dilatation of the ventricles | 1208
raised intracranial pressure | 1208
hydrocephalus | 1208
intubated and ventilated | 1208
external ventricular drain insertion | 1208
ICP monitoring | 1208
gradual recovery | 4032
discharged home | 4032