11-year-old | 0
Hispanic male | 0
Maple Syrup Urine Disease (MSUD) | 0
newborn metabolic screen | -105,840
blood amino acids confirmation | -105,840
congenital nystagmus | -105,840
exotropia surgery | -105,840
growth along the 10th percentile | -105,840
two significant episodes of severe metabolic decompensation before age 7 | -105,840
one episode complicated by cerebral edema | -105,840
intensive care unit stay | -105,840
mannitol use | -105,840
baseline learning issues | -105,840
behavioral issues | -105,840
attention deficit hyperactivity disorder (ADHD) | -105,840
good dietary compliance | -105,840
stable blood amino acids | -105,840
normal growth velocity | -105,840
presented in septic shock | 0
metabolic crisis | 0
cerebral edema | 0
intubation | 0
hemodialysis | 0
insulin continuous infusion | 0
pancreatitis | 0
pneumonia | 0
cavitary Group A Streptococcus infection | 0
trophic feeds of BCAA free formula | 0
dextrose supplementation | 0
intravenous lipid supplementation | 0
BCAA free total parental nutrition | 0
natural protein restriction | 0
elevated leucine levels | 0
prolonged restriction leading to negative amino acid balance | 0
pulmonary thrombosis | 168
renal infarction | 168
hypercoagulable state | 168
normal renal function | 168
three doses of dexamethasone | 168
neurologic stabilization | 168
metabolic stabilization | 168
transfer to pediatric progressive care unit | 168
antibiotics course completion | 168
resumption of home feeds | 168
weaning off intravenous fluids | 168
leucine levels remaining high | 168
natural protein restriction to 3.5–4 g/day | 168
weight decrease by 1.1 kg | 168
increased work of breathing | 240
biphasic stridor | 240
tracheal tugging | 240
subglottic stenosis | 240
tracheal stenosis | 240
transfer back to PICU | 240
laryngoscopy preparation | 240
intervention under anesthesia | 240
increased IV fluids to twice maintenance | 240
D10W+0.9%NS infusion | 240
operating room on June 5th | 288
70% sub-subglottic stenosis | 288
tracheostomy | 288
nasogastric tube placement | 288
BCAA free formula administration | 288
high risk for decannulation | 288
sedation requirement | 288
muscle relaxation requirement | 288
natural protein of 4 g/day | 288
valine supplementation | 288
isoleucine supplementation | 288
intralipids resumed | 288
glucose infusion rate maintained | 288
amino acid monitoring | 288
trended up amino acids | 384
continuous insulin infusion started | 384
increased dextrose to 8 mg/kg/min | 384
hemodynamically stable | 384
continuous airway pressure support | 384
no end organ dysfunction | 384
elevated leucine (1050 nmol/mL) | 432
metabolic acidosis (pH 7.23) | 432
anion gap of 15 | 432
altered mental status | 432
decreased ability to follow commands | 432
dialysis consideration | 432
growth hormone course started | 432
natural protein increased to 7 g/day | 432
normalization of anion gap | 456
normalization of metabolic acidosis | 456
improved ability to follow commands | 456
stabilized leucine levels | 456
trach change on June 12th | 456
sedation weaning | 456
paralysis weaning | 456
BCAA free formula held | 456
natural protein decreased to 3.5 g/day | 456
increased activity level | 480
BCAA down trending | 480
leucine remaining close to 1000 nmol/mL | 480
BCAA levels rising again | 576
lethargy | 600
leucine level 1322 nmol/mL | 600
concern for infection | 600
elevated white blood cells | 600
elevated platelets | 600
red and white blood cells in urine | 600
Enterobacter cloacae urine culture | 600
IV antibiotics treatment | 600
elevated ESR | 600
elevated CRP | 600
down trending ESR and CRP | 600
normal renal ultrasound | 600
normal serum creatinine | 600
dialysis discussion | 600
second growth hormone course started | 600
physical therapy initiation | 600
BCAA stabilization | 672
BCAA down trending (leucine 519, isoleucine 70, valine 169) | 672
natural protein increased to 7 g/day | 672
modified barium swallow study passed | 672
transition to home MSUD formula | 672
solids foods introduction | 672
protein count goal | 672
enteral formula supplementation | 672
insulin weaning | 672
dextrose weaning | 672
BCAA normalization by June 24th | 864
tolerating home nutrition | 864
supplement regimen tolerance | 864
regained admission weight | 864
weight gain along 50-60th percentile | 864
prolonged admission for tracheostomy training | 864
physical rehabilitation | 864
increased natural protein tolerance | 864
discharged on 12 g/day natural protein | 864
natural protein prescription decreased to 8 g/day over twelve months | 864
muscle wasting correction | 864
puberty onset | 864
scheduled laryngoscopy for laryngotracheal reconstruction | 864
parental consent for case report publication | 864
