32 years old | 0
    female | 0
    cystic fibrosis | 0
    bronchiectasis | 0
    recurrent hemoptysis | 0
    pancreatic insufficiency | 0
    malnutrition | 0
    admitted for massive hemoptysis | 0
    treated with broad-spectrum antibiotics | 0
    CF exacerbation | 0
    computed tomography angiogram | 0
    centrilobular ground-glass opacities | 0
    left lower lobe | 0
    pulmonary hemorrhage | 0
    referred to interventional radiology | 0
    bronchial artery embolization | 0
    right common femoral artery access | 0
    left bronchial arteriogram | 0
    microcatheter used | 0
    left bronchial artery embolized | 0
    embospheres | 0
    post-embolization arteriogram | 0
    resolution of hemoptysis | 0
    discharged | 0
    re-presented with recurrent massive hemoptysis | 3
    inhaled tranexamic acid | 3
    admitted to MICU | 3
    repeat embolization | 3
    repeat CTA | 3
    enlarging left upper lobe pseudoaneurysm | 3
    systemic to pulmonary arterial fistulae | 3
    electively intubated | 3
    diagnostic bronchoscopy | 3
    pulmonary and systemic arterial angiography | 3
    embolization | 3
    left pulmonary artery angiogram | 3
    supreme intercostal artery angiogram | 3
    embolization of supreme intercostal artery | 3
    left thyrocervical trunk angiogram | 3
    embolization of thyrocervical trunk | 3
    post-embolization angiogram | 3
    transferred back to MICU | 3
    hemoptysis improved | 24
    extubated | 24
    septic shock | 24
    Burkholderia cepacian complex | 24
    weaned off vasopressors | 24
    transferred out of MICU | 24
    hemoptysis-free for 11 days | 24
    isolated hemoptysis recurrence | 264
    transferred back to MICU | 264
    repeat CTA | 264
    enhancement of pseudoaneurysm | 264
    multidisciplinary decision | 264
    recurrent massive hemoptysis | 408
    intubation | 408
    repeat CTA | 408
    pseudoaneurysm altered morphology | 408
    repeat embolization | 408
    pulmonary artery angiogram | 408
    pseudoaneurysm opacification | 408
    microcatheter advanced | 408
    coil embolization | 408
    post-embolization angiogram | 408
    clinical deterioration | 408
    comfort measures | 408
    expired | 408
    acute respiratory failure | 408
    Burkholderia cepacian infection | 408
