51 years old | 0
male | 0
high-grade intermittent fever | -360
cough with expectoration | -360
breathlessness | -24
hypertension | unknown
childhood onset bronchial asthma | unknown
chronic steroid therapy | unknown
nebulized bronchodilators | -360
steroids | -360
quinolones | -360
tachycardia | 0
tachypnea | 0
bilateral crepitations | 0
wheeze | 0
respiratory distress | 0
eschar on left chest | 0
noninvasive ventilatory support | 0
azithromycin | 0
doxycycline | 0
oseltamivir | 0
throat swab for H1N1 | 0
sepsis workup | 0
intubation | 0
meropenem | 0
teicoplanin | 0
CT scan of brain | 0
CT scan of thorax | 0
CT scan of abdomen | 0
bilateral multifocal patchy consolidation | 0
minimal right-sided pleural effusion | 0
collapse of left lung fields | 0
consolidation of left lung | 0
Gram stain showing Nocardia species | 0
acid-fast stain positive | 0
cotrimoxazole | 0
imipenem | 0
tracheal aspirate cultures | 0
Nocardia otitidiscaviarum identification | 0
resistant to cotrimoxazole | 0
resistant to amoxicillin-clavulanate | 0
susceptible to amikacin | 0
susceptible to ciprofloxacin | 0
susceptible to linezolid | 0
susceptible to imipenem | 0
susceptible to ceftriaxone | 0
negative acid-fast stain for Mycobacteria | 0
negative HIV antibodies | 0
negative H1N1 RT-PCR | 0
high WBC count | 0
neutrophilic predominance | 0
progressive thrombocytopenia | 0
positive scrub typhus IgM antibodies | 0
ventilatory support | 0
transient hemodynamic improvement | 0
deterioration with increasing inotropic requirement | 0
blood cultures with yeast-like cells | 120
caspofungin | 120
Candida tropicalis | 168
deranged renal parameters | 168
deranged liver function test | 168
deranged coagulation profile | 168
anuria | 168
worsening metabolic acidosis | 168
renal replacement therapy | 168
bradycardia | 168
asystole | 168
death | 168
sepsis | 168
septic shock | 168
multiorgan dysfunction | 168
community-acquired pneumonia | 168
nocardiosis | 168
scrub typhus | 168
candidemia | 168
