58 years old | 0
male | 0
Caucasian | 0
admitted to the hospital | 0
shock | 0
diffuse ST-elevation at the electrocardiogram | 0
fever | -168
persistent cough | -168
nasopharyngeal swab test performed | -48
SARS-CoV-2 infection | -48
levofloxacin | -120
current smoker | 0
hypothyroidism | 0
chest X-ray | -2160
pneumological consultant | -2160
interstitial lung disease | -2160
high-resolution lung computed tomography (CT) scan | -2160
mass in the right lung suspected for cancer | -2160
endobronchial ultrasound-guided transbronchial needle aspiration | -2160
severe hypotension | -12
asthenia | -12
emergency service called | -12
electrocardiogram revealed a diffuse ST-elevation | 0
blood pressure 80/40 mmHg | 0
heart rate 110 bpm | 0
oxygen saturation 88% on room air | 0
body temperature 37.5°C | 0
emergency coronary angiography | 0
absence of a coronary artery disease | 0
normal left ventricular function | 0
admitted to the COVID-19 ward | 0
high inflammatory markers | 0
increased liver enzymes | 0
normal troponin values | 0
arterial blood gas analysis | 0
respiratory alkalosis with hyperlactatemia | 0
bedside focused ultrasound | 0
lung ultrasound showed an interstitial syndrome | 0
bilateral B lines | 0
small sub-pleural consolidations | 0
bilateral pleural effusion | 0
echocardiography highlighted the presence of diffuse pericardial effusion | 0
swinging heart | 0
inferior caval vein of 2.2 cm with no respiratory excursion | 0
global left ventricular ejection fraction of 50% | 0
blood pressure values increased after fluid therapy | 12
pericardiocentesis was not performed | 12
oxygen saturation rapidly deteriorated | 12
high flow oxygen therapy | 12
diagnosis of pericarditis | 12
corticosteroids and colchicine were started | 12
heparin prophylaxis was started | 12
high dose aspirin was avoided | 12
empiric antibiotic therapy was administrated | 12
second nasopharyngeal swab tested negative for SARS-CoV-2 infection | 48
third nasopharyngeal swab tested negative for SARS-CoV-2 infection | 96
enzyme-linked immunosorbent assay based test resulted positive for IgM and IgG antibodies for SARS-CoV-2 | 96
total body CT was performed | 120
locally advanced lung cancer of 8.5 cm with subclavian artery and vein and thoracic lymph nodes involvement | 120
pleural and pericardial effusion | 120
histological examination confirmed the diagnosis of lung adenocarcinoma | 120
oncologic evaluation | 168
moved to the oncologic clinic | 168
died for rapidly worsening of the respiratory failure | 168