35 years old | 0
    female | 0
    gravida 5 | 0
    para 2022 | 0
    presented to tertiary care hospital | 0
    at 36 weeks and 2 days gestation | 0
    new-onset vaginal bleeding | 0
    five-day history of fevers | -120
    headache | -120
    neck stiffness | -120
    altered mental status | -120
    dog bite | -72
    prenatal history significant for IUGR | 0
    IUGR diagnosed at 32w5d | -2712
    fetus weighing 1477g | -2712
    past medical history significant for motor vehicular accident | 0
    splenectomy | 0
    diffuse axonal brain injury | 0
    loss of short-term memory | 0
    secondary seizure disorder | 0
    cesarean delivery due to unstable pelvis | 0
    tremulous chills | -72
    fevers to 102.7°F | -72
    husband noted off-balance | -72
    slurring words | -72
    endorsed new-onset significant fatigue | -72
    persistent headache | -72
    transient spotting across bilateral visual fields | -72
    new bright red vaginal bleeding | -72
    symptoms prompted hospital visit | -72
    wound on index finger | 0
    well-healing | 0
    no erythema | 0
    no swelling | 0
    no tenderness to palpation | 0
    category 2 fetal heart tracing | 0
    placental abruption | 0
    underwent emergent repeat cesarean section | 0
    neonate admitted to NICU | 0
    respiratory failure necessitating intubation | 0
    core temperature lability | 0
    platelet count 8×109/L | 0
    repeat testing confirmed | 0
    transfused with 2 units of platelets | 0
    platelet count increased to 55×109/L | 0
    post-operative platelet count decreased to 16×109/L | 0
    thrombophilia | 0
    baseline platelet count 400×109/L | 0
    concern for ITP | 0
    concern for TTP | 0
    hematologic emergency requiring plasmapheresis | 0
    infectious etiology considered | 0
    splenic platelet sequestration | 0
    hematology evaluation negative for schistocytes | 0
    normal ADAMST13 level | 0
    excluded TTP | 0
    sepsis considered | 0
    DIC ruled out | 0
    normal fibrinogen | 0
    normal PT | 0
    normal PTT | 0
    sepsis syndromes | 0
    profound thrombocytopenia | 0
    remote history of platelet count 14×109/L | -43824
    ITP considered | 0
    unresponsive to transfusion | 0
    started on clindamycin | 0
    started on gentamicin | 0
    started on metronidazole | 0
    concern for infectious process | 0
    immunocompromised due to asplenia | 0
    susceptible to encapsulated organisms | 0
    dog bite risk of infection | 0
    bacteremia with Capnocytophaga | 0
    mortality risk 25-60% | 0
    rabies considered | 0
    dog fully vaccinated | 0
    dog quarantine | 0
    no evidence of rabies | 0
    rabies prophylaxis deferred | -72
    infectious disease consultation | 0
    x-ray of finger unremarkable | 0
    started on meropenem | 0
    tick bite exposure | -8760
    contact with goat placenta | -8760
    Coxiella burnetii exposure | -8760
    started on doxycycline | 0
    neck stiffness | 0
    fluctuating mental status | 0
    intracranial component considered | 0
    platelet count <70×109/L | 0
    lumbar puncture deferred | 0
    encephalopathy considered | 0
    altered mental status | 0
    MRI of brain with contrast | 0
    no encephalitis | 0
    no acute intracranial processes | 0
    chronic changes from prior brain injury | 0
    blood cultures positive for gram negative bacilli | 0
    Capnocytophaga species preliminarily identified | 0
    converted to IV ertapenem | 0
    10-day course | 0
    Capnocytophaga canimorsus isolated | 0
    bacterial identification via MALDI-TOF | 0
    16S rRNA sequencing | 0
    neonate intubated | 0
    respiratory distress | 0
    discharged to newborn nursery | 144
    neonate blood cultures negative | 0
    platelet count recovered to 278×109/L | 24
    thrombocytopenia attributed to infection | 0
    discharged on sixth hospital day | 144
    completed IV ertapenem outpatient | 144
    asplenia | 0
    thrombocytopenia | 0
    fevers | 0
    altered mental status | 0
    zoonotic exposures | 0
    IUGR | 0
    preterm labor | 0
    preterm delivery | 0
    delay in antibiotic treatment | -72
    fetal distress | 0
    vaginal bleeding | 0
    neonatal respiratory distress | 0
    favorable outcomes | 0