63 years old | 0
male | 0
dentist | 0
employed | 0
experienced systemic reaction | 0
acute and diffuse urticaria | 0
recurrent loss of consciousness | 0
treated with steroids | 0
treated with epinephrine | 0
anaphylactic shock suspected | 0
referred two episodes of transitory loss of consciousness | -8760
attributed to laryngeal hyper-reactivity | -8760
evaluated at the Allergy Unit | 72
determination of Immuno-CAP | 72
chlorhexidine-specific IgE | 72
total IgE | 72
Basophil Activation Test | 72
exposed to chlorhexidine via inhalation | -672
sanitation procedures | -672
daily cleaning and disinfection | -672
aerosol products containing antiseptic/disinfectant | -672
positive CD63 expression | 72
SI=6.0 | 72
tested a mouthwash containing chlorhexidine | 72
CD63=9.6% | 72
SI=4.0 | 72
disinfectant containing chlorhexidine | -672
2.0% solution chlorhexidine digluconate | -672
mixed with other components | -672
anaphylaxis | 0
allergic contact dermatitis | 0
urticaria | 0
photodermatitis | 0
drug-related skin eruptions | 0
facial flushing | 0
swelling | 0
paresthesia | 0
generalized urticaria | 0
itching | 0
difficulty in breathing | 0
reduced blood pressure | 0
adrenaline | 0
anaphylactic reactions | 0
occupational activity impaired | 0
systematic review | 0
CARE checklist | 0
PRISMA guidelines | 0
search strategy | 0
inclusion criteria | 0
exclusion criteria | 0
target journals | 0
hand-searched | 0
characteristics of cases | 0
occupational allergic reactions | 0
health-care workers | 0
allergic history | 0
type of exposure | 0
clinical picture | 0
diagnosis | 0
management/treatment | 0
health outcome | 0
Nagendran et al. | 0
Toholka and Nixon | 0
Waclawaski et al. | 0
Wittczak et al. | 0
Vu et al. | 0
IgE-mediated reactions | 0
immediate-type hypersensitivity | 0
delayed-type hypersensitivity | 0
skin prick tests | 0
specific IgE | 0
basophil activation test | 0
sIgE | 0
BAT | 0
CD63 | 0
SI | 0
anaphylactic reaction | 0
severe anaphylaxis | 0
occupational anaphylaxis | 0
chlorhexidine-induced anaphylaxis | 0
hypersensitivity reaction | 0
allergic sensitization | 0
antiseptics/disinfectants | 0
health-care settings | 0
exposure | 0
risk factors | 0
prevention strategies | 0
health surveillance programs | 0
life-threatening events | 0
medical community | 0
side effects | 0
severe adverse reactions | 0
conflict of interest | 0
acknowledgment | 0
Dr. Bernard Patrick | 0
English manuscript | 0
discharged | 24