5 years old | 0  
    diagnosed with Crohn's disease | -105120  
    older brother with Crohn's disease | -105120  
    bronchiolitis episodes | -105120  
    anti-tumor necrosis factor drug (infliximab) | -2928  
    protein-losing enteropathy | -2928  
    recurrent intestinal pseudo-obstruction | -2928  
    admitted to hospital | 0  
    abdominal pain | 0  
    bloody stool | 0  
    gangrenous bowel | 0  
    ascending colon removed | 0  
    developed pneumonia | 24  
    ARDS | 24  
    PaO2/FiO2 <100 | 24  
    ventilated | 24  
    lung protective ventilation strategy | 24  
    fever | 24  
    hypotension | 24  
    tachycardia | 24  
    tachypnea | 24  
    bilateral crackles | 24  
    arterial blood pH: 7.10 | 24  
    pCO2: 55 | 24  
    pO2: 95 | 24  
    HCO3: 17 | 24  
    BE: −7 | 24  
    O2 saturation: 98% | 24  
    lactate: 6.8 | 24  
    hemoglobin: 9.9 g/dL | 24  
    white blood cell count: 19,300/mm3 | 24  
    platelets: 61,000/mm3 | 24  
    increased neutrophil band count | 24  
    CRP: 10 mg/dL | 24  
    procalsitonin: 100 ng/mL | 24  
    chest radiography diffuse infiltration | 24  
    chest radiography consolidation | 24  
    antibiotics initiated | 24  
    vasopressors initiated | 24  
    Pseudomonas aeruginosa in tracheal culture | 24  
    Pseudomonas aeruginosa in blood culture | 24  
    oliguric renal failure | 24  
    continuous venovenous hemodialysis | 24  
    fever subsided | 264  
    laboratory findings back to normal | 264  
    CRP not back to normal | 264  
    cultures sterile | 264  
    general well-being | 264  
    weaning attempt failed | 336  
    re-intubated | 336  
    restrictive pattern with low compliance | 336  
    HRCT interlobular septal thickening | 336  
    HRCT air bronchograms | 336  
    HRCT consolidated areas | 336  
    HRCT bronchiectasia | 336  
    HRCT ground glass opacities | 336  
    neutrophilic infiltration in tracheal aspirates | 336  
    negative mycobacterium tuberculosis | 336  
    negative viral respiratory organisms | 336  
    normal immunological profile | 336  
    tracheostomy performed | 552  
    prednisolone initiated | 552  
    clinical condition improved | 648  
    pulmonary functions improved | 648  
    CRP returned to normal | 648  
    discharged from PICU | 768  
    no mechanical ventilator support | 768  
    tracheostomy present | 768  
    bronchiolitis episodes in past | -105120  
    no PFT applied | -105120  
    no BHR determined | -105120  
    no subclinical alterations detected | -105120  
    no histopathological examination | 336  
    parental disapproval for bronchoscopy | 336  
    no conflicts of interest | 0  
    

  Final Answer

5 years old | 0  
diagnosed with Crohn's disease | -105120  
older brother with Crohn's disease | -105120  
bronchiolitis episodes | -105120  
anti-tumor necrosis factor drug (infliximab) | -2928  
protein-losing enteropathy | -2928  
recurrent intestinal pseudo-obstruction | -2928  
admitted to hospital | 0  
abdominal pain | 0  
bloody stool | 0  
gangrenous bowel | 0  
ascending colon removed | 0  
developed pneumonia | 24  
ARDS | 24  
PaO2/FiO2 <100 | 24  
ventilated | 24  
lung protective ventilation strategy | 24  
fever | 24  
hypotension | 24  
tachycardia | 24  
tachypnea | 24  
bilateral crackles | 24  
arterial blood pH: 7.10 | 24  
pCO2: 55 | 24  
pO2: 95 | 24  
HCO3: 17 | 24  
BE: −7 | 24  
O2 saturation: 98% | 24  
lactate: 6.8 | 24  
hemoglobin: 9.9 g/dL | 24  
white blood cell count: 19,300/mm3 | 24  
platelets: 61,000/mm3 | 24  
increased neutrophil band count | 24  
CRP: 10 mg/dL | 24  
procalcitoni