65 years old| 0
male | 0
admitted to the hospital | 0
cough | -24
greenish expectoration | -24
chest pain | -24
asthenia | -24
weight loss | -24
valvuloplasty | -25920
aortic valve replacement | -25920
Warfarin 5 mg once a day | -25920
Carvedilol 12.5 mg in the morning | -25920
Carvedilol 6.25 mg in the afternoon | -25920
left anterior hemiblock | 0
acute respiratory failure | 0
admitted to the ICU | 0
poor ventilatory mechanics | 0
inadequate management of secretions | 0
use of accessory muscles | 0
mixed acidosis | 0
orotracheal intubation | 0
invasive mechanical ventilation | 0
systolic blood pressure 104/54 mmHg | 0
partial oxygen saturation 80% | 0
respiratory rate 36 rpm | 0
heart rate 120 beats/min | 0
left pneumothorax | 0
thoracic drainage tube placed | 0
IMV support | 0
sedation with Propofol | 0
analgesia with fentanyl | 0
metabolic acidosis | 0
shock caused by dehydration | 0
severe hemodynamic compromise | 0
tension pneumothorax | 0
central venous catheter | 0
nasogastric tube | 0
bladder catheter | 0
chest tube to drain pneumothorax | 0
pneumonia due to non-specific microorganisms | 0
tree-like infiltrate | 0
consolidations in the upper lobe | 0
consolidations in the lower right | 0
consolidations in the upper left lobe | 0
pleural effusion on the right side | 0
left pneumothorax with chest tube insertion | 0
leukocytes 14200 mm3 | 0
hemoglobin 8.9 g/dl | 0
hematocrit 28.9% | 0
mean corpuscular volume 77 fl/red cell | 0
mean concentration of hemoglobin 23.7 picograms/cell | 0
mean cell hemoglobin concentration 30.6 grams/deciliter | 0
red blood cell count 374 mm3 | 0
platelets 166000 mm3 | 0
monocytes 3.2% | 0
eosinophils 1.4% | 0
lymphocytes 3.9% | 0
neutrophils 91.3% | 0
basophils 0.2% | 0
glucose 114.3 mg/dl | 0
sodium 141 meq/L | 0
potassium 3.2 meq/L | 0
chlorine 111 meq/L | 0
calcium 7.9 meq/L | 0
BUN 15 mg/dl | 0
creatinine 0.9 g/dl | 0
treatment with ampicillin/sulbactam | 0
treatment with clarithromycin | 0
antifimic treatment with rifampicin-isoniazid | 0
antifimic treatment with pyrazinamide | 0
antifimic treatment with ethambutol | 0
bronchoscopy | 24
pale palate mucosa | 24
erythematous stippling | 24
cavitary image in the right upper lobe | 24
bronchioloalveolar lavage | 24
bronchial brushing | 24
cultures for mycobacteria | 24
cultures for fungi | 24
Pseudomonas aeruginosa | 28
Klebsiella pneumoniae | 28
KPC producing strains | 28
Mycobacterium tuberculosis detected | 28
no resistance to rifampicin | 28
Ziehl-Neelsen staining positive | 28
Löwenstein-Jensen culture positive | 672
Colistin 300 mg initial dose | 28
Colistin 100 mg every 8 hours | 28
nebulized amikacin 500 mg every 12 hours | 28
complete resolution of pneumothorax | 240
interstitial pattern | 240
left pulmonary cavern | 240
pleural effusion | 240
bilateral right predominance | 240
hemodynamic instability | 312
increased dose of vasopressor | 312
inotropic support with norepinephrine | 312
inotropic support with dobutamine | 312
atrial fibrillation | 312
rapid reverse ventricular response | 312
death | 312
