31 years old| 0
male | 0
admitted to the ICU | 0
gunshot wound to the abdomen | -672
gunshot wound to the chest | -672
exploratory laparotomy | -672
right thoracotomy | -672
left arm injury | -672
left elbow fracture | -672
open reduction internal fixation | -672
septic shock | -672
acute kidney injury | -672
chest infection | 0
infected laparotomy wound | 0
empiric piperacillin/tazobactam therapy | 0
prolonged ICU stay (56 days) | 0
received several antibiotics | 0
continuous fever | 0
leukocytosis | 0
persistent source of infection (abdominal wound) | 0
persistent source of infection (left-hand ORIF site wound) | 0
frequent dressing | 0
debridement | 0
carbapenem-resistant P. stuartii isolate in sputum | 528
resistant to ciprofloxacin | 528
resistant to trimethoprim/sulfamethoxazole | 528
resistant to gentamicin | 528
resistant to imipenem | 528
resistant to meropenem | 528
sensitive to amikacin | 528
unremarkable chest X-ray | 528
highly febrile | 720
piperacillin/tazobactam every 6 hours | 720
persistent fever | 768
increasing leukocytes | 768
septic screening (tracheal aspirate, urine, wound, blood) | 768
piperacillin/tazobactam changed to meropenem | 768
septic screening results | 840
P. stuartii in urine | 840
P. stuartii in wound | 840
P. stuartii in blood | 840
carbapenem-resistant K. pneumoniae in urine | 840
carbapenem-resistant K. pneumoniae in wound | 840
carbapenem-resistant K. pneumoniae in blood | 840
tracheal aspirate culture report | 888
carbapenem-resistant P. stuartii | 888
carbapenem-resistant K. pneumoniae | 888
resistant to amikacin | 888
resistant to ciprofloxacin | 888
resistant to trimethoprim/sulfamethoxazole | 888
resistant to gentamicin | 888
resistant to imipenem | 888
intermediate to meropenem | 888
meropenem dosing regimen changed to 2g every 8 hours with extended infusion | 888
colistin added | 888
colistin loading dose | 888
colistin maintenance dose | 888
follow-up septic screen | 1056
MDR Acinetobacter baumannii in left-hand ORIF site wound | 1056
MDR Acinetobacter baumannii in tracheal aspirate | 1056
unremarkable chest X-ray | 1056
meropenem discontinued | 1128
colistin discontinued | 1128
transferred to ward | 1344
stable with no signs of infection | 1344
received multiple antibiotics | 0
completed prolonged courses of colistin | 0
completed prolonged courses of tigecycline | 0
completed prolonged courses of imipenem | 0
hospital-acquired pneumonia caused by carbapenem-resistant P. stuartii and K. pneumoniae | 0
