45 years old | 0
female | 0
fall from 18 feet height | -504
difficulty in breathing | -48
past history of pulmonary tuberculosis | -8760
completely treated | -8760
conscious | 0
oriented | 0
respiratory rate 30/min | 0
heart rate 120/min | 0
blood pressure 112/68 mm Hg | 0
reduced air entry on the left side of the chest | 0
tenderness in the epigastrium | 0
bowel sounds were present | 0
X-ray chest posteroanterior view | 0
large air-fluid level in left hemithorax | 0
collapsed underlying lung | 0
obliteration of cardiophrenic angle | 0
rightwards shift of the mediastinum | 0
infiltrates and scarring in upper zones bilaterally | 0
plain computerised tomography scan chest | 0
hydropneumothorax | 0
lung collapse | 0
ultrasonography of abdomen | -168
no evidence of solid organ injury | -168
no free fluid in the abdominal cavity | -168
provisional diagnosis of traumatic hydropneumothorax | 0
intercostal drain tube insertion | 0
50 ml seropurulent fluid drained out | 0
gastric contents appeared in the intercostal drainage system | 2
nasogastric tube insertion | 2
repeat chest X-ray | 2
Ryle's tube in the area of left hydropneumothorax | 2
diagnosis revised as TDH | 2
iatrogenic perforation of stomach | 2
surgical repair planned | 2
tachypnoeic | 2
respiratory rate 36/min | 2
SpO2: 92% on oxygen | 2
heart rate 118/min | 2
blood pressure 130/78 mm Hg | 2
blood gas analysis | 2
PaO2 64 mm Hg | 2
PaCO2 39 mm Hg | 2
pH 7.38 | 2
vital parameters monitoring | 2
electrocardiogram | 2
non-invasive blood pressure | 2
SpO2 monitoring | 2
rapid sequence induction | 2
injection thiopentone 250 mg | 2
succinylcholine 100 mg | 2
tracheal intubation | 2
intermittent positive pressure ventilation | 2
anaesthesia maintenance | 2
thoracic epidural catheter placement | 2
injection bupivacaine 0.25% 8 ml | 2
surgical exploration of the abdomen | 2
large diaphragmatic rent | 2
stomach and spleen herniating into the thoracic cavity | 2
reduction of hernia | 2
diaphragmatic tear repair | 2
fresh ICT insertion | 2
feeding gastrostomy | 2
stable intraoperatively | 2
shifted to intensive care unit | 2
mechanical ventilation | 2
reduced air entry on the left side of the chest | 2
chest X-ray | 2
extensive infiltrates in the left lung | 2
arterial blood gases | 2
hypercarbia | 2
PaCO2 58 mm Hg | 2
culture and sensitivity of pleural fluid | 48
growth of enterobacter species | 48
sensitive to meropenem and amikacin | 48
early weaning from the ventilator | 48
tracheostomy | 336
nutrition maintenance | 48
enteral feeds through gastrostomy | 48
minimal ventilatory support | 48
high grade fever | 48
leucocytosis | 48
tachycardia | 48
systemic inflammatory response syndrome | 48
infection under control | 672
left lung expanded | 672
gases exchange improved | 672
haemodynamic stability | 672
ICT removal | 672
transferred to the surgical department | 720
tracheostomy | 720
gastrostomy | 720