24 years old | 0
male | 0
Nepalese | 0
admitted to the Emergency Department | 0
fever | -72
cough | -72
fatigue | -72
disoriented to place and time | 0
blood in the nasopharynx | 0
no oral injury | 0
no urinary or bowel incontinence | 0
no neck stiffness | 0
vomited coffee ground emesis | 0
maintaining 99% oxygen saturation on room air | 0
blood pressure 126/84 mmHg | 0
temperature 39.4°C | 0
intubated | 0
portable chest X-ray revealed normal lung parenchyma | 0
severe deranged liver function | 0
SARS-CoV-2 positive | 0
started on SARS-CoV-2 treatment | 0
started on liver support | 0
acetylcysteine infusion | 0
lactulose | 0
vitamin K | 0
rifaximin | 0
intravenous pantoprazole | 0
4-factor prothrombin complex concentrate | 0
fresh frozen plasma | 0
fibrinogen | 0
sustained low-efficiency dialysis | 0
computed tomography of the Head | 0
no evidence of intra- or extra-axial intracranial hemorrhage | 0
abdominal ultrasound | 0
liver normal in size | 0
coarse parenchymal echotexture | 0
spleen normal in size | 0
both kidneys normal in size | 0
body temperature fluctuating | 24
ventilatory settings | 24
repeat RT-PCR for SARS-CoV-2 positive | 168
developed disseminated intravascular coagulation | 168
bleeding from the intravenous site and endotracheal tube | 168
died on the 10th day of admission | 240
multiorgan failure | 240
acute liver failure | 240
acute renal failure | 240
disseminated intravascular coagulation | 240
fulminant hepatitis B infection | 0
hepatitis B viral count >17 million | 0
cytokine storm | 0
altered immune response | 0
severe COVID-19 | 0
marked activation of coagulative and fibrinolytic system | 0
lower platelet count | 0
higher ratio of neutrophil count to lymphocyte count | 0
H score 172 | 0
hemophagocytic syndrome | 0
COVID-19-induced cytokine storm | 0
immunosuppression | 0
severe hepatitis B infection | 0
severe spontaneous hypothermia | 0
poor outcome | 0
inverse neutrophil to lymphocyte count ratio | 0