35 years old | 0
    woman | 0
    previously healthy | 0
    abrupt onset of dyspnea | -72
    loss of consciousness for 5 minutes | -72
    received illegal hyaluronic acid injection into the dermis of the forehead | -72
    received illegal hyaluronic acid injection into the dermis of the right cheek area | -72
    body temperature 36.8℃ | 0
    blood pressure 150/110 mm Hg | 0
    pulse rate 127/min | 0
    respiratory rate 28/min | 0
    confused mental state | 0
    crackles in both lower lung fields | 0
    normal liver function test | 0
    normal renal function test | 0
    white blood cells 21,080/µL (neutrophils 91%) | 0
    hemoglobin 11 g/dL | 0
    platelets 240,000/µL | 0
    troponin I 0.16 ng/mL | 0
    CK-MB 0.6 ng/mL | 0
    C-reactive protein 5.307 mg/dL | 0
    D-dimer 1.278 µg/mL | 0
    N-terminal prohormone brain natriuretic peptide 9,177 pg/mL | 0
    arterial blood gas pH 7.505 | 0
    arterial blood gas PCO2 28.6 mm Hg | 0
    arterial blood gas PO2 66.1 mm Hg | 0
    arterial blood gas HCO3- 22.4 mmol/L | 0
    plain chest radiography ground glass opacity | 0
    plain chest radiography consolidation in both lung fields | 0
    contrast-enhanced chest CT diffuse ground glass opacity in both lungs | 0
    contrast-enhanced chest CT dilatation of the pulmonary artery | 0
    contrast-enhanced chest CT right ventricle dilatation | 0
    admitted to intensive care unit | 0
    mechanical ventilation due to worsening hypoxemia | 0
    hemorrhagic eruptions in anterior chest area | 24
    administered antibiotics | 24
    administered corticosteroids | 24
    administered diuretics | 24
    hypoxemia improved | 120
    initial blood culture no growth | 120
    no evidence of fever | 120
    excluded septic embolism | 120
    discontinued antibiotics | 120
    weaned from mechanical ventilation | 168
    discharged | 192
    completely improved after one month | 720
    follow-up chest CT improvement of pulmonary lesion without fibrosis | 720