71 years old | 0
African American | 0
female | 0
type 2 diabetes mellitus | 0
chronic kidney disease stage IV | 0
hypertension | 0
heart failure with preserved ejection fraction | 0
chronic obstructive pulmonary disease | 0
gout | 0
admitted to the burn intensive care unit | 0
maculopapular rash | -168
allopurinol | -168
erosive rash | 0
ocular involvement | 0
oropharyngeal involvement | 0
skin biopsies | 0
SJS/TEN | 0
SCORTEN score 4 | 0
IV corticosteroids | 0
IVIG therapy | 0
respiratory failure | 24
intubation | 24
septic shock | 24
ileus | 24
oliguric renal failure | 24
continuous renal replacement therapy | 24
bloody diarrhea | 504
drop in hemoglobin | 504
infectious workup | 504
Clostridium difficile assay | 504
upper endoscopy | 504
antral gastritis | 504
colonoscopy | 504
perianal skin breakdown | 504
epidermal SJS lesions | 504
ulcers of the cecum and ileocecal valve | 504
ulcerated, edematous mucosa | 504
histologic examination | 504
hematochezia | 504
transfusion-dependent anemia | 504
colonoscopy | 672
radiologic guided embolization | 672
ileocecectomy recommended | 672
high-dose steroid therapy | 672
IV dexamethasone | 672
IV methylprednisolone | 672
prednisone taper | 672
multidisciplinary conference | 672
infliximab therapy | 672
septic shock refractory to vasopressors | 1728
death | 1728