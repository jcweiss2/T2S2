77 years old | 0
    woman | 0
    menopause at 52 years | 0
    adenocarcinoma | 0
    endometrial cytology | 0
    MRI revealed primary malignant tumor in uterine cervix | 0
    MRI showed small amount of fluid accumulation in uterine cavity | 0
    cervical biopsy | 0
    diagnosed with Stage IIB cervical cancer | 0
    CCRT with cisplatin | 0
    whole-pelvis irradiation | 0
    brachytherapy | 0
    MRI before brachytherapy showed primary tumor shrunk | 0
    MRI before brachytherapy showed fluid retention in uterine cavity increasing | 0
    no signs of infection | 0
    WBC 1400/µL | 0
    neutrophils 868/µL | 0
    lymphocytes 448/µL | 0
    CRP 0.41 mg/dL | 0
    fifth cycle of cisplatin administered | 24
    presented with fever 38.8°C | 72
    presented with malaise | 72
    COVID-19 negative | 72
    discharged from outpatient clinic | 72
    came to emergency department | 96
    decreased consciousness | 96
    worsening general condition | 96
    fever 37.9°C | 96
    GCS score 13 points | 96
    WBC 2300/µL | 96
    neutrophils 2254/µL | 96
    lymphocytes 56/µL | 96
    CRP 1.39 mg/dL | 96
    CT revealed extensive pyometra | 96
    CT revealed small inflammation of small intestine | 96
    consciousness worsened to GCS score 7 points | 96
    left conjugate eye deviation | 96
    suspected right paralysis | 96
    no nuchal rigidity | 96
    head CT showed subacute cerebral infarction | 96
    head MRI showed subacute cerebral infarction | 96
    pyometra considered predominant site of infection | 96
    transcervical drainage performed | 96
    intrauterine purulent material reddish-yellow | 96
    suspected sepsis | 96
    intravenous meropenem administered | 96
    general condition worsened | 96
    respiratory condition unstable | 96
    frequent seizures | 96
    tracheal intubation performed | 96
    anti-epileptic levetiracetam administered | 96
    L. monocytogenes detected in pyometra material | 168
    L. monocytogenes detected in blood culture | 168
    administration of ampicillin and gentamicin initiated | 168
    lumbar puncture performed | 168
    CSF pressure 18 cmH2O | 168
    CSF gross findings showed sunshine dust | 168
    CSF polynuclear cell count increased | 168
    CSF total protein increased | 168
    FilmArray detected L. monocytogenes | 168
    FilmArray detected cytomegalovirus | 168
    diagnosed with L. monocytogenes meningitis | 168
    diagnosed with cytomegalovirus | 168
    intravenous ampicillin continued | 168
    intravenous gentamicin continued | 168
    ganciclovir initiated | 168
    vital signs improved | 576
    blood test results improved | 576
    moved to general bed | 576
    able to open eyes spontaneously | 2880
    state of consciousness stable | 2880
    GCS score 8 points | 2880
    grade 2 leukopenia | 0
    grade 3 neutropenia | 0
    grade 4 lymphopenia | 0
    no complaint of abdominal pain | 96
    no intra-abdominal free space on CT | 96
    leukopenia | 0
    neutropenia | 0
    lymphopenia | 0
    no abdominal pain | 96
    no uterine perforation | 96
    meropenem initiated | 96
    vancomycin initiated | 96
    frequent seizures continued | 96
    tracheal intubation | 96
    levetiracetam administered | 96
    seizures frequent | 96
    CSF pressure 18 cmH2O | 168
    CSF sunshine dust | 168
    CSF polynuclear 1157 cells/µL | 168
    CSF total protein 455 mg/dL | 168
    FilmArray detected L. monocytogenes | 168
    FilmArray detected cytomegalovirus | 168
    intravenous ampicillin | 168
    intravenous gentamicin | 168
    ganciclovir | 168
    moved from ICU to general bed | 576
    four months after admission | 2880
    opened eyes spontaneously | 2880
    consciousness stable | 2880
    GCS 8 points | 2880
    E4 | 2880
    VT | 2880
    M4 | 2880
    no nuchal rigidity | 96
    no abdominal pain | 96
    no intra-abdominal free space | 96
    no uterine perforation | 96
    grade 2 leukopenia | 0
    grade 3 neutropenia | 0
    grade 4 lymphopenia | 0
    CCRT with brachytherapy | 0
    fifth cycle cisplatin | 24
    fifth administration cisplatin | 24
    three days after brachytherapy | 72
    two days after fifth cisplatin | 72
    three days after brachytherapy | 72
    following day after outpatient clinic | 96
    day after brachytherapy | 24
    third day after hospitalization | 168
    fourth month after admission | 2880
    24th day of hospitalization | 576
    first admission | 0
    four months after first admission | 2880
    administration of CCRT | 0
    during CCRT | 0
    after CCRT | 0
    during brachytherapy | 0
    before brachytherapy | 0
    after brachytherapy | 0
    during hospitalization | 0
    after hospitalization | 0
    after diagnosis | 0
    after drainage | 0
    after treatment | 0
    after meningitis diagnosis | 0
    after ampicillin initiation | 0
    after gentamicin initiation | 0
    after ganciclovir initiation | 0
    after ICU | 0
    after general bed | 0
    after four months | 2880
    after first admission | 0
    after lumbar puncture | 0
    after CSF analysis | 0
    after FilmArray | 0
    after tracheal intubation | 0
    after seizures | 0
    after meropenem | 0
    after vancomycin | 0
    after levetiracetam | 0
    after consciousness deterioration | 96
    after emergency department | 96
    after CT scan | 96
    after MRI scan | 96
    after transcervical drainage | 96
    after purulent material drainage | 96
    after L. monocytogenes detection | 168
    after blood culture | 168
    after ampicillin and gentamicin | 168
    after lumbar puncture | 168
    after CSF findings | 168
    after meningitis diagnosis | 168
    after cytomegalovirus diagnosis | 168
    after moving to general bed | 576
    after four months | 2880
    after eye opening | 2880
    after consciousness stabilization | 2880
    after GCS improvement | 2880
    no COVID-19 | 72
    no uterine perforation | 96
    no abdominal pain | 96
    no intra-abdominal free space | 96
    no nuchal rigidity | 96
    no relationship to cerebral infarction | 96
    no obvious GPR in endometrial fluid | 168
    GPR in blood culture | 168
    L. monocytogenes detected in both specimens | 168
    increased fluid accumulation in uterine cavity | 0
    uterine cavity fluid accumulation | 0
    cervical tumor shrunk | 0
    applicators inserted into uterine cavity | 0
    uterine cavity manipulation | 0
    immunocompromised state | 0
    high risk of infection | 0
    sepsis | 96
    meningitis | 168
    uterine perforation risk | 96
    peritonitis risk | 96
    septic shock risk | 96
    neurological sequelae risk | 0
    mortality risk | 0
    hematogenous spread | 0
    ascending route unlikely | 0
    immunosuppression | 0
    malignancy | 0
    age risk | 0
    leukopenia risk | 0
    neutropenia risk | 0
    lymphopenia risk | 0
    CCRT risk | 0
    brachytherapy risk | 0
    uterine cavity infection | 0
    intrauterine infection | 0
    L. monocytogenes infection | 168
    cytomegalovirus infection | 168
    Gram-positive rods | 168
    Gram-stained images | 168
    fluid accumulation increased | 0
    tumor shrunk | 0
    fluid retention increased | 0
    purulent fluid | 96
    reddish-yellow purulent material | 96
    sunshine dust in CSF | 168
    increased polynuclear cells | 168
    increased total protein | 168
    E3 | 96
    V4 | 96
    M6 | 96
    E2 | 96
    V1 | 96
    M4 | 96
    E4 | 2880
    VT | 2880
    M4 | 2880
    frequent seizures | 96
    respiratory instability | 96
    consciousness deterioration | 96
    general condition worsening | 96
    fever 38.8°C | 72
    fever 37.9°C | 96
    malaise | 72
    decreased consciousness | 96
    paralysis suspected | 96
    eye deviation | 96
    seizures frequent | 96
    vital signs improvement | 576
    blood improvement | 576
    eye opening | 2880
    consciousness stability | 2880
    GCS improvement | 2880
    antibiotic switch | 168
    empiric antibiotics | 96
    definitive antibiotics | 168
    appropriate antibiotics | 168
    risk factors identified | 0
    predisposing factors | 0
    immune compromise | 0
    treatment-induced leukopenia | 0
    high mortality risk | 0
    neurological sequelae | 0
    improved vital signs | 576
    improved blood tests | 576
    moved to general bed | 576
    spontaneous eye opening | 2880
    stable consciousness | 2880
    GCS 8 points | 2880
    written consent obtained | 0
    consent available | 0
    no competing interests | 0
    acknowledgments | 0

