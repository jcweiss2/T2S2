65 years old | 0 | 0 
male | 0 | 0 
admitted to the hospital | 0 | 0 
multiple blisters | -432 | 0 
erosions | -432 | 0 
superadded maggot infection | -432 | 0 
previous episodes of lesions | -720 | -168 
treatment with steroids | -720 | -168 
unknown generic medications | -720 | -168 
lesions all over the body | -168 | 0 
febrile | 0 | 0 
flaccid blisters | 0 | 0 
erosions | 0 | 0 
Nikolsky sign positive | 0 | 0 
diagnosis of PV | 0 | 0 
skin biopsy | 0 | 0 
tzanck smear | 0 | 0 
intravenous dexamethasone pulse | 0 | 72 
supportive care | 0 | 72 
intravenous antibiotics | 0 | 72 
isolation intensive care unit | 0 | 0 
oozing from skin ulcerations | 0 | 168 
hemorrhagic excoriation | 0 | 168 
peeling of skin | 0 | 168 
oral methyl prednisolone | 72 | 168 
hypoproteinemia | 168 | 168 
pleural effusion | 168 | 168 
blood culture showed enterobacter | 168 | 168 
pus culture showed Staphylococcus aureus | 168 | 168 
pus culture showed Proteus mirabilis | 168 | 168 
intravenous Tigecycline | 168 | 240 
intravenous vancomycin | 168 | 240 
sepsis | 168 | 240 
high grade fever | 168 | 240 
albumin levels fell | 168 | 240 
TPE | 240 | 360 
TPE cycle | 240 | 360 
Nikolsky sign negative | 288 | 288 
no new lesions | 288 | 288 
exudation from lesions reduced | 288 | 360 
dressings dry | 288 | 360 
lesions showed re-epithelization | 288 | 360 
lesions showed healing | 288 | 360 
oral lesions healed | 360 | 360 
erosions on back | 360 | 360 
erosions on thigh | 360 | 360 
erosions on buttocks | 360 | 360 
IV methyl prednisolone pulse | 360 | 432 
cyclophosphamide | 360 | 432 
discharged | 432 | 432 
monthly IV dexamethasone pulse | 432 | 0 
daily oral prednisolone | 432 | 0