70 years old | 0
female | 0
admitted to the hospital | 0
hypertension | -8760
heart failure with recovered ejection fraction | -8760
non-ischaemic cardiomyopathy | -8760
paroxysmal atrial fibrillation | -8760
remote cardiac arrest | -8760
ventricular fibrillation | -8760
cardiac resynchronization therapy defibrillator | -4380
ICD | -2190
fever | 0
altered mental status | 0
jugular venous distention | 0
soft systolic murmur | 0
white blood cell count of 10 880/μL | 0
haemoglobin 7900 g/dL | 0
glomerular filtration rate of 78 mL/min/1.73 m2 | 0
lumbar puncture | 0
cerebrospinal fluid cultures grew S.pneumoniae | 0
chest radiograph | 0
right-sided consolidation | 0
pleural effusion | 0
pleural fluid cultures grew S.pneumoniae | 0
blood cultures grew S.pneumoniae | 0
transthoracic echocardiogram | 0
TV mass | 0
moderate tricuspid regurgitation | 0
estimated left ventricular EF of 45% | 0
transoesophageal echocardiogram | 24
mobile mass with independent motion on TV | 24
mobile echodensity on the ICD pacing wire | 24
endocarditis | 0
CIED-related infection | 0
Austrian syndrome | 0
IV vancomycin | 0
ceftriaxone | 0
prophylactic anticoagulation | 0
ICD extraction | 120
intracardiac echocardiography | 120
lead extraction | 120
AngioVac-assisted extraction of the TV mass | 192
near-complete removal of TV mass | 192
discharged | 264
wearable cardioverter defibrillator | 264
IV ceftriaxone | 264
ICD replacement | 720
ventricular fibrillation | -720
defibrillation | -720
alcoholism | -8760
immunodeficiency | -8760
intrinsic lung disease | -8760
Osler’s triad | 0
pneumonia | 0
meningitis | 0
septic emboli | 0
pericardial effusion | 120
embolic complication | 120
valve replacement | -8760
valve repair | -8760
valvectomy | -8760
percutaneous thrombectomy | 192
AngioVac device | 192
TV debulking | 192
PTVD | 192
surgical intervention | -8760
medical management | 0
antibiotic therapy | 0
cerebrospinal penetration | 0
mortality | -8760
surgical candidacy | 0
rehabilitation | 264
cardioverter defibrillator | -2190
cardiac arrest | -8760
cardiomyopathy | -8760
atrial fibrillation | -8760
cardiac resynchronization therapy | -4380
CRT-D | -4380
single-chamber ICD | -2190
battery exchange | -2190
EF recovered | -2190
non-pacing QRS | -2190
narrow QRS | -2190
arrhythmic events | -2190
device upgrade | -720
device interrogation | -720
septal leaflet | 24
tricuspid valve | 0
right atrium | 192
venous drainage | 192
venous return | 192
bypass pump | 192
filter | 192
extracorporeal system | 192
thrombotic material | 192
venous circulation | 192
TV surgery | -8760
PTVD cohort | -8760
sicker overall | -8760
co-morbidities | -8760
surgical intervention | -8760
mortality rate | -8760
length of stay | 264
blood transfusion | 264
operative approach | 192
valvular disease | -8760
interventional services | -8760
infectious disease | 0
collaboration | 0
case report | 0
images | 0
text | 0
consent | 0
COPE guidance | 0
European Heart Journal | 0
Case Reports Consent Form | 0
financial support | 0
research | 0
authorship | 0
publication | 0
manuscript | 0
resident physician | -8760
Internal Medicine | -8760
Rush University Medical Center | -8760
fellow physician | -8760
Pulmonology | -8760
Critical Care | -8760
Cleveland Clinic | -8760
health equity | -8760
discrimination | -8760
health care | -8760
hiker | -8760
outdoors | -8760
Supplementary material | 0
European Heart Journal—Case Reports | 0