61 years old | 0
woman | 0
admitted to the hospital | 0
general weakness | 0
fall at home | 0
infected heel pressure ulcer | 0
admitted to the Department of General Surgery | 0
urinary tract infection | 0
thyroid dysfunction | 0
hemodynamic instability | 6
loss of consciousness | 6
admitted to the intensive care unit | 6
intubated | 6
unconscious | 6
hypothermic | 6
temperature 35.8°C | 6
hypotensive | 6
systolic blood pressure 75 mm Hg | 6
bradycardic | 6
heart rate 45 beats per min | 6
obese | 6
body mass index of 36 | 6
generalized subcutaneous edema | 6
marked in the lower limbs | 6
large areas of macerated skin | 6
extensive heel pressure ulcer | 6
surgical revision | 6
soft abdomen | 6
inaudible peristalsis | 6
irreducible ventral hernia | 6
no features of occlusion | 6
hypercapnia | 6
compensated respiratory acidosis | 6
arterial blood pH of 7.36 | 6
elevated serum bicarbonate | 6
HCO3 32 mEq/L | 6
hypomagnesemia | 6
0.5 mmol/L | 6
hypophosphatemia | 6
0.4 mmol/L | 6
severe hypoalbuminemia | 6
20 g/L | 6
CRP level of 34 mg/L | 6
WBC count of 5.7 × 109 cells/L | 6
thyroxine T4 1.0 nmol/L | 6
TSH >100 mU/L | 6
extreme thyroid insufficiency | 6
myxedema | 6
fluid resuscitation | 6
inotropic support | 6
hormonal substitution | 6
intravenous T4 500 μg | 6
T4 100 μg/day | 6
intravenous triiodothyronine T3 5 μg × 3/day | 6
suspected sepsis | 6
urinary tract infection | 6
heel pressure ulcer | 6
initial empirical intravenous piperacillin/tazobactam therapy | 6
4 g × 3/day | 6
replaced with cefuroxime | 144
1.5 g × 3/day | 144
metronidazole | 144
500 mg × 3/day | 144
metronidazole withdrawn | 168
urine culture | 168
lower limb wound | 168
Escherichia coli | 168
Corynobacterium | 168
hemodynamic stabilization | 168
intravenous hormonal medication reduced | 168
oral T4 | 168
serum thyroid hormones normalized | 168
extubated | 168
gradual increase in CRP level | 168
CRP 156 ng/L | 168
emergence of clinical signs of pneumonia | 168
radiological signs of pneumonia | 168
cefuroxime replaced with piperacillin/tazobactam | 168
CRP increased to 206 ng/L | 192
no fever | 192
no increase in WBC count | 192
abdomen still silent | 192
moderately distended | 192
no signs of bowel movement | 192
enteral nutrition | 192
computed tomography | 192
considerable amount of fecal content in the colon and rectum | 192
significant expansion up to 9 cm in diameter | 192
enhancement and edema of sigmoid and rectal wall | 192
bowel obstruction | 192
enemas | 192
violent and abundant diarrhea | 192
CDI | 192
diagnosis of CDI confirmed | 480
PCR test | 480
BD MAX Cdiff assay | 480
GeneXpert | 480
enteral vancomycin | 480
250 mg × 4/day | 480
persistent diarrhea | 480
replaced with metronidazole | 528
500 mg × 3/day | 528
enteral fidaxomicin | 528
200 mg × 2/day | 528
intravenous tigecycline | 528
100 mg initially | 528
50 mg × 2/day | 528
piperacillin/tazobactam stopped | 528
no clinical improvement | 528
lack of response to treatment | 528
colonoscopy findings | 528
extensive swelling of the mucous membrane | 528
no pseudomembranous formations | 528
fecal microbiota transplant | 528
frozen stool from healthy donor | 528
donor screened for pathogens | 528
fecal microbiota transplantation procedure | 528
500 mL liquid suspension | 528
5 enema portions | 528
diarrhea disappeared | 528
no adverse effects | 528
rapid decrease in CRP levels | 528
recovery from myxedema | 528
no problems from digestive tract | 528
discharged to ordinary ward | 1560
65 days in ICU | 1560
