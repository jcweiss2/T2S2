history of nonalcoholic steatohepatitis | -10000
history of alpha 1 antitrypsin deficiency | -10000
orthotopic liver transplant | 0
incarcerated inguinal hernia | 1
inguinal hernia repair | 1
cytomegalovirus viremia | 2
treatment with valganciclovir | 2
discharge | 4
encephalopathy | 30
increasing home oxygen requirements | 32
arrival at hospital | 35
require 4L nasal cannula | 35
oxygen saturation >92% | 35
encephalopathy characterized by sparse speech and disorientation | 35
nonfocal neurologic examination | 35
white blood cell count 9.3 × 10^9/L | 35
creatinine 2.12 mg/dL | 35
blood urea nitrogen 53 mg/dL | 35
arterial ammonia 204 µmol/L | 35
induction dosing of intravenous ganciclovir | 35
empiric antibiotic coverage with vancomycin, meropenem, micafungin | 35
intravenous micronutrient supplementation for B1, B6, and levocarnitine | 35
lumbar puncture | 36
opening pressure 8 cmH2O | 36
Gram stain revealed encapsulated yeast suspicious for Cryptococcus | 36
start of liposomal amphotericin B and flucytosine | 36
start of continuous renal replacement therapy (CRRT) | 36
start of rifaximin, zinc, and lactulose | 36
ammonia level 692 µmol/L | 48
neurological deterioration | 48
mechanical ventilation | 48
empiric intravenous doxycycline | 48
ammonia level <100 µmol/L | 84
cryptococcal serum and cerebrospinal fluid (CSF) antigen titers >1:2560 | 84
cultures from bronchoalveolar lavage, CSF, and blood revealed cryptococcal growth | 84
repeat lumbar punctures | 96
opening pressures greater than 45 cmH2O | 96
large volume drainage every 48 hours | 96
thrombocytopenia | 96
nadir of 16 × 10^3/µL | 96
mental status transiently improved | 120
tracheostomy | 120
culture clearance | 168
complications of cryptococcal infection | 168
persistent hydrocephalus | 168
oliguric renal failure | 168
progressive splenic infarcts with necrosis | 168
splenectomy | 168
sepsis | 168
duodenal leak | 168
persisting renal failure | 168
failure to thrive | 168
move to comfort care in hospice | 240
urea cycle disorder screening studies | 240
low urine orotic level | 240
normal serum citrulline and arginine level | 240