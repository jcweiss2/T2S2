28 years old | 0
man | 0
iron deficiency anemia | 0
unknown cause | 0
referred to the local hospital | 0
elective esophagogastroduodenoscopy | 0
intermittent diarrhea | -48
rectal bleeding | -48
computed tomography scan | -48
cirrhotic appearance of the liver | -48
splenomegaly | -48
gastric varices | -48
lesions consistent with gastric varices | 0
glue injection | 0
Histoacryl | 0
lipiodol | 0
exsanguinating hemorrhage | 0
admission to the intensive care unit | 0
resuscitation | 0
hemodynamic stability | 0
loose stools | -17520
occasional blood | -17520
heavy drinking | -17520
no regular alcohol drinking | 0
no family history of liver diseases | 0
iatrogenic upper gastrointestinal hemorrhage | 0
variceal bleeding | 0
portal hypertension | 0
cirrhosis | 0
uncertain etiology | 0
repeated esophagogastroduodenoscopy | 24
general anesthesia | 24
Sengstaken-Blakemore tube insertion | 24
CT angiogram | 24
no active bleeding | 24
provisional diagnosis of portal hypertension | 24
provisional diagnosis of cirrhosis | 24
transjugular intrahepatic portosystemic shunt | 48
removal of Sengstaken-Blakemore tube | 72
postoperative melena | 96
further admission to the intensive care unit | 96
third esophagogastroduodenoscopy | 96
oozing gastric varices | 96
multiple bandings | 96
further glue injections | 96
further attacks of melena | 144
Doppler ultrasonography | 144
repeat CT angiography | 144
inconclusive TIPS patency | 144
high United Kingdom Model for End-Stage Liver Disease score | 144
transfer to regional liver transplantation unit | 144
TIPS venogram | 168
migration of glue | 168
afferent system | 168
efferent system | 168
inferior vena cava | 168
right atrium | 168
pulmonary embolization risk | 168
repeat CT scan | 168
good TIPS patency | 168
glue cast distribution | 168
mobile glue cast in right atrium | 168
embolized pieces in pulmonary arteries | 168
transthoracic echocardiography | 168
mobile echogenic structures within right atrium | 168
normal biventricular size | 168
normal biventricular function | 168
consulted cardiology team | 192
unsuccessful snaring | 192
risk of breaking glue into pieces | 192
interventional radiology opinion | 192
cardiopulmonary bypass risk | 192
liver failure | 192
open heart removal not supported | 192
anticoagulation with low-molecular-weight heparin | 192
magnetic resonance cholangiopancreatography | 216
sigmoidoscopy | 216
final diagnosis of cirrhosis | 216
primary sclerosing cholangitis | 216
overlapping ulcerative colitis | 216
migration of glue | 216
liver transplantation candidate | 216
multidisciplinary discussion | 240
IR approach | 240
standby rescue cardiothoracic team | 240
fluoroscopy | 240
mobile glue cast no longer visible | 240
echocardiogram confirmed glue cast | 240
lipiodol dissolved | 240
radiolucent Histoacryl in right atrium | 240
IR option not feasible | 240
multidisciplinary meeting | 264
direct atrial extraction | 264
liver transplantation surgery | 264
cardiopulmonary bypass support | 264
Histoacryl polymerization | 264
complications | 264
portal vein thrombosis | 264
splenic vein thrombosis | 264
sepsis | 264
embolization | 264
anticoagulation management | 264
waiting list for liver transplantation | 264
planned glue cast removal | 264
cardiothoracic unit extraction | 264
migration of cyanoacrylate glue | 264
severe complication | 264
conservative management | 264
minimally invasive | 264
invasive management | 264
multidisciplinary approach | 264
