46 years old | 0
male | 0
Caucasian | 0
admitted to the hospital | 0
sudden pain | -24
redness | -24
hardening | -24
subfebrile fever | -24
pneumonia | -2160
relapse of pneumonia | -2160
osteomyelitis | -168
recurrent episodes of pain | -168
swelling | -168
lateral side of left thigh | -168
right thigh pain | -504
pathological fractures | -504
Anaerococcus prevotii | -504
abscessotomy | 0
active wash | 0
antibiotics | 0
debridement surgery | 0
external osteosynthesis | 504
femoral trepanation | 504
external AO fixation | 504
pathologic fracture of the left femoral diaphysis | 504
osteomyelitis of the left femur | 504
osteomyelitis of the right femur | 504
sequester | 504
fistulogram | 504
contrast flow | 504
femoral region | 504
X-Ray | 504
CT scans | 504
MRI scans | 504
abscess | 504
intramedullary space | 504
fistulas | 504
air inserts | 504
interfascial spaces | 504
bone destruction | 504
purulent discharge | 504
Ilizarov’s apparatus | 1008
intramedullary osteosynthesis | 1008
silver-plated intramedullary nail | 1008
left knee remodeling | 1008
passive knee motion machine | 1008
femoral resection | 1008
shortening of the left limb | 1008
screw migration | 1512
abscessotomy | 1512
biopsy | 1512
pathological examination | 1512
debridement | 1512
external fixation | 1512
amputation of the left femur | 1812
sepsis | 1812
intensive care unit | 1812
stump debridement | 1812
Meropenem | 1812
Colistin | 1812
right femur healed | 2592
signs of osteomyelitis disappeared | 2592
left thigh healed | 2592
rehabilitation treatment | 2592
outpatient treatment | 2592
follow-up | 2592
osteomyelitis | 0
haematogenous osteomyelitis | 0
pathological fractures | 0
Anaerococcus prevotii | 0
anaerobic bacterium | 0
pneumonia | -2160
lung infection | -2160
purulent processes | -2160
molars | -2160
infection | 0
immunosuppression | 0
diabetes | 0
peripheral vascular disease | 0
drug abuse | 0
surgical implants | 0
immunodeficiencies | 0
bacteria | 0
bloodstream | 0
bone grafts | 0
tissue flaps | 0
antibiotic-impregnated material | 0
hardware | 0
antibiotic therapy | 0
one-stage approach | 0
debridement | 0
re-implantation | 0
hardware | 0
infection | 0
osteomyelitis | 0
femur | 0
pathological fracture | 0
displacement | 0
osteosynthesis | 0
bone healing | 0
knee contracture | 0
amputation | 1812
broad-spectrum antibiotic therapy | 1812
informed consent | 0
conflict-of-interest statement | 0
CARE Checklist | 0
manuscript source | 0
corresponding author | 0
peer-review | 0
scientific quality classification | 0
P-Reviewer | 0
S-Editor | 0
L-Editor | 0
P-Editor | 0