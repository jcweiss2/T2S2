62 years old | 0
    male | 0
    referred to critical care medicine department | 0
    severe acute pancreatitis | -192
    respiratory distress | -48
    chronic cough since childhood | -40320
    heart rate 122/min | 0
    blood pressure 114/66 mm Hg | 0
    respiratory rate 32/min | 0
    predominantly thoracic respiration | 0
    distended abdomen | 0
    tense abdomen | 0
    absent bowel sounds | 0
    Hb 10.2 gm/dl | 0
    total leukocyte count 17,900 cell/cmm | 0
    serum creatinine 1.9 mg/dl | 0
    serum amylase 2897 U/l | 0
    CECT abdomen findings | 0
    endotracheal intubation | 0
    mechanical ventilation | 0
    invasive hemodynamic monitoring | 0
    intra-abdominal pressure 24 mm Hg | 0
    nasogastric tube free drainage | 0
    decrease in intra-abdominal pressure to 17 mm Hg | 72
    nasogastric feeding started | 72
    severe cough | 72
    feed visible in endotracheal tube | 72
    aspiration suspected | 72
    endotracheal tube upsized to 9.0 mm | 72
    cuff applied | 72
    thorough tracheal toileting | 72
    recurrent distention of nasogastric drainage bag with air | 72
    gastric content in respiratory tract | 72
    communication between respiratory tract and esophagus suspected | 72
    bedside bronchoscopy | 72
    gastric contents regurgitating into right main bronchus | 72
    right broncho-esophageal fistula diagnosed | 72
    septic shock | 72
    severe acute respiratory distress syndrome | 72
    high ventilator support required | 72
    vasopressor support required | 72
    chest X-ray bilateral lung infiltrates | 72
    right lung predominant involvement | 72
    death | 120
    