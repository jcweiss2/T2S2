77 years old | 0 | 0 | Factual
female | 0 | 0 | Factual
breast cancer | -10080 | -10080 | Factual
chemotherapy | -10080 | -10080 | Factual
radiation to the chest | -10080 | -10080 | Factual
severe aortic stenosis | 0 | 0 | Factual
coronary artery disease | 0 | 0 | Factual
90% occlusion of the left anterior descending artery | 0 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
tissue aortic valve replacement | 0 | 0 | Factual
saphenous vein graft bypass | 0 | 0 | Factual
midline sternotomy | 0 | 0 | Factual
induction of anesthesia | 0 | 0 | Factual
intubation | 0 | 0 | Factual
left internal mammary artery dissected | 0 | 0 | Factual
left internal mammary artery atretic | 0 | 0 | Factual
greater saphenous vein small | 0 | 0 | Factual
cardiopulmonary bypass | 0 | 0 | Factual
decline in cerebral head saturations | 0 | 0 | Factual
reduced mean arterial perfusion | 0 | 0 | Factual
reduced cerebral artery perfusion | 0 | 0 | Factual
use of vasopressors | 0 | 0 | Factual
extubated | 2 | 2 | Factual
postoperative course complicated | 0 | 0 | Factual
persistent lactic acidosis | 0 | 0 | Factual
high-dose vasopressor support | 0 | 0 | Factual
mixed cardiogenic and vasoplegic shock | 0 | 0 | Factual
lethargic | 15 | 15 | Factual
leftward gaze | 15 | 15 | Factual
right upper extremity weakness | 15 | 15 | Factual
symptoms resolved | 15 | 15 | Factual
bilateral tongue ecchymoses | 15 | 15 | Factual
tongue numbness | 15 | 15 | Factual
dysgeusia | 15 | 15 | Factual
CT scan of head | 15 | 15 | Factual
no acute hemorrhage | 15 | 15 | Factual
CT angiogram of brain and neck | 15 | 15 | Factual
no large vessel occlusion | 15 | 15 | Factual
mild calcification at bifurcation of right common carotid artery | 15 | 15 | Factual
50% focal stenosis of distal left common carotid artery | 15 | 15 | Factual
right lingual artery completely occluded | 15 | 15 | Factual
mild distal collateral flow | 15 | 15 | Factual
left lingual artery multifocal irregularities | 15 | 15 | Factual
postoperative platelet count normal | 15 | 15 | Factual
prothrombin time normal | 15 | 15 | Factual
international normalized ratio normal | 15 | 15 | Factual
fibrinogen normal | 15 | 15 | Factual
no prior history of vasculitic disease | 0 | 0 | Factual
ADAMTS13 inhibitor screen normal | 15 | 15 | Factual
volume resuscitation | 15 | 15 | Factual
low-dose epinephrine | 15 | 15 | Factual
high-dose norepinephrine | 15 | 15 | Factual
high-dose vasopressin | 15 | 15 | Factual
systemic vascular resistance improved | 48 | 48 | Factual
otolaryngology service consulted | 15 | 15 | Factual
serial examinations of tongue | 15 | 48 | Factual
flexible bronchoscopes | 15 | 48 | Factual
persistent tongue numbness | 15 | 1440 | Factual
persistent dysgeusia | 15 | 1440 | Factual
supportive therapy | 15 | 1440 | Factual
tongue sensation returned to baseline | 1440 | 1440 | Factual
taste returned to baseline | 1440 | 1440 | Factual
discharged | 1440 | 1440 | Factual