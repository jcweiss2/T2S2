63 years old | 0 | 0 
female | 0 | 0 
168 cm height | 0 | 0 
53 kg weight | 0 | 0 
papillary thyroid carcinoma | -9936 | -9936 
resection | -9936 | -9936 
radiotherapy | -9936 | -9936 
stenosis of the esophagus | -6720 | -6720 
repeated aspiration | -6720 | -6720 
respiratory insufficiency | -6720 | -6720 
pneumonia | -6720 | -6720 
purulent pleurisy | -6720 | -6720 
pleurectomy | -6720 | -6720 
restrictive ventilation pattern | -6720 | -6720 
recurrent nerve palsy | -6720 | -6720 
percutaneous endoscopic gastrostomy | -6720 | -6720 
tracheostoma | -6720 | -6720 
home ventilation | -6720 | 0 
mobility decreased | -8760 | 0 
secondary depression | -8760 | 0 
never left the bed or nursing chair | -8760 | 0 
stopped talking | -8760 | 0 
mandible nearly fixed | -8760 | 0 
could not open her mouth over 20 degrees | -8760 | 0 
left axis vertebralis stented | -4380 | -4380 
stenosis of the internal axis carotis | -4380 | -4380 
arterial hypertension | -4380 | -4380 
secondary lactase deficiency | -4380 | -4380 
esophageal stenosis dilated | -168 | -168 
decreasing general condition | -24 | -24 
fistula between the esophagus and tracheal membrane | -24 | -24 
referred to the University of Erlangen | -24 | -24 
examined by several chiefs and consultants | -24 | -24 
deemed too unstable for open surgery | -24 | -24 
inability to open the mouth | -24 | -24 
recurrent nerve palsy | -24 | -24 
minimal invasive orthograde approach impossible | -24 | -24 
referred to our hospital | 0 | 0 
suffering from pneumonia | 0 | 0 
4-multiresistente gramnegative Pseudomonas aeruginosa | 0 | 0 
put on veno-venous extracorporeal membrane oxygenation | 0 | 0 
partial thromboplastin time of 60 seconds | 0 | 0 
preseptic status | 0 | 0 
ventilated through a tracheostoma | 0 | 0 
low ventilation forces | 0 | 0 
thoracic computed tomography | 24 | 24 
big fistula of the tracheal membrane | 24 | 24 
tracheal cannula ended shortly beneath the lower limit of the mediastinal fistula | 24 | 24 
decision to try endobronchial stenting | 48 | 48 
plan to close the fistula with a pedicled omentum majus replacement | 48 | 48 
surgical plastic needed an abutment and a secured continuous airway replacement | 48 | 48 
procedure performed | 72 | 72 
vv-ECMO began to be partly ineffective | 72 | 72 
rising septical issues | 72 | 72 
high volume input of physiological saline | 72 | 72 
oral approach would only allow a small flexible bronchoscope | 72 | 72 
approach for this upper part of the trachea had to be performed through the percutaneous tracheostoma | 72 | 72 
retrograde manner | 72 | 72 
trying different Dumon and one-hybrid self expandable metalic y-stent | 72 | 72 
plan was to changeover to a more floppy Freitag stent | 72 | 72 
whole procedure was accompanied by a mandatory additional ventilation | 72 | 72 
nasal jet catheter or a special double-lumen endotracheal tube exchange catheter | 72 | 72 
ventilation line was introduced either orally or through the tracheostoma | 72 | 72 
placed distally below the main carina | 72 | 72 
successful retrograde stenting was performed in four steps | 72 | 96 
Step I | 72 | 80 
manually compressed “y” of the FS was successfully pushed downward on the main carina | 72 | 80 
Step II | 80 | 88 
frontal surface of the stent was cut with at least 1 cm opening in the longitudinal axis | 80 | 88 
stent surface was reduced ~40% in the sagittal axis | 80 | 88 
new stoma for a regular tracheal cannula was created | 80 | 88 
lower new edge of this stoma was fixed subcutaneously | 80 | 88 
Step III | 88 | 92 
jagwire was introduced through the mouth into the trachea | 88 | 92 
jagwire was running out of the new FS stoma | 88 | 92 
leaving the dorsal membrane of the cut FS behind | 88 | 92 
soft-tip stiff DLET was introduced for more stability | 88 | 92 
dragged out of the new stoma of the cut FS | 88 | 92 
distal jagwire was introduced into the oral orifice of the FS | 88 | 92 
bending up a curve | 88 | 92 
oral part of the FS was still outside the body | 88 | 92 
bending the FS outward at the level of percutaneous stoma | 88 | 92 
pulling the jagwire at both ends | 88 | 92 
FS flipped with its upper part over the soft-tip stiff DLET into the upper third of the trachea | 88 | 92 
whole fistula was bridged by the FS up to the level of the vocal cords | 88 | 92 
upper edge of the new FS stoma was fixed subcutaneously | 88 | 92 
Step IV | 92 | 96 
regular tracheal cannula was introduced for ventilation | 92 | 96 
lungs were not aerated at that point of time | 96 | 96 
spontaneous breathing work increased | 96 | 240 
vv-ECMO support was reduced | 96 | 240 
lungs became re-aerated again | 96 | 240 
patient woke up again | 96 | 240 
could communicate with her family by writing and her eyes | 96 | 240 
infections continued to be very severe | 240 | 240 
spontaneous work of breathing never exceeded a tidal ventilation of 170 mL per breath | 240 | 240 
reduction of intravenous saline injection was limited | 240 | 240 
mandatory but reduced vv-ECMO support | 240 | 240 
patient along with her family decided actively to reduce the vv-ECMO support | 240 | 240 
died on 18 November 2016 | 240 | 240 
pulmonary infection | 240 | 240