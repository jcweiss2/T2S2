62 years old|0
    male|0
    hypertension|0
    hyperlipidaemia|0
    dizziness|-168
    fatigue|-168
    nausea|-168
    vomiting|-168
    transported to the emergency department|-168
    evaluated|-168
    discharged home|-168
    syncope|0
    ECG obtained en route|0
    anterior ST-segment elevations|0
    ventricular fibrillation|0
    cardiac defibrillation|0
    endotracheal intubation|0
    ventricular fibrillation recurred|0
    resuscitative efforts|0
    restored sinus rhythm|0
    spontaneous circulation|0
    heart rate 77 bpm|0
    regular rhythm|0
    hypotension|0
    no appreciable murmurs|0
    no lower extremity edema|0
    extremities cool to touch|0
    mechanical ventilation|0
    rate 28|0
    tidal volume 500 mL|0
    FiO2 100%|0
    positive end-expiratory pressure 8 cmH2O|0
    breath sounds present bilaterally|0
    ECG wide complex rhythm|0
    slow ventricular tachycardia|0
    right bundle branch block morphology|0
    left axis deviation|0
    high suspicion for acute coronary syndrome|0
    received aspirin|0
    received ticagrelor|0
    received heparin|0
    epinephrine infusion started|0
    bradycardia|0
    hypotension|0
    emergently taken to catheterization lab|0
    coronary angiography|0
    no coronary stenosis|0
    right heart catheterization|0
    elevated right atrial pressure|0
    pulmonary artery pressure 61/28 (39) mmHg|0
    pulmonary capillary wedge pressure 15 mmHg|0
    Fick cardiac index 2.6 L/min/m2|0
    point-of-care echocardiogram performed|0
    dilated right ventricle|0
    severely reduced function|0
    concern for pulmonary embolism|0
    immediate pulmonary angiography performed|0
    large bilateral pulmonary emboli|0
    EkoSonic thrombolysis catheters advanced|0
    tissue plasminogen activator delivered|0
    fibrinogen monitoring|0
    Doppler ultrasounds obtained|0
    no evidence of venous thrombosis|0
    formal transthoracic echocardiogram|0
    depressed right ventricular function|0
    CT chest|0
    bilateral peripheral ground-glass opacities|0
    wedge-shaped opacities in right lung|0
    pulmonary infarctions|0
    refractory hypotension|0
    vasopressors started|0
    broad-spectrum antibiotics|0
    viral respiratory panel negative|0
    tracheal aspirate culture positive|0
    methicillin-resistant Staphylococcus aureus|0
    completion of catheter-directed thrombolysis|0
    repeat ECG|0
    sinus rhythm|24
    first-degree AV block|24
    left axis deviation|24
    incomplete right bundle branch block|24
    prolonged QTc interval 498 ms|24
    developed anaemia|96
    CT chest|96
    CT abdomen|96
    CT pelvis|96
    mediastinal haematoma|96
    persistent ground-glass opacities|96
    tested for SARS-CoV-2|96
    COVID-19 positive|96
    transferred to COVID@-@19 ICU|96
    enhanced contact precautions|96
    supportive care|96
    extubated|192
    inpatient rehabilitation facility|192
    discharged home|672
    lifelong apixaban 5 mg twice daily|672
    mild exertional dyspnoea|672
    transthoracic echocardiogram|672
    improvement of right ventricular dilation|672
    improvement of systolic function|672
    lactic acid 19 mmol/L|0
    troponin I initial 77 ng/L|0
    troponin I peak 6424 ng/L|0
    brain natriuretic peptide 127 pg/mL|0
    prothrombin time 18.2 s|0
    international normalized ratio 1.51|0
    partial thromboplastin time 28 s|0
    fibrinogen 193 mg/dL|0
    D@-@dimer >20000 ng/mL|0
    COVID-19|0
    coagulopathy|0
    increased thrombo-embolic events|0
    right ventricular strain|0
    pulmonary embolism|0
    syncope|0
    out-of-hospital cardiac arrest|0
    ST-elevations in anterior leads|0
    slow wide complex tachycardia|0
    concern for acute coronary syndrome|0
    depressed right ventricular function|0
    bilateral pulmonary emboli|0
    catheter-directed thrombolysis administered|0
    ground-glass opacities|0
    positive COVID-19 test|96
    extubated|192
    discharged home|672
    lifelong anticoagulation|672
    no shortness of breath|0
    denies chest pain|0
    no venous thrombosis|0
    mediastinal haematoma|96
    persistent ground-glass opacities|96
    improved right ventricular function|672
    improved systolic function|672
    negative viral respiratory panel|0
    positive tracheal aspirate culture|0
    methicillin-resistant Staphylococcus aureus|0
    COVID@-@19 ICU admission|96
    enhanced contact precautions|96
    supportive care|96
    inpatient rehabilitation|192
    discharged home|672
    mild exertional dyspnoea|672
    improving dyspnoea|672
    <|eot_id|>