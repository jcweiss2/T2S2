40 years old | 0
    male | 0
    admitted to the emergency department | 0
    persistent frontal headache | -168
    throbbing headache | -168
    over-the-counter painkillers (paracetamol and NSAID) | -168
    chronic lower back pain | -168
    lumbar disc herniation | -168
    NSAID use (intermittent) | -168
    headache recurrence | -168
    fever sensation | 24
    diarrhoea | 24
    temperature of 38.1°C | 24
    pulsatile, fronto-parietal headache | 24
    lumbar puncture | 24
    neutrophilic meningitis | 24
    elevated protein levels | 24
    hypoglycorrhachia | 24
    CSF bacterial culture negative | 24
    multiplex PCR assay negative | 24
    contrast-enhanced computed brain tomography negative | 24
    empirical treatment (dexamethasone and ceftriaxone) | 24
    treatment discontinuation | 24
    morphine administration | 24
    pain relief | 24
    discharge with diagnosis of aseptic meningitis | 24
    paracetamol, ibuprofen, tramadol prescribed | 24
    headache recurrence | 48
    fever | 48
    gradual deterioration of general condition | 48
    neck pain | 48
    photophobia | 48
    phonophobia | 48
    loss of appetite | 48
    fatigue | 48
    temperature of 38.6°C | 48
    slight psychomotor deceleration | 48
    neck stiffness | 48
    hospitalisation | 48
    second lumbar puncture | 96
    lymphocytic predominance (78%) | 96
    high protein levels | 96
    slightly lower blood glucose | 96
    empirical treatment (acyclovir, amoxicillin, ceftriaxone) | 96
    CSF culture negative | 96
    multiplex PCR assay negative | 96
    eubacterial PCR negative | 96
    panfungal PCR negative | 96
    tuberculosis enzyme-linked immunospot assay positive | 96
    CSF direct examination negative | 96
    CSF PCR for Mycobacterium tuberculosis complex negative | 96
    CSF mycobacterial culture sterile | 96
    HIV test negative | 96
    syphilis screening negative | 96
    tick-borne encephalitis serology weakly positive IgG | 96
    Borrelia burgdorferi serology positive IgM | 96
    immunoblot test negative | 96
    CSF PCR for B. burgdorferi negative | 96
    lymphocytic choriomeningitis serology negative | 96
    West Nile serology negative | 96
    Toscana virus serology negative | 96
    mumps IgG serology positive | 96
    fever | 96
    headache persistence | 96
    discontinued anti-infective therapies | 96
    temporal relationship between ibuprofen use and symptom worsening | 96
    ibuprofen suspension | 96
    morphine administration | 96
    symptoms of meningeal syndrome for 8 days | 96
    fever waning after 2 days | 168
    complete resolution of symptoms after 6 days | 216
    investigations for auto-immune diseases suspended | 216
    no headache recurrence | 216
    no neurological sequela | 216
    diagnosis of ibuprofen-induced meningitis | 216

