15 years old | 0\
female | 0\
acute myelogenous leukemia | 0\
induction treatment | -336\
ciprofloxacin | -336\
linezolid | -336\
meropenem | -336\
tobramycin | -336\
liposomal amphotericin | -336\
pancytopenia | -336\
tachycardia | -72\
hypotension | -72\
lactic acidosis | -72\
admitted to the pediatric intensive care unit | 0\
severely impaired left ventricular ejection fraction | 0\
sinus tachycardia | 0\
incomplete right bundle branch block | 0\
NT-proBNP | 0\
high-sensitive troponin T | 0\
fluid therapy | 0\
noradrenaline | 0\
dobutamine | 0\
milrinone | 0\
deep sedation | 0\
mechanical ventilation | 0\
respiratory insufficiency | 0\
va-ECMO | 0\
cannulation of the left femoral artery and vein | 0\
distal leg perfusion | 0\
va-ECMO blood flow | 0\
pre-oxygenator membrane pressure | 0\
mean arterial pressure | 0\
noradrenaline | 0\
vasopressin | 0\
levosimendan | 0\
hydrocortisone | 0\
residual LVEF | 0\
CVVHDF | 0\
anti-infective therapy | 0\
meropenem | 0\
ciprofloxacin | 0\
metronidazole | 0\
cotrimoxazole | 0\
liposomal amphotericin B | 0\
acyclovir | 0\
linezolid | 0\
vancomycin | 0\
PCT | 0\
CRP | 0\
leukocytes | 0\
high-sensitive troponin T | 0\
creatine kinase MB | 0\
total creatine kinase | 0\
microbial specimens | 0\
viral myocarditis | 0\
myocardial biopsy | 0\
mean arterial blood pressure | 24\
LVEF | 24\
noradrenaline | 24\
vasopressin | 24\
levosimendan | 24\
acute ischemic injury | 24\
Dacron conduit | 24\
second arterial cannula | 24\
ECMO circuit | 24\
ECBF | 24\
MAP | 24\
venous drainage pressures | 24\
lactate levels | 24\
PCT | 48\
Hickman catheter | 48\
broad-complex tachycardia | 48\
esmolol | 48\
metoprolol | 48\
left ventricular function | 48\
aortic valve | 48\
pulmonary edema | 48\
intracardiac clot formation | 48\
second venous cannula | 48\
left atrium | 48\
catheter-based atrioseptostomy | 48\
ECMO circuit | 48\
ECBF | 48\
venous drainage | 48\
lactate levels | 48\
MAP | 48\
cerebral oximetry | 48\
regional oxygen saturation | 48\
left ventricle | 48\
therapeutic anticoagulation | 48\
unfractionated heparin | 48\
partial thrombin time | 48\
PCT | 72\
CRP | 72\
leukocytes | 72\
high-sensitive troponin T | 72\
creatine kinase MB | 72\
total creatine kinase | 72\
microbial specimens | 72\
cardiac systolic function | 120\
ECMO cannulas | 120\
LVEF | 168\
mean arterial pressures | 168\
CVVHDF | 168\
renal function | 168\
leucocyte count | 312\
respirator weaning | 792\
allogenic stem cell transplantation | 1008\
LVEF | 1512\
ventricular dilatation | 1512\
discharged | 2160