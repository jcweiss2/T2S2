57 years old | 0
female | 0
alpha-1 antitrypsin deficiency | 0
chronic obstructive pulmonary disease | 0
polysubstance use disorder | 0
severe malnutrition | 0
hemicolectomy/colostomy | -8760
admitted to the hospital | 0
acute abdominal pain | -72
vomiting | -72
constipation | -72
generalized weakness | -72
slurred speech | -72
black stools | -672
tobacco use | 0
assistance with some activities of daily living | 0
clonidine | 0
paroxetine | 0
buprenorphine/naloxone | 0
albuterol/ipratropium inhaler | 0
temperature of 36.6 °C | 0
heart rate of 122 beats per minute | 0
respiratory rate of 22 breaths per minute | 0
blood pressure of 155/109 mmHg | 0
oxygen saturation of 100% on 3 L/minute O2 | 0
severely cachectic | 0
body mass index (BMI) 14 kg/m2 | 0
abdomen was exquisitely tender to light palpation | 0
ostomy output was black appearing | 0
peripheral white blood cell count of 27.1 × 10^9 cells/L | 0
lactate of 3.7 mmol/L | 0
urine toxicology was positive for cocaine | 0
urine toxicology was positive for buprenorphine | 0
fecal occult blood test was negative | 0
computed tomography (CT) scan of the abdomen and pelvis with contrast | 0
diffuse small bowel dilatation suspicious for a small bowel obstruction (SBO) | 0
managed non-operatively | 0
initial improvement over the first three days | 72
WBC had decreased to 13.6 × 10^9 cells/L | 72
increasing clinical deterioration | 96
WBC count had increased to 22.4 × 10^9 cells/L | 120
repeat CT abdomen and pelvis with contrast | 120
pelvic abscess measuring 8.2 × 14.0 × 16.3 cm | 120
persistent SBO | 120
percutaneous transgluteal pigtail catheter was placed within the pelvic abscess | 120
280 mL of purulent, malodorous fluid was immediately removed | 120
abscess cultures grew mixed flora | 120
abscess cultures grew Enterococcus faecium | 120
abscess cultures grew Candida dubliniensis | 120
given ampicillin/sulbactam 3 g IV q6h | 120
given micafungin 100 mg IV q24h | 120
repeat CT abdomen/pelvis | 192
drainage catheter within the abscess | 192
bowel rupture as the underlying cause of the abscess | 192
transgluteal drain was upsized to improve drainage | 192
became confused | 192
hypothermic | 192
tachycardic | 192
tachypneic | 192
transferred to the intensive care unit (ICU) | 192
concern for sepsis | 192
blood cultures drawn | 192
blood cultures were positive for Dietzia cinnamea | 192
same antimicrobials were continued | 192
improved | 240
repeat blood cultures were negative | 240
taken to the operating room (OR) | 336
jejunal enterotomy | 336
jejunojejunal anastomosis | 336
ileocolic anastomosis | 336
abdominal washout | 336
removal of the transgluteal drain | 336
cultures obtained in the OR of soft tissue and the abscess revealed mixed organisms | 336
post-operative course was complicated by confusion | 336
post-operative course was complicated by deconditioning | 336
post-operative course was complicated by ongoing malnutrition | 336
completed antimicrobials | 1008
subsequent imaging showed resolution of the abscess | 1008
discharged | 1008