74 years old | 0
male | 0
obstructive sleep apnea | -672
interstitial lung disease | -672
morbid obesity | -672
hypertension | -672
atrial fibrillation | -672
diabetes mellitus | -672
admitted to the hospital | 0
epigastric abdominal pain | 0
abdominal distension | 0
poor appetite | 0
nausea | 0
belching | 0
constipation | 0
cardiac workup | 0
CT of the abdomen and pelvis | 0
moderate colonic stool | 0
enlarged pelvic lymph nodes | 0
enlarged mediastinal lymph nodes | 0
enlarged retroperitoneal lymph nodes | 0
bronchoscopy | -672
fine-needle aspiration | -672
flow cytometry analysis | -672
discharged | 24
presented to the Emergency Department | 24
no improvement in pain | 24
worsening abdominal distension | 24
using baseline oxygen via nasal cannula | 24
vital signs within normal limits | 24
abdomen soft | 24
mildly distended | 24
non-tender to palpation | 24
no rebound tenderness | 24
no guarding | 24
admission laboratory values | 24
CT of the chest | 24
abdomen and pelvis adenopathy | 24
aortoiliac atherosclerotic disease | 24
right upper-quadrant ultrasound | 24
heterogeneous and coarsened echotexture of the hepatic parenchyma | 24
no biliary tree or gallbladder disease | 24
concern for acute mesenteric ischemia | 24
CT angiography of the abdomen | 24
extensive atherosclerosis of the superior mesenteric artery | 24
moderate stenosis at the ostium | 24
endoscopy | 24
non-obstructing Schatzki ring | 24
gastric ulcer with oozing hemorrhage | 24
bipolar cautery | 24
serum immunofixation | 24
M spike | 24
polyclonal gammopathy | 24
IgM kappa | 24
quantitative IgM mildly elevated | 24
free light chain ratio normal | 24
flow cytometry of peripheral blood | 24
no increased blast proliferation | 24
no lymphoproliferative disease | 24
declined bone marrow biopsy | 24
worsening abdominal pain | 192
altered mental status | 192
asterixis | 192
afebrile | 192
vitals within normal range | 192
oxygen saturation at 94% | 192
white blood cell count elevated | 192
platelets decreased | 192
ALT elevated | 192
AST elevated | 192
lactic acid elevated | 192
total bilirubin elevated | 192
direct bilirubin elevated | 192
INR elevated | 192
ammonia level elevated | 192
repeat CT of the abdomen and pelvis | 192
no acute findings | 192
transferred to the progressive care unit | 192
IV N-acetylcysteine drip | 192
lactulose | 192
IV vitamin K | 192
CT head | 192
no acute abnormalities | 192
EEG abnormal | 192
diffuse slowing | 192
serology negative | 192
tick panel negative | 192
anti-smooth muscle antibodies negative | 192
continued to worsen clinically | 216
respiratory status decompensated | 216
bilateral ground-glass opacities | 216
concerning for pneumonia | 216
broad-spectrum antibiotics | 216
more lethargic | 240
tachypneic | 240
ABG | 240
pH 7.46 | 240
pCO2 34 mmHg | 240
HCO3 24 mEq/L | 240
bilevel-positive airway pressure | 240
admitted to the intensive care unit | 264
unresponsive | 264
comatose | 264
hypotensive | 264
worsening markers of septic shock | 264
increasing lactic acidosis | 264
increasing total bilirubin | 264
direct bilirubin elevated | 264
ALT elevated | 264
AST elevated | 264
reduced hemoglobin | 264
critical thrombocytopenia | 264
prolonged INR | 264
intubated | 264
gram-negative bacteremia | 264
evidence of septic shock | 264
IV fluids | 264
vasopressors | 264
ventricular tachycardia | 288
defibrillated | 288
returned to atrial fibrillation | 288
rapid ventricular response | 288
acute respiratory distress syndrome | 288
deteriorated | 288
initiated comfort care | 288
palliative extubation | 288
died | 336
autopsy findings | 336
diffuse large B-cell lymphoma | 336
involving multiple organs | 336
liver | 336
lung | 336
bone marrow | 336
multiple lymph nodes | 336
lymphadenopathy | 336
right cervical | 336
peri-bronchial | 336
subcarinal | 336
pelvic lymph nodes | 336
large mass | 336
matted lymph nodes | 336
right lung hilum | 336
enlarged liver | 336
multiple ill-defined pale-yellow nodules | 336
infiltration of medium-to-large atypical lymphoid cells | 336
vesicular chromatin | 336
prominent nucleoli | 336
scant-to-moderate amount of cytoplasm | 336
immunohistochemical staining | 336
CD20 positive | 336
CD10 positive | 336
BCL-2 positive | 336
cyclin D1 negative | 336
CD5 negative | 336
CD138 negative | 336
MUM1 negative | 336
CD21 negative | 336
CD3 negative | 336
BCL6 negative | 336
sections of the liver | 336
areas of necrosis | 336
nodular and diffuse infiltrate | 336
atypical medium-to-large CD20+ cells | 336
bone marrow sections | 336
greater than 90% involvement | 336
diffuse large B-cell lymphoma | 336