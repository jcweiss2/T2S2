67 years old | 0
female | 0
admitted to the hospital | 0
backache | -672
calculi in both kidneys | -672
ureteral calculi | -672
HLL | -0.5
double J catheterization | -0.5
purulent urine | -0.5
fever | 0
chill | 0
low blood pressure | 0
imipenem and Cilastatin sodium | 0
fluid resuscitation | 0
Norepinephrine | 0
Hydrocortisone sodium succinate | 0
anuria | 48
ARDS | 48
invasive ventilatory support | 48
CRRT | 48
transfer to ICU | 48
sedated state | 48
cold, clammy extremities | 48
loud bubbling sound in the lung | 48
lactic acid 10.6 mmol/L | 48
bicarbonate 10.8 mmol/L | 48
central venous pressure 20 cmH20 | 48
diffuse dysfunction | 48
LVEF 20.3% | 48
sinus tachycardia | 48
broad ST depression | 48
elevated troponin I | 48
elevated amino-terminal brain natriuretic peptide precursor | 48
creatinine 356 μmol/L | 48
VA-ECMO | 48
CRRT | 48
imipenem and Cilastatin sodium | 48
Vancomycin | 48
lactic acid level declined | 50
vasoactive drugs stopped | 58
arterial blood lactate level normal | 60
extended-spectrum β-lactamase-positive Escherichia coli | 48
inflammatory indices diminished | 72
anti-infection regimen continued | 72
minimum serum trough concentration of Vancomycin | 72
LVEF 35% | 120
black and necrotic skin | 120
weaned from ECMO | 144
renal function scaled as acute kidney injury grade 3 | 144
CRRT discontinued | 144
urinating | 144
vascular ultrasonography | 168
computed tomography angiography | 168
vascular surgery consultation | 168
necrotic tissues amputated | 168
spontaneous breathing | 120
trachea opened | 240
anti-infective therapy replaced | 240
Cefoperazone sodium and Sulbactam sodium | 240
physical rehabilitation | 240
weaned from ventilator | 480
tracheotomy tube sealed | 600
discharged | 768
intermittent hemodialysis | 768
follow-up | 1296