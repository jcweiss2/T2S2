90 years old | 0
female | 0
low back pain | -672
nonsteroidal anti-inflammatory medications | -672
hypertension | -672
hematemesis | -120
Mallory Weiss tear | -120
Forrest 1a ulcer | -120
esophagogastroduodenoscopy | -120
hemoclips | -120
intravenous proton pump inhibitor | -120
hemodynamic instability | -72
drop in hemoglobin | -72
second OGD | -72
slow active bleeding | -72
additional hemoclips | -72
adrenaline injection | -72
melena | -288
repeat OGD | -288
friable tissue | -288
active bleeding | -288
computed tomography mesenteric angiogram | -288
no evidence of bleeding | -288
no signs of pancreatitis | -288
empirical GDA embolization | 0
super selective angiograms | 0
GDA embolization | 0
Nester microcoils | 0
severe epigastric pain | 0
hematemesis | 0
urgent OGD | 0
fresh blood | 0
large blood clot | 0
increased serum amylase | 0
increased serum lipase | 0
exploratory laparotomy | 0
pyloromyoduodenotomy | 0
gastrojejunal bypass | 0
edematous pancreas | 0
generalized bruising | 0
fat saponification | 0
hemorrhagic pancreatitis | 0
pseudomonas septicemia | 72
atrial fibrillation | 72
CT scan | 168
acute focal pancreatitis | 168
loculated peripancreatic collection | 168
multiorgan failure | 216
death | 216