45 years old | 0
male | 0
admitted to the hospital | 0
fever | -168
cough | -48
generalized weakness | -48
loose motions | -48
altered sensorium | -48
herpetiform rash | -168
petechiae | -48
ecchymotic patch | -48
disoriented | 0
irritable | 0
not obeying verbal commands | 0
moving all limbs | 0
no lymphadenopathy | 0
no eschar | 0
chronic alcoholism | 0
heavy smoking | 0
thrombocytopenia | 0
raised urea | 0
raised creatinine | 0
raised liver enzymes | 0
increased serum bilirubin | 0
increased lactate | 0
increased ammonia | 0
normal coagulation parameters | 0
oropharyngeal bleeding | 0
platelets transfused | 0
arterial blood gas analysis | 0
severe metabolic acidosis | 0
fluid resuscitation | 0
improved urine output | 0
broad spectrum antibiotics | 0
intubated | 0
mechanical ventilator support | 0
neurologic deterioration | 0
hemodynamic deterioration | 0
respiratory deterioration | 0
magnetic resonance imaging brain | 0
normal magnetic resonance imaging brain | 0
retiform purpuric rash | 0
purpura fulminans | 0
high grade fever | 0
hypotension | 0
blood negative for malaria parasite | 0
dengue serology negative | 0
Leptospira serology negative | 0
presumptive diagnosis of meningococcemia | 0
Gram stains of the skin biopsy | 0
negative Gram stains | 0
serum/urine Neisseria meningitidis Ag detection | 0
negative serum/urine Neisseria meningitidis Ag detection | 0
lumbar puncture not performed | 0
low platelet count | 0
venereal disease research laboratory | 0
negative venereal disease research laboratory | 0
CARBOGEN | 0
negative CARBOGEN | 0
rapid plasma reagin card test | 0
negative rapid plasma reagin card test | 0
acute hepatitis profile | 0
negative acute hepatitis profile | 0
hepatitis C virus antibodies | 0
negative hepatitis C virus antibodies | 0
vasculitis workup | 0
negative vasculitis workup | 0
blood cultures drawn | 0
sterile blood cultures | 0
urine culture | 0
sterile urine culture | 0
Weil-Felix test | 0
positive Weil-Felix test | 0
doxycycline | 0
bullous eruptions | 24
skin biopsy | 24
mildly hyperkeratotic and flattened epidermis | 24
widespread separation of the epidermis and dermis | 24
direct immunofluorescence study | 24
negative direct immunofluorescence study | 24
extubated | 48
shifted out of ICU | 48
improved neurologically | 48
improved hemodynamically | 48
serum creatinine improved | 48
liver enzymes still elevated | 48
serum bilirubin decreased | 48
retiform rash started to fade | 48
discharged | 336
total 14 days of doxycycline treatment | 336