28 years old | 0
    male | 0
    insulin-dependent diabetes mellitus | 0
    presented to ED | 0
    urinary incontinence | -8760
    dysuria | -8760
    worsening shortness of breath | -8760
    cachexia | 0
    suprapubic tenderness | 0
    diffuse lung crackles | 0
    decreased breath sounds on the right | 0
    blood pressure 150/91 | 0
    pulse 84 | 0
    temperature 97.5 | 0
    respiratory rate 16 | 0
    urinalysis white blood cells | 0
    leukocyte esterase | 0
    blood in urine | 0
    glucose 10,000 mg/dL | 0
    admitted to ICU | 0
    chest CT multiple bilateral densities and nodules | 0
    consolidated cavitated mass in right lung | 0
    abdominal CT bilateral hydroureteronephrosis | 0
    fluid collection at bladder base | 0
    post-renal obstructive nephropathy | 0
    bronchoalveolar lavage grew Coccidioides immitus | 0
    urine culture grew Coccidioides immitus | 0
    Coccidioidal serology reactive IgG and IgM | 0
    complement fixation titer 1:128 | 0
    severe disseminated coccidioidal infection | 0
    intravenous amphotericin B | 0
    CT-guided drainage of prostatic abscess | 0
    drained pus cultured C. immitis | 0
    monitored in ICU | 336
    follow up CT resolution of abscess | 336
    downtrending serum creatinine | 336
    symptomatic improvement | 336
    transferred to medicine wards | 336
    amphotericin B completed | 336
    symptoms resolved | 336
    discharged | 336
    