62 years old | 0
male | 0
uncontrolled diabetes mellitus | 0
septic shock | 0
epigastric pain | -72
shortness of breath | -72
septic | 0
tachypnoeic | 0
tachycardic | 0
hypotensive | 0
temperature spiked to 38 °C | 0
blood sugar was 20 mmol/L | 0
intravenous insulin | 0
bilateral lung base crepitations | 0
abdomen was distended with crepitus | 0
crepitus at the right lumbar region | 0
crepitus extended down to the patient's scrotum | 0
cardiopulmonary resuscitation | 0
intubated | 0
inotropic support | 0
white cell count of 70 | 0
thrombocytopaenia of 14 | 0
C-reactive protein of 248 | 0
deranged renal profile | 0
serum creatinine of 578 | 0
urea of 47.6 | 0
coagulopathy | 0
mild transaminitis | 0
severe metabolic acidosis | 0
absence of the right kidney | 0
gas production in the renal parenchyma | 0
air locules extended from anterior/posterior liver space | 0
air locules extended to retroperitoneum | 0
air locules extended to lateral abdominal muscle | 0
air locules extended to pelvis | 0
air locules extended to scrotum | 0
fluid resuscitation | 0
antibiotic therapy | 0
renal-adjusted antibiotic dosage | 0
IV Meropenem | 0
cultures grew Gram-negative bacilli | 24
Klebsiella pneumonia | 24
image-guided pigtail | 24
placed into the right renal collection | 24
surgical intervention | 504
extraperitoneal approach | 504
nephrectomy | 504
histological diagnosis | 504
acute pyelonephritis | 504
emphysematous pyelonephritis | 504
good clinical recovery | 720
discharged | 720