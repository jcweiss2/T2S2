20 years old | 0
male | 0
schizophrenia | -7200
cannabis use disorder | -7200
social anxiety disorder | -7200
delusional belief | -7200
oral risperidone | -8760
risperidone 2 mg daily | -8760
paliperidone palmitate | -6240
paliperidone palmitate 100 mg monthly | -6240
quetiapine | -4320
quetiapine 1000 mg daily | -4320
weight gain 35 kg | -4320
clozapine | -1560
clozapine 175 mg | -1560
CGI-S score 3 | -780
cannabis use disorder in remission | -780
social activities | -780
weight gain 10 kg | -780
sertraline | -1170
sertraline 100 mg | -1170
muscular pain | -504
CK levels 7499 U/L | -504
low intensity weight training | -504
clozapine dose increase | -504
clozapine 200 mg | -504
benztropine | 0
aggressive fluid therapy | 0
rhabdomyolysis | 0
CK levels 45564 U/L | 72
myocarditis ruled out | 0
NMS ruled out | 0
recreational drug screening negative | 0
discharge | 336
sertraline discontinued | 336
aripiprazole | 336
lorazepam | 336
CGI-S score 6 | 840
visual hallucinations | 840
auditory hallucinations | 840
clozapine rechallenge | 1008
CK levels monitored | 1008
liver enzymes monitored | 1008
CK levels 2218 U/L | 1512
light workout | 1512
CK levels normalized | 1519
weight training | 2016
CK levels 4734 U/L | 2016
CK levels normalized | 2023
clozapine 200 mg daily | 3024
CGI-S score 3 | 3024
planning on resuming school | 3024