58 years old | 0
female | 0
internal haemorrhoids | 0
RBL | 0
osteoporosis | 0
dyslipidemia | 0
depression | 0
pelvic pain | 48
dysuria | 48
empirical intravenous antibiotics | 48
ciprofloxacin | 48
metronidazole | 48
increased WBC count | 48
transfer to referral centre | 72
exploration of surgical site | 72
band removal | 72
superficial abscess drainage | 72
CT scan of abdomen and pelvis | 72
rectosigmoiditis | 72
moderate to severe ascites | 72
exploratory laparoscopy | 96
serous ascites | 96
SIRS | 96
transfer to tertiary care centre | 120
ischaemic colitis | 120
hemodynamic deterioration | 120
respiratory deterioration | 120
ventilator support | 120
ARDS | 120
antibiotics broadened to carbapenem | 120
colonoscopy | 144
superficially necrotic segment in lower rectum | 144
inotropic support | 144
volemic resuscitation | 144
ventilator support | 144
antibiotics | 144
modest improvement | 216
WBC count decrease | 216
repeat abdominopelvic CT scan | 240
circumferential thickening of rectosigmoid colon | 240
state of shock subsided | 240
extubation | 360
transfer to floor | 360
discharge from hospital | 432
recovery from intensive care unit myopathy | 720
recovery from prolonged intubation | 720
intensive rehabilitation | 720
follow-up appointments | 720
muscular weakness | 720
poor exercise tolerance | 720
colonoscopy | 26280
normal colonoscopy | 26280
follow-up with respirologist | 26280
persistent dyspnea | 26280
severe deconditioning | 26280
no residual cardiorespiratory injury | 26280