50 years old | 0
male | 0
admitted to the hospital | 0
cough with phlegm | -168
fever | -96
shortness of breath | -96
sore throat | -168
white sticky phlegm | -168
cold | -168
yellow phlegm | -96
chest tightness | -96
dizziness | -96
no chills | -96
no chest pain | -96
no hemoptysis | -96
no abdominal pain | -96
no diarrhea | -96
emergency treatment | 0
routine blood test | 0
white blood cell count | 0
neutrophil ratio | 0
high-sensitivity C-reactive protein | 0
procalcitonin | 0
interleukin 6 | 0
biochemistry profile | 0
creatinine kinase | 0
lactate dehydrogenase | 0
glutamic oxaloacetic transaminase | 0
glutamic-pyruvic transaminase | 0
emergency chest computed tomography | 0
right lower lung infection | 0
heterogeneous right lobe of the thyroid | 0
black loose stools | 0
increased frequency of urination | 0
urgency | 0
no significant changes in body weight | 0
history of thyroid enlargement | -8760
unknown Chinese medicine | -8760
government employee | 0
market surveillance | 0
denied recent exposure to poultry | 0
family history unremarkable | 0
vital signs | 0
body temperature | 0
pulse | 0
breathing | 0
blood pressure | 0
saturated oxygen in arterial blood | 0
fractional inspired oxygen concentration | 0
alert | 0
collaborated during physical examination | 0
pupils equal | 0
round | 0
reactive to light | 0
enlarged thyroid | 0
pharyngeal swelling | 0
no tonsillar swelling | 0
coarse breath sounds | 0
scattered wet rales | 0
heart rate | 0
normal rhythm | 0
no pathological murmurs | 0
no abdominal tenderness | 0
no rebound tenderness | 0
no edema | 0
sepsis | 0
severe pneumonia | 0
multiple organ dysfunction | 0
respiratory failure | 0
myocardial damage | 0
impaired liver function | 0
gastrointestinal bleeding | 0
enlarged right thyroid | 0
hypokalemia | 0
hyponatremia | 0
hypochloremia | 0
blood gas analysis | 0
platelet count | 0
neutrophil ratio | 0
biochemistry profile | 0
blood urea nitrogen | 0
creatinine | 0
high-sensitivity C-reactive protein | 0
procalcitonin | 0
lactate dehydrogenase | 0
glutamic oxaloacetic transaminase | 0
glutamic-pyruvic transaminase | 0
routine urine test | 0
urinary protein | 0
red blood cell count | 0
coagulation function | 0
hepatitis B surface antigen | 0
syphilis antibody | 0
HIV antibody | 0
hepatitis C antibody | 0
throat swab | 0
influenza virus antigen | 0
bird flu nucleic acid | 0
smears stained for bacteria | 0
smears stained for fungi | 0
smears stained for acid-resistant bacteria | 0
bronchoscopy | 72
sputum smear | 72
multiple blood cultures | 0
urine culture test | 0
Mycoplasma pneumoniae antibody | 0
Streptococcus pneumoniae antigen | 0
galactomannan test | 0
1-3-β-D-dextran test | 0
cryptococcal antigen | 0
blood tuberculosis immunoassay | 0
TORCH panel | 0
rubella virus IgG antibody | 0
cytomegalovirus IgG antibody | 0
toxoplasma IgG | 0
IgM antibody | 0
rubella virus IgM antibody | 0
cytomegalovirus IgM antibody | 0
herpes simplex virus IgM | 0
quantification of blood CMV nucleic acid | 0
fecal occult blood test | 0
chest radiograph | 0
right lung infection | 0
right pleural effusion | 0
endotracheal intubation | 17
mechanical ventilation | 17
imipenem/cilastatin | 17
linezolid | 17
oseltamivir | 17
methylprednisolone | 17
respiratory failure | 48
myocardial damage | 48
impaired liver function | 48
acute renal failure | 48
NGS | 120
C. psittaci | 120
meropenem | 120
doxycycline | 120
ceftazidime | 240
weaned off mechanical ventilation | 264
tracheal intubation removed | 264
oral doxycycline | 264
chest CT | 336
vague patchy shadows | 336
pleural effusion | 336
repeated biochemistry profile | 336
discharged | 504