55 years old | 0
male | 0
admitted to the hospital | 0
weakness | -120
light-headedness | -120
muscle aches | -120
non-productive cough | -120
wheeze | -120
frequent shivering | -120
no shortness of breath | -120
no chest pain | -120
previous evaluation at the ED | -48
discharged from previous ED visit | -48
intravenous hydration | -48
Penicillin V prescription | -48
asthma | 0
hypertension | 0
diet-controlled type 2 diabetes | 0
lisinopril | 0
hydrochlorothiazide | 0
25 pack-year smoking history | 0
quit smoking 16 years ago | 0
syncope | 0
blood pressure 109/87 mmHg | 0
no pulsus paradoxus | 0
heart rate 109 beats per minute | 0
respiratory rate of 24 breaths per minute | 0
temperature of 36.5°C | 0
oxygen saturation 100% on room air | 0
mottling | 0
cyanosis | 0
no jugular venous distension | 0
no lymphadenopathy | 0
clear lungs | 0
no distant cardiac sounds | 0
regular heart rate and rhythm | 0
normal S1/S2 | 0
no heart murmur | 0
unremarkable abdomen and extremities | 0
portable chest radiograph | 0
right upper lobe infiltrate | 0
borderline enlarged cardiac silhouette | 0
electrocardiogram | 0
sinus tachycardia | 0
no tall QRS complex | 0
no electrical alternans | 0
white blood cell count 16.6 103/µL | 0
hemoglobin 13.4 g/dL | 0
sodium 129 mmol/L | 0
potassium 4.2 mmol/L | 0
carbon dioxide 21 mEq/L | 0
creatinine 1.0 mg/dL | 0
glucose 152 mg/dL | 0
cardiac enzymes normal | 0
B-natriuretic peptide 915 pg/mL | 0
lactic acid level 3.8 mmol/L | 0
antibiotics started | 0
fluid resuscitation initiated | 0
three liters of normal saline | 0
no improvement in symptoms | 0
no change in blood pressure | 0
no change in heart rate | 0
no change in dusky mottling | 0
no jugular venous distention after fluid resuscitation | 0
intensivist consulted | 0
bedside ultrasound performed | 0
pericardial effusion | 0
diastolic collapse of the right atrium | 0
diastolic collapse of the right ventricle | 0
normal ejection fraction | 0
subcostal view suboptimal | 0
syncopal episode | 0
bedside pericardiocentesis | 0
200 milliliters of bloody pericardial fluid drained | 0
symptoms improved | 0
cyanosis improved | 0
open pericardiotomy | 12
pericardial window placement | 12
repeat chest radiograph | 12
smaller cardiac silhouette | 12
repeat electrocardiogram | 12
slightly increased voltage of QRS complexes | 12
CT scan | 12
pericardial drainage tube well positioned | 12
trace pericardial effusion | 12
right upper pneumonic infiltrate | 12
small bilateral pleural effusion | 12
pericardial biopsy | 12
pericardial effusion fluid analysis | 12
adenocarcinoma | 12
pulmonary primary source | 12
bronchial brushing and washing | 12
negative blood cultures | 12
negative urine cultures | 12
negative bronchial-alveolar washing cultures | 12
discharged | 24