17 years old | 0
female | 0
admitted to the hospital | 0
sudden deterioration of mental status | 0
disoriented | 0
dizzy | 0
high-grade fever | 0
infective endocarditis | -72
intravenous antibiotics | -72
Staphylococcus aureus | -72
vegetations in mitral valve leaflet | -72
intracranial abscess | 0
mycotic aneurysm of the right cerebral hemisphere | 0
CT scan of the brain | 0
ill-defined hypodense lesion | 0
perilesional edema | 0
peripherally enhancing lesion | 0
intracerebral abscess | 0
ill-defined hyperdense lesion | 0
focal contrast filled out-pouching | 0
conservative treatment | 0
neurosurgical consultation | 24
discharge | 24 
informed consent | 24