67 years old | 0 | 0 | Factual
male | 0 | 0 | Factual
admitted to the hospital | 0 | 0 | Factual
left leg swelling | -72 | 0 | Factual
cactus plant injury | -168 | -168 | Factual
Primary Sclerosing Cholangitis | 0 | 0 | Factual
mild Ulcerative Colitis | 0 | 0 | Factual
deranged liver function tests | 0 | 0 | Factual
progressive left leg swelling | -48 | 0 | Factual
worsening of erythema | -48 | 0 | Factual
pain | -48 | 0 | Factual
felt generally unwell | -48 | 0 | Factual
paramedic assistance | -24 | -24 | Factual
presentation to ED | 0 | 0 | Factual
Blood Pressure (BP): 71/41mmHg | 0 | 0 | Factual
Mean Arterial Pressure (MAP): 48mmHg | 0 | 0 | Factual
Respiratory Rate: 36 breaths per minute | 0 | 0 | Factual
Heart Rate (HR): 125 beats per minute | 0 | 0 | Factual
sinus tachycardia | 0 | 0 | Factual
Temperature: 39°C | 0 | 0 | Factual
Oxygen Saturation: 86% with 0.21 FiO2 | 0 | 0 | Factual
admitted to the intensive care unit (ICU) | 0 | 0 | Factual
pH 7.15 | 0 | 0 | Factual
PO2 84 | 0 | 0 | Factual
HCO3 15 | 0 | 0 | Factual
Lactate 7.6 | 0 | 0 | Factual
Sodium (Na) 134 | 0 | 0 | Factual
Urea 7.6 | 0 | 0 | Factual
Creatinine (sCr) 173 | 0 | 0 | Factual
eGFR 27 | 0 | 0 | Factual
White Cell Count (WCC) 13.8 | 0 | 0 | Factual
C-reactive protein (CRP) 22 | 0 | 0 | Factual
Hemoglobin (Hb) 114 | 0 | 0 | Factual
Platelet (Plt) 81 | 0 | 0 | Factual
Liver Function Test (LFT)- Total Bilirubin (Bili) 99 | 0 | 0 | Factual
Alanine transaminase (ALT) 61 | 0 | 0 | Factual
Aspartate aminotransferase (AST) 83 | 0 | 0 | Factual
Alkaline Phosphatase (ALP) 96 | 0 | 0 | Factual
Triple vasopressor support initiated | 0 | 0 | Factual
Noradrenaline 20mcg/min | 0 | 24 | Factual
Adrenaline 20mcg/min | 0 | 24 | Factual
Vasopressin 0.04units/min | 0 | 24 | Factual
Piperacillin-Tazobactam IV 4.5g | 0 | 0 | Factual
Meropenem IV 2g | 0 | 168 | Factual
Lincomycin IV 600mg | 0 | 168 | Factual
Vancomycin IV 2g | 0 | 120 | Factual
Emergency left lower limb fasciotomy | 0 | 0 | Factual
debridement | 0 | 0 | Factual
below knee amputation | 0 | 0 | Factual
LRINEC Score of 5 | 0 | 0 | Factual
extensive left foot and below knee tissue necrosis | 0 | 0 | Factual
dishwasher fluid | 0 | 0 | Factual
liquefied fat | 0 | 0 | Factual
unviable skin and muscle | 0 | 0 | Factual
Histopathology | 0 | 0 | Factual
oliguria | 24 | 192 | Factual
blood gas showed severe acidosis | 24 | 24 | Factual
left internal jugular vascath insertion | 24 | 24 | Factual
continuous renal replacement therapy (CRRT) | 24 | 192 | Factual
Group B Streptococcus pneumoniae (GBSPn) | 24 | 24 | Factual
Ventilation sedation | 24 | 120 | Factual
Propofol 170mg/hr | 24 | 120 | Factual
Fentanyl 40mcg/hr | 24 | 120 | Factual
CRRT (Day 1) | 24 | 24 | Factual
heparin circuit | 24 | 24 | Factual
Renal dose | 24 | 24 | Factual
Triple vasopressor support continued | 24 | 120 | Factual
Noradrenaline 23mcg/min | 24 | 120 | Factual
Adrenaline 18mcg/min | 24 | 120 | Factual
Vasopressin 0.04units/min | 24 | 120 | Factual
Intravenous Immunoglobin G (IVIgG) therapy | 24 | 24 | Factual
Rapid Atrial Fibrillation (RAF) | 48 | 192 | Factual
HR 110bpm | 48 | 48 | Factual
oliguric | 48 | 192 | Factual
pH 7.40 | 48 | 48 | Factual
Lactate 3.9 | 48 | 48 | Factual
Sodium (Na) 131 | 48 | 48 | Factual
sCr 116 | 48 | 48 | Factual
WCC 26 | 48 | 48 | Factual
CRP 105 | 48 | 48 | Factual
Procalcitonin (PCT) 21.18 μg/L | 48 | 48 | Factual
Hb 83 | 48 | 48 | Factual
Plt 63 | 48 | 48 | Factual
INR 3.1 | 48 | 48 | Factual
Fibrinogen 2.4 | 48 | 48 | Factual
Echocardiography | 48 | 48 | Factual
Moderate segmental left ventricular dysfunction | 48 | 48 | Factual
Ejection Fraction 40-45% | 48 | 48 | Factual
Dilated atria bilaterally | 48 | 48 | Factual
Raised Right Atrial Pressure | 48 | 48 | Factual
Amiodarone loading dose | 48 | 48 | Factual
Amiodarone maintenance dose | 48 | 72 | Factual
CRRT (Day 2) | 48 | 48 | Factual
AN69 anti-inflammatory heparin laden adsorbing filter | 48 | 48 | Factual
Citrate based anticoagulation circuit | 48 | 48 | Factual
Sepsis Induced Coagulopathy (ISTH -SIC criteria) | 72 | 72 | Factual
bedside surgical debridement | 72 | 72 | Factual
pH 7.31 | 72 | 72 | Factual
Lactate 2.4 | 72 | 72 | Factual
Sodium (Na) 135 | 72 | 72 | Factual
sCr 79 | 72 | 72 | Factual
WCC 27 | 72 | 72 | Factual
CRP 127 | 72 | 72 | Factual
Hb 78 | 72 | 72 | Factual
Plt 50 | 72 | 72 | Factual
INR 2.0 | 72 | 72 | Factual
Histopathology consistent with NF | 72 | 72 | Factual
Wound culture for microscopy culture and sensitivity (MCS) | 72 | 72 | Factual
medium growth of GBSPn | 72 | 72 | Factual
Tissue culture (intraoperatively) | 72 | 72 | Factual
medium growth of GBSPn | 72 | 72 | Factual
Vasopressor support - weaning | 72 | 120 | Factual
Noradrenaline 20mcg/min | 72 | 120 | Factual
Adrenaline weaned off | 72 | 72 | Factual
Vasopressin 2.4units/min | 72 | 120 | Factual
oliguric | 96 | 192 | Factual
purpura over the right forearm | 96 | 96 | Factual
multiple weeping skin tears on right upper thigh | 96 | 96 | Factual
RAF HR 130 | 96 | 192 | Factual
pH 7.36 | 96 | 96 | Factual
Lactate 1.5 | 96 | 96 | Factual
Sodium (Na) 130 | 96 | 96 | Factual
sCr 116 | 96 | 96 | Factual
WCC 33 | 96 | 96 | Factual
CRP 103 | 96 | 96 | Factual
PCT 15.37 | 96 | 96 | Factual
Hb 91 | 96 | 96 | Factual
Plt 53 | 96 | 96 | Factual
INR 1.7 | 96 | 96 | Factual
LFT - Bili 131 | 96 | 96 | Factual
AST 127 | 96 | 96 | Factual
ALP 121 | 96 | 96 | Factual
Double inotropic support | 96 | 120 | Factual
Noradrenaline 20mcg/min | 96 | 120 | Factual
Vasopressin 2.4units/min | 96 | 120 | Factual
fulminant hepatic failure/ encephalopathy | 120 | 120 | Factual
refractory oliguria | 120 | 192 | Factual
pH 7.39 | 120 | 120 | Factual
Lactate 1.2 | 120 | 120 | Factual
Sodium (Na) 134 | 120 | 120 | Factual
sCr 124 | 120 | 120 | Factual
WCC 39.5 | 120 | 120 | Factual
CRP 74 | 120 | 120 | Factual
Hb 116 | 120 | 120 | Factual
Plt 49 | 120 | 120 | Factual
INR 1.5 | 120 | 120 | Factual
LFT- Bili 139 | 120 | 120 | Factual
AST 69 | 120 | 120 | Factual
ALT 97 | 120 | 120 | Factual
ALP 140 | 120 | 120 | Factual
Dual inotropic support | 120 | 120 | Factual
Noradrenaline 20mcg/min | 120 | 120 | Factual
Vasopressin weaned off | 120 | 120 | Factual
ICU acquired weakness | 144 | 144 | Factual
unarousable | 144 | 192 | Factual
no response to noxious stimuli | 144 | 192 | Factual
Pressure Support Ventilation | 144 | 192 | Factual
refractory oliguria | 144 | 192 | Factual
pH 7.44 | 144 | 144 | Factual
Lactate 1.1 | 144 | 144 | Factual
WCC 43.5 | 144 | 144 | Factual
CRP 109 | 144 | 144 | Factual
Hb 90 | 144 | 144 | Factual
Plt 57 | 144 | 144 | Factual
INR 1.5 | 144 | 144 | Factual
LFT - Bili 150 | 144 | 144 | Factual
AST 95 | 144 | 144 | Factual
ALP 154 | 144 | 144 | Factual
Sedation weaned off | 144 | 144 | Factual
off vasopressor | 144 | 144 | Factual
Noradrenaline weaned off | 144 | 144 | Factual
Antibiotic de-escalation | 144 | 144 | Factual
Lincomycin and Vancomycin ceased | 144 | 144 | Factual
Meropenem IV 2g TDS continued | 144 | 192 | Factual
CRRT (Day 6) | 144 | 144 | Factual
Hyper-Ammonium Therapy initiated | 144 | 144 | Factual
Rifaximin NGT 550mg BD | 144 | 192 | Factual
Lactulose NGT 20ml TDS | 144 | 192 | Factual
2 units of PRBCs transfusion | 144 | 144 | Factual
jaundice | 168 | 168 | Factual
Hypoactive delirium | 168 | 192 | Factual
deeply sedated | 168 | 192 | Factual
RASS -5 | 168 | 192 | Factual
new onset lateralizing signs to the left | 168 | 168 | Factual
CT Brain | 168 | 168 | Factual
No acute intracranial pathology | 168 | 168 | Factual
Ultrasound abdomen | 168 | 168 | Factual
Acute Calculous Cholecystitis | 168 | 168 | Factual
pH 7.44 | 168 | 168 | Factual
Lactate 1.1 | 168 | 168 | Factual
WCC 44.3 | 168 | 168 | Factual
CRP 109 | 168 | 168 | Factual
Hb 129 | 168 | 168 | Factual
Plt 66 | 168 | 168 | Factual
INR 1.3 | 168 | 168 | Factual
LFT - Bili 235 | 168 | 168 | Factual
AST 75 | 168 | 168 | Factual
ALP 175 | 168 | 168 | Factual
Conjugated Bilirubin 142 | 168 | 168 | Factual
Anuria | 192 | 192 | Factual
Hypotensive BP 71/33 | 192 | 192 | Factual
MAP 51mmHg | 192 | 192 | Factual
Febrile 39°C | 192 | 192 | Factual
RAF HR 160 | 192 | 192 | Factual
palliative care pathway | 192 | 192 | Factual
deceased | 192 | 192 | Factual
Troponin 616 | 192 | 192 | Factual
Ammonia 158 | 192 | 192 | Factual
LFT - Bili 352 | 192 | 192 | Factual
AST 100 | 192 | 192 | Factual
ALP 299 | 192 | 192 | Factual
CRRT (Day 8) | 192 | 192 | Factual
Renal recovery assessment | 192 | 192 | Factual
Furosemide IV 250mg | 192 | 192 | Factual
Acetazolamide IV 500mg | 192 | 192 | Factual
Vasopressor support | 192 | 192 | Factual
Noradrenaline 2.5mcg/min | 192 | 192 | Factual
Lincomycin IV 600mg TDS | 192 | 192 | Factual
Meropenem IV 2g TDS | 192 | 192 | Factual
Digoxin IV 500mcg | 192 | 192 | Factual
Metoprolol IV 15mg | 192 | 192 | Factual