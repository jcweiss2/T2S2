1-year-old | 0
male | 0
10 kg | 0
admitted to Accident and Emergency department | 0
irritable | 0
drowsy | 0
Glasgow Coma Score = 7 | 0
mild right-sided weakness | 0
unequal pupils | 0
right pupil 5+ | 0
left pupil 3+ | 0
no external injuries | 0
intra-osseous needle placed in right tibia | 0
intubated | 0
fentanyl 2 mcg/kg administered | 0
propofol 2 mg/kg administered | 0
rocuronium 0.8 mg/kg administered | 0
hand ventilated | 0
normal end-tidal carbon dioxide | 0
head computed tomography scan conducted | 0
acute right-sided subdural hematoma | 0
significant midline shift | 0
transferred to operating theater | 0
systolic blood pressure 98 mmHg | 0
good pulses | 0
peripheries mottled | 0
pale blue skin | 0
venous access gained through left femoral triple lumen central line | 0
arterial pressure monitoring established | 0
tympanic membrane temperature 36.0°C | 0
received 30 ml/kg of 3% hypertonic saline | -1
hypertonic saline overdose | -1
surgery commenced | 0
anesthesia maintained with O2/N2O and sevoflurane | 0
positive pressure ventilation | 0
passed large volume of urine | 0
Hartmann's solution infused | 0
blood loss moderate | 0
no transfusion required | 0
arterial blood gas recorded | 1
mixed respiratory acidosis | 1
pH 7.08 | 1
PCO2 9.2 KPa | 1
PO2 31.6 KPa | 1
Na+ 154 mmol/L | 1
K+ 3.0 mmol/L | 1
Cl 129 mmol/L | 1
Ca++ 1.36 mmol/L | 1
glucose 14.1 mmol/L | 1
lactate 0.8 mmol/L | 1
hemoglobin 10.0 g/L | 1
base excess 9.8 | 1
highest serum sodium 158 mmol/L | 2
Hb 8.0 g/dl | 2
right fronto-occipital hematoma evacuated | 2
transported to pediatric Intensive Care Unit | 2
ventilated | 2
sedated with midazolam | 2
sedated with morphine | 2
extubated | 4
postoperative fluid intake maintained | 4
good urine output | 4
SaO2 98%–100% | 4
self-ventilating room air | 4
respiratory rate 24–28 bpm | 4
no respiratory distress | 4
heart rate 140/min | 4
blood pressure 112/66 mmHg | 4
pupils equal | 4
pupils reacted to light | 4
awake and alert | 4
electrolytes showed normal Na+ | 24
electrolytes showed lower and normalizing K+ | 24
developed temperature spike to 38.8°C | 24
temperature spike resolved with paracetamol | 24
discharged | 168
follow-up after 1 month | 720