45 years old | 0
male | 0
suspected snake bite on left foot | -48
swelling of left leg | -48
anasarca | -48
pain at bite site | -48
suspected snake bite | -48
non-venomous snake bite | 0
shortness of breath | 0
altered sensorium | 0
inability to speak | 0
weakness of bilateral lower limbs | 0
swelling of left leg (documented on admission) | 0
non-tender left foot | 0
raised temperature at left foot | 0
minimally conscious | 0
reduced alertness | 0
non-cooperative | 0
disoriented | 0
blood pressure 106/60 mmHg | 0
heart rate 102 bpm | 0
respiratory rate 20 breaths/min | 0
body temperature 37.2°C | 0
SpO2 91% | 0
bilateral crepitations on chest | 0
pitting edema over left foot | 0
two rows of teeth marks | 0
no fang marks | 0
hemoglobin 15 g/dl | 0
total leukocyte count 24.37×10^9/L | 0
neutrophils 89% | 0
lymphocytes 6% | 0
platelet count 19,000/mm³ | 0
blood urea 122 mg/dl | 0
serum creatinine 5.01 mg/dl | 0
serum sodium 117 mEq/L | 0
serum potassium 5.1 mEq/L | 0
no deep vein thrombosis | 0
bilateral raised renal cortical echogenicity | 0
normal coagulation profile | 0
prothrombin time 12.7 s | 0
INR 1.03 | 0
serum procalcitonin 0.27 ng/ml | 0
normal left ventricular function | 0
bilateral multiple B lines on lung USG | 0
intubated | 0
admitted to ICU | 0
provisional diagnosis: snake bite with cellulitis | 0
sepsis | 0
AKI | 0
DIC | 0
IV piperacillin/tazobactam started | 0
IV clindamycin started | 0
magnesium sulphate dressing | 0
RDP transfused | 0
CRRT started | 24
IV metoclopramide started | 0
oral calcium polystyrene sulfonate started | 0
IV glucose-insulin drip started | 0
oral pantoprazole started | 0
IV vitamin K started | 0
IV magnesium sulphate started | 0
oral conjugated estrogen started | 0
persistent bilateral chest crepitations | 168
body temperature 37.8-38.9°C | 168
blood glucose 70100 mg/dl | 168
total leukocyte count 31.65×10^9/L (day 7) | 168
Klebsiella pneumoniae infection (transtracheal aspirate) | 192
piperacillin/tazobactam discontinued | 192
clindamycin discontinued | 192
tigecycline started (100 mg LD, 50 mg every 12h) | 192
reduction in swelling | 192
serum procalcitonin fall | 192
body temperature normalized | 192
blood glucose above normal | 192
hypoglycemic episode (47 mg/dl) | 240
severe palpitations | 240
tremors | 240
sweating | 240
25% dextrose administered | 240
blood glucose 83 mg/dl | 240
hypoglycemic episode (49 mg/dl) | 264
hyperventilation | 264
profuse sweating | 264
palpitations | 264
25% dextrose administered | 264
blood glucose 86 mg/dl | 264
hypoglycemic episodes (days 11 and 13) | 264 and 312
tigecycline stopped | 360
IV meropenem started | 360
IV clindamycin restarted | 360
IV polymyxin B started | 360
blood glucose below or lower end of normal | 360
CRRT stopped | 456
serum creatinine normal | 456
serum urea normal | 456
electrolytes normal | 456
sepsis recurrence | 648
Enterobacter spp. infection (transtracheal aspirate) | 696
meropenem discontinued | 696
polymyxin B discontinued | 696
tigecycline restarted (100 mg LD, 50 mg every 12h) | 696
hypoglycemic episodes (25 mg/dl) | 720, 744, 768
50% dextrose administered | 720, 744, 768
tigecycline discontinued (second time) | 744
oral minocycline started | 744
IV cefoperazone/sulbactam started | 744
blood glucose low or slightly below normal | 744
gradual improvement | 744
discharged from ICU | 912
transferred to general ward | 912
