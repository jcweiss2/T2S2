81 years old | 0
male | 0
admitted to the hospital | 0
lower abdominal pain | -72
bloody diarrhea | -72
abdominal computed tomography | -72
thickness of the descending colon wall | -72
intravenous hydration | -72
antibiotic therapy | -72
cefotiam | -72
levofloxacin | -72
diagnosis of ischemic colitis | -72
follow-up abdominal computed tomography | -48
ascites | -48
thickness of the entire colon wall | -48
renal dysfunction | -24
convulsion | -24
transferred to our hospital | 0
slightly clouded consciousness | 0
temperature 38.0°C | 0
blood pressure 140/92 mm Hg | 0
heart rate 95/min | 0
skin cold and moist | 0
abdomen distended and tympanic | 0
generalized tenderness | 0
severe inflammation | 0
anemia | 0
low platelet count | 0
renal dysfunction | 0
hypoxemia | 0
metabolic acidosis | 0
low CO2 level | 0
tachypnea | 0
colonoscopy | 0
diffuse mucosal edema | 0
ulcer formation | 0
bleeding from the rectum to the ascending colon | 0
no evidence of free air | 0
whole colon wall markedly thickened | 0
huge ascites | 0
vital signs deteriorated | 12
blood pressure 60/40 mm Hg | 12
heart rate 115/min | 12
severe disturbance of consciousness | 12
generalized cyanosis | 12
diagnosed as having necrotic ischemic colitis | 12
septic shock | 12
emergency surgery | 12
operative findings | 12
large amount of ascites | 12
colon wall markedly edematous and sclerotic | 12
inflammation of the transverse colon extended to the greater omentum with necrosis | 12
extended right hemicolectomy | 12
ileostomy | 12
resected specimen showed hemorrhagic necrosis of the transverse colon | 12
pathological findings | 12
mucosal hemorrhagic necrosis | 12
submucosal edema | 12
venous dilatation | 12
congestion of blood | 12
ischemic colitis | 12
stool culture | 12
O157 | 12
verotoxin | 12
diagnosed as hemorrhagic colitis | 12
HUS | 12
acute encephalopathy | 12
O157 infection | 12
treated in the intensive care unit | 12
ventilation | 12
delayed emergence from anesthesia | 12
encephalopathy | 12
poor oxygenation | 12
intensive care | 12
HUS improved | 120
encephalopathy improved | 120
without dialysis | 120
discharged | 768