84 years old | 0
female | 0
admitted to the hospital | 0
hip joint endoprosthesis | 0
increased bleeding | 0
postoperative anemia | 0
hemodynamic instability | 0
received packed red blood cells | 0
fever | 312
antibiosis with piperacillin-tazobactam | 312
diarrhea | 336
septic shock | 432
circulatory failure | 432
lactic acidosis | 432
blood smear | 432
high concentration of plasmodia | 432
rapid test positive for Plasmodium falciparum | 432
artesunate | 432
ventilation | 456
hemodynamic support | 456
death | 480
no travel history | 0
plasmodia transmitted by packed red blood cells | 480
look back process | 480
donor traveled to endemic area | -720
donor contracted malaria | -720
donor did not mention recent return from endemic area | -336
donor did not give information on malaria prophylaxis | -336
donor released to donate whole blood | -336
donor had general symptoms of illness and fever | -168
donor did not report symptoms | -168
donor diagnosed with malaria | 0
donor took malaria prophylaxis | -720
negligent manslaughter | 480
donor sentenced to criminal fine | 720
donor sued for damages | 720
donor convicted under civil law | 720
donor must pay bereavement compensation and funeral expenses | 720