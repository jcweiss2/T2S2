3-year-old girl | 0
fever | 0
respiratory distress | 0
admitted to intensive care unit | 0
no known disease | 0
secondary parental consanguinity | 0
sibling died from fever | -24
cousin died | -24
upper respiratory tract infection | 0
ampicillin-sulbactam | 0
azithromycin | 0
COVID-19 PCR negative | 0
poor general status | 0
low consciousness level | 0
confusion | 0
blood pressure 170/78 mmHg | 0
heart rate 110/min | 0
body temperature 39°C | 0
SpO2 88% | 0
weight 13 kg | 0
height 104 cm | 0
crackles in both lungs | 0
left lung crackles | 0
normoactive deep tendon reflexes | 0
normal light reflex | 0
COVID PCR positive | 168
hydroxychloroquine | 168
favipiravir | 168
increased respiratory distress | 72
deep respiratory acidosis | 72
pH 6.96 | 72
pCO2 91 mmHg | 72
HCO3 22 mEq/l | 72
intubated | 72
SIMV-PC ventilation | 72
hemoglobin 6.5 g/dl | 72
white blood cell count 16,160/mm3 | 72
platelet count 503,000/mm3 | 72
blood urea nitrogen 44 mg/dl | 72
creatinine 0.8 mg/dl | 72
AST 65 U/l | 72
ALT 57 U/l | 72
total bilirubin 0.68 mg/dl | 72
sedimentation rate 60 mm/hour | 72
D-dimer 5820 µg/l | 72
bilateral pleural effusion | 0
atelectasis | 0
consolidation areas | 72
ground glass opacities | 72
persistent fever | 72
teicoplanin | 72
cefotaxime | 72
decreased urine output | 96
amlodipine | 96
hypertension | 96
refractory hypertension | 96
enalapril | 96
esmolol infusion | 96
furosemide infusion | 96
albumin transfusion | 96
peripheral blood smear | 72
clustered platelets | 72
anisocytosis | 72
microcytosis | 72
hypochromia | 72
polychromatic young lymphocytes | 72
bone marrow aspiration | 72
LDH 1162 U/l | 72
ferritin 1512 ng/ml | 72
D-Dimer 7840 ng/ml | 72
triglyceride 247 | 72
normocellular bone marrow | 72
no dyserythropoiesis | 72
no dysplasia | 72
no storage cells | 72
no hemophagocytosis | 72
normal renal size | 72
normal renal echogenicity | 72
normal renal vasculature | 72
left ventricular hypertrophy | 72
mitral insufficiency | 72
azithromycin stopped | 120
meropenem | 120
IVIG 1 g/kg | 168
repeated erythrocyte transfusions | 168
anuria | 240
progressive thrombocytopenia | 240
microangiopathic hemolytic anemia | 240
creatinine 1.9 mg/dl | 240
undetectable haptoglobin | 240
reticulocytosis 8% | 240
LDH 2540 U/l | 240
negative direct Coombs test | 240
schistocytes | 240
HUS diagnosis | 240
normal ADAMTS-13 | 240
ruled out DIC | 240
TMA triggered by COVID-19 | 240
aHUS type | 240
fresh frozen plasma | 240
hemodialysis | 240
extubated | 336
urine output 0.9 cc/kg/hour | 360
LDH decrease | 360
blood pressure reduction | 360
platelet count rise | 360
esmolol discontinued | 360
oral antihypertensive continued | 360
asymptomatic | 672
hemodynamic normalization | 672
Hg 11.6 g/dl | 672
platelet 192,000/µl | 672
CRP 3 mg/l | 672
creatinine 0.6 mg/dl | 672
LDH 230 U/l | 672
D-Dimer 140 ng/ml | 672
discharged | 672
oral antihypertensive discontinued | 1008
no genetic mutations | 672
sequel pleuroparenchymal shrinkages | 672
ground glass densities | 672
regression of findings | 672
