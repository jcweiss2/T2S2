30 years old | 0
female | 0
admitted to private nursing home | -192
severe pain in abdomen | -192
fever | -192
giddiness | -192
gaping of episiotomy wound | -192
resuturing of episiotomy wound | -192
evaluation for fever | -192
platelet count of 50,000/cumm | -192
worsening fever | -168
breathlessness | -168
hypotensive | -168
conservative management | -168
shifted to hospital | -168
severely tachypneic | 0
severe hypotension | 0
inotropic supports | 0
intubated | 0
mechanically ventilated | 0
platelet count of 40,000/cumm | 0
deranged liver function tests | 0
creatinine of 4.1 mg/dl | 0
coagulopathy | 0
international normalized ratio of 4.3 | 0
bilateral chest infiltrates | 0
arterial blood gas showed a PaO2/FiO2 of <100 | 0
severe ARDS | 0
ultrasonography abdomen and pelvis | 0
two-dimensional echocardiography | 0
provisional diagnosis of acute febrile illness | 0
severe sepsis | 0
septic shock | 0
polymerase chain reaction for leptospira | 0
dengue IgM | 0
malaria smear | 0
IgM antibodies for hantavirus | 0
falling platelet count | 24
coagulopathy | 24
blood component transfusion | 24
severe ARDS | 24
lung protective ventilation | 24
renal dysfunction | 24
renal replacement therapy | 24
septic shock | 24
broad-spectrum antibiotics | 24
inotropic support | 24
progressively worsening chest X-ray | 48
alveolar hemorrhage | 48
worsening lung function | 48
ribavirin | 48
expired | 240
multiorgan dysfunction | 240