87 years old | 0
male | 0
admitted to the hospital | 0
atrial fibrillation | -720
heart failure with preserved ejection fraction | -720
hypertension | -720
dabigatran etexilate 150 mg orally twice-daily | -720
weakness | 0
decreased oral intake | 0
mild cough | 0
increased lower extremity edema | -168
atrial fibrillation with rapid ventricular response | -168
serum creatinine 1.20 mg/dL | -168
eGFR 57 mL/min/1.73 m2 | -168
verapamil 120 mg daily | -168
metoprolol 25 mg daily | -168
furosemide 40 mg daily | -168
verapamil 240 mg daily | -48
metoprolol 100 mg daily | -48
furosemide 60 mg daily | -48
fell while getting out of bed | -48
vomited three times | 0
axillary temperature 95.7 °F | 0
blood pressure 102/48 mmHg | 0
ventricular rate 36 beats/min | 0
oxygen saturation 96% | 0
jugular venous distension | 0
hepatojugular reflux | 0
bibasilar crackles | 0
bradycardic, irregular rhythm | 0
systolic murmur | 0
3+ pitting edema | 0
IV normal saline 2 L | 0
IV glucagon 1 mg | 0
chest X-ray | 0
right lower lobe infiltrate | 0
ceftriaxone | 0
levofloxacin | 0
acute renal failure | 0
hepatic dysfunction | 0
septic shock | 0
pneumonia | 0
electrolyte disturbances | 0
elevated serum lactate | 0
coagulopathy | 0
IV insulin 10 units | 0
IV dextrose 50 g | 0
IV calcium gluconate 2 g | 0
IV sodium bicarbonate 50 mEq | 0
computed tomography of head, neck, and cervical spine | 0
no acute hemorrhage or fracture | 0
FFP 2 units | 0
vitamin K 5 mg orally | 0
Profilnine 5,020 IU | 24
FFP 2 units | 24
vitamin K 10 mg IV | 24
unfractionated heparin infusion | 120
warfarin | 168
discharged | 456
PT 54.4 s | 0
PTT 100.6 s | 0
INR 6.0 | 0
fibrinogen 279 mg/dL | 0
diluted TT 125.0 s | 24
diluted TT 113.1 s | 26
ALT 546 U/L | 0
AST 422 U/L | 0
alkaline phosphatase 111 U/L | 0
total bilirubin 1.4 mg/dL | 0
direct bilirubin 0.5 mg/dL | 0
CK 170 U/L | 0
CKMB 5.9 ng/mL | 0
troponin T 0.08 ng/mL | 0
NT-proBNP 3,695 pg/mL | 0
white blood cell count 18.52 K/μL | 0
hemoglobin 14.0 g/dL | 0
hematocrit 43.5% | 0
platelet count 214 K/μL | 0
coagulopathy correction | 24
renal function improvement | 120
hepatic function improvement | 120
INR 1.8 | 120
PTT 46.9 s | 120
warfarin therapy | 168
discharge | 456