72 years old | 0
    woman | 0
    treated diabetes | 0
    hypertension | 0
    hyperlipidemia | 0
    candidiasis | -432
    HIV-1 diagnosis | -432
    CD4+ T-lymphocyte count 32 cells/μL | -432
    VL 16,600 copies/mL | -432
    ART initiation with ABC, 3TC, RAL | -432
    CD4 cell count recovery to 265 cells/μL | -288
    VL controlled below detection limit | -288
    abdominal pain | -360
    vomiting | -360
    decreased level of consciousness | -360
    emergency transport | -360
    blood pressure 102/58 mmHg | -360
    tachycardia | -360
    labored polypnea | -360
    Glasgow Coma Scale score 13 | -360
    metabolic acidosis (pH 7.0) | -360
    hyperlactacidemia 199 mg/dL | -360
    abdominal CT showing gas in mesenteric and portal veins | -360
    intramural emphysema of the colon | -360
    diagnosis of intestinal ischemia | -360
    ART suspension | -360
    emergency laparotomy | -360
    jejunum to colon necrosis | -360
    mesentery normal blood flow | -360
    NOMI diagnosis | -360
    subtotal small bowel resection | -360
    jejunostomy | -360
    preserved 70 cm jejunum | -360
    preserved 95 cm small intestine | -360
    complete large intestine resection | -360
    lactic acidosis resolution | 0
    CD4 cell count 163 cells/μL | 504
    VL 49,600 copies/mL | 504
    HIV-1 subtype B identification | 504
    no drug-resistant mutations | 504
    R5 tropism | 504
    single-dose ARV administration tests | 504
    DRV 400 mg | 504
    RTV 100 mg | 504
    LPV 400 mg | 504
    ETR 100 mg | 504
    MVC 150 mg | 504
    RAL 400 mg | 504
    omeprazole co-administration | 504
    Cmax LPV <0.01 μg/mL | 504
    Cmax RTV <0.01 μg/mL | 504
    MVC Cmax 0.580 μg/mL at 2 hours | 504
    RAL Cmax 0.566 μg/mL at 2 hours | 504
    DRV Cmax 2.18 μg/mL at 3 hours | 504
    ETR Cmax 2.09 μg/mL at 3 hours | 504
    ART resumption with DRV, RTV, ETR, MVC | 600
    MVC Cmin 0.45 μg/mL | 600
    DRV Cmin 1.72 μg/mL | 600
    ETR Cmin <0.01 μg/mL | 600
    3TC addition | 600
    tube feeding initiation | 672
    Cmin MVC 0.128 μg/mL | 672
    Cmax DRV 1.1 μg/mL | 672
    DRV Cmin <0.01 μg/mL | 672
    ETR discontinuation | 672
    RTV discontinuation | 672
    ART dose interval adjustments | 672
    VL decrease to 32 copies/mL | 2016
    sepsis development | 2568
    catheter-related bloodstream infection | 2568
    death | 2568
    