10-year-old| 0
    male | 0
    admitted to the hospital | 0
    born by cesarean section at 38 weeks gestation | -984
    weight 3200 g | -984
    length 52 cm | -984
    APGAR score 9-9 | -984
    perioral cyanosis | -984
    neonatal sepsis | -984
    patent ductus arteriosus | -984
    newborn screening normal | -984
    discharged after 11 days | -984
    recurrent pulmonary infections | -984
    multiple hospital admissions | -984
    severe gastroesophageal reflux | -984
    breast milk intolerance | -984
    Nissen fundoplication | -936
    gastrostomy | -936
    atonic seizures | -936
    childhood spasms | -936
    valproic acid | -936
    Fanconi syndrome | -936
    oxcarbazepine | -936
    severe hyponatremia | -936
    phenobarbital | -936
    phenytoin | -936
    atomoxetine | -936
    aripiprazole | -936
    quetiapine fumarate | -936
    haloperidol | -936
    sertraline | -936
    pregabalin | -936
    olanzapine | -936
    topiramate | -936
    levetiracetam | -936
    mirtazapine | -936
    ethyl loflazepate | -936
    lacosamide | 0
    clobazam | 0
    brivaracetam | 0
    acetazolamide | 0
    hypokalemia | 0
    potassium supplementation | 0
    weight below third percentile | 0
    height below third percentile | 0
    head circumference below third percentile | 0
    subclinical hypothyroidism | 0
    selective immunodeficiency of IgG and IgA | 0
    nephrocalcinosis | 0
    microcephaly | 0
    elongated eyelid fissures | 0
    eversion of the outer third of the lower eyelid | 0
    arched eyebrows | 0
    broad eyebrows | 0
    depressed nasal tip | 0
    short columella | 0
    small teeth | 0
    spaced teeth | 0
    micrognathia | 0
    large cup-shaped ears | 0
    low implantation of ears | 0
    bilateral retroauricular pits | 0
    polydactyly of the right hand | 0
    polydactyly of the left foot | 0
    bilateral palmar aberrant folds | 0
    sacral dimple | 0
    Kabuki syndrome | 0
    KMT2D gene sequencing ruled out | 0
    exome sequencing | 0
    homozygous variant OTUD6B c.433C>T | 0
    pathogenic variant | 0
    weight 24 kg | 0
    height 1.24 m | 0
    delayed head support | 0
    delayed sitting with support | 0
    no gait development | 0
    emits sounds | 0
    obeys simple commands | 0
    solid foods orally | 0
    liquids by gastrostomy | 0
    levothyroxine | 0
    gamma globulin | 0
    insulin resistance | 0
    allergic colitis | 0
    facial features | 0
    hand features | 0
    severe intellectual disability | 0
    seizures | 0
    dysmorphic features | 0
    craniofacial dysmorphism | 0
    recurrent respiratory infections | 0
    chronic constipation | 0
    congenital heart disease | 0
    hypothyroidism | 0
    hypogammaglobulinemia | 0
    allergic colitis | 0
    insulin resistance | 0
    abnormal corpus callosum | 0
    mTOR pathway involvement | 0
    difficult to control seizures | 0
    severe mental retardation | 0
    genetic panel including Kabuki syndrome | 0
    genetic panel including Rubinstein-Taybi syndrome | 0
    genetic panel including DiGeorge syndrome | 0
    diagnostic odyssey shortened | 0
    adverse reactions to medications | 0
    irritability | 0
    insomnia | 0
    tremors | 0
    hallucinations | 0
    seizures decreased to 5 events/month | 0
    discharge after initial admission | 24
    patient's current age | 120
    <|eot_id|>
    