62 years old | 0
male | 0
referred to the critical care medicine department | 0
sever acute pancreatitis | -192
respiratory distress | -48
heart rate was 122/min | 0
blood pressure was 114/66 mm of Hg | 0
respiratory rate was 32/min | 0
abdomen was distended and tense | 0
bowel sounds were absent | 0
Hb 10.2 gm/dl | 0
total leukocyte count 17,900 cell/cmm | 0
serum creatinine 1.9 mg/dl | 0
serum amylase of 2897 U/l | 0
chronic cough since childhood | -62400
endotracheal intubation | 0
mechanical ventilation | 0
invasive hemodynamic monitoring | 0
intra abdominal pressure (IAP) was high (24 mm of Hg) | 0
nasogastric tube was kept on free drainage | 0
decrease in IAP (17 mm of Hg) | 72
nasogastric feeding was started | 72
severe cough with feed visible in the endotracheal tube | 72
endotracheal tube was upsized to size 9.0 mm with cuff | 72
thorough tracheal toileting was done | 72
nasogastric tube was kept on free drainage | 72
recurrent distention of nasogastric drainage bag with air | 72
gastric content in the respiratory tract | 72
communication between respiratory tract and esophagus | 72
bed side bronchoscopy | 72
gastric contents regurgitating into the right main bronchus | 72
diagnosis of right broncho-esophageal fistula (BEF) | 72
aspiration | 72
septic shock | 72
sever acute respiratory distress syndrome (ARDS) | 72
high ventilator and vasopressor support | 72
bilateral lungs infiltrate with predominant involvement of right lungs | 72
death | 120
right broncho-esophageal fistula (BEF) | -62400 
congenital BEF | -62400 
severe acute pancreatitis | -192 
massive aspiration | 72 
raised IAP | 0 
nasogastric feed | 72 
massive aspiration through the BEF | 72 
increase in the mean airway pressure | 72 
air to leak from tracheal to esophageal lumen | 72 
repeated filling of the nasogastric drainage bag with air | 72 
conventional barium esophagography | 0 
surgical closure | 0 
severe hemodynamic instability | 72 
high ventilator support | 72 
recurrent cough since childhood | -62400 
early diagnosis | 0 
management | 0 
prevention of life threatening complications | 0