75 years old | 0
    male | 0
    presented with painful right scrotal swelling | -48
    scrotal swelling | -48
    pain (right scrotal) | -48
    scrotal pain increased gradually over 2 days | -48
    fever | -48
    rigor | -48
    history of diabetes mellitus | 0
    medications for diabetes | 0
    dietary modifications for diabetes | 0
    pulse rate 110 beats/minute | 0
    blood pressure 100/60 mmHg | 0
    temperature 39° Celsius | 0
    central abdominal tenderness | 0
    suprapubic tenderness | 0
    scrotal redness | 0
    scrotal tenderness | 0
    increased scrotal temperature | 0
    clinical findings consistent with epididymo-orchitis | 0
    elevated white blood cells count (20000 cells per microliter) | 0
    neutrophils predominant | 0
    scrotal ultrasound showed normal testis | 0
    thick fluid collection around the testis | 0
    diagnosis of infective process | 0
    received parenteral antibiotics | 0
    little improvement | 0
    developed anorexia | 96
    developed nausea | 96
    developed severe abdominal pain | 96
    developed backache | 96
    fever (recurrence) | 96
    rigor (recurrence) | 96
    abdominal tenderness | 96
    abdominal guarding | 96
    abdominal X-ray showed mild bilateral pleural effusions | 96
    abdominal X-ray showed dilated loops of the small bowel | 96
    abdominal ultrasound showed fluid collection at the pelvic cavity | 96
    normal serum amylase | 96
    normal serum lipase | 96
    CT scan showed large amount of air in retroperitoneal space | 96
    CT scan showed displacement of right kidney toward midline | 96
    CT scan showed air extending to the right scrotum | 96
    CT scan with oral contrast showed tracking to retroperitoneum | 96
    CT scan with oral contrast showed extension to right scrotum | 96
    laparotomy done through midline abdominal incision | 96
    thin pus in peritoneal cavity | 96
    air collection in retroperitoneal space | 96
    fluid collection in retroperitoneal space | 96
    initial intraoperative evaluation of small bowel showed no abnormality | 96
    initial intraoperative evaluation of large bowel showed no abnormality | 96
    lesser sac opened | 96
    posterior wall of the stomach intact | 96
    mobilization of the duodenum | 96
    perforation in posterior wall of the duodenum | 96
    suturing of perforation | 96
    peritoneal cavity washed with warm normal saline | 96
    2 drains left in abdomen | 96
    admitted to intensive care unit | 96
    clinical condition improved | 96
    drains removed on 5th day | 168
    developed complete abdominal dehiscence | 192
    developed right scrotal abscess | 192
    another surgery done | 192
    abdomen closed with tension sutures | 192
    drainage of scrotal abscess | 192
    general clinical situation improved | 240
    discharged after 10 days | 240
    tension sutures removed after 3 weeks | 672
    improvement of clinical studies | 672
    improvement of imaging studies | 672