50 years old | 0
male | 0
admitted to the hospital | 0
distortion of the oral commissure | -72
dizziness | -72
headache | -72
malaise | -72
vomiting | -72
shallow nasolabial sulcus on the left side | -72
weakness in closing the left eye | -72
diagnosis of acute upper respiratory tract infection | -72
diagnosis of peripheral facial neuritis | -72
tuberculosis | -14016
cured tuberculosis | -14016
no immunodeficiency | 0
no major trauma | 0
no toxic exposure | 0
no smoking | 0
no alcoholism | 0
no drug abuse | 0
no hereditary disease | 0
no unpasteurized buttermilk consumption | 0
blood pressure 135/85 mmHg | 0
temperature 36.5°C | 0
pulse rate 85 bpm | 0
increased white blood cell count | 0
increased fasting blood glucose level | 0
increased glycosylated hemoglobin level | 0
normal serum creatinine level | 0
normal cholesterol level | 0
normal C-reactive protein level | 0
normal creatine kinase level | 0
normal procalcitonin level | 0
normal blood coagulation parameters | 0
negative test for human immunodeficiency virus | 0
negative test for Treponema pallidum | 0
emergency head CT showed no apparent abnormalities | 0
chest CT showed chronic-appearing fibrotic streaks in both lungs | 0
dexamethasone administration | 0
head CT re-examination showed no apparent abnormality | 72
headache | 72
dysdipsia | 72
malaise | 72
fever | 72
neck stiffness | 72
slowness of the pharyngeal reflex | 72
peripheral facial paralysis | 72
somnolence | 96
aphagia | 96
slurred speech | 96
brain MRI showed multiple abnormal foci in the brainstem | 96
increased cerebrospinal fluid opening pressure | 96
increased white blood cell count in cerebrospinal fluid | 96
biochemical cerebrospinal fluid examination showed increased potassium concentration | 96
biochemical cerebrospinal fluid examination showed increased chloride concentration | 96
biochemical cerebrospinal fluid examination showed decreased glucose concentration | 96
biochemical cerebrospinal fluid examination showed increased microprotein concentration | 96
negative Gram staining | 96
negative India ink staining | 96
negative acid-fast staining | 96
transfer to intensive care unit | 96
physical cooling using an ice blanket and ice cap | 96
anti-infective and antiviral medications | 96
intracranial decompression using mannitol | 96
symptomatic and supportive treatment | 96
negative test for influenza A and B viral antigens | 120
negative test for anti-Toxoplasma antibodies | 120
isolation of L. monocytogenes from blood culture | 120
identification of L. monocytogenes by time-of-flight mass spectrometry | 120
genetic identification of cerebrospinal fluid pathogens by high-throughput genome sequencing | 120
respiratory failure | 144
mechanical ventilation | 144
administration of ampicillin, amikacin, and meropenem | 144
transfer from intensive care unit to standard medical ward | 144
ability to walk and eat normally | 2880
central respiratory insufficiency | 2880
intermittent mechanical ventilation | 2880
satisfaction with treatment and recovery | 2880