32 years old | 0
    male | 0
    sudden onset shortness of breath | 0
    syncope | 0
    seizure | 0
    chest pain | 0
    flu-like symptoms | -72
    developmental delay | 0
    sedentary house-bound lifestyle | 0
    hypertension | 0
    tachycardia (110 b.p.m.) | 0
    hypotension (90/52 mmHg) | 0
    hypoxia (oxygen saturation 92% on room air) | 0
    clear chest auscultation | 0
    normal heart sounds | 0
    T wave inversions in leads II, III, aVF | 0
    dilated right ventricle | 0
    mobile thrombus in right atrium | 0
    mobile thrombus in right ventricle | 0
    thrombus passing through PFO into left atrium | 0
    elevated urea (10.6 mmol/L) | 0
    elevated creatinine (144 μmol/L) | 0
    high haemoglobin (168 g/L) | 0
    high haematocrit (55.9%) | 0
    elevated lactate (2 mmol/L) | 0
    elevated D-Dimer (3.84 μg/mL) | 0
    elevated troponin (2.28 μg/L) | 0
    haemodynamic instability | 0
    emergency pulmonary embolectomy | 0
    extensive clot in right atrium | 0
    extensive clot in right ventricle | 0
    clot passing through PFO to left atrium | 0
    D-shaped septum | 0
    fresh clots in pulmonary tree | 0
    fresh clots in right atrium | 0
    fresh clots in left atrium | 0
    fresh clots in right ventricle | 0
    severe tricuspid valve regurgitation | 0
    clot removal | 0
    PFO closure with bovine pericardial patch | 0
    tricuspid valve annuloplasty | 0
    epinephrine infusion | 0
    severe right ventricular dysfunction | 0
    ECMO initiation | 0
    weaned off cardiopulmonary bypass | 0
    full ECMO support | 0
    continuous venovenous haemodiafiltration | 0
    intravenous sildenafil | 0
    weaned off ECMO | 144
    sepsis | 192
    acute kidney injury | 192
    critical illness neuropathy | 192
    percutaneous tracheostomy | 480
    weaned from ventilator | 672
    IV heparin anticoagulation | 0
    warfarin anticoagulation | 192
    oral tildenafil | 192
    haematemesis | 672
    traumatic ulcer clipped | 672
    tracheostomy decannulation | 888
    discharged home | 1032
    complete recovery of functional status | 2016
    normalization of ventricular function | 2016
    no evidence of acute brain ischemia | 0
    no predisposing factors for PE | 0
    no evidence of Bechet’s disease | 0
    no evidence of underlying malignancy | 0
    negative antinuclear antibodies | 0
    negative factor V Leiden mutation | 0
    negative anticardiolipin antibodies | 0
    negative double-stranded DNA antibodies | 0
    negative beta-2 glycoprotein-1 antibodies | 0
    clear chest CT scan | 0
    clear bronchoscopy cytology | 0
    <|eot_id|>
    